`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PzeNb3leAkgZimhqkyozRRAgbJiPXymdEE1jNp1q5XDVmD4HXpOX1L3u1cAQ25oF
MpV1Kezp9HfZ70i9jJ0K3XMf6k08JI8mXDlOadbBb0MuIb2g2X98+NSqzGET3Ex7
9SI4/cjAz9lDzs0lXYi31yjU6VDzWULaj6I3RVJhZu19q5VUwI2kiG6qf4Lb4kjG
11zgunFEO91w17UzIl8fqk7J0yuxDhVv9bfrvK3bhp3Ll0NyjmK9QTEVbRQNtjm7
tEwtnMbX46cEBJCoFAUnOw/bcv5U3WOVNF7WChAkMEgckTq+bjk58wh9E5QzFyhk
IXpB1wI+ZPIhdvrL1Z+rBJgsUQt9VmiZR8gRhZNe6qjUKkbM+BlHxcEpvToAGdRv
yqmISik+gqZPDTDEKHlAtoHFEz70gwoH+50ltLtX0xCBEUpJXYkkq+nGqvbiGI52
ZWAlDcowbj7tQCSQUXnOs0+TiTsbRm5q9LeQMm1DVaZR6LRGWLNtkpVZDZE1BOUl
PosDfgOJHLdi8VswVj3WEhbpiDnMlqcRiTKR67eCD7GlgeMG3PWpV9Yt33ZZFu24
3ojfCcSTG6IvWcjeYp8aIsWX7LVWEZlRY6d4zI0z6yoqbvzCz3Q8uFz4+qnDxOqY
VWxaMiyqw3gSVeojupQJbH/oAWzQqi24+NSRY8aoSvbsuoC25N6aFYFlcwObWQvJ
y2PsMOMXgZyVV0hjVo9LkYbh/OzhL6MdL/JT99SMDUFgcIweglBk5q+VgC8+CvQX
MlnOxzkv0KDxVQ9m38WJYKuPXu/NTcb13BU3zhPDVBfPZ4Vd3Ea73nHXKqlnAPwZ
qHdpKJZi2EQbxTwXq75U0/PA950yU+Ga6krz59Htx0ilQWQtuKAemdLChETbCIxX
CCUW3lMrzwuIXcQeZRLC8uOPtP1VyuHnDLhZKzv6YfY+cWuO2W170kAZo7RtpQUU
4t2epAeV8/Hm5TsmEiH/lFeYrHVqX59bKMl3tvXEftMseJhPc4Yhj28yWejbNkfS
B5mFxIdYPHSraAbN3GfAaNwm8cZ2u8KBTqFQHfROBkVAi38tWBDOxMpNDMi8jplo
y9tRphi4epTWuvM2n8OSyeZtC3fmqfhhb3fqq3N6eijfctB3GgEOfL5HZt9b2AhX
JuZYoxUt+DYdlgXzGxx3CNoilMXv+W5KeP9/IXCZYBsN6mLm9s9We7XKU8Pqagbl
lt+av8XoEV9nvnutJyd//+q4+hgvvQvMI1Xx713/iwzt3gB/CAb8QFR6bwvt5RBG
wq0Agj/Hj/bJtxGZdQBWTckIhl5NzsmkvDXjhY/OybNMfIJZP9nUUdD/oBPHlSSC
RknOhtm3zZa5z0KIRJWQu5lVjug2W1kAc1FEgNJgWNkHYf+QKYTXUkC5+2kUux3l
cxPEnuBkOImPewZDDl9k/4yjKR11CiL2pGQ2gSWPkA2nyWl0lpM6hzMTk3V6KgpW
ifSiG7Twf/QH24cTlUsWPBNCMxvDyeqvdiMSqR0uTSo9+U89IULaki+RsNGJa6DB
xrhcTsVAewKZ2mJovdJBv4kPqfbPJmx5RpbqcyDCHb3erwhuo6pFzXYMfRg80Fnw
TSAbh+oT/i+EDP6v1wwO09x0RvuHrqaGkc56aX6f8ZLcv+jchre5NgLQVY7MPpjt
bpucu9DQeoKxVdgyW9BoIv0MVRa2IQSOcJ6TwL1PYUAqqQZ4z7nL7PZMm4jsSFmT
7fUBkKW/wH1yiK/arLZqFTsi7EPEgW8rI0x9pk3UyEtGviVy92ZilMkHkjFIzszK
4uQrpWy1cp2wjiQ8DNmMG9srTec2ENHlB9iWa9vT3gaLIxYpFjLL8+t9v0WmCoUU
CgHvRAQVeClkL7H6Z8mWq/N1CYtag31FyUXFC5anI9xlZmSZXqDV1owep8kamjkc
iLaygav0VrWW3NaFROivEYENHgyef4tGJzGIMGtDILJioY6UZJRWsU1qCyXvSPDD
3OPixEugzKQn3TA88Mnckk+3oxVbEVWLLafVaGkuZF8//QOjB0C7nEtl2rDeATbr
ZyhinfCbfP1FQVWzohnhELvvsPzK0jxh47tidFmTGVvfMZzzIUu7G0QYPd+uLBXa
TtEiURdHyP2WkuWlx+nmFIk3IiaV9InviJ+5nGB1F4qJ2xy+OxU6PtQloHncugWZ
OC0sUq0w27YSWabmPa5UOwlC1VlquvxE2BNbDL9doBFu6tf24HoUZ+hTS6ioe0j+
jqsBOH6mHpweZih7lSFQLn5mf715R0w8Kf7LuNsZsh/oOjYVMfycdjPdhfQ97iiM
noixIXNQnPFnCyCUToEfiBX8I0yo9yrFmr/EFk5yJzI3nYAKMDo/nR5IJdfgscfq
7rEj6MiaDC5aJaNByquvLtLzTTveK0ZRThSxx1LGsr1Mj3ciFHbAMx1u6lDvfTrV
Pnco7XU5cln009UUd62VthUTn9r4Mf64ZryW4uxJSvqPV5iNrkePbxUxw6CivNO+
0Sl+K6/lsRtXWGCmHYeCVLJ5dI2iyMCGS2vE6R47Dlp3xf+PDSgoY7VdZfbRf4VE
UcQyyDzAX0LdZdlgQFYDyiP0klKLc+qmy3Pj9MMq19w3Cszs3VGf15Gq5GGEsDsW
vYtiz8Jpbh+qz5p9ieejy0n4Kx5uhS/Aa5seduA9wFqMU7h0SppC53tNwkF+Ql63
4QUwr6DHP3ZQ9xE7ll3P0Rc+u1Nj+FeK3YFxM10X9oGuCt+uUpmQmXIUg7ESprcc
8bckinuRDk8blACsa9wrDzikEYiwQ5ERQH2iYxp1GMh/RwPd44dJlof4DeR8diNs
dsJVNxMkNuZNSuryQ+7boK3d3Ix6WXJsRKrHBEZNRVPwxvcAS6w1BWzqx7zNSipJ
auKVZ6sK+scUYSbppfZzlF6G7qllY0H7dQYpS8ZqmMCVdvRbey8nQUAX311LR9mM
grU/Zx+XiqoNtTs5eLP4OvH+MOQJI1l7mW3VAy7rK+wCm+2/CZz9kO8d/ImO9b9m
rlDbWVFJuzmwmuAg6km44i8n5RTqfPkUzXMy1rWP2QlsO4WtnCuRib3PGlNNYH/L
+W1MGtI3xCwOpAMU/03/l92oSX50TwwmPjXs4Utom3CEQrbIq6akB8mmw6doTwaL
V01Zs3WBpbT4g4M2snptxxwGIF7rU2cV8kAW9FzYLOJm1w8+jsis2XO7Gai1iHNl
a7X6AvsyYIxUT6XeS//AzNkueG2EBYPuTuu+XxldMmjtw4FfkWm7Bd2LEDxodymN
xF66+huQl7lXu653l+G77CeNHSNc1HGohdICJ+ifOHl+b2OU+ZmhtmbrUfbpMNR2
Pg0c8MRGFj2m3nU8NjoBNCSz3G4LChHxxgUBZPFILtgEtgdUpKJvnUcToAyV+YQx
ZYtKoOnYYBsP4r9mblfQc5/fy0i/KOKdeISk01FxYOSkgKBby4XCrrKm6AkQA1i+
A0T3hzodvMXTmIBsTLRd6i3tPuaaaiJwhRRY8NIOs6mWgxtgLN5Ltj8MnHSiWmrc
gKmFJKDdDezsASMDkkiCQfU5MwLOnNR2rOiG02tvPsHa7nSUAsNvQ96cOa3Z3G+F
UuCNnq9EWAOBmH0nTE7R5Z5WAT3Kk1exk/P6lA1n0QdL+Kyp1+N0xhHxJcgMu1Aj
kjfyX/nWqXfB3UKxniMW49tJln29gMFEXGUSZT1hzNmxxGc19gJ+hl8lldxwihXB
NuIwVhwkFsQVcQsbp9BTDA4HXSExfwu5wd3nXcfj8LfIc0fOJLYlIojFecIiU1jS
ZGcKgrO0JArJRCMgtJTC2qaW/kRCX4SyDB00sXCSNtopLrj2nxDxNdACvLQkz/Od
8rnfyKR4HaVq04kCLxJ5K2hVRw57p87a1tMMf7xtXV4w0DSRUt5vq/M9Q8O39+1k
pYl+oZZiKc5X6BDG0pltSGOH0NemgXWBnsxzxrVT3Zzcp+LCX15PMrX4AtHV/JwV
eunOW9GOHoihxz9qqSAc65/W8tNqyeVWQGsk8TEJ/hU3j+1CrdIGjkvGLrSIbs+0
0Cw2LqLHujRc0IRrIhvMVXf7qDMcejb57NM33k6wuRvYBQeJXn8AHiKbRbjFCExL
ji/FSfo1uoHie3Xizy6sDhlLBHTh+8AWUtmvj22kOv5Yc9RDxO4e3r3SpwrKm+Su
aDuhJaxCKzZZ/pttgti1KRWmiESX2GizhN1vfQlyZ6lbBh3NZVPaTZg8aZd/IRWn
FI1q3E4y2hFkc4AVq0b4AgTGALw38Bwep3ShhshXmV+AWx5GPCho6qzIoyRV0w3+
e0N8LEBLG9CegLYANIfpZNVN2o7v4bKz056ndn5PUV/1anlRZTfMUJ9N/cTHkSch
rqJ6JM6BjsYu8tU2Lm5QHUiLQ98/XMdKgeR/zbBTqN8n4Ugr7A/EVZnP4FK/mLIU
lNhKY9o+yHdS1o/liFEPbBuTcjBZS2INKk+DPBx8Fanfk177CBGrG3nGBV3yOFTH
YQ4U0+Gr7nbxcPKJNXuI1MxkVQzHU36LLe+5K6q5x/BX44aRHII9wZPe7a2OeqoH
iFfovLhU6O7/EtrNCGQkVx5cSOkVa4s15+r7WKvoLD0APRqXzWocY2j0oXhNX2/D
1szx3zfUayCAAk8qefw2d0fGwdkINpA4kZvXgNbS0i3GJzjNer1PGhjGjq6nLHu+
GcwrGX8YCE4eprWTNphb1SAW5h8RMYP23YmpOclP1LAZ4gv46dMoIBop8+IKGvaw
IHIncKfK8OAVgx+3bZFkiZusvkVBPgsinjx+ThOHEnTsbXq9eeh1W05BCBx8+cNE
QhnVjnm+61zDZ8EmizgsQkeAwPtDJ2Ap66MTlutPoIR+UPjZCjJUcaxAwxk2Qdyv
DLkMmHtRY9HeZxcyjmDIjVDGQ1AjBAOj1NRVs0fL8GuZ1NYUyNKKaTcYdn0kBiOt
NjDeZogRrbWFQUF4mkbeVFvK2hYhWhiljkasfjoZ5IEYu6YVmW+Yyl/L1jlj5wHt
3OnVmFNiL9qlJen8e2TxR6BYTujLsOnB7gsipZNOhD02Iut+sGDEuPg6/wWhcCY5
vD45t7ADLbZJmGF1sGqhNglZUbO7C1B/PW9NSssMzN0NapNwOxxwnpvCGGw0HCld
BkMmZ//1tycFQu+hfExaNpFgmdsqHR5zoWnbiiBM66+mX99JQB0d+Qm3NTrUEXuF
m8FDQUkYkgCbr0Q6JXlUfihqQQ/lyS2PHASqEM+pP1SIaN0o85VggIhszGX97dj+
ZxNlfmm2VGy2WaZBp7NTLK8SFiezqQGBA4oC9K5opftnm8Pr2BZLR5gyHlbhCcLT
m9OOaoCvXLAc8076xA7tSY9IuNbkEfUTKBYdBkuwNIrBkw+XGYIvDXIFm423SSoI
MCKLUfTcH9wV9j/wG+OEnqK9c+1n/4SeLu66VIHdF/nXux+XvTbEa3JqDSTaoXCI
lD/AxgYuG//ss6BNfO05LZuZbf9FPKUR9xu23a0EtYzPOOIFUJufty9uN9juMV+/
O34acKtdBWRgxjpuM9V9Chmh3QAj51J2TiJ/qnK84MWKlwFlOV44HChnsyDaUurN
ecN5njmrudVGk4/vfD6sSxIXF8jK5TPyaOrQ0Ix8yhoroMalSnvYPl6UC3nO/Hmr
KvtyyLyWHLm5j56FY+F/c5keyveAV7lPQoV58U5kRY4HPvHVAPxbdRho+X+i6XED
YzrkOU11Q8TcsgFYAfrI8AP34e+DE8W2++N0cB1P7bSA4FUixi6oIvhsYwmyaHtu
fPiNeBpednVw6AcCBV6XV7Tf+oAuNIg8E+YNSwsTcp33m2+mIEhMkozT5HS0gWy5
WB1/S0J6iKU6DqM2I4I61pU8XR9j47n4LTqbA0Zn/zlFt7BHw8phY7b2AmNm7JxY
Z9ndfvFLnv9MHY2NWNz+wLloQvqfRJq2uIHwTC74dm5wPWmWBMqx5K8My86uMuhz
9nzrGK+pRv8m9ED0Eqy66uEEY6scEjMErOn9WEXU+YMD0hBgjmDUD09s3sWOoWls
6ahYI0ohXU6b3t+rHeE7lQOCVUuCP0RMY3QdnQorSt53tvmwoUnanWvLxWCvkDgQ
ll+PJ//7NeW/Fm4b/wYIRaDZIhiCMzTFmYOgapM3KA08BfT9OTlO0MFbagzzKyf2
uPJM9SfnoB77xWIaIO1uIg+6O6TiLeGM3yulC5t1uBCZm2MIcBzQtPgnZGzt6GKQ
0ek6kDPFbJrES0DUfRf+GOmMUt9YwRgqcSS3hHlUbTUvj9nck3QzZAGyeWm6A9+k
gH8Efw/Tet2XRhnOuAOna1/alNHdWL+vHKeshzERN0fGD2sohHYykII1raCdJnbb
uHiRdL92jc6PI0oMkvmm2fEfB9165Jmd+Y+iEfUNURmYMOH+DsN5gMJ/qcWYN/DM
oNFu/Wqk3L7Fp6MZXku/ciJpnIJ8yiaqc4C063UKA7JJwzJodmqhhj3O4Uu+pz4m
R06gHkY2C1VwH9jWYdKEddRNnYi7kIb4tGzOI6dhg9AklYk1oeepYrBvLqQE7wrJ
BBsLX32aK5Emhqje9J416bzQLYccbbGgUzRPe7atLFZUWErxX7bOML/pl4FfF7Ks
fdAhuYF3OvsDIqeUcBXu47H/tyeQF+ruczxD6O3CRf6wZYfZwzGEyoxxhf+NvzUF
JIm16mN04bRMH11XcxOiZDeJAgLqL/ocJIOHTXzWVvHbe8lr3jlKTWc2KDzJDOrr
u9wcgT0tLWy4O44cH6L5D5pccilCiTk5u1/ya8O1ezjvscKS3LNjo3vC/pAxxNVL
XyzLBIz+ARAvZA4TXAnra3rR33a497aP2E4oHIrgoZDV5r1LDgK87KxuaIkcpirW
q03HLghWcyKZY/RUOhV5r/UOVVOagNs12pPbKLqIoOBny5H67i4R4lT7B6/X9HqB
v4sbUZW4shawJS/mpTenA7L7PFjyPcwuI1NSnZ5/t2NuGntOa//UuKdq/prfqq4N
lyHVRCn5sK8l5pUIf9YhJTqzn234iaQ13hTNpsHHmX/6MdefMaJfUj2qLR/HGpUp
jQwn22lLUSE8zRsl4E9A7/84gYyLQz71AdxOCh0plmIDHPmJptd8z9mSZYW9ez5E
i9EFjR/r2MVJMvzLBZ3dJ8KHuu5jGBu4CbpzF1tFq5butbyR9CKcbkePojbcs5DK
M4HTDBQ8Kg5EOS1kxb9TH5+CNQKaaKF5U5SZ0/q+sTOOImFnsjld0I2A/ZUvzFYf
UFPNFWF/PPRfW1ObZkstUvzwK+Ql9DXHIi/bBajoHyYlRSiiFpIJbupUMbjL7Ful
UPNwxscEVwVr2MMG8oMS+A/xRpNAcG4EhcTsOlSh1PBvpkVO06sIpxXgo7nGJbaA
tPzxO9IrlXQSRbbFtMiSimwvcGfvADvdYRy1zSS86sFId5/aYczXm7w1VaSIiom2
r2W1L/UN2gYXAZ20eXmeVeUq3bzRxNsThXFezH4H4oPL5y4fuNsvXSOplcHVkSo+
xEAW1Sp/O5rMPzMizh2wAq81XWcFUafQF3qkXEtHHFK3QcPOFqhjFz1xA4qNDQ6J
VXqrjZxaDf89VMT/x8bbH25bVlo9O2ZCnfIqbfuRZNJCt9zq70W+gw3qgy7lPld7
T1AYPDy1+fwU7A4KJaOboBiCYvw488QGzVUUYzpcVi0J+SOgPoKcFxOg2eFyNUnQ
hKK9lLuQQu6i5LIP9WRc2eRNFON5tSCLUfwwg/VZ0f4qBWPC52goqAUPsQ7goTdw
jXGq0sLf7W+5QgqvEcW/PJLzHfuQnGyTCKcK3+vkukywNA+kBK2xUfMHKp+wxswH
Vv+kws3+dtxFb5Viw7bRsrynhDjV3AJvc82nNTCPHHqREYtZfecDmM7Hs3biSKDZ
M1rBqb4t0KxSHb8BX3EuPHSZl9F9KxVN4FAaYUlASV2i6fSrOx8qERw2wVQv9CnE
9kmLfIjSF7F9IUDkXQhzl94Xb61E8S+JYmoDV+spEU5npT23F4RKzl/IxXYcirJz
tZgClxXqHQChdGAP6yIY+JQ7bheeVFFbXX13Jf67B53HWYK9FDb4U3bLYrnpAfwx
Nfd8zev+XjvH1qqD9vQl6TpuSElYNKXGPcVH3Jt0jcJSZ2aZAK+N5+PQYLEDbL1F
d5+3qLUXZsq5YaFLrTWsYUj8/03anb4pkylfDsZNXlZUXGlAQxw0PVoG8uwPjtPL
0gHjOPV6dSNstDHJwKMmYW55KiaYCsiQ4YHdZUVnUAAk0/BQznWFxy+Wx9MUuyjC
aZNCcZydpeKOobT5+VMqyxSUfwDW7/f/ePGTEJOreQJUstQqy+VabrO2itR9NyFq
ypE3WLPcfkIBE2q0EwrA+wQCpkxeR/oB4U9hK+LOCxnYmVHWxKlzXoIIc3x74utc
VVQneV8kEn5jmLbAgjm6b7FppJMHOGQxWOlJAhQJn10W9y30xM/1RL10naWC+ueG
HuRy2Scnp6Z0OD+VIPkfvidQz2HTc9piXk+4T6t/gAIs+OKsXgadcJcssucxGRbM
v6o7tlG9/mKh8n0owui3CzccjSk+EDLGP0nV2rQlwOSf58Ltmeg7DHAcB5jnUJqA
BPnF7zfyNm5a3UltkLd0HNMarbuPNhs0dVu6gaVL9ppb0UYJdV9FFnXKjzDEF7ez
C8pN3AELk6ZdH1W2gvvu7ndhdAkff2ED6PydX8ObJJA2YVIKyzow1O4TWTZxSvZm
OA5wHxm1+IL2ZRKU1jczCocFFCfPD62FrbXJVE06iXWWfkTW37cN7QhAepgAkbVB
I3IAugW2xSQU8yFpy3K1UYpS8Q6+Fb8nY3PW7s01UsX0EcOJl5asO+v3lfLpFb6r
QrqBujofWx9TsuLVW03u7zSro6sFNBhrrnxGFuaBGNMhVic52ufEZ4It8wWSc5xL
puUbMQNV6TUm3Cyv8X1UaF30JmOiFT30KJJDR5/a6YmCIlF1dGdJPhewXyxh57uB
hYIC0OZCiricodiYzucIuLvKfX4M36bSpaFBurb+vTIE6yBJpVELo7iuNJEdEd8l
9xzh/iN6sgW8I5NS5MWrDXmGz/TkycvqTxtRb/WpNaBfClRO20wLCuzKSbqK491W
SHD8hF5QfNF9k33HqD9sB4LpZV7/dPRIb/RX/uwgtfznNJ+7zGypL1Vzn/mdguzF
sP80/J0Viwl3KeJIVmmJHXVEO17rRn8QrCn1scVsVwaXrmhgtbEVsx27fo4FwlKz
JTr/sh3+SK9sr6SPhQDciMGz4tFe4k3me0Ui+ocMUX+02KuOz9qZ2OjKbqBVGWY5
ZnYWrrE011KjIUMppwo1oRKOthbmGgaacvdQkuiUKbAb0qsQRqk7Z6ec0SJEPj1Q
/uA+hcZ94CWwZ0mp388CHuDtmJAumI3iVkjd4QFfpCvVUWSKvIlB45ZS1bU1cvY8
ePFjtFXqSjAGCgN2E6gpxY6uVdBI8/rREKxBgm0GdgHNQMHmK+yAEzxd9DT+Ha+F
V4aRdFPNlUCmxOVh9Fo8g4eYVkJpjBr9OVMHztd3duw1ONSD7j8sZbdYGaRW7gZy
2ftTLVyZB6Xfuhy2XEej0HeqqQHtQb3GUMO5YgCWJgZxtM6+bhAQZIf06iGQwjHZ
oz6CVO+0wqytGZ7hEEhhwrNcJF1EoqUGIuyCX9jBwPVgtrTMIkmQ+LfOMrPcu/7V
zaiiAptBD8POiub3hDjPGFXjAYAIv0PALe2+vrf1yrQQT/nnxG2hZ6P1mly1bGsQ
UyaC0UNxJb4/KkwNIC5lZA/zNOVRnnoEpdLAMSiYhQiXyX1V64QdStzq9qoG+Wxg
qEyGgNRXC/HEMJVvkpBnIpvPx7D16gCnenp5arBWFQP/4yJD+gVvK7WZVJDB9EBC
ZQvADFZJIVIYZRDobPvdcH32wLgeYFCWZnycVV/5SkK482S9MZFxwDluRj0DfPUw
BaAz3jEO0zpVL5d705QXfAELffo7/qheky+VWTjfHAJI8pQtoEtoiZ1SHcwqHpG1
AcdENTvXny4bAbKhJhQdYu8XZGg76O4wNYDfv8eeIhirAx6nzt2YjRQyAKJPXgYk
wyU3o/YEj/JFVPuNyKpwW27rW7rDDxKH+P/i4JGyHYz+uVdqkT9/il866sArpmJA
FUUqxQoPH3c1vu3CpmJRbDGfBKABm8LCAmZaHWLk15iB9GFtdW4RePrPAJZdnU39
pzL2Ug8kwTWorUXaaTNexDyVushfYuJv0aEKBdvVOkJSmnmcB6R4726w9LoSyRnw
srxrIGppyhBJZz/Gci978QHylhrEZPrUmFoV1pY5fXgqGyq1KhQfUi1x4+zOok7x
4I9dXJEiyI1lujHYSrW9RxASV647AOyRaZtFkjhwVlt6mwXXcC3OfyDn/mya2kJB
710am8yOFy66n23EUIFR68jeFkFc1upa94rj/TnisZcuUDaKDLhRcT1XI5Y6cAp4
Igjmw3d6dEW5UL8mlg27LP98IxIyqKr61wDVUNnQtcnlfcwCd/r2vGntE4erjHa/
odAF6CGsOWh6nAmJyaEIT/0UVqFDIIguhmeXR796mlChvvnGxxiEMaiCQEaK21hL
yLnKKvMCJ7i/CrRaLVFDOhX9ku9OYJvG+eOUK6kBUnzfHl2+3Qe9zQHSa9BzXPXJ
uDaKS96P/tQuhhGzQGMUGlY4GF0F4VIUTfnJ6jXd0p2A30LXfucgF5NhtS3gBftW
bq9QO3Ve3vA4CzNIN6XTwZR9SimB3otozuc2R7o7o0Mmi2vE+EyAulq4G3t50jS2
OzlG75nAYL4SPhtW0p/CmGZF6rbt5naaZid9/ubMl5TPv5/UY5tCRs9lUoDjn4Lj
S90xaSHXcgNVRXzotf+kgwl0M17aaalnZG2iz+75eC5J8upFv0E6S6rZ//dL8Mnl
Uk2Jj5pO9CWcbpWRZA83ZkxeN8iy6zP0jT2/zHTQE/eXDdhJWOLxBNtPGHmZgUcR
HMGEKAQdUCc2phhvz19rEC5qeDHpv/4xdobLozRgdEuKlGp1Q0pjGRAyk4UusTFU
wkV3EEhWXgnFg/fidSJs8e7mT0i+OnX4VYF5F9ILmdZfFcKHmc2SQOK3S7QBjCuA
fcz7JtMLddnSZIBwl46lYO83nb+qjcvf5epLrKuBYjF7r8ILAHTCN+LtgPfo4yXq
ZNWXEyytb4qbNhrBhXPxD3Or1rnpS6/btssa9bZvzTJxxD4bqn73FNR0vYi8gyb/
CCkiDJ/VDfqdJKI5zkubhEKn9JISR6OAWkoSZIE9WrjRGQ/4xWRIFwAO45omASfw
WPJQFKJIu2AN43qXG1vZADa111/7ILXG4sQ+eLVbkKP1amUyxZqplHRnBt+KKX9p
+DVQO2XkRlRNOauB2sGH8DZsB3Dy1NDgpB1OJmC7ntPSuBfZr8+CBpp7VUFgxTuI
hUf6dGudMh4PRa20Exm1mKeyX9WfaRpfev9AAWr5/BZk2iaSrY2Gog05tgV8Rq32
Q/qYXyYBWiN25RjBXxBGzMk/g3JWC5bW0hVsAEwQf+BGLuFzC8szNNHbGC5/NS+c
HhJsM3pnBfCguzsccYnqZQ6mTiwto8O/ExwrdRv37gccWJI/QtSY2pBXyg26wZek
ph2e/LQiqmCqzs6F4CA/7nV8JS1cvjbBvBU9QVN2jNStvL1my7U59sk82PheVjZ3
ZteYRLobUf6KFf7U+KroG8qzlKGAlp+3qK+IO8rESyCs2eB5OriCYqGkzJIgOsYL
f2xKFgWGPKuOR05tHtOUH5Vfd1KRPR27SgvSLFgwOilVl262fM/9ltcu+dOTWQw8
8tk0A72syujmm06CRcuCDTTSlfApkb3E3lLxuzG5MxQCRikefdOZJI13FFU8WJB8
dm7bdnWlUaQfrSG7jVd+rivrT9Rm7cJPXkigbj7IcM2yU0BuRaJT1aPRgMvUS0rG
pI22GeE38674Lgn08Xr4VLFC8LkFli4ZvGODF2Eun+/WQJtpUMEXS7rgsBBgXaYS
+4tSByMKcPx478XXrK49jt4pI/O/v/uTI6HkEdxwUwDxRrLDNVcaowO1/eyawvZ9
z8o68NCBh+9I6pTqWf33uCtjK4HOOLIi/A59h65gVivv8AiM4zL5QfGe9SJ2ZLHE
KoioxRsL3Q4hx4lhJXu/IWWxD139WbJrMHNYCKcrFeIT3HZFHZYGZznD85Dl0O9s
pXK2kMZh3RZrEpF4y3XbUw2wheXTZ6GYXzuKwpk3tKrLcJjGqw9onUUAUKTUUfi3
AkXevw7GwoD/ZmZPP+MW/f1gZvxS/yxXAXfKpQsc92VDXMiOs7czTMC0BFcDjv2+
8/pWRPySgjlewrwmb7BS3qKW5h2QUidUNTvsH9OYpI4YLqr+2z69rSKb+TfkcSJt
LcZ26H0S9PzcQRGjxSoeAlIuI3jHkeCNnkZNCZBw6u42FG7KABa3UmDa7IaF/QDH
fo3GampjZTFuCBsTCzPo48Lzhda2h5Y+tCwrlg4yI0HEzaeiTriheO3u6F113PmM
TjtcoGEzvotxeT8l6avdfNET2CRm/PyY2NRIxD9o9kBNB+aT7RI+CA5pzxVrxCAi
2i+7oY7Ez6zWMZF+g+cRreOUmZAewjmBd6ZI4FE3/OX2LUFJum4NRbN14QyScbSh
vCfJe4aFrNwKDljBJfk4ujfVslQsTnVLNgt4XclcGkbM6gViBrm2Y5oV0znguKZQ
+FPsHShlvUxaBZ6BX28C78eZbrOwyjzGWfZXw3bhf9Xlvk3Y3kuXKfL0chMjgjCo
9TtM/tIz6rwXoSfyIA2XXqjIMyuZwqRDb3m/WiatP49nVfW86tUiw2qRM7x8CeD5
6UKCuILtqztXpwecCL/4nScr+YqsKd5LkDSFiqveCXBjEExybkMItn+m778gpspG
cqkf+CDXyaCLIReiRbqBwHGbnJBFbqVToKh9EobdyVjIdRUeiH2R1Z8yJxzrXi8X
IVxkrYu0QJ7/GqLvKcCDMbk5Y7KYuzsvmO9jIiI1KsflHcURNRuJ3yEs3UEyGAxp
VF2X7x7nib1StsEfAPROOyLCZn67B079TiOMM4qYa5+0IoSRsT+7jCJj7a9M1mD0
JoDHO37VHVuatNNm2ouq9oM7Idr/ZeOUJQRPrN+Lar8wpivYxskdekZyFSEyJgkO
xifhLXjTVuSYgR+Zgda+PqTeXfK5qTUQ5h7BK7aPpyRfRQMoeTkIaLkCNcjiEbaf
MbiIIkpQYCbBAMn73OqBozid0WYynhLQFhBwzmMkZjuFex6czGLLbS+AJ9Rp+aX+
oa6hGc+uyQQW6S7Br8RWq7YeQDD0dPyBIU31sZu6VtkUK1TGQ/nMUO7hJ06cO+B1
h0zq/8MCYZ3pg4Coqk5dvBN0KSNpqb/Hh7iWv1ocY+A0j5wswzBiQWVEh6w+p2GR
lKGspXP09pKK+yAJoiWvTNKXfoHLiIRRrmAmfO711znnCKqfNXjnH9km4S6Eq77v
zqMNFpJ9D23xuLMQ9B4HADyhGGvVb4FnHQsBxT2ITjg4ruFbC+a3jIYgSAgUy1rD
2SFTxirJaripK4V7YvlrPgtCzh2rq2vyKCO/SNocHLLdGoOryCoqtfURWrzqkgxB
P4O3hBn9PXnZ7EV12ipnYnVa78lruYmqvvPy7BnbxQZuSEETTvqIoUmJUsgLz38i
wyGkYLOdiyfpYdZYuikWX/bYrUBqAjezLMGU32bO0gSkREhJpm8i/RmC2TBCUyBQ
B1Io4EuwqjSi2Pi4nF7W/DvsRoqV9wgO9NlJieuWUuGOt7hwDknSbIU1jr6VClOg
lIHn5sxm3mQxYkGyR45mPUQxF6ZP+egnqS9EizJd8uukcVuLR0iP5yeu3YMueSEF
38S1DZ3HaV6uMQNHE0sEnhEXEIoS025uY1zhGBI9ZK35Xx7P/wdRxSvTcIh3XEej
PRaS9TgEeIruXHRiRy0lAlRyctzwp267GCIRP0WFhws1t6sX2xVVrk9OOYiKA3SF
UJoUvOONHaFWBl0YSch6peEFshKvdONJmmEEo+cxzBieMjmPMb2UzCahIBo8vfUb
/iqVy/j8ZQpjf4D8scJiQgIniDHw/nMXFbUQdtfEA3YftSCzJVHjG8cH5MJUFn2k
LgNXoh2EnO+xOpuBzO+dRhZO2CcMrxx5CnW95xXrTBjqaocsksh8VVpT4jFz/M2r
Jl5W83LnQ6/bDZs3nasygU11zOQB2zNoEMQvlDqnMKIEgXnjxNJV9GGkoMtY/9+Q
bJl+azHsW7VyQ3iRkqPL0fo1+S9aYbMUhsJ+ACrz6oN6xE95gOuOzyrm7S8VYj0x
UVcvc8oD8m/jtPDqj0hF8Dvc7Fj4acTQcHXzfMzsfYYYDmVxlfJhlVFmON03Eq5l
ccYMpi4lVeOBGuzqjeC9aaGYywWJntdV8hpec2R7XvLJYrnMyVUcj28Bd0//ukfp
MyVSANKIj7/zeJKXA+ucZInqG+83U+jv7rjakqfGdCnHh0QCGgdCYqKAMXyZHCmo
BBHYuMjLIveQBFFPzH7N7JekAn7rEOT5fFF6VZgM11UIEfUyjhXjcbelg7sDGpuY
7eWcSLNL1tGm2HpLjCU8R9+KhPdaQTAePEdJ9SyqPawoBqekT8hCV4MSNNtXfmEK
r9OiZiSKs5vNgn910ErxVvzpsAwThOT2TcH2caMS1zsxHeV39SklTm1LTVE9EB16
+Tg0zibCiObjqtdyE1UK/zgK+5uDZ6N6HsS07xOH0sV39Y0XPiLBX/ATz9XCEEED
q4ybsPfe4Mh8vvv/+7dpAAM68eXafcTVHxnBWFAB1eL1t2CCf82352Qy3dDLisrb
sRC1kO1g3Zu9p06eEDsE5nIdkIFiRbAH+f+7Mv8cYhkWgU/3n0GthWbH7V7a7tOt
gH+Uq3q8+5srKLVYSU3rH298VuRrFih7CmhKm1vgEhGVNXCy5rB05Ol2m9SA080v
365gn5BpuPPJSDaUZ08GMOA4X/IuOGaFahiEF1haB8t4JV+PxzxDAI/VfoS79EYK
y6lcP5Q95283Zk67twot81tyEliDhxh3786TdVnXFLGhohYX3SEDAbh3li9dcXDC
kzlZVnVQB1y/dRjOIqG0cbtEfP3xCSzE4j1DTcIOeQuvAKu6qSkzCwmx4t3P3Pyp
XAxtUEmGq9v6hHlOkmKoWYr2fEnFCPPJHa6M5LbD4nVU5zZpQ9IpAB0lKkW2GgKJ
kOXp+9oYlhBnKxWIGwzmwow6fUoa2u4PWH76rEt6iTgYqs8UfidqneOIX97zescE
+6NLKCm71wWrBCNGssRv9qvSXuwh4SmJOaa0L3aH/wdtsmUi36tS+dVPLCPVVpH5
Ea+HuD7Nt1HjsNW/6EvtcXOm1R/j2yov6QVpEgdG+0U9yXa4/sGeWoq6BI+Svkax
XeJhFwyrdV50lEYYOVYhdLRJ27a3h5h6D/oOOaP0LRDruUuAYo0dJKq0v57/ioAv
VSjY3QfSmbIPpcbBQcz0QpWWFEwU2tF7YW7nvit1+VCHJ2aKzyOoQAjUXBzNTRya
YSxlNgEAClKuP2jZuBXCUoQLOjKgeHKFh+DD2ot+A4S13A/jOREMv3YRlk6PmR6F
85/MToU+elSauiMJj6ZYq3Yh3bnsp85rovpcSVcesiuuon8oD2FFhGdwHkaY1E6i
Oa0wEfnxTf4SKawOVgLoag3mKKJSYFt+itTH7/Pd+RDtAPISSbxAHuj2F9nOGzJk
Yhc+Wr9YySEKsjtgcjhCdFT5W+sMznvNCPUXVhdRAMfJz3vTz/0+VSl4g4m1wyt2
+rdZoWWlL/wkeZN/KBkc7abl4iDTNTJgEd6ZKngyioaccOmhXkbgTLcl4IEGM6X3
4/4ZcME2goKkvXjRyUlQNcyJ8D/p22y33bWusD51BBXL6x1idUsRBLLK0TyG9Qbj
wsRhb+vnqIPC5xlZdHS/T/UilwWC0N6E6LXiUXxUD3DC21tvWLVQ6C5RGOfvPD2h
I6EvI1aynsEQkNvax4zC/mi0vALYgq2i+Scb+C+RnC6qDGvWyiU5n1cUFnvywnrX
ofbY7Pwxig5vjH11tr2cOdsAozy5C35DBODFPOLeWEL6PkmJha06c/YkpQEyu4eL
rXG2mJJWywQj9e3H3cZBSPh/vp4il8D+FEK6LhnexDXHQL2mDA2+U7giQDAkfKi6
lnPtZd9N8Rfc30DJk3ofCtcs0PebCxXkBrLbcPGCqdbLlu3eVfVbJNFZO/vrtMMJ
2KJO9x7QpKkarrApdfl1KnQ/d21F8MShUK87b578nZi7oPWMwjLpA6jy58fanslX
67t2rcKWbwfsazICpQFZByY6NLJADN4iN45KfJ0itrHPm4f+mSbPifY7BhrHiiDR
F2QEfP8jfAHO3iXSj3k1n/zd0kOmbhO+3uMDeHnw5BBbM5z/w6VsUd+/Wrrlc0yG
R01s/jUjCTx+CL0Dh2T3WS7tTLfIvuEyrC44WKh6cN51tVEpHmUr0835Kz3PHrJs
FPh2Fhnoo9k5COn7yFOCQ/XldoaUHhij7CQQCzVMsKOdftfAFW+hgvB8jm9gSza8
OBZfPv+Uofd3PWf6LBZXX+IQd67aXHnxDM9dO7doxmrTDj9WL4NisLRjJtThKlcv
qxIDjPX+Re7siN6t95Ak9etr2fRJAV7H6epJCsEQfgCG6lFkkDZNH33R7ouq9WSk
IYwPpMOmL3GOJ7ZZWEkacNRdVQmNokje83O9kvQJeg8tppMgFFOn9ewM48sdvU1n
b6Pem0h/olF/L5vvnsgwsFctqe0ddNgmcO1I+UkUdlR6Y/U7pFb0Q61IJpUqdRtW
Bdn72JsNdAQSmE1jpr5HGN0RfKxFandmz+aFVwHoR/sJw5l0xhJnCnJeQqD9OdiW
POAGwr6PW31wlBEckTt+WnEzOo2nthmPkmRDlp/2v+ZB3uiUVoyyHIc/S1H4PunV
4JgCc5L4LVUH3brb5p8BHhuJ2R1vz/jB9ayr+lVEajtF+2nOIYdE8xjpNSZIZlWP
NMVo2MvkSkL5cTAlMVdDArs/qoyRz4sVpy8T3w9kzNDplXBdvHMVPnu7aQOkEDp9
JLbse9QPzFlIuRx8txQsH9PiwTvXHDSmbPVASCCzIErSUc3xGAQygs/69m3VGinu
pmgIz4C9qolp+odWXjwwdeXCMdw4kf6pefmBWd10VhwDRFh00HDeZV/Q0L0/r0vw
VtqcJIup9TRPgWbQ3Cs/10QTyEPQOTYpjnu6EY1pSAvBrVmX29DltheaSZM39LTb
RnD417zU0kLriMunaB/6cbL+NLNoJCmABpqF/UJ/l/ZFPJJLjcD43s+X97Apt5nm
YPHi0hxNPc3KH5d5R12D1MQJQTjt/etVSAIJt+fo+RD0VRzFMlMToa4fvwu1NJdi
6fsgI2R/s7ffHnrpe5j1OBg6u9zzooCqOTBZPM91WgkPPVgjeuGakyCuCN0fIHnL
QiUOnCc30Q5FLk6BwoqGo9abqGMUSqMHdvOAQSZSFlL3e8vTS2+5uwhhZ0ZLvLjm
SSh6BYTO33/9U/rmP7zwcqLVMNXn+nQ/StL8e30KCRbTUkgC7HFWRyoE4yLh8z+F
rcS9q4ynf1vl+o8F7IeVNK4HByBzBIinpQKqefanxDNKoyHRkuphZlvsh9n2gRQa
ypLvsO/+GwUB9WTuh8vCAzKPOt5FthyZ1jQnXRD3k9zuAaYrrANEnT1O+bhihHnL
HlsO08dkn0YyGwu/02v9kILPmD/WBOVuLT0oND4+cZEEFcoOwkA2U5QP1su/+ygn
TFlEils0yenbkEmslDEi3/QdRD2dyNt8ZfDucxGJzHRgLliTplinJ5DjrBBubrwu
XgwiYBRNLcujLAvkjiWwbuk0usBsrQTN0eJwHUfhWZ4wUbWkHtthvQhIsMte/6Qj
oNEHE+aRTud1vCP33xwzuO8/FxUNUfUPnWV4k1RLCvnhdtyuQ2mi2HVP7HHgGDb7
8AlP+NLlu8V4BPG/fAUb1VuINL3Fk3Fl+f7DYLOy+mnKruk9oyTYfFPmWpfdEvKl
rQvkqWTquOicDR7F1UuiZV8ai0Wb376i+9OGXq/9pkqTu80DVu+FXfFRwX3Fk0NT
qC22DUzR14vU9vlSCLlyE0lC+NUr3kvGKVkrHFcThufTSENDKRU6BdHQUE7CXws4
ViRYEcoQkcHBYAXl5rvAddh0gg+Ir9JrQgZ2aTOE8ZSbdVsgf90rOJwz+WWwj7s/
lVKVljTUz7UhS+/QMXYyM73f3/uftq+8gyt8yAsFi23crFUIMK53pLyfwehchcOH
M7vfOOXWeuspylXa2+gQkSyygIEmPg6o4JyUdS+UJ4hXjp6Pzp4h9aPobYon6VrJ
5OHo0ZZ2GHuW72/HrwBUzegJulxP6bfHkWrTqq67L+0k94VQj0neH8lzhrALO7bR
+AMyKjHxE5cv+o411zbpA5f7auZafqCOAx1u6xHXAGI7XwPj/WaeCeTGbl09LXgN
ZfgRd6vIfjULmxF8eQVZIe4jYfD5lPaZBhdqJWJ3+5oOuvKaRu9BPnRR0rytUQzb
AGQx+unv2ozvBSFbIJB8v3ixBLMuCP7n5qU4wTqTevCJeNGxWGLwsUMdJJB4FULN
qfDbHpqLbmLA15osB3MmJXJaZwrOw1n8idT4VropLhrPBcpAlPNmuygKWCeyuwQ9
F3F7e7OICPEWNEZjJ9E70lSR8pcMssulbrXqYFrcKCY+aaxEnbIJST/m9U01QrI2
+dWrQogm+eLl8tcA0rfxvrQYtQajb9d55OqPSKCfvPkOS91acTLlW7jHaRqWxgJk
XX6UAAieLBt/lHSNaBnGRcf4F33cKfi1+sW8rHyTjp5WnUi/Z4rV9jKs/aJ9xVuI
`protect END_PROTECTED
