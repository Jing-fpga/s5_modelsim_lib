`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZiY4D2010tRx04j7b2d4stRuL0qS8HCFie4OlJgeaRVNdIuGzsIYenlSUjhFsjxF
aPlJknpCdEXpl9EbPC35YM7QQVId5ARuQzhTEz+/LSef/d+NFUjbtO9Jqvck03Yb
D078aaANhqNsh+gPzTUFikov5YqkMhwWwdYY936WGpKipFQCjRjI1ANdgAjNRS7j
gsgPgstH3fgO1vysQdZg1scD2xzdrfDyYus8Lth/1+6JO2B+2NgBYrv8JiuvOxVn
uW9XOz7os4A5SVNQRWlTLotm8Dyl+U/BatLYzklvQ8tihXqf+wTnX07eht77B2Zx
sUNPRl9zNANFrOIPXMlriDlpBQb7FdsgRcUm69O0IVS/WXoQFTXveya2oKjnU2yg
p3cUJUdykcJpb2od5WwSYfS4BE3JHCYOOPFD09/KsFKG74CCDapPUXLKWcKj0Mzb
xYE4nsGeP8ueMt0JKg2ObOq3YD6mpM442zQlqb88+eMDqI+2TJTb4/FnnvgRYm/Q
4qqrRzAXO11vCiOns+CJYJVVv+vCO6LejBlVoP5rxUOWhVguV2pY2vmadtLGhMQA
uNXJRvMtRPvYRUSIxJ5vvymlfrZpqSKt9rnIrQiY048iTPqLdexNTBdBDZp4ixo/
onYSNRQrKfP2BNy0xcOLaskg7d3mYJrMV9dkWbSso7DfS4mSMFXbH0OzAtvk9Yfx
vqK3ERBg7GJmwpVMOiVAZA==
`protect END_PROTECTED
