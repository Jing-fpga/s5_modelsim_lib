`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6+Wk/3i5bet4CQxBOIAmuedJ/pnI7wDIDjSrB698TX3dY5J6GqMw2OVfDLRl+Oiz
uMY0UsjQdgxpMYv0MRLo0G04ULCTEdG4ChtKtlxyN1nSzeK5b0A/tJjECIBdQQq5
y3ED9HAgDO+Pb8iXg/z1Zq5Trg8jgwJj+bp37I66AWEJOT1qezdBLTDIXTs5u6xp
yxJqD6Lcx9YMS9XfNwo2oZ2ucI5MmP0cLuMPcygI2TlssayZC3nE2+q1B8Z34yAO
gES9vH8ygHNMLbY7XLg3qGvDBztfrgbJFj2xJ4BVRtoZ54UybuFJUkPZlcbZ0fhZ
Zo0JRyPuLYSIOBUMSTSXHmb3TONwFTbCIOfX0LuEYiVBFNqsbQX03l9/9y6N8txT
9U+w2mfGiZKk4ptd1IgohC0g5RYhplxyzMvyWEXyqx0awa6VG4ylo64XO5xY0KfM
Qw8uc60mIDGO30oeHqm+1sODTfDnJjbqtOBw9o7Ua/wc6QoYPu/mH88r91noFNWF
MxwOFgvSvqM6/gcfoEMfSUozePwE+i2rc+gQKo9lkPYqOMl7Gjh+LzUSRQp2/MOm
KK/C94UcMi3wJd6+BDWGOzi7OOl9xFNL6B/GLZf4Il+ZnRS8okyDF3TDtrnJfQXx
lXNdW4But/P1VD50VSXzm9v8qf8WuABg9t7RYeJgFJ3f8R/jRk0FK3AJts/sA0r/
FKX5bWeQk8UdYQeNNrHX+aIIc/hPmMSsscKsW3Ohanj9TMl2ifY3WWuHQG2VssmH
mnrjEZ+v90uPyMV38t6hrKzVMrG1ALHtg8H/Ye19mJSihhJk/CNiAPykLlzb6hDZ
Kp/DKbytxMk2ZIWV7n5y3il5aeCqbREcurJGi9LMPctl4eUZ5kKLUgSpjufNcIIv
SYPQIvZTZWcqoDCegQS3Di4T8SNr9h7boY8FLsiH6Yy5UmMIqgScZ/UseXLt384+
witMajYzr4YIzsWAV0c+ljN4XslwstP33pBRBSLT3VwOQqH1/ABCYK5Qw5TZeUyV
gAdI0lYTqNCwDo4AbY3i14yG0wYDWWaxVFFt4DQ8iVaz9xKOGEIDmJrn5T4UpE6Y
YhQATxYThHujSYxp/26MSn67HN5Wv20tRclfR9guCRxUzY0bmeZkwIhTh6qG19X0
GwPJlD7leJ37wTO6j49bc5RP8IaMgqVVYlQ6XM7p6TFKFhtVEdlBDygMzwMugW7Q
N0GlulmCH4Y53MCrT7lt+GI/x/cYDe5xZ3VzOZRvWuV5HOq5RsoTxcdt+UA1FbxN
9f1na56vJWIGLhvDf/lx0EaJ+/UV61AyVexxgQeRfThO3Bk9stRbWP7qmiv965/A
2ooF17ghuOsmDMQLDZ24u7OpWyR6RXlAz/T9K67W+gmb9qFKcHbaGaH4EiBJegSI
KmdMGuJhnAfV6rOJ/G4naCcNmnPyIQOsJxgFoH6cF50zmlgfdxzHhA30z71lExAR
GjjSrIQaKCQZyEqvmRP/Q1pC3o5gL0d5oCsfajzWAIJP/pjN31GsqEntdbL29jst
t40ltbsj6zR8hke9gHHtFw==
`protect END_PROTECTED
