`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/02lsHbwSlKUMp7jNHJ1eOtQE1lY9GyIVAOIGcM4beciELFpHEKZrIIbItKx6NER
M6DzEnCR7kX560+L4DYR2dS6+EDS2TbV0D96jEqE1WMdwpnDzHMLzAdILScOXapL
6smI3pAg7vMrNq5lCjEeRDngezylNiqM2dH4C3B//MOSFY+k8Zt8GqCtgk2aRPqf
tsw4gy7SyZWiWJedxeEucKAJRdKfIy7QpyjZoO/UHaNh3EJ8mA/gCvCYnRKcqNxz
w0QZFXtfw66OW5IV3BGDJoke3U7VAAv37rliqJiVpED08f0pHW6NQIy4vC/juRNN
CzscSIy/+BYTAobPX7vBDt40W1xdw45Zw2SmCTWFd9VWFTVcWVxZ9OovPOFSUXqc
37HVIhBWIgIJKNbXz/5A+mJhQSEjw6Q+J6b6JkRou9q9QmFV0JfOrUAivlzedMxf
VZWM+2gTpI6ga0K9pIwPkf/rQqmA1x17oYg3+mGmfUwCxhd1nliCkl77dOBHIXPn
THFIqbeL2Q3+gc1xWRLqN4Iu2IpCU5NhgF7hPHSGnaFjHfDWAsXm8YCkOYOaWgi7
S1Px9ir7pQY1+yzxSzfWiyEekNgIIPSde9iX5ENM2nmkRZEpSEvfhQlu9mYFKuAU
RoOoVjwzzmSFyoO7G+xPKdMadCKNp87bf3eGNTuX9RsydlrqbpPCloO3nbat5jAq
9YKfAwSsy7jP12F8xoe2prhbRMjtFm2ddwsddOil/Zs9rqYBsfL8ug6PHVONqjsb
EvJfRRlkUrljc4gJraJhy95bkjQ8OnqoT28u8cqFG7qdzAcGoYJFvdiZbsUhju2k
6uIJnWMp6fOZDYf4wBsHtVlZwR2WsgYBNA1bRZHzvdxd5eO0Nh4k+zCbU77Gi5zi
AbAJBbPHApuMISqZgRK0qBcIs0q3Tt8FTfsE02eFrCG4HU0GALOn0EzA83VLllTS
VPYYBFzNjso7C2CGWhviPGBrUAcaibOdNICT3HOC3GikzKDDSjQdkdolSPdth13+
ZLP3TCvwN3zAUE217G+SGDpGW7sZnWXLSPaJD2/9zcpCdf50BzjzapLInXz1WW8+
3f5P2Br2HkDYBMmJExBRDbTZyo8m8FV1OlVxFxkBnhphkdu1qPHD0YCtagVRXlLW
6GInsnaNHRbtsNIZjOGOsgpSTTdN+bf2cZRmRA3qz9cx9wTjVY7hNJJC+FPwiIzl
rdc7W1A8HPoxn3ogDYOgzCbmQm6+NR5SB9MDX6XVcPKV5/OCVPzcqHD1dDFJpZPx
CmeSCZsabmKXw0BvXFsFBEF86LhrQh78kTGHOCqdxARA6EYs18o4Xwnuwo09D1Oh
DEb+66N7+7Uhun9i3Z0pHZ+dKQUMyyH7NkAY42cMy1BmaBd5fel4KFPMO4Qqu8WG
aTxtDmM/6K5GuEUdxvwD9uBPVpv+iDmVCYhkIYw88X4=
`protect END_PROTECTED
