`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sstEtWQJ+XCH+xvV+y2wN627j41t2hQRfFGrlGRRSFSHVpDEuDD8Y3O9Fb5P8Q68
2k2SU5PwhhWZp8dh93nP0SPWKU8+WlGM7qKcLTAZVe0n+EkWaSBfIq7FmhFTOIfh
wAuwaKtKPrciIVbFqXemvC+Ii/ihZHn+L31JjV4GVNx16ine0HG1e7NR2LPXuDIF
aHJR03ISaf6XPKVeLibDamOALfVl+WFUZRy5mFcDQbvAp4PNr2fRxnWzhgGDroyU
7m9/6UDKhGkRzU1Y7cUV04FH4Cn/wjRN0M+0hA7VBg7x4G29qEBJw/d0Sy9S2KEZ
B3ByGGjXiChvknjv3GSAnxJkQkIO0J7N8PHKdkuPSRXjCYQ6ZxeTcW+SKiIMIQm6
OYldM5HYkFqfc4b6G0niZx+A92D2CXQ+lSYVAe3fIaa+pd3Nsw55mvx1g+QbcOt3
SnWORRqR8Wy0HpK9bDDJ0EqXOEseoFAYnhpCKg5Z4vHFmAVAuFoytNKV8rnKsgJ6
S5RkLGxxmOCM75xRR0z3zYA5fQv5m//wv7wiT0x+QBa07osigCbyxYq3qp0GSmf1
+wtRgtOIhaAHLck9fUawO8vA0fm7RY+2ZHhpNmIkwBQtAN+61O6qCHZNRwrKfuKq
sxdMOUevpM6B1Gs9RKj1xHv8ETWuEMX1k3HmsTJBcz94fhw209ZjvjGtB3YK/KB0
8eXPcjPX8ErKwUe2wj5pl0krOVss5oTbrD7DYdkG4guIVdW7gXK6F9rU96xNUr2L
FpT4H4vGxjt/uaMlLeRYpvUDmh8WOsFsrEIArhqZEMFeeHC5lMAbUO9LbWZa6+qD
wkphF7LAl9jcjxs1eTMrsou6QcjpV+u8YFJwL9rfTQF8pObmq87s/K/sK8bQUDIS
PAnQfF7ZhP6B+Ge3OKm6p/HTuvqXs31vI7PaEX0aRRaHWbq/dG7xLelQJOlKY2QO
jNb7psjB73K5ovtJzu9gT6h8OLnOi+BjipL7P67XMlrpna+7ETCc3WcE6copiMPB
xuqraeke7DQJc6YYjOJ07VwhtxzAQzFBeU7u5SietmhdomzjtTqubKoQHJvOcg8b
EShLLOvTnN66lOuBxhXaxqrj9/MnaKAm8plOkx2bj9XE9oXmb4pGiVFSS7hP+rQ3
zaAekNA8EfRTzyquorrnRPPt5Att2TLvDz+5QMfb1tPgPXNFeQQ+QvAyNw9cC4Cq
2tNuA+gTNH+24mHSBydwcYrZwPMaG/23+NArIkfCSg/ESu/kca8IbCmzSe5CetPl
pbddPqFNjb1Bg5Kysxr4Vfp4kXj5gXU148L8v9DKv/lUqCsXZAtR2t7ucYMe9pR9
OYCJ+D9eER9TE5A+QRBzZ6JDwbGgW2XEQOnG4zNHm9BXYdF1BY8C2I2mX4yDpG+d
KcJ/ocNshj1KbauSQT4OsXZNDBu/eoN/psSlLYINiMas9z33rstrryLGHJzGCafr
u2ogHf9Jo+ecVpD4Jy+UOBArLZ/NNFEAJNrxRBmM9oUnqn2LLsVyQv1Q7uFzFbhh
Jb/313inJt5lebTiOH6NY5PoFA2AvFtbaVGQCjUc5YI6qqO2GFp/aItjKZ1cirrN
xerboIvWwzCSRz65/65d9GjDrnxzjSFdYGJig9KRdpMZdUsM6hAmJAZvghrS6yqb
ClDqYo60QnofNaVT1w9bflbnKL3lAOpDNxi7DtIL4VyFVlG9M+XHyK+6dSWCW7e4
yiZRrdKMHmkBbD1u3wubo+5YWL+ioyknQahsI9bIwcwekEtAR493XnStt+ySkFlT
sefyVv26j1mZ2KargZS9/UlFcMnhxWJBjjYc6q+PmZAVJMtXg6/yMRdUDsMFuMk3
mw2jtwyCAFkQkSJH+oaQnhkSOWegih+fonBcbWlxjTxIeIyotQSLil0vrAutSw3S
4iUv9+BtwhYSqfAw4UcVc0unG73NfmhD+Wy715AWf1TOhbwwdvaRLaeWvCw8Uu3i
+yEEod+m5JDjVQNe7BPZWqmmLM5zX0HQJQOFq5jQ9Gz7kfw5il9Rm+QO47+Y/xPb
auWgRWd94P14YIMvrq59tStkg8ZXqJva77Mkb58yeh+RUrG5TsIFYf1/LWApML+t
fP04taVzQnZ5mmlL0HWunYC9vVEiBCt+e3UdyYj8I2lj0elga4X13foPbr5w3W92
DvMsXIWgriX/tFmPtJ+m4NwU2ui6QiJRmxHAgklTv1ygbMXTzBe4GaH8N9qiraJB
ekzeL6IrB6znmaZaU7j66LKJELUFGlkka611ESgQU7TYkX3bxi2GI9o77KYC/JlE
+oef1MPFbyUMLjFazcaVx9UjYTIU+J4d1tHv6QYvUkNcVOUz2tmvOzWLpmTYAi7d
c/Bg1kXw2f8+o7xagrwRgspJuie5+oy8St/qJO3W+DfLtvKkbu4vJxV9h4sgNCBd
JLxMZcTLBlCmBiJqj632/ysy4Mj9EXae4fmeCbKI2jcAk0sl9QFw98ZP5wNrd0oV
i9+Ti2C+Xoinb97SaqGLTk1DP7b9b1B4OTjh9JEfbGj4ysXYqL1D9RWjjIrFK8mx
5pYGesHwvRucAqwL79OWY/HW74FqUIjj4UDVtl3wERO1H8aRFDyzrbR6o6LZ71yW
KGcWoIuGTMrnJqmBeW7stm/telugt6S657qoST4y0oSU5LpbKKqUGbIWSYKLFWRz
aiBiq/DZqyXz+f47npBEDUGqEMiTJIRg0OYt1G224aORQ6kucXxcW5Ngcma10BId
/UHLMw2L5ILfq6TsntvzrvUHfYmL8QEnygWNIhV9+bwhAhFqU52cZ1t4wbGsEEBN
lY1/q2oHEcjDXoSENq9botfL9itpwsE/4O6eGKnFcnfVMgLGiKEoQAgfmAG0+JV7
eDkKqif8h6FV9HU+I5WcP9CaiU9NxZzc5HAxfxJ7jz9SUv/1fJkxGd3b4UXTMoiy
sYA5Q5I7SWtr2duzHxxKwbEzWyGkCRCr1S4jpFKhOqSRbjrGPIqLhcsr1bchFIW8
j2AreA4JyjgPALWf8k1WjCfQuNNSlnMGD3mY5LgaQDvUFMJKhLFb3cwkeMxAuSyt
21AI1A/dJ/Hae3x/t0zEPzGX1wsOBBn1hzNGkyzJDMY82Ii8uD8A/zCEQlgV72pf
0k3BxpgX4DwfudGnJG7EqsgTAskI/ybwUNDt5oh3ZOwnheyDdSifABKCvgnzAt5j
JHUOj09S/WQiVnObWOodB8QoC0b347IEkPNdIRzKfc/Boc6SAhTHXhpvxBRokt/C
XnM0eBm4EtXsPBgnG3p0U8pAAKKtqhzagsnGE5UnTcrpTmo1IUWzSXBOVs049OyI
flmMm8i+Z3sOb7ims146L+dB8EIAjqv6w7r0Z3qeWiAXDc0GHQ8rR+FG4nu0fVPK
5+0vPVSR1PSVjaofPrjJjIP5WTKwNQeg8XwopLVCP5pr0DfLEXAqTxEl6dZ5Z/QY
xc78RSUDpEBh6uZ6nlmyQDdCcq+zn65IJpj3XatsBLxiuHAZw0v7dwaAfUW8YGcx
MgKyDbdixwkK+y24vI1KL9b4mOqMJkVuB1KWOscVSYLoUHOYcyzkKbm0dyV6+2Uc
frubEP+XCb3d0oO5655lsbmuCLMxTZjr9ZSUGvo31tRqCBhJnPtpn64ooeJZyuf1
n8NuGYggIFrwq5cfChQOdQ0K8c4L1e0/y7jpWvY3O4rVGg0+mO/iMq0kuKrDAztF
yrQFYYBQ18WTAzENtXl6paOkF/pBa9W9Xh4sc96XZ98GGG5gRNTCHnWZb3iqMbL8
6UNf2HmLWn7EgOrsX7dfP3SGilYSogyTBv4hDcNo+rdrhfX9CtVftiEt8ERJrvJu
bqR5PZwxwRXlOK7V8JQ0jOPWls7oW+P8HrBe9Sl70LhFxn/foFtnx6QRCKm70VRP
C9spM5Ji+WV0SDhRDQqqCZcU1XhhCOGp9SRobhg398LMTC+P9RS1bGPgs3pWvcFG
Mvfc8sf1SnybYZqNll1RFzwFY+SklfiEeXMOIa7aR7ILyf3Bt6YrhucujDUlyqu2
4trunxKhWNueo3y09ALnV6GT0J9WMrGms7t8G2IxyLiQL62MOGUODwT7bmSF9+hW
DHez1R7dUlAQUfrLIHkL6Hia5Yci+mRmcIXcHw/HnJou9pOlxK4O3XEDVYz470N0
In/txL1gYtCVmgJ042kn4p8TTzL08RwDLQPKnPxZAz+4R6BtOVrbJsBOzVtYK45F
wROGYZO56Ovapu1PWCOb//JuzQgFuXMMzZYdsYXRRzSg4UUO3P8bwJQyZMXtAMqZ
QiyaRnjxoVzAekUMWmaxiQBqbayXPD4vZTHAbJjw1JH5ZVY1oOfnG9KW4G22xIky
EvW9DiKNOVgiE2UhM3R9ewqsJ7VRGDBv9m3JI2f/Gim263fRVnyFS08kdzkUf6pC
bzFHAElyAwrU908n9aQg29jYdGm6OGPn1+M9YFMuA4RovL80IGKLJK1kNApRQ1jP
AjqTcI2pgvXnRpFlvQLsYx/Tpnw6KK323Rnm6FMVtlaQ4CahbLt5CIpgxeqmKqbk
/K/97Cvr3zgE/RTvWX/ndlc7qCY6tJCcirzeidyWxXe8CBdyrY2zIDoBNWO61IKk
yqy58a6jskCEBsLUnjoBR7sZg4Becu4PH+DrB8Ee7O3axxPoXivpeyU4FcGjjRqn
qMPwIAC86L40iPRrUqux5buLPhlF8uehD4yHSKhzvB90TG3vnBijLWtKYiyWC9Cm
0A9QXeQlS8pIRY/1gIDmCLX4Vcykk7d8JNn+08qg/Qj9ecZQx+4WVJhhGLSixD0s
O8vSjJOyLa+0qYPdNPNmVApRQDyu9bo7hVViQ/Cs3/XWqOCFm0n5MvkTccYvkIkL
jSCbXkcbtg6rA1VUNp+11CAAx8/BkNl23/7DDSYcgvby7RGFLW7pgmMrzvWWf6ml
p6xNAXsUA60bqJ1Jg593BGXLNNetIau4Vn7NQkrsrkFrKTtwMDHVTnqCSd6WNwFU
rZAaePmOM3LaPDyUp4Lp4q7kJ3vKHwLjJluoWkaO6xy6UEAGGI5KdRuDwHZoFnVh
Ky+SUPGfNtwrxpgTpofkvz4Ld7jU47FUzsyjqrMVpDuAV5904IDVSi7yU8aA2rRh
mu/TPHgH7gLYSE5lKAJa3v1UzvJLfSfdXJ8tis/ha5l2yOe6sa2rW3IO2OOX914O
78VENevpBSsqmaADud5amEh/ifA301tDB73HsXz62eGCcA8y2CX7yN4sMOmjuYMc
HJdU/bFVhQoNQR1RXi6YQS/dlG6I5ujHiLbjpvCtmXD7Dv0/jRMp6NNzWlbyNDje
wnN/p79VYGbDyoy/zCgrQZPlR4CIxRoVJcqvqcaZvvIMm92vVMdeVNdhfH2Un/5y
BiYm+Y+M2WDMX++gsx5+3ptmZEUqnqMvHfI0E7Rovd0dvD1vaHc9ZeGIISvcHjCL
WPKFCRqLY0K1vXLO9dVnLSy1fTmedljFYgklDewufprThRy7xc/4GdOHR6ov91xq
+EUTpdybclKsr1neYq26URa8Mbo4Z2j2GZg/IUhhCqEZmErQR1Oy6m96Go57yaKF
yp+JlpmypIAN+sfGNlc68VxArCfaZSkz8nPVxTWpsyRrn5+3y1sRyLxpdJ3u87CS
JiX0gaKWrgQ601JrIKUrhDMLEyWG/9GjRVWqiXSVLZMuBCDffmBaCB6TEkkX3UR8
7Vvrz5sKxXvSZH60zc47/2SypcPqkJWbfougaZVvE3/wwWAkY74jdPYiyybmKYx1
+NuHrBbi4tczV15+w7nSJlfMUrF70CtxN8LkbG1ke9rIwerkYSuXZKxM3T3MAdoh
u+40TLTBJvv31BKrxZd3lsXu1i/bp7g7bSjzg2f4h2SfAIPCsWHEur5+kUX1T1oy
KObMkcU7liTsifDEufFVkztldleh3bDgIJR0S/dj7mccoK24kkrQ+RCPnNpSd21D
KWs0LSmMRCcxiXAZ0+7ZUJZpxr91B0+i/VwAY/CZyu3zdKxxpAFgAVTNvmtGOcLN
xsvIABWaKLgS7MAfPQhu4YUPKZ8dLVd5HPB582+NTukeIsJRLUUKpgCxiRNIID/G
ZwciM+IZUjsovkkuOmxmIozJD7wt7yOzezL6M/WO/4QH40g5Q4L1NXtXkvzG0rbA
Y3ELtRI2jgNhwjHQnxfpBu04z+45oMrTiWeKfzkKXdpVjWbUwToLPL1Dp0TpBViu
hkJ3wXqNEVpC9L5Qfj/C8GqSxcfA9qTas0PbztuwUFfZQDzHTls6ALlD84DeP+eq
YcejlRz0J7N2HEG4eZFdoBGMnPfFcwjTknY9TKlaQQ/+7QP1jIBth2NjAVWCwe37
tbaj07CUkpA2QIvMmAjLywZQsLN5upaQ7fR49W9We287X7pD6FvOdNX6oNengo6Z
r3c+8VKlVCgNW0OzMz6NzVzpi6EHK2cG0tk2iCOJXmSpQgw+WjZk0F2szm9PJjvc
6qF6Z96wl1M0PDpY+Svs5az8xq/15ofPXdGUNXZbbtDLwylVUmdOuaAczv1KVQPA
/oMSbAo+gmshz/1OAj8TyFoMUYFyDjwIXS6j8LwuLvGZ1YM7meig/O3IpnPqHcUb
0ffPUawTcTC8dCUAFnvP2zFlyUa+SUsdLaFerz2QP4jt4YYaSBV5igwdwbeuLF9j
n5msrDG1ALez2QUz+GcaQ+MgmL9bJcPBdETXBspm74MbHK06Kgtoe/C4PjwePiNL
Ft7OeqV3YuF5NmY0B0U8aaaDIjRGJiqgqrDdIA/nP7uzR/CsYcrzBhMAxZ65dMNO
fFZFARTcecDrVZLjwjAfRWZn3odQvrvUCZylxrrgAGvQekrND0766B6UqaoUIvND
OTZYLJjHj92hEZIuOS1Ax7YXsxqDkfGunF6V63gj2zjshGin141oork62V7hmIlL
vxdCmuXCUOllXhL3vnNGjoQRjiueXR+2u0kHjaJzxbMsYpnj6UZu5Xhe2giyLa62
LzJjMfRbt/lKiwbBCyGg0Evh4W12Q5K5ePKuRg5eC6BoIDhYZgzWRIcEOC3lo/Ha
m/LFZXwihtPuxUb/JA/FKUxpS1eDor8ASDwxz03xpqJLByxBGleoMd2dMYhfbtSq
u1QIhetapWZGs1acthYoeExj2Ru2Or6IqNYFE7uYbkoTdvQd+etBPtZXtyyIWx0k
Lp2ss5z9RMnKdH4+oXCVP4K0GRJ2t0+k1nLKSRxf5cKsWswwdS8IifYf8/3U8iKv
luQJfhlv9hNHiTemStMq2e8PoU90Q++fo+vtqOWoftys1Yag7pjWdUeq8gRQFlAD
AvnUqz9E0+FklsN0wvPFwHJwTSBGdPqY7s/pijkHBo0l73/Fz+AFHAdBKb7qaZgI
gVFFtKJw4g0up3pQ39ZTh5bKkJ1mxSeYE8iJrFtPw0RrWRzjMEhFUWzH+y8A47Rj
+UeYFRREyzE9UGaXypEBspaXfXyS04vsqsOBIAqXYbElF1mBvOSKsCh3s92N8/du
C8IDX8kVragBTdP64Ybrlu+sq0tLX3pdjgZQCWUCgSmWYEff7g6xkozeC9VenovS
OBc0nP3B0yt178aSq1ZuwCJkhjSfEw5HdgKd8nb2BPli3fCzDWJXX2bT7fIfoLoK
PIJAQHaPZz9UOlpLntDHLs7y65E6fz3rIhhMrMdXprtN8ZeuaWcumLfj42lf2Wpo
k0C1anabBZlXRKnyVOw0RVC0T3pZeoYKDI/Mr1p2tVW4OGeu0JNX40wHVeLn52L1
K8VT0PYA1mR0JpltKMHP3aSeVKYqcu+plsoZ/xOilh6OsZcpgQqFXj23SBwInlRp
rT2vLvW39FkAXoiiCkPHtLvvctp7PMVTm9ssKbSCaas/lKtQ1iAw8w1oYjVHAb1s
CSWlPy2hYnB65dp7KSG+UOBLEsRUh8YJKmEUzB4W6OqOslTFhylva6vp5QTlrZOk
cI7ynU7whxdtkYR93RLU861UWJkzBzn+btfbfZ6dhAQGoa9Nf7ILQMtZKA+TKuZ6
54ARgi1pwZdE2RGeYNzlVTNn/vt8oOkpMZH0fI2n5z0qHatglvA+mkRpeVU02AaL
qlyvzEHxRfWz72Ak35mMx8wJAZ8VujFqr4uw/BI6qWYqzbnRKn3sWgCWo5pc9te5
urhG0fgRiPbwZrFLu3ioDrgoKOlSp7CpZTMQHoyeQKWMy4knxoqlBp+OVxTzR2wK
prq0GnEEavWeP6Nl+6DdZKzEXRhtqwX6N2NdTSnC5B2W6B41XDF4opnqEeD9LKaA
EWRcE6gkyLCY0oh5ZyI9kmSo6zpUI46NXr8XsVp5QR/kzNfG9dSlstqbIZIKBS/6
+K0BtxPYlgJu/2p/1uqXkFfdNkPx8K1Sjxc5lMwZrm0IX9Y3tiNOL15RLGKTl+A8
T3trhl6JlpFceEkz70eP1nYFre341ZDQmki2rqH/R7zlOua/3hP7srKZj6OO4B5G
+L/1VpXKJ/Goc5rjs0R1SkEhYqoHmVP5kLeSKN6+8YKkDwLjz4qLrS3oMrIkNiJH
u/To/5GM2TxTYMTyRNVgPP31vWDdBBaT76Qp/24jQZpASwUbmFXpmn4kskrbSThd
EAyDeoQeygGmquyBFKDQcTdtBaqoMRISCYJjW74asp8Ziqvnvp2C3pR2vYlHcMkH
S41QTHGbvkj0u7uQgV07wZXkKn4hW9rtw3SM1J70n+KpsJJnoYs5/QY176EbwfY8
wEBZwZ5I7FiLDVfspZ/GnWESAn5DOYd477YkzqeGGRtYFu3+PUAOLBICMmIm43GB
tmtDwVTkR90IbRWfPH2sGLNpWZvpUK2eJ44Gxk2TCdLUSufxF5+Tab65mtfJbLhJ
nCB2SYpr2Uogp+0EbpROUH8oZ5HziOFjh5ncKCYf3L8TLtkbIE11uVf8ctpMsq8b
OEIjVmA033dK7J3TiWF/Q6ty2GiqJk/zpWhWNPzIDFKeeYXlgGfMw4hAUhf8fZWX
Xl5N71bc589G4ou64K0d0Thl9o4B6EM81gWu4wAd/oO3ObH9JlPOURIzIZ0spBld
zZkSJGo/SCTGoOayRIt/fjXqS53jADWHfoEFKHSyiy0C2WgCcki8jUubWettM6IN
MA8EBSTPWgPfia1Q3jUVMVz6lrnqwXgNYGGnvx1WaD2KAtnRWJSB9sHHLlyAHpZe
PEBVsb6ejO8u+P/VjMknxfkPpXHBc5WakB/V9mhE78jBSgCPb6ClkhXz8wiXKicN
E5Rsncgyfcw2eE4+6xpvkUG8mV6CnPIfDtbVLOIzV42r1Eu+msj5r8qY1rgeWjof
iuC+F7S4q868iTsxq3teoxNssoBz0eqwsIpeTnxSxJ60R3V+KfGjoDZRiDU6pc00
iwZUWo3FZdhzqKBWZfCdS69OCkIwdUPDKW/7lt/Wo2O6oWBuRUbJG7YOD2Azf8Ve
A2mUQ+ST5D22RVp7M/agrrznMLoFi7cEK1JMJDtBlLQIEzIV8QMPg3BB8uxREJ2g
/Tujn7PSRx1hqJPFozUBl9azL3K5hR3/JMnVslf4arrouSr6/rNFa2lxFQZ7aDYh
aMh3ynSPl28BVmUpuVC2LlaiDR7y8tQTTLEKh0ixkdva6wfiYCW0y5HRXert9A6B
DJHwYyojc63/bDX8qKK8+VPRQyA2gKfPKo6Qvi+vBEn2Hx/B5Ck5REKFebi2KIT2
qu22iKS8zLAWVc0ecmcPiRTFw5s9DoSqkUCnKr+ZSCxhuSz5h5O+XE3R4fdgz3WH
FwUsfMadQkYiq9slgIXIupQWHNSvH97opuCcFtgckxW9inUkDC6SKWmKSFYKtoVM
BK22LEeHcSI9r4wiwZ6QjJmpIUZ5mURxPBLg8mTaXxbOtGsLSqjoLGdLvf7hDua1
Du2jVSdGLnp1rBjGU0uAbr3pTfWhXJGtEZ04pIwv5A73QMxBq3WRvDiRKIbf7AxS
s2HQxQYNPbhez5aI/wqmmyShXWcyUskr7IueAJi0a++tfppCfg1Q74+VCf4l8eLw
5weBSrhFlaAXWPMkMP0ADboUz6vxaL0my4OCyp3YEmts9ElSoLSNfj/vK1C0SEjg
ql9vO88fjm3XXJmLxST7VS+yT7QGAQouPI2YL7fVgW4llj3X+3k052UC0x4f4Ylo
Iut6sHN0L65JL8Y6MmV2WD4hDqLt5J9rmUOGhB7Mqh8oBk+j4E/SfIqHTSg/6PJg
0jI8qlqva7tHwRwvs923KJVSi+Ta3M9tOkonyiX6ulU0OYvBDSgHzZHamsUPu1gM
qMaKzXNFFp9B/x64NWgMT0Am79BbT1WrB6pKd+d3+3G3TEjqrJ+CzuziNRkZLVId
mx5ifbo7mFy7o/59yVEnRW+TyjRDBQwXALjpwrmS/lY1IRtvrI2APTEb6RNfjda+
EBlpXB6gbi7f1EeeaBi01jCP+CRUv/ENhw/sk7onpFBPxGjzjRj73arYarp+L+8P
7BkHiSw1VzaGvqa8OOepiLeOwrhcrioAIuO+cVwTc/LHNrCNFKQqaS2/aHsGOQb2
ahHDJFVmNnOp16d5YIo2tEvGmks9BC3s9PNPuBqNlRuiJSmfCeNAEhH0HXF8Q0Iv
Eqnj/35wKIgk65Vv0hVW80Bu0tFM2sXMFhVGoFaGHgPmZDMoI2FzIbUCLu6Pg6NE
sn9AnoHc/EGWo8JkcIszecbLidKkzdZn72w0qb03jyoHB+eP5Feyl0zhWJ2yVkf9
QLUH+pj7P1izctgtvRR7BFG/dfaaEPgdIeS0d/RRvIVHlTKk44J5yFV7cwJq/YJM
dSc2ujYpgjhrsn2QqTn9ksNRjSdqwBaTo4rlYQgxTyM2TEq8ytTxF62/5bSEbvlY
75hv1PJvboeAQQz9vE0xxyO1mUWMj1ia1x4G9IZmP0NUMyAVs9/F7YeCvltgiEFe
2dBec5BHK32iE8lu0uIyPqV/5iV5LmeWfgGXREHmAaEcas2BEd4Q/V2j3q1T0ldF
z8aLfxwBAHueUh/YvWlewjJEPfEyfpeNGBGsrMmsBkiOvkM/fkirGsBx+79IFidh
ilECI0avZ/sXxgt7pxDsbUGAt7YDfgv+4/9FHqBjcCF/TqEJ2XcJO9pMcBiRs+PF
wpD8wFj2h45pKX3w10HdoyZjIl1f21/+dYLapO6MldzgUxHMNMMY4L9Y38W7l+I3
AZHAny5c7Jgs/CxuIvZ2CF2HgGGtcHNpgnEX+KenMvcV45ld8XY09Ovl+XCHftgx
NuyAK+WsyOi+Km8GvcKqSI2cs/3GKqHo9jJlGzUfnLiYG9RP851Jh2dWUksqUX0T
2lS6hrD0YelPbHXWIWm+QVo90z5ouzRs1ClQsSjrFH1FSBG5cELDWxSI/iQNjGjs
Yb4W2LEwlEHrtfZ+f146l8A24NIb0cQuw5G5gn41ywp7FlMUlcDlSMwzw2o3Nfe5
K/Y3CKLh1RZvcvbIJ6xxJ34piVdJezuZwyqBq19qV4spMU37psYjDVZro4W8vTIS
MnszwyS0nNI9OchvVYCMnoXcNxoEqcZWrqHeIbbybXPEvLmCas/nu4AvV/BbfFX1
y+dCqkTBhjLsy0foBIJhW975JGSw/bTNjFTz5lrEY35hfrtthANKgmrzOrpuaRX7
SuAfqzKJtgJRxt7iUr9vj5N3xpOOFlw/L0MyjAgerC9CgVykPIEGf5JVF8Y+MhsF
DbpieRHhEH6aTc9pb9GtyXzfdZyy5/ZR88IKXUiEhln5CXvv84/EvP0wxSuNUbCb
/lRMy/aXJHuVmQBEnut/eXfk2vPFsUclaIWojKrfWIuyupmUNG7p7PgEGuAHIO+w
dPJhVOHaVXDJG6PQmEO8oRK0yvecx6NJPUVnPMg7vp1wZkWal1TS8G9kV6kUj8ww
ww3C65ew+l3vNLbGE5t91QlUSD0Zxo8uJfsH+kwV38L2KtOov39UbmWW6mKazqZ9
ka2rmWqMGUGBptt9hMRMmD+T2TZE1ovKwQqbsz41ljrLG3jRoZ7KYXb2OlLAUmHe
hgZ/G018JGhFbHz8cNssuzgsdBWt32zn1EAhZRVgQrsLIeZGcAV7Y7CEL0YzGqYo
pgX3e7zc/udqgY5R4zgN9oQFW7SQzQpLQOOQvDmmHruDQiio1jgv+Q9i7pe4Il6a
ZQJ8nClNVNm3bQ2PeW5i/+O+GCfJOZx4WO3BR8W4RWnvHd/G65t3Do/+olHtr+U4
qALki4+5Ibn8rY7KXmgOJWCw0izuK1e+1CRNcRf8aIdN914qWvv2A5P46mSm2b2m
WkesHs5L6ErSv86+E8PlLJCAPTbhtffzAuVfDVBTJOo=
`protect END_PROTECTED
