`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bVBbOt38BlZKdRZC3mf+8Wq9fm13H58tQ/YaM55lLWpc17uR4SSOgU21rMQ005yK
gegnK2DrseZl9qOE3IuBjjDzlTfr/tP11mQUi7GKjEOjU27wSkHxL1SNahvKkooP
2fAjmz1kjJOG7rlo8d90Ma+e3CMEFROdbdSoTbyBQvC/zMaj4M+KttwcV9+w0Xuq
iMkr0ShZLcxn3V3b16BOUFH6A+5/2pXp9nXB4Q/W+ZSxqcLKEtbd10vtU5H7XRCr
HyPjWp+saMyvDHEIG88cs5DbzkVzjkp6ZZFt3uhQlNMvTZROJ1tGqhrcRZ5p2Qi7
IGXo84bx2EYXP9adbxc+ZPlE+rYhFTE0PtGIzJ/0p0boQfH65/cMdynWvIHxDtLY
06iOxmO153qGGi2NocpuvgIAqM2zDbVwl2G8g4bJTfB5mj+Z6Dgrlf4S7/hObr1U
TeOfTkrmJVqvwgFFpgShbopAP0+hPPgEvvVZnCPZtTiYoM8hQYfyeSLSLHAhKSc1
BtucmXH0WbxNScG/wZbqHCaS36y1eQ7M4bQCSQHD36KwCnZMfdnbR/roM8Uo9Cvo
2wsik2MwW+jk+SmFZQi/PxWpeMPeUU+Etrc/3VoQbdVplD58umA3EhdV5KtyGLOe
/VT6MHP0DCLKVg9NVUdkRGyyQxbJtMZdI/YCrJ9kbvMbfmA0aJ1Biep2bzTuQHfn
SiHj7c839CzXzCrOqRzNL/6ufdAA7BFaV5HvDtHTeR2/j5gWyjQsknBY+9FHqoF1
8x0pc27nqDkidb0DPmOj40Iilt7oVjMuS6Vrl+2iR1zJBYU11zmnE0ips4Hnf5VA
KVpuKQyrqN6ss+PCizeFlMtiCJ1EuvNfd2nruGtW2WShYeTMDNsSAv1qq+xSrpr3
JtLS3NqE807+ZQ9yQpJsLm+Btd4uvIpd2TnggcbNpp8XicuDgEmro9EWPcG6pQR7
eu1yNL1r2GuV/Hw/58um2K7Nw6/favgW6TUrULbhiUkRjwqjiva7XcBcFsEkkjaY
ov584TdidijSHOICeI3HtyIM7GxGzsh3dHLoXCSLuNrFXC5/S+JyUvdOEqomnyE1
4QMGkyfgltkyBpDmU6nBoxvw83CLmuB3bjGoW6DWMfFXKuCVOp6+X5oSysLKtm5r
PyBnKXoohYPoJGxmIck2+4n1B1sfl2XTjTaGN8rfjGUusm1Xu9qpKMh0F6vXKIJK
4hBWzxTzXZmZ4rbUBZJ4mUznekWEF5RS/Nht8rx8Y4VgCLqQypWN30mvlEezfppE
w29rGfln7DiSLwh7Pf6Penp+9rIf/u5AJD7TG6jn4kcIe+WwSkjxWVmBIeSB0MN7
ZIae2ibalBGQEWI7Dp3PT1dOpwu+rPX90Kb0PvlIo3dQzDrtYkzq9It+cjcuchru
wV3rsJP3y/+D5AO19EYFvnEsB0/bdJzHevxmvl+GJ2evHnMPHCJ7uvatCPYqNbLT
pQeyVDyqwyR45Vki5K/WigOM23ZDSANx+QoM5aoK/ahqZpLiXLghcH1zklPlIE/W
UfEwolId/f7/L+yAZWopyxywMw/PMXUqaHQ0gRfjUA5NrsV+RbiPqEAl5c5dq9Fr
ET/r/2MgOJTeQwOZ2ON1e+WUL25Yq43rROPNErd07oDiGcwqv1PQbQTr1qUMslXm
W6tbgb9KFEh9xtEpisMgYWQIRT9NxyQUWvDoyvhncANUnLYxq5t02Zpdi9jSfqiG
nTfR+M+4m/doLnOVdrTXGcTKfZBkEUm0Z6Dj/yq7M08N25awHdRh8n57DAlgFz98
+KIh6o3m8vI/v4vyH1X1OuX6aELezla+hZ8/ulaxDSux+3cbHn3Y03bSmVd7NQ7g
Uqi1v7Lrf3I/A7vjHNlp813n1eexpl87N8OEm14XtSUyY4CfCnDgPjFDmJGfYlOO
53RIbn8urB8Rx9AyhMKk7x8sBnwSNW1MOFZj5v2DmDORSECtMFBCAmzYGk+mN3R+
0JU65J4ezVSsaGlrnQN8dJT9w3dGah9HcEw9oyx0ofB4ufuTHfSUPS/YIyxFWucf
TB5LUHLGT3KXCCDEqKpk44kbByOtGDV+qV7l1l5WW3KNj5E7c8qX0TX0sOJik1HH
lzQrc1Fu8rMCvOe5LWhLYWyzEN2RoEpitlkNHU7/mc/ijAusC6ijIEg3nN4CuJpQ
2FImneWdmYJI9IBmLzcXrcWRUcLe3wUgBMVLN9QTQi7mbFbMsHSXu1ZKw/gqqR0p
xJpoebNpgiCMt7PIrnf1wiYJsqhm14IVuYf5HnNAdkKm1ft1f/Vm0FwJB7V6H2Hi
EktAqHuOGZHxqTEnzVgQciPCCy8J6k6U5173+o4kxhfCKVl3+RSIVYuTgjfwE6wF
jDE2eRx6WNqg4b4zlXw5SK7wbnGqun5EZ087DsNdsRqD4dxiEL3WbEF5kqXoIonk
eDLP8nsCIhvykSbU1kpKeiKKR8YJCef9GQupnJIdGdTbCgxrv2cGxcVOY55XyyvI
09ikTGX7QPwmj2ODQKGXfDjltUceVj42qZq8dQlWY4XcY7d2B0wjDjLVvOIwle7u
riy0m+M1gEhcTuzcnhxWqP2gMmFOiix/F1nQucnlHaRPl1YCIL1LRgFB6FCWcWUN
KgYO/y6R6dW6lQHnCg5WPCi1u7PSbQbMH/kxRskDLXsTYyGD+Ry/67AXasijYtGq
oVELokGr8+Uk1i7Dz9ACc90acmTDavJLz5jy8pY7kyRdpRL+Ws05BV3v/C7Gkyms
9+luzVvlCm1uHiOS2JGYb8y7STeU4KCM3u88tnfSKYDUX8A6Spww9LvvNcWQ7uvN
vA9j6sQF7tK0kXDUKYO+S/pqukOjuEMl73RkOoophr4B7+6SS6UO2rbSFGa4fAUO
O6QYq7fdNIVS2LchETIMQeLBvgSIYet0+ACgm9lGlnBcQNx9Vbe1cDG+plPUwjO+
FqBUExL3NB0iSTHM5wjSihfwUcQP92xoPlWPKtyHD9zKC1bqGa5cFf2gEShLdoO8
GrHftsWK6WLQ0KhUEBuNbuvTTf4Wzt6OtIPhu58l6Z+/YeBEuZytPm154B9JRfqT
x/mUeWWSUzG6rKM84aM+l2lHPNFu3JElTeRcekOnvIl5FywZ0E7moURE9HLcyqWx
wgH0abp594VIDaVyt+2Qid5DABr9Q2+QfCXLvnBCyQSjpzQdsjWju0vccAXumdI8
ozUQlcr5DTQxn8zm2Mj4U/DQI1LX6k3sLTU4PwXjxe/qX8ma6L14zsHQpYwx//hM
yirXbv5mlb8HvuEr6z1yuq5/cQ0r7Xzb/Bkjnj+t8dQVWww5NrFG/VJuL/hNfo4x
Z5oDfAhn2yjJT4YjUw1D+GPgTlduKT0II9Vf7QEF8PLE9HyMGCJgbyiMVQY1UEmE
kUju6DZieh8Vx4vUOz4k3TwOhxBPvDJqgdWEnDYeebYfNoWwz0G9kVWvleYLe5a8
3mt3ajZAkEEHBqzpaQuAeORE/YpNhFAHibe8a180U8X6fi7o1/3LZtQPuRYna6jV
tkN98I3klxt8IGslaRUg9636TMVcw+/7q/bSm/J1EetVTlpC9/Qg0lwnW/PRlmvZ
q6uZdT66FNILhlateE1hVr99BVoMicvEjFhbYNpqdJ2z8Sk/0qT/pm01+y9wm2M/
+NY6Fl2NEiXjSkylkf1tG7PY006it+Llqx8cm/C7GHHNCG00jNYRVB+Beg2kmvhy
35b6U3G1hxIhSdiGFbaz8tb8uzkgJJbky4ArD/UKDyTwq13kDbLCEMoTBm1jM+eQ
h3c1c0Ir9HzBGoNzTjNZGdENfiBXz64+AMQGfuFet0AuZynP2526JPxOg6lcmSxg
JO2yOTKzWMvvvB8JqW2ngt5Itm1oflLzP/ktLSlP6ZOfYA2dzZTTA4GYd4znWHXr
THfUKox1ey9T4ZWaGbANxPDGjGUujSp7p0ZgszZlTouRoT2mnKt4MD/1Q14seHhr
9iVUKFeFfhmLJ288C1x0wA7rJZue1cz/PD0Y+UtDSR5/pBT8Icq1yVRMzKpYCnaN
wDfwjG2GcPHBsAoRbCAR8UkTCH395gSora68fHbWVs9tjccwMPTGWCAVZg1Lkn0Q
hdQzhiwAA7QOalyLRPmqrR2Q21/Uh8iN6lwdBVUpJbfvAE7PMBSvHz/J+UBOd7bs
t2nST4GpuD28YGDiCwjRJLuGTSUfC5W9uff2K+VyV9yretbSqP940Gvh+mF1aqjZ
LQepKG40dmusRnNFZcQTJ2Q3/uR3XT+OwoDByIi5OHO4HxFrOfuwL0klleX3GPhQ
yziTM3kzoSoCPFiifOHSyeAn4I0iC+rnWCZAIyCAf1udnMroJWYbW8iKiCJ4ACER
2/BQevEosSwnMnk1nFpY9fvHpGjyG20d+r/vTrtRoX6rBRBld0+7yiNPiow+X2SE
P1qqsyW4SPJ6yG2HetOUDvXJvL6FihWKrqw3hbqJPwF2Na5MRfetIfGfOxAinubc
j62/M9zFNhtMaTPgpnnz5NWYlSg27Z1IDdg8de4dRwLDbxLXj/ObWyAGvrfs9/jW
UQJ9vrCFoXeGMQfRSYCZdKOw1IK41cLmdS7rb/f5yf8p7L4lBflTInT09IXdMgqm
NMRRtI6IukEiEzp/h+b0zyNVitSh1XWtKWHtm36qFOJayktzwLLhYZioHvl9ofP2
cL5t1ig5Id+WGu5xm+yDb7sFVwB2bMg3sE0wCaYpk6QFIBAq043YQCEGDBW7KRQz
DPCZNfnxhJkF45RX/ndgAsXHbG6H4EdHTZNcOAX4yk36bosnMDFLvVG6/q7r2jEy
fLQ73WrX2v4oIMuHA1c2DPu1aGTq9ePQoDhfu9KCfMlTysivQDHqcCMcBQPNWAGe
cYYhmB6VTOovXbbID64Y0y6a5h7OjEfYDbMqLF6g4U+D1ABHUEfMdYhZvKk597xE
zobwquQ/G5jXmSVldYoTdpoxmb8SNiMjOm+O4YN+zvBnHxtjmUdzI3nkWDkVNsKa
ift0uJuthiOJsinFGumBQ0R6k1hMBCoec+DET4kCcRq02gTJeetHldmRKAdOh1yF
4alaatnwU+VkXvSCUn1hmMnsTXkecykVlf7UnX4mh8ctwffdtLpVTX04zjfyrMP/
BFZrlRzcY9TyHfupt8QxPK6tOZPFiZwyIfNoWl+zBkaM4/KplJfHL6mwkmSj1giP
rVARMDQJDEbghCqJJKkSVlC+Xj7eqAbYMxoN/S8nK9qLgeS433qVz9RwpeQdEPjk
2+nPIZDqYyQxsHp+lVlkAT2vBx5vzC7DSSYuv3XWyGL1OeTVeQTNjoD3mdkHTCQq
1nUkjUzGvUt9svGn3LHnKSpKuH0/isgLLVPzIojGr+J7RuGYVOmY7cnkcoqVvEe/
yVK6SdtxoS5wHyoLEaHL58QEjYlV7nfrr7QnM77DxK8hD2yO5rvcBmCVIhUoBX6r
jw1SjfaMPohZI4fMm9TFwHE78xNkgYk1uwAwtgctOocHT+P8QuSmEF5F/ydqhP/2
G2KcgTg9ESHrbx0kdBxcSBTTB/hm/DYzfAAZQPkHVcpvVforUjNNytkq2iOtruF5
hOiGzzHizLdqptFa06Z57o2se53qA9XWRWWVpCyxMnJUZ8j6m/5VwkydnVcIbpWG
AXcCT2tELt7SZtQ7w4cQMiTN3R1VwDQMIfiWR9WliPv49A79S7SzWcGAjo1iUgDa
Scc/4UQM/pytVK0lIUbM/RM73LD8Pfp1Xm28Tjy3e+k=
`protect END_PROTECTED
