`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CaXvybP7wijMvxJ7wU8Dupp6n7Bd6HtMwg4vDR8mPrdwN4yPJORbR0YHCnFNzQbG
Arc4wWvcz8EwhEF5S2GMS6wVIhAxp2k5qbuWF3U3tIBiksbqfjDmYkcSerYm7S6g
s1YIzObKzk4Fbb4r1dk7zE8Nu/nu7AQ7eTmHLhTSq+WrhCrhVzPp3Bb8I34VN4BA
wcvtZLLli5gNZ8Ypyj4V8tFL7wSjTGIsJpn6p/jkAzCoI7lsMvVNgBh7qR8ZAxd0
FBOxLaFpEBEmnqW5MWTKLs8HOJSUtvWt0dwnR6WMMnPmJU8DIT8QLbhw9+eL5eKm
6iZKqkNKtZ0xsIkV7uMOIMRahR4tbtt3Unn+UV8kn+csuJ1RKnil/X92g34h47Sg
172R8Fm9d1qumDSMJvd7+5CAEpLIuUWbujczK+JD3dL5uphcXFrGG5TEzAbH+Xxs
nn1XJjNmetcWTplz9dWFaPxk9nXuPyrhX0mqtbIFlNhM1VNFK+NDzyAgEd0/tutn
+LJA35MZx1MpyYut6YSrvFubBPRtsv2NQwyD9loAdxtVQBipK++nQGzdJMyraG+Z
uAOEijICLsPau3qYMA1UPmUdj8BNeQvHEHQGU435UkqqCftiamGJH5avdBn3iJ6D
C3+r1tkTU9Wojm/ynBsaxJP0gtcskikHsv6RmIJHyvCt4ne998dYdsYtCCTw6597
oTQE6UkSmC1g3Zog3FC80ZMl2GRNZK7RH3ftxMXEl93l3pgVdMp0u87OLkzegtba
Z/8ganK38rPO2aIHTeyhArXERnDIskKUxa499GD7zMpVqrGJGY7sacCTtwf9GmpY
Nrfk+5nWS8aDmfUyoZMwOMCVNdOFtBPhnEohOyntSozAO78AcWsmH2lWMP4pMkmL
JTs09oGBoVQYgv54QdJe519JFoj+rx/NGAb1JQYWBtcox95ccON5Rfqh3E10Kbb0
fGqj0p3D68zllAlD822yPLyhKOFPmyqzqsvRVg3GCyI44gOgXUSPPftwndhWrj7R
0RsDiotWAKXz4ND83UPpb9m/mHdAMWbO4sXnZ7DM9CSuV4ZV95Ct8OCn5tMSUFYo
sBEO/pHw6ahtLEJG0KpsKSmfqFp/r4cqoFNhc3Dwsw5N9WkOu+GMDgJRsQe33m+8
BPZmM2b31RHjsx6/j66dUztA+QjUaI37HdxJcnIi3iQE3O0m8rq3Ecge3jg8v3zA
FYhSM9RbCcHxdlz2kcQ7QjVoMv7Ic18+1tp7AypXkg+x46Cwe4U31hrzjiYHjTQZ
ZmyQRdtyM3JDTT0PpJ0W7+EMaDglpUr1PyFAY68bXTmWXxSLtlQ7ON7lrRhgmWI2
2JUo8ZNLnRNR13PIe2N1iuORwdmqBxXppqArB5qUp00iUdpEj4MfdaJfrTB06cTM
3a/VKcvfpR23v0CAm0JfejBBkXK6dNooPrnJEO7L8+L2yo12VlSw0siz6XUdSfBo
p4Qavt20N8KrHXr5lYLCWZBj3y7CTruzqFmEkGqyDsf0TQW4GrMiZ+hDgyJgoxDN
1KydfsEAfooQe0oqB5M3b7vSsWuA2oELi6pdeTuHVygd6f4nA4PlxbADMaoGo6gP
uciwM59rqMDNjG+ntAoevHnCnWqMMe6lPARTr9HpkqaqKRUDnVuQUSpO8kkUVMIa
LEGBQyE5Fa3fkTm3DUqHIvVNcscMBanLhFfzEZ9kgi0acu0C1jQNiM/kOLy9dywF
xo3K5EBniwFqOgb7PkK1nNFeQG3rIFTV3FhDOBRvsfRd8cDaYv5rcr1CcZye5lle
+bRJKajJi2nJj57raFoFjUyHmNrDEG0IlXPY22RYX5NxJBAsshQQKG6bjfLrXtK/
mEk7nT3SKBTNPXWEI1jd3WGLopMOyLGfu5mEBO5jB/03dlO+ck4ePSZgiqIjUNd0
Lm/uvRocrVzFbrX/EHb2tqpYx9CWDFnnDx1f7ZOZjHFrQUdhEC2+LFmQrsV4fHtj
wwC3iqKgBuQ1de/ZP0yydo77GwPZf84DBAvuVhqNUTaWL7FiLcTgUP+havK1Q2Re
efe2zH3EBFt75EgtY39L3Ms+OGxGeAysWsYyfpYM+hRxJqiE2zIYWca2XGdPMcGy
kk+byfhlXyvMtlyTlTTCVmoa/uJbrcoPmaNjTPxQ60kXVdByhU8Bel01OjJ/ihQ+
4Ixxk8gfYlkQaqBMw9dfJ+sMmysw+B6fvNVZ10HOPto8PUQequhbrgGC7ih7X70G
TBj7rgZhr06IXJeNDRb5UeHf5QzP60UxCZdRE/bx+joQK2T+WQTP4Id2+0XzIr+j
buSczK++rI3Kvr/d1ykb8IEguUGcWv2cs2hvTTy1xdTejUnV/RfJf6Rs2Z3uoG84
ksLN3osuRHBTwBau/7iVABs+J/9+2poMTd8s7bJmHaW+sD5ehJtSf25kCuGY/FkW
BPWRwvfhrM0PZgSUmEJNREZIBuw1Dxry3ce/312adluS+v61P+ryqcJ+5FiqTMqY
p6pEGIIamVrPtwSr3y/c5e7VeH0+sLJW1faaS1qoKUld2PkJRdEHZx/hk85odOiw
AtRTCNOo1k8OSoSR51k67/krH5kyek1URRinbP9lGDgqQavWhhgXKeVPCbg+FnPy
JxH3Gsy7CmLpf78U/G1fZ/O4151GSV5Wi1AJAQ5ATW3SqqwPza++yzSLxmu4+gPM
UdBO0ggG1RkYZ4X5RgdMty3tAZwocbiW5lUgdgSIJyhB0IAcY7bgfUJVyKtQnZNL
8jnyJXeSqcvxZH/dqTt+GfmA8GWO4NHN1kPS39QtyVjFwTBOb9KE3IPzTN041HsH
K5vr2fQPFXF3peu1t8q1yRw+efS83oOShEhrSx5MOKxPaoYKoNbpIcl5dzTVFjmr
RQi460cqiX4r2IUb560JMV+LWh0AkqmWvcC70VA61W8OdEp3p4HcdTEJf7YT3RH9
qY1hmTmYv4aOYW6Cci6Zyqp5TT5hTawq9Ady+4sXwQPB4+9a9BUrgstyDTVRofkk
TmVBYBlSuB3EEcwyEz2z17yOT/lZb5JOGxNBsS/YpljWt3wwyBr2tiLD1nyXhzb3
50KjnJPmxZpTg/v/0zvCL1l22kVKRXPt3nVXKbvixh1kyCc6bXky72zlUsCaQyqU
mJULDhl8MJkyvo00Pt1RrYOPsow9Q1VMX/1j5q49b/UnYKK/B+C6D65NJP8c6hFt
mQeDcuYkkQO5rU112azvpJRwKcOM+5fDojL3mTclYneG9zj1t4hmB+xBj/onrfG0
fvFBRqXk98ljbdC4GRvTd+944HyFC4zAQPJ+5wSO9J8doJtXO5nOzyby5JGcFscb
PthrjfMD/NW2y52o8Jm0gy1ueia49TgWrC4Sae5lAN69eZs3CgjAhLUHkTkE1HME
yQgTZhoLvmCP6DjjzNJNrCJln7ksUcULFHQMvgCTP+1QzkHGiXOQxxb+Q9RrmEy7
mlaP/5yAV4RbS+H7K0k63FAdJPbiCk3Ev/WJtsvxHs1L1xSBGqM5wb5YTF5oN3eD
yMrmWkKDKsF+e0gZ4kD0jpSR+TH0L7mifVw2V+/CWKu2Nj63iw3Lfe73PPE60zn5
/TWcP3/roV144ueey9y3O516MH7zOF1yFXrnbB8i5TrnqB4Pn7y59QmPAmUakbNA
sYyjJWzjq4+qWDiv4f0ipNgDb50TsXl9D3+tBNALsyBJITsvMfGxh5ru7OTLCc2Z
yTL2Gj9DA/4XQhHgaodq6g5WPr9jivUuh5FyDdKoP4IODXcDV0Ey8/HqRju3sgnq
Po1z8w1dl4oV122cFQf2P2yhhwN+z1Rk+tWnyNKJJl3moFWZg9+DeLy21oklphFG
iuBuHayPWsDE9RyEckzbmcfJkRlqW+lyDe1PythCj5slZi8d+/Ou7yD+hAw709U6
BShe25jGXM9+uFfn3OC9+76pSiao7lxRYgVHZR55XbweDTWUphbGrRA/L5i0gpJD
aWWkKGOLU5PWgTiDwNtTs0TWYW8/gqSFWbOnDOoOdGz9gu6nNa21Qck13a5w75Ly
elZrWuJdk/nPohBE4pHCjOGHSaEkP1B+hwJxSLxAaiCva4EJTHYosdnGKJFNO21O
5tqr5uzxe0voehVapUSXtOGm97AmRTcPj+XciohvUeA5e5ZPaPoOzZR1/zcRnHDO
jTAW14IHmXh/Sox/IOTzqLSxqqarOvklsWoC337BlbPIZP+UUj/aVJp8qjP27ibA
RUEUn8T4PEgMoUmQnM9rCumdI5j+qz6Tug2Gy0yOphiV0IedDDvUbUTY9L1kIBCR
gR0TStPQLkKeu8Tng+gL6RmXvbS08otWadYWVjlRgPeetmHvRaLwb5MVsk8S6Uwf
wb5xFXTV7JA7/wxybuk2IiMh7vcw9gGmCaZxwd3UHZjz4+GMiUWKVDK7Nurhj3Re
sEXrARjwOmnsatbAhthl4WPtpjp96vIkIqe0EIcalwyKrjBfrYWCUunvqeNloR7g
3EyC1HenegFIGkv3H9gpMYAHivTr9aptNnZBPZnjHk9xL4FBUPTekkYT++HmJN1F
qVOKh48RX8HZNGHnmTkAv/ghc28/yRN0SJwvi+FIg5E4TNTHuATnvGIje0e2tl70
FjIXOkpKcc97tqaCDFTKkBi4e+6VgJ6J8MgB2bGhVIo/Z31j+UdjHBDVlRFQjnuX
BJhcpqFrl1rCKRWcIx3KRk3+4fqSKJ9LDcSVn6j+roQI8rAwBF2Dur/g2giOuyVa
PQDKhPyGX417IkhH13oAij03ZwmhDt5KkPMXdZpzm/s4NmC/b5rMZinaN88w844u
bEmInkpzKRXfEc6Y6l4valdStYpnGq9bP3F4BosGeGWFI0toxrZN+nt7b35bIWjO
vh1jW6pemvvSqAZh41J1PtXH+Kpgf6Fxl+5h7B67C/OOVpLLQRe4oNUZ4WpfuKO9
3jKvQvPzoRNIepsO7xn20NmRvcpwf1WJ6acYlDNiZI9uj2ULACvz+b92EX2R/ufr
aJVmkhrVySll4cc8pWxhASbSmn27+HejYnSqdjRxuR0sWjjlED5RJWm9FxHSboMV
NYwpt9rOCGFCXw8JTYk7ZU1Tik09kHdGAjhgp3ShXmUKnSsi3Npdywsk2wQsHb1Z
vmFE8N35lITdDTtxE7wX/A9eEBs/EFu5pPztTyezp2qHr9WeBlENUXgIJ+d/URYT
kBoPADBHvOa109Lbmg5mnM561jGGoHPfDQs+EXHTx4Li2GwqA0gw3Niyzsw9a1p3
uu5w/j8dHG3YrHONXrIzb1IFfhmW68aYkU7jlL+nYVzkK+nSl6ZAAdxL1mKIzqc0
IkkgMcirZ5NlVhg5ZDtII24NBvJ0W4eazFhAlshTZkDjsC6Wg/hslIjjX6RfnTmx
CfDcEEi9ns1alFD/wYnk+z/HgIt1LBEVzWGFIjN5h0rSgtT6CvCYmASJRbZDl6oT
ABQ9H9V856NrNwl8Xa37lCetKtJ747lpacm6uoWcj/bUmyWbPAsfdSWNFpoAR4/o
PXzVe8mL/3bLGkT3UGJZQV/IGiXmDiUgdQqTaeQvvl+G7Jhg4LM/aQBlLwfocAze
2GZtu1OMCfsA+MWcS3nK+b+ffi7kQ3Je86AyQYEU0PlOcLEo8V+VFsKyP9fDNRWR
5kh1xYLs9YIz1OJx1YLegQiMwhFeksdCaoU8saGYGaWp1K++D7sI/Vm51KKzB0Hn
LDg4EftuTqgL/MsdWEiUANN9K1UbETqN2ai99zWkkbuFJnO8wpFu87OqE16xbpGg
rVfYs/A23Oqf86J1ps0AbGBdW4whA/J346ootqSJzjElRPpehzFiiKghi80CvqqW
uPQF3LGyiscny+Ey0HBMmNpb5K6SdTX+GqCTU9MwdU6EBZwqymTap2oyywDUkjCu
y+LewQ+90UBZWrDZL/l+7qki35k5T59hn8cVcIN8H61URRK/EvW+3AGFHQEbWjXj
azPaAc61B1420eVVRtwmghsmVsVAD3AlDIomWFafbYrivoOd7dHmdLAFAx1jPSyo
Dcy+EsLQresz/xrlhHATWdnWA3W1KvLI5AqaEVYJitab+gHVDiVpcco29FnqmFFZ
0imgiqc/3rnNWN2Hvlb8TbYPJ7H4IHBGA5xmOT28EuqEiMTErruyUWQESr4U62Bg
Nra6bqjQuMNOH+n43FE6AgCbO00DLCPoGqz2id1sK5e0O8uS6N3U4R/FW01Zg7Uq
jGv7Hwg6Gz8p9l5/Ef7YhAbQWiAWj1p7e0y5a8QHiTMsfrksmsP+Uu3do9mt46cn
wpnTJxGlcRORQfjSU0q+XoRFv7233nhpR9JzmySQlxLJjPl8yzncCeAugfWYKM3T
jSU4drDPlBbmlRnwddq2dlpBK1wP7x2XV2rQygHBcSHv9aAj6ar2NS8CeGOULqs6
1NDYnecjoKKkVSLTiDAwm/JXIyXPn5FNdEkPmh5uLZ4MpnfEyJ+lmiOrztmnWh87
mZY3F03DdDqjfaxqr3asrYga5aK+mCAAPIDp3p+fhtdPvKtiE3X7DyYQa9BY9gnd
umo7K7pzFqHsT5ayaPLAptQYYmQrD0k3k+HDktFuuJkgTa9xOn8SiwUIGEKaUW6X
etogH9b4Zd7+IM3kaJbQ8lnEwj+mErBFACUZ1meb4GDO7Wg73kkebUI/N5r66EH6
bSbyf/C6okJt3lSfBozKKxxmSL1Q3yVXVrvK1pJOzI+aViRgEGuZ6CNUcGRA372m
a9tAVi9+cRb57InDJxCF5BP9zCq/R9VkOKaebFO8Jyfoes9tMJp3S+b763g9Tciw
rMvnRRZQHAa4wRmW0YBwrYaCBrvZkscVrYr4Vhf1IdOuQnt2/J5u2cbHe026NLMJ
o4MpvtRGowPCgHNNmf7JF5FbgNmwTOF4cXwMWm3ib2ieOFjQoyL9Bdl5cJKmpaIx
EWXaTwTV7HolbZYtBMSeNOTFNj5UlUuIww8y9YZpnH5F9Aerzq75bJDPZFdYQWHG
peFeXhNq7hbkNrsgFnz5OHuDWYMQfwI8BtPJyTp2Em3lMv8PTFA4F+y3jG6lTTRL
Quet0TDu1R5eSe5gPsNYZwjHu3sJt2FoB0WJnvU1haUNsNd+F03kp7N5kkRNS/GI
8S/cvDAi/SB0hD3LqC9DlcKYgpYbtZjC4cGYVQiPi56AYpOdtqmjDrZ6BeHeYRX2
7mXBxBPZKSu1i6pn6gj1c7OkPxmmx/RGPLUsa83cHkaN/+aHGfSWf8+rRbRuNvoe
/osgyvvAz5SluRkkzAFjBP96bNcE9s1oCKpcH+xS4qVJEK+sR3DFxTpGAWG5A4HH
7xLqvgbS1lDVop0T2iGsZkv/A+aneNim3oDycXrP2dVCmh7VGQ28d1THE5R5+re1
scQfwN2bfzwhty6SerS90Bcoj/XF+mujW2ERPoEQ13jozA6zuWQEmuB2e/BmEx0e
AdBoAlVGdoY/U1DczxxDYHge0bUKCoAE6b7yhhvWl4BjVuPSr749rN3MjXKUC7fO
1SffUvH5LVYNPSkUji5ldP1Hkj/VLUneACDC8XgT2rFvAvttj2GIjrrMpTHXvwTB
rbIWyTde0jr3gUYr8Ww/7qnlqFpJNROJBLvFg+4uO1oxllHATsJfSKi/R3joBFf0
8TTrLyMGb/VwcKGXIAum1nZ2GLpYAbeu+bGR6ZOcTstqEsOxllTSdLoz++esr/Si
ICmZc4F/b8x5SjzHnI9aj3VyNs52Ujivnc5ByV5tu+672ujvF//KbRUh7oXrsExh
CAYCbkNwRzldcLjubnIUsNe+bNCIXfLiOsm7xRHuEknhJk4v4oRfNZnVzwazrEpD
XNvddeRAIOvQv1rFr9s7WMcNeXzhaSeEcyGvvXd2MX6cHJqVG7tlCr4vF1A2uPVN
7m4zSMDLmIxMUTFwUrbuv+Y+9dqQ4zbD8JiUjpUWSeKkccnEbT4yLljgJ55PZHBI
46cMnXYdFsspmPBes8n+aMXZYPpWNmnZRH12RuvzDLjOb7708/AJqPbrjJ4tKBAh
x96LQ/fQ2v66b5LwmNhbCAx6qwI61sDDEgc/zjctHwNtcgrjxEw9uswIOyd7LToI
Zft+GF8aAH9sUo+RPnoN0CQEOW9+VreMPvin0o4GTmeoxGaGoN4TJwE5wotfPlLa
tDNOlXd8KsEZ//NTs/JsTeK0VzpSyS5prukphCqb61e6EV592e80gz/ZPYuPROdn
lRhWpYJS0/2okudZJi5sGlpcwPEt9ro6TvhrEXwGo/XpaWAVTwLy0IE3Y+C4ZGT/
/GO6EJi2dlPh8Ugd3H9cgYjeeZlwbVDwf0RpBXgjpbgbb0F4EYfmaqTWl/SxI8Th
SDJT1039To5mLdCQvrgnZ5zgEnmve5yMA4JUcKpHJPGqwPlxszNhBh5/GU+lIYf/
gzzDF/2Zz+ru8tYCKzevxkmKdwQrIhNcLwYAfKyXyL4jttXMA50GYkbKs9vY3bNm
nLz9yQlACgytC8L4e8mPD0SZNDusC678mdpUmS8unCDa9gqVHte7c1LCkrPvt47b
rF+lZSI8W32FN0tc2uRO89R4MBWvB0lJLy8Z5Cc7fJeJQvbzNApqLSXQAnNxE9Rk
sucVnYaJgsq626FWF+tOm4hgY2X9aHOaElxxoJ/rhzPA5i4nrWXumAf9VuBbXETU
9tMAa49jz68C0K6f0MOTGdbn9a//p/9miHckXf23pIrnboaUHaGYsXRAZjYAIQF3
m9FrvtH8NK+gpsKiIG0nE4CL/bOLyQ9uu3RiTGcs+1CvTf/Sgd2I5kRccj8JP+LS
2FxEQMSzFwss3ItElc69SetDQQrgmCFdOgWXRUEuNt4BTUJ7aa0RonsO0/Gsi2n0
nolphI4DWZJRmrZPmBSubFPwujE3JmUni62Ibh+EQvSf+R1u4RqI7S0su4eThwiL
NuTnoxoTNmetshSoMItgkFuz1DxDW0Q5hSyI5ZMBLcuGsyqOOQj7D1njbD62Q2Dc
yB1w+r3v3dp7QGEwwOk60N2XtOOoZ3qaLcaKascPyMkj0gjv+v3ukpyh2raEsczP
nRJfhZuXujcV+UhmW8aALxq5v0waxUefjULmqlvZn3AYV1D21uJv5qd4OLYR0ZM7
S4iY1V3RIhHpSelWSA01uF0YB7pfjZDy4V5TcvYoKAMshSu027Ju9O61JZgvAq6s
6Sm7RYKjdo2Jh9kZx0VuYAWWfsZo28QVU8V11iI3C7LqejmyIREtQiz3tqoXTaEb
o26KiyTJ4l+zt5EecW+ebZ13hdMpItyDMe8qhyV0+S1AOiijDqobayVaTNr28yxc
rG6Q4KeQ4jvquCkTk3FDQBmRoeSB534b2GqG5ztVfCPccUEZCL6Atb4OXE2/Bmg6
VyliAyzzK/7iT3+wj9kvTTcazDi7xuE5r26CuSmNw5GAtaVngo5K72rjgpYa3CWY
O6sOqU+CEJtubsY0vQuD5AkEj/o+gffeqM1pijLnaY06yNZAo5AazGufXIiNFMdn
M8RFKDgQc2Yt28N0rid+G3eqBliqODkI4gTzaprcutgSHWPP1UKY4tUX9cACEqj/
lxJ9r3rhkC3NMRZ+Jg8QeaI3GTFK0tYGLU+q2wM0O4OtzKfKWas4x5GQ4Mnuj7c9
4fXnNrEYwtLiOXTB2vrOFANds5Gdy1AfafuCimtHkMDgWKElr45JMkTQRVR+8s82
K3bA9tEbYGVBmaTmW7Mx11rsmvLd55UeBXjnh7rJ00gOC4ssawsiN04llb6jHXs8
VefkwIBCH55cJ7OG6PQoyexd0LqqYCG42diwiQ2EsnPk6ouE6op5e95vCylAGmPk
qcp61kSPHN5SCS/tDxjAtVxRVT88oWHAjGeE1Y/qSpPd1hfDpc2SVJb1ps/NOIyk
16td7VDLLhBrcSyYQbybGK5D3+2YHj9qDpHA9owlDpqsaG6vb/Hv2M9aSkc3DIJ1
aMfB8Ms5aNTNTEETO3xl3fkin9f5byxFJAutxT5ohwt4V5yDZMKJQzCwD5/fyjdt
pbPnaLCshoR8mWhOfAz7iuPY1Poi+NOOOPi8GQnJiUveeh82wm2uelmSYCsnUWZ7
u0G2jhX+r0t1FB5xjkJeqt8kkwglyaBfHEh9+rm7H43wtFQsGE45+vcUoHgifjaw
PzZDgQtggv9pvBkIJXKNzJkPP/hmvn+XXhwZWwvNrCcq6iQpGNfLTZD44xD9E1So
sdGNVIqlJB00zc1HHTF2kLDb/m6SlOb44UdWIGO+3BU0zxm4r20utoyr8/QPJRT6
vQqwh7N9aPWxPb+iEgSrdee4UL1cipo0ZRzEWIOt6OhPHinOieoATgMHR5lMfG9F
xDD6CeIeojJvpoauyXQ/HCDMh/Fy9LMKCjOXO/S1hrgUYZkHlMD/QEF36UjdjG/v
BXmnh4MCqkobhHSZF+szDZAU1onXsGOgLeF60TFnkDQfCej5EbmLRRBezsDoP/MV
TWEKjrS95l+rFH34Rx9801x+R4HstWdlOKgUF0cJS86rrtjB846BDRKtWwsXycy3
08C8EzniLaT6FOws+TpUnPe6fZBmxQCY8FX7JzL8CPTXyAmPdQea4jiHAPOO2zi8
I1ZBKYtSpMKZTv6RV9baYMe9xmaBsmskshL4Z17nYzSW/fGYKQyvGIsRHNvK3v0F
rRtTV8fWRJaQSo0TtlZ+n+XABLcbEhHoo6dW3XHqPPoiERC6OcF/QZXoL2wwEzzY
kEJokZo7lxhTqwcLH14DH5UlW2xsmqvF4LvniQuLccoGjc7830Ek2IB4e2t30DQv
rYA7u7jaf8FaKvsovoLi+KO2vOTa5+YWdGed9f94eY4xdzgZBPvV4offlhTEQWDd
C9mMivdMJyrk6GVSyjapOMLiMN/VfBXLXqGvqJ04aTPRxCo4wBBOKnbudAWAyqRM
pCed8BomHKN5t4YO1yxZo4d9GUJ+rfO0hzlR9pp3j4GqwVIRgdUWwLLykVR0iTgu
7G31IbTEY/qz2Fxdn4poRDMvmNbetJqaMYn5W8DUijKab8ZIWrrHZoN2MdV3doyR
bpcDM5ZzRwrhgWqHN95RoUh1mx7SDvV5G0te1RVRdVX0WpT2q2yys/0Ck/yasx72
RuuXuLLjY7G3wKAwIbhYs4BT6wEVKod4VZeFY8Kyawn44EbRqXlOgJqT7j/3JdxE
5wBtAwK7lRBwkrzLvpjzZmHm90XCCoU+nqlrFSM/pxjNk6l1ZJXMTgvxOs7300Mn
Du7lPoO713+dQBziWcpriEkLm33IDHwjR9nU22gG1S5+ToneedyEzMQh7bFYPzI9
c2wZjWr7i/FxCebDTa6vCkcUv5T9pPsMc+6VU97rYQyNRIDKLkA7We/kvBouPPfr
aqux941ePmlqQ0/RmO30l0GORCQ3xe34vXXpn8QbtCdQKqcyy4fiayeI7fzJrX/n
BZg0hqbrRO1lSQ4pnLQgRF7NtieM6Dj8abAHKUBB4EDEjVyEON39buGi+C1wqGXQ
FJmh1DnFfB+4UcDDxuBgMO+iEGaEAwnh/Kzh+g3WM0QvARf84qoDOyYOwYxQMWFw
Ir7gy9dTCwUfXw3VSFerA/Hg348jcwd5y2lEX9IChnAa/1l9grg9XQSGUOMsLI72
7IICZA8+lYBeetTkn+lEZVjmRAxJib5d3N5GHEO5cNNwlIJDzSKnOTUoVBn5sq6I
dWRIilYSlijhlBqOKG93sssxhDk9u51MLdqloiUI3BVSycpw35lNQXYF7NsJ9dex
R8r6iXB95OHEU817dx0GtMqWdMqK1U0VPfCRBihwa3n14SDo/cMrn0QftlOTS5Rv
iuqHOr+T4SztdxUU0frW94cfPZk9XAH92gzPlu5XOA3TSOtyPFbP4kRXO1sgxuER
PJ2NjGD0O4gDK/BuuI4kk5eGECHVLO9hUHTrNliu2Oo685zdvkctDZK6mjbZ1s0x
Zqa2Cd+WcNjKnreNzlgU4HXtgTLHjLIpt9T+kbWAUdDsQ2+fWReEq5cMnY7E2dWl
KEQ9+T3Rs2ddk5qEfrdO/6WOJRoA8oP67I/h6bMO8o+UUCaIkEh/kGbkBbpKO+cP
pLUJT4CZGwX5TAdi5bgwHIUWV+fHgDWa/rBQWibfbO7QRRrre/0pbr0sIlae903C
0NkaaFP/zW83fUKTxuxxLsZYrHwywDvESNMSI9qCdgjkerUja3ksUOFnsT7/8zQ5
PiC+AsE2F6k2isgwZP9EFp5a2pAWkDoGYUNZvKNhWFTDru1gae0SDgH1XmN0A1cZ
d63+j+qCNHZ8EzY9JMBMePEUey4aWsmK1sojomw4fqC3CFr+xfKMT33Z5aSnMkTS
uc5IR/Mu6cXFVaTaK9WEoxCamTITe6x3a9ADgPkoS3sg1dsqeXHESNwLroWfHMLa
oYbTaAktIN76uOWQMK4j2rxPIjyodtgfMf7M3IhKfKNBJlRDJ1itmX7IIQX3C++p
s7d2vlNHg2T30tCH14/rTsp00qVR9RBqdLKylnsliN7rldShbrPrT5dL+E4o9Tek
UaxZPVjeHoNsBboR1ymRF7imLSBX4Ww0R0elhc9WCyoS9c5fnWmD8qHFlzhHtxco
/tp4GUjsoDW52tgb9uVyFvyW/rln7eIK2XLiAS9Z6hppfBf27bTUyYCAqznag3TX
zFDPVvaWiC9COVQ5AbJXVRsFkn12/7aySHta+Ohl45jV76FCbRa5eTlYPWAvzMGn
yrVRqU3Il5BcDGRN6p2gDK+sQw1Dc7DoeMB672QT2nHLAzNuat2ElZBEKKIIEMha
2Es77BvYGBOJdkajhIWFE4pcPtYhfWSVZlWIbk3RmZGpDZYmFe3A7SfDrhWseTOb
vVCfxfH9mfNfFe2L71Qc18pDlc4dsDpR9kXMj+T7jqxKbprIultkUfF/vhktIxZC
l0XbpdbizW3DjRPMVLTeGXIgQShy7qxiMbzjxbG8dYxM0SUT18OH1xxBWwa1KjwD
I1hw0uMubBrWImUIwtBJkNzkkDr6bzVf1+lBOY3zyZGbN7DCU+r82nM38Nnl1aY1
r3dZWw4bK7NPrh4pp8D1C412n+BLjGdr3KgQOgfkWyJ9IUB3YjoS6Db7Q+qn5ilQ
xnjmlqlw1ZOC9Il2MJHfs8AuBHayVrlQSUH9feqnXRju22CKiCN4M1eXRr1FG0Rv
SV9Yaxovt7MwCuzqD83b4ew4KohnUPA3sk5mdNU/fdtazT7QR7o+X+DMFloyqPpF
bfVePmlGuTRZHmYbNMqyazGjoo/DL90e3NUKFfoByRun56OW01Dret2mSDD44UMn
CA7ps9tQ2/n3PwXqIIJFqFFX2AqRtBfNh5LVHWi7/3gp/v5OdobzViFKRYd5TY2C
Y035dxxT12KuZIkjiEN4SvCddkki10uI9KY+FCNu0iXkYNYb0M0mtiUlbqTcrsxy
chJsUtMnPi2Z4BuxXnMQZCLe8fyipXChQyp3qsdUzdIGY2+IVvVSZM01DRcAp4WE
Qde3ipRilspfK0dhDBOgzF7wzRQSzrmiBfek0PWcDpmeoIVdXU1vfsHEOUXW45b+
ADWz/x0+srXW8YTRBYjJuOmDyMCNQrogZt3NmyxZth/P+g6gQqI/3Xr44C6/pXFz
+ywstOtzcfnztRcPB5V1Q+NfF7RCTsmiFioK2ey5/jWwc2uPNlozBB3G829HRKrP
lx2RbdEerKH7LH55pW8mqANF81OHCbClIa9O6VmogWpOv+8n7nl9Qxb46L1cP47s
Vig3Te/dR96e2jN8h6o5IBWfytIEVEBexY2xGUaOAbvV/uFCT38oMVX5dJBeHF6l
NxS5d1H42nSkztj2VxPF7tT/HVRWyjBTP/7cwOppIh3GX4sjyBdrvNwuFFAWOpw0
CcvU5Lu0GqFE0K4hYnhu+6cd0kbws09Dar/1TQCCE75tk6IGqcowzr2dsUgjB7L0
kitwZ1WIOgowyZNHHEs+LF/V6bX8cPYAS7o1lvNC5klRVaNeHt9xAmjPqiy0rk78
U53t6U8umsf3btFR2UMmildkF2236+4RR2v4Y0k9RoouYwCWNl8ZY2rq2n7kAGj4
7RzjWXXK835YB1pZgylmh3godK4ZUvNPmqkYBiPNP44RX5/ppcbkS7X3uytXQoQV
lrLSUsBqfDsUl/WhjRlC138ThgKYUjGopueDAmVkcCQkdY+bq1TfoGnzAJU20ZRp
pq35/e29dH6eQxZK5QBybPcRhHGY/KCW29zJLQJ47urozCV7T4byk8CMtd/az3zx
dvCFiDkDGowM2ekQNxuwi2B6YNQNP5ly6zqGR4xAoAIy+ZqoLQ5prZYSxU8MdMzR
ML/NgRq8HALf4oihmulqg80wISJB+CbtrherEmLQlN02203aoZefSMlGNyPv3l8h
wfgusAhxIN5NvCHOTxe9y974jFMcffaI8Mqu5XhWeysLG1e5kgQ/iU/qmBN8qxyu
Cmdsw/Eehgnnb7n9FfyA5mYTE+Ahkw7FXCicI8KdbjeJ+Ql4IqVv+49Oz9/umucw
3IAN4Eu9Y3rL1e0oCPnp7ewElvsUG1ed30E2c3stQ4l4epD0XxkryHsFSQWIuxbg
8dZBAFHcWM+XghUTHtgirtpleK7Whg0DHfULXvkkFlDG7wxq0y0voieEtNskgStc
LA74R61Vc7eOzt758EKYyYQIJVFYfuLhTXINM9opeIURCG5+BYVAt8D/MitV0OJh
aktBSXMzO74v0KV1fu6yFfRZCE1lTzunK4nzMmQ/6+aebmOeFHoJZacWZ2F4OwVx
fIDPRgYXgbrYOn2AgrG7jmksQqSyvsZvVkBBuoHWrS4AAN0PmjsEUSOOrQu/pVVU
A11nm1fjSswP7jfdsJ+lRXGz2um0kgbMRwpVlUwI+zfPSlHpAGgDU6zdY7idzHdl
g3YCwwk3bf2G+rov9ySlkbG2LxrN/XiBXlYfbSrN6CXIc1lUvlP8RgA127CcvOT5
jN9HlhcHdR6HBuWAawBJ7F7LQe6ZEV8Ntuv5ED2APbuBBhPIbvsM6WnF4VKXrcPW
UyEvJB/ffl9HK0J/mQEDGWYi3/f84yK+8yDK8g7aUGtom+pNO1awWuvodZjZMy2/
vo1Q98NpIjgtNq4wqf7RTQ8jKgqQsctSsTRR+4fRazVDxYTd19/hvLc+k/MqpnWx
7t/ETztfeV/QQIvLWHZ/WIxgJ6AIXK89AQwHU9RnmcPWrtIuW6/vwOkHB9Ll5gKG
h5vuJwuYkdcr3kTQ12WE42EyPXYYWAsLwnWTMrSIGUdkURZf6Tmlugtc4Z/7swTC
nVaEediHHZZZ/m6JVM0BvybBDU/2DE9Y4HLkJBWc+DXVI44pBWUY5U6tmfd2caSd
3snZm8+5D0WPfWoF0DVnaxulE9zeHV9m3lA3HwfZ2gqu1Pk62hkCUKbGZBlN9BG4
mwAtmESFBt0mnAf+U05w/l8tGTKrBFfqWxU6/C7Mn5vQE7mHfu+CfUvyO7eLCQia
BAJ6XCcJmrpcJxO64n4fLNn8cvhVB5VfKXVN0Ib8JlCyCJNokOkERMdrjw9G2PYq
3XhqH/8etq9IltZTORkz/Jo0g7uWfj4UguPDKteT3dmyKZbMQqWnAaGQ+7StLcNT
W1GgND1rRZQuTCsvmO6oOa+leGvmSo60KcOOSPrZgHmGh/ufkvXW9uflbxtRnJ7w
K7rTRzcuOil+vzvpugBJ/bpV3dmXmsmF2ObSGxzBaJBSkPhteUlPOWeFDTjpbdJN
Xgpvy8nuM7oyfg7ebgOErRZ/DbJ+jEHeIJLF5aG3kXQ6SbIN7JH6eO0aMC6UF0Q9
ynKY7mGtUjdY2kcdqdh59/VN11BcxyAWomCeKCxC/ZcKGjKJOKDAjzKc7kA3pepx
E/ncx+JXzaqscD/rYnsWtkr0QZiFMfuMPmuw4hh4himSkKso8ZdebSWvZXCWIrkb
HjkrobRcTYNupSLFs4ezPBbiEFf8elBPJa4YhDJ970HrcN5Mc5K536s0/KYzsdvi
DYQy7ajkqu/pSfFBL8DAUFM1odeRGv8xTaEpTMt/po2HV9JRhxldgHcROTB5dy/W
EMQfKYpeWFBeCHoLBIv7YDVRSkIpvjBSIK2Y1JYMI2rrm2Rc7VpJjt+HSrRzJ39p
VuR5bWM5D80/T6a28N1M1qZ85aZBLv1tZR7TUR74LwLcPLacPt4SX5+oZZID9QcS
4r5k4ntep+Km2slijqtAUCNTWh64aYgDawk10c30J3cKVJv6P0Tpa2WKn6HvMZYO
cv2OhIBOmKPBgK73gddghKh8FgNSM0uPzRs55YhoxQCCNm5u0MLxGvvHOgjR5lwq
i5fFK9JdzSw7JSDwX9SDbvcFeNthIZfU27n8DDtAptYHRx1kxRtFlvPVUah01P/s
pt/GGMfxLBuRNW7YiEYfd47zzguWvLn1b781Rgk+qCvkrLGIh2WLGQNc+FmXSCeU
KulxV0I7bp4mklaGzIvFgdzcSSfcFvKE+Bve0qV4P5mu0C5iCuHA5aNs8zdwGWYN
7cVNBerthW7DLknio9pKO0ITDFsFHDhEbkEXgXQL5XPH4V1Lf4Xqz/R4nZp/MBTf
kxdTQKOtuIaGkeZrLcMyGn+iyT0PGYcsF2sFAi38K857NvJWdB9VOnWH3IqYMtDD
QLwIk2h68aJTkhDNFu0QQ/eaAhswOfizqqcVVEpoGJxYlkzZhFU8Lbjdmql0jQLZ
99bgUJRX9gBM2TbIfkmyBR4e2ro6LGYrFAWnD3c15390AKCWsyFuye8COZLLsdsz
8Bnyez4IB9+uiAg8SEWVQaxtHOpC+c/EceOq+C9/n8c8imW6Si6AcsE1mSPRLg/z
T7uUCkNYft4TIRk8fMQs1ekpwdYUv8U4pOx6TTHcgQrwa8dD2/wjkF8dEfW33VvQ
qY3cO/+sYIudmqCRx7mEXtGIgAqpk7AAolrrVstCGTNjsF+H5L9aMk9aENUslC67
X6BtbwMMZka6j966fGzjgnh/G0+xolr7O8fL9eiwlWWmGSiayMLxj0Zj0w7ynYW1
+f1wXeGNEwDh3H52x5RsGlqhZRKyTp4P4iP0lvnoyNoy3hSt5zXzSz65CAyouIHK
CRJS4rCAM5Ur9h3+OR6xibbnJDBwdrcYEjwLEgpiemXNS/JjIVz+xNRdm6PRbOyw
UWB1Kb7u/4bgPa3YWVv5chZQNl5AmCmVULYFBH/aC3q5sQat3PQdO9xeEiKyyZv1
M44Kv34B9YxxZNhHAXLdRA==
`protect END_PROTECTED
