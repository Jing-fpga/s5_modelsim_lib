`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jl+XDt+HU+piaLwG6jqRvDXAHXsJGPdhZbP7thRcfdHUBoKl8+mt+nUduVzVxbHu
6jyBvGZWn0MdnSFsdo+eayVUpGHVHyNTqHeUemCs3aTb6v2Jp0ZkyQcgsjgcCT03
mqIQOTnTx2bWmnW/WdOdehCAf907KL2bWvFuusA924DLW/cA5l8PKgx4mA1+mha/
tCqV4E2TFt529MdfsNGsIKEF0+BT6Cxj0OgGq36XgSkKszhPpllVkvp4izbSaDY7
Coogdu4OYu2ZtipSxGd6fUtEB+QUQUe3DWxl7n/dQOzadxyVQmznyUvLjoaBcq/q
NZNceIuVFYB8Tofk//qWyNu7j+5VjiHg8cdpwkbn4HNm6fgq6ya9JpSlEh2ITTJz
77AZyJrNCc20VPFt/0FexQCqbPtLkNwK/Ah7/95qEiQzcVtl5xqAkqvTW+dN6i8j
mGaFuqEcMSBaTwieNV7p2BbeOA+baWVH1QZRIW7UtSvtya9/wV5g/dqsNh88dht4
9Ha/OgxE06xpfXvZZR/z+fxZfJO3NVPEf1PApHq67vSPxnQ5ra19BL2BpKylAdHg
jwStdx5cMOTrMd6ngxg0w8g8XmLeRelBpc7IXfAXT3uilfG7J5n12Olg2F6O0QYN
l/BBuUNsADpf/OKXmFSyNbKvwX+axibUAFU+wY1W17fym4aHjHtwocVlBEUfREvJ
iGkwzS1dXPCO/oFfXrKQIDqjdq9GJuiYiGKXgcmJ29XvsU56JTPEhXrhXhzr+NdG
zrpWRpUhOcNLYbc7owWqKhcI3OYN3BTUp9WzAz+IJlNjq9gfYNZHltLMKd7QHrxs
I+9j3e6udmxBvfyFd8C/SiIL/ED8JE3GNJ70EZKammzQ9xksffkKmx9gbyRPh1Nj
lj4gWELQFhsf1ZtjmbiEOQW/etElLsyCJRL6OuEepLF+bIeEqiGRxYm90IWYsDT5
em5yPr5c7Uv/TNVuccw/hf37jXkGrqSgrfFqexoArGbhkLa8l6Dh4NZQT0e6csCY
VN4YcqiNMYfNvofMTPPYq8aKghs2PbZ9/iff1437tn7o4vBaBhHtbdkIV1nla06a
elv/saL2SbEv6O3TgHhCQ4+nKawbyyjWkB3paPEaRv7jZERMVJLA9EBpByYPz+NG
GW9hxe60h/itQzCWQ1kJjthid7/4Xu16NTHLsCAxWbv/NRsIf7pY6bUtVnV9NbUY
leCmIC6oNc9CdUUj0cDmrpITyAa+hiGM6mF83ygfdwTCRr9HCCWHKz9XErULbZb3
Qmo8G8EjWhIbMqwfknJgOuvTy1qMURk+xMa7WrhuvbE9KUQRBY5ttaMB8t2GQ1r2
H+i6kn9sASt93t5UpmqKeYa51FdKZLMkhvMPcbQFiDFex5VkHyzkeNpD3GRZERVA
kxEFTsoII2/VFg117MBNhDL2k1xHkl9RU1R9S8i102efcMbDHP0dgXJqEe+KCSyZ
slXf3uMd9oRr7sFJ3EuvmGSuoaevA1R9JNn3UNVfa4VQ8tzfWznsuPmlZMejTYF4
CbRwQk4kKevKS2pBMygWnQLN18y2nm0MBUtwTsQLykP7Q23BDJRTf0GF5CXaz3Gz
0MdaeTAli3oiW8Jx+4xRHyNlWrsQNk8hJ22TOPLptVsqJrXoe4rLgRrC49YyvSMo
mBteDcTa9yDNwR03Cnbom2ldM+BFWrW8ykwbjKMZqweHoxgM4SClLP1F+PL5zNd/
vB7xUCFMOj5DJSi8xhRwmdP3GdeAKv5eVd7JS9UC+UpsTNcnSLEK29NU1fbArOIB
DdBSMYuM5nLIiHebvr0QyrqlZHvsMQ3S0Wim6iloIKS4GSN4gXClCQ5TTkC0zLJo
1b7sXEZfcXS5yqQ5PX1wbwYCn7naZwwL2DbfoBPT0VYUPrM8zYjBNHIjjstc9RvT
VetrKBTc1wEMFr08cGhpJR6sFwUJ94pa3yZoJW9lDvfrBk30tOjt6h7wRy+mr7w+
2WgM8TRF6i6nWxVqqjjbSQJkNb4fR2tCrYyDaVhOQ2h4mvsCP8b7EdTvZxq2jSwy
k1R8z1QecqKvd63uyULi9d1q6o5NTMTKAE2dITBBlNSLC1J91GXVGmYSfG5zt0X1
QfWI5KaEDbc7SClnW3W21WkVnR+iuy79pjV2HDBjdrWFvSC83U5Nw0BtQ/jBDrzm
ovSpD1n9vnbeS2aZP2QNv2lBSWJx86rbgl8jDLpDTsg+nRvs/nnnN3GcMG62kYGO
KNG6nFK2xTIe0yEQumGEOAXwCq5dazDqM4yfu+Ym9SttSkbI76fxmnEPtnPOmgZt
BJrd2BYlHMnpg+sP4SftjIGwc5Iy+fYXCNzEDJOtfkrdKtzjYuET22+dobmoHMmf
E0ID1TSotrVgDGCDyQGjgRVv+l++GDWji5ioax8jsTIB0YG8vjCkfUUSFjBUAWqI
epsB9xvWVYS8pePAeN5igVPMXO6zsKuIQaozsjYbXr5I9LxHugCRlPxUowfFryZA
taJkNidbwjaFg+tnerX9kK1b3mmqIeRZcB+/ZYa4l7BAXhLGgRHfSCKHc4dT67Q/
UBS1ie1hC0cI05Y5Waa2LwHY4aPm1w9iaPvyHwyeEHjcVk4UlRofDDtHSPt94vfE
iC+m18BvDe0FauOAd1BUf9fecIkQYNp2OUedqFezDR89T7+SpA67T/4j9K36wJ1v
AJWRGcto23FJK3Joe6gg0WmLrhuix/iMmh2+WQSfwa3kpoEn0htoBWvOT1h/gTp8
TpBgpbN1yVJ17Zfn1lCvHurnjoAo5MI8usWHd9gQDlFuEOaByMLLQCu0iimnQe6b
aU5v+TPR0O+44bnouLJb2UY2YAE6LQr4b1LMwdUBfTB5UuoAltPE6dgEbYph9cTb
IQkCEXKRklwcqcW+Kgpf3YfT5Ay0kA0edRVYlwAIDQbGIXdIzi1RDdrVoZQJ+AZk
Uv1wgrXTmUoluZgBUhkHCI3p9XC9Aq/cSwdkrHil74lqyn28mycgGQgN4DlB4YVd
kla5i/0Hdg+W/9FFUHeGiKCvHwiI+Hwlb0sFSx26q3PMIbtOzznycwPPnpeVk3DW
AlmkifY52U5nLpJiato3mO3MRMaShjVmGmBkHdcCsnCDHIhn9vvP3Um4mcu+oTPX
4HvZZbJSk/GacRLaz3yfONgcI3lB6Ja4HJSTpO8xZ/9ikNXtbMOYMepmTSPi/9bi
4VVkifD+d1+wuZJPUnkjQFHFbLgJHcPLEDh5wMR8eqkQuEUpmiE34xr9neZTNtXC
aqddNL5zyZoY/7lZoWTs3qrITQZU2LAqEmqcbm/R+HouYCmUVaOLfY+jCiDU5LHy
eUFN75L1hXaFaVkq6vqGK1AGODwNHOqwONye7i54xIx663WZsOBXEI2onLVBIuBE
`protect END_PROTECTED
