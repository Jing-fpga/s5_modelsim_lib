`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BS0nA6fGeNpeXibvygxUv89PwC5YXCIucHCV1i43tTGazLPR53f07ikxLySINrUN
zi/pfy2q2E+iacpw6QJI+iX8JBttkZ+G/M83E8gGts91+xCDvI+9iVkCjUoAywZj
HUKYb62ZczfPW8LPBbh6npwNv/k5Py9MHtMQOKWvuGtWa05BjmJS8wp3jqTbonYy
+zsn6PsxLOuRUdTIbuEgC9jLvNhG8Zwdg3eBJahkDnHwMd9Fz7MCvkiI/CxnJZs2
eFxf+XqbBNf3zkMk8oDAXLlLzLiQhrHPp7xDbBIDoPPq4tWI06fu2CwkDYu7uSo+
IW/TMd++qPRyeixGKpoWTyENsS7QYOfdpPe270FdAmnfkFsIJ/d70xXqb8a3WliI
e4R/5/AbFsbv7Hes7stIOkbxrLvDbR3z35QJX7Dds9cpiTaUn/Ew8vmog451KToX
fjEo1vOMK9y0cZwkDEgBJBYUfojvrgIQheUtpD7Pv3B1Vv5Sj3K8et2hoI/H4b+u
2LnLRi8y5rSjlznuboyhq9NgHVUi+CTJshIH9tFmjlZkaA8EuwpqbqTJ3R/ynqBy
5fR84DidE12cnJL4RfKDCTKpBQsLb2fVBkO7TLd8agGt/dBPOUuq//F/HVr10jh3
EnsHma6Vv5j6ol9a0Ry0OfFFcoMOGFs7qDj0AVZhNr3/Fyv/6L5A6vm+x9v7kyL9
PFbIFZAdUJ9VpLZZKCgxV4H4vjI9wWfJL2Mxc0URFC5dGuVLlX/3P98LbtGvPEn5
FJGqNI+l4kXXApAFE5tv+WFp0BrN+K69Tp9CU44nwseZvC5F/FN431kAFHzGbCgl
TZm3zkwiZUSAq8eOX5hgd4JkmCbeabl7lQ0VKjaBu8mV7LDQAB15B9phumJMfeXk
Q8Jy+lajJp5GbIifxOH7TeGdkZiQ0QQqRvUG3VvhLcwl+gFtW+w3+akHFss/GsAf
/6OYKC5RFLufYuITceXVIV6gXjtFynlR3eX+HjdKMkB1CJWG0g4Eo9Vw1ZA9BZ0/
ItJWuvEKXweKbDPmgPZiJvqDAiho8atpBM/oPPDGlh2jzeYJU2ZNeG+p/8/sEv1K
CrJ7i0zawksOmlKWw6rRLGXFLzLEViCMZ9bizhPYbuCx+4acaXUFZhUsL3vFH95o
BGMydL6kYa6hHc4HBMKB543jrw+N4lD/oXbjK3jesTfAv7WASzD4RZRn2LYO1FLO
LMAcqSjqVHSDiXZwADJ7bRe8YfrEiWPNFT6BcRAbItp+6oLfGzKzhHABTMrn8bd8
eAOEgfvJNO8ybOkRAp8v2biagKCH7Afg8NJZA/vimtwUkvAmmp9coscqrgyNBp6N
EjRBXaTY1M2YNgMjMH9rz7NhHd59N0RANkLDCogL7Ov6Jd8rvHBV9cg4C547F1Nt
0m0LVpO5ZvAdz/NTfZMDt8XvAPWF78nggI2/uDS+aIUWwxQjkBqOEslLkExTjavJ
484YEg9f5DkMG+YoTe7trblVpjGBgpjipzRhf2HvbM/ysdfGFicLZf8SwzCDcSe1
c9Iz0YxM5XtcYer4sZ+CGSflnSDaT8tkmON8ol0Ci54EH8WK2fJMUw1/U/cTgP5r
x4G5nkUs2EGAjXdEEvb+bcW6nQ+aVIEyH0fGfPKZxLLoQOtA8+fLjJrmUW5Xi2La
M7uVoQVxMf8HshXl83dht7z+Lara664okj2BMblpqlsJvXeDdvPPO9/IjBJ5iMzY
XgRbSliI9KfrT7BISBXBIgAMM3Xb/iF4bESmayrhPksopdipBjgw4NZC+Bw+AK5g
2VSWFuUtZK+AC2Sq9hBwCsJ7dx1vdmKZp1PQFOos90goexpJj2uNmNtHUSuSF0Yx
238wUjqqMqjDOl/sl+veggpfpojXVnsO6Z4X6nl8+0WmPwRBp0Z28yH0KtytI0Pq
K2MIgpLCYAx5kAWuxZf69zzMZS7tMNefmnwpXxbxPJzoTkmWmIXR/M6hC0lP5OBs
TDJWkZvesdyXzCh6LjsKCv5EH1Yvvd5ST8OPzgOHQ8iW0EbM3Nedryt8HGEOjtN2
DqhlRicFV/INz5VLcToJ0ws72bUVgP1dxvAbHFHPEbQt1TyKJTR3gLUoiWyRstKZ
NPLDrtUv/Of32HKkXGcv1Nb8bXWu8CiOyYH9RJDr+3tmS7fITGhJsHGPgIDlDoay
+SsQBHYE4lgF6foUh9zZT7vWVQqFMafLB2CRdfmTBc10qkXR5mnypdYF1ZRlOCr7
RS1XYKhQgwkyThFJfwLNYVPT6PmAkvnkYpvb44VsvpkrWVGeQcb6aack+bPpudJA
NNlSqnYeqEmI+5ggrZo2fA==
`protect END_PROTECTED
