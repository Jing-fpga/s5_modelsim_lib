`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z2auXKp1RdLvwZVP1vikIE3ZnN9EDj5B+KxZQ0usI5PrP1AGBrR7DyCdEdKhjFTo
k+7OKCyI6KVAnWJJ4QUledEkZB9fLMYEsS1CLOjKK5WgiI1jj4rr1Dq8jmou3XOH
BgO48eMCmeUbzGdu/56eKsvK+Cyf31YMe2J263MupWPfPEbfUldLPN30lNTEXHyY
hjKj+nJbxJqxzWmAPpy0m7N1lifRmTYlq48f+TnbSeZ9+e03b9ABOb5c+ChRYBNB
1AA1uks9gzrczo5qx2EQlH+xoCrL1VxqWVM8rS1mblSfzJ6fvw+0d3xi0SEz7Cxj
N/qMUEEYPLam2qYEEOLILWfDVIT+GCmGNhNdixATt8z7U8mjB88lPz50uB/TM63s
MeSlhAz8KKR1x6V0b7ofEniKzufwONmTFwNNjWcD3MXtFqJvk+UpDp7u1t4Bp+J1
Ya/M2vbQBA6qId7rEAmbv7qBLhfNRst/8PICKOKWvqQQFr42OIt49lgVc/OqM5GO
40j0jBwL/+MwxKYsjGIM3zIrBMbQcX9OcWheQFEVrzX7MLIZAz8fiacHepneBJb9
pIwIXbGRlWpNZsG01aBFg1MQgFMJFRdjK6dE+h6IWWJVhhV5tLbpnKXFyS6eBgEu
0phtGOrbjQADJP/PiKorfvJRkReXudL4dVj6tyqMXx2KHEiJH31T5AnRtpp1Znu4
qF5A7R0tBiInKwrA3Alqo0OOwMBNpRcRPjRy6+uhZN0MrpeWTzY04+nrbtCsWwOg
9aiHRegtqxc8Y9LfOKjOBeMHEJXUoWOqZpUrNwf38yjucVXoPkpfBdgdX9p5ZxHz
g4A+4DBvULbYRK7ZS7jM51J8PotOAEbYqAbx+fe91QKi+BQAgmr4jpyMYN9Yg/e9
O2znyqKmOFeV9/Q8YghxIyhwYDlYnqah/r0Xd0M8Zc8ubYjV9Tqv2SbE9Cul+6KX
Ib5sCjYgsC9RYpXjfNeUwUo1ULNktc+FuNIKBjhUvt/U/l1mIerT21hbJBkpoDFr
Zz0W+DcotMS13ugSoEQPCnlmI4JixDRs3ifHAn3oGtiJxLqwurXGuH3cIhMEdSQr
S1a1/cJR3eWj3IkyQS0MByKakWfx++VU5lFcRTDJRhVVI87jFKbRjUPcvTZzrHMG
3xABABL1t3GKF2vTgQy14CkV2j7dJXbzr3xiAEjkGf1Cnu4d/I2TpBhtH2ySPIu7
kusLB5g9pK2Y3E7zAiNAqDAGiJWVLgCARANtNaZCLRGAc5aWAaVziDHEdRVk/M3Y
vlBms1+AK1ZENj8bU7DBDyjqu5MyrlCnPKM4zuqaii9FTSG9oagfnbs/B30Y8XuS
hSD1/PhDwqdE2w46Q+xo8SKo8insksDmQvPMMP29/1Or3kRhYzJtUStMjelZI+wG
YuOLRQWMMxYRAZqyf1bCjyA/0pRPq7QdhIzodM6l7oAUCYuxxrB3MLB4DlKEg7u0
3G8I/8Wnv7b/d7ZwR4RnfDLRFBbnA4UyZI0ZO3jH3ixkxN08OZOAahJaXtdrRwgF
95PPMaAHQ4Qk5hvlvSXhiDjuxc8j8l7pYhncKpPTopKeaNtDwf3pBP1Gu587JxEx
uBzReDlBX9/TckFeqRXQ+5Wqj0Z3rW5gObgoyqER3E7ZrOz5CTPnzUrPQoqi9WEh
e6qOyeEebZF2OXykGrrCugboxPKXUmMfMo4Kg4mf9unrQbAwP63R9gWFiboVa+e+
Eu5YNgXnqwrnDCJ3O4FbK+5K/dVMClpk8w+jV/2dg9d6t8egUZbfFP5MsrD5exwi
8+VhD73OzuXtvYSniHDhobRIrlzCMxbvyoOoUm//b5aQ2bzxbcKM5kljXbL0c/Uf
d/HS8eEpNBFEJI6YUttvoQkUK/3ZLoB1RJCeITwO/zCc48MaHgPSxe37zWbM6io5
4olUnWX5OqgITM+2WRhrlsgN1hqXEMSwjKA6iroswLMgRz5ZHwAMQC7KS256QpfD
SvM0Lha+tz9P8aZeNH2qBFuqibNXJrEfjnqSEk/VI2eMcG0KKvLKpcDafNAhS0G3
c1KJASTQVcPW/1FwYBEKPRKg0coW2p6Yvih110nGangev6U3VgZ7tiGRV0ANxdKR
+j86ECuw3qeSb7WAUm0WSpgooY2j0v8W1lujM7FhbQ0p5iBOdJ+lk2r26or05PyV
jpZSw5iIcx4WsgkePt6raRKLEV0yUb9fBE+eCU8NXCKti9/I6m8AfeaKQUN8I6km
dTcAs1R1Bj0aQcEoIC9SOx4g6EQUHaug72T4v2rNseGc/5RCCxCJHIXfcKvKwujI
SxFpOHBnDT12fZaBQdnvkMZ0gk2NoZNH5aNgPcOjntyP8ziAROgz7yOLMOSfo/eM
jrt2+8WSc9FbnuKHIaUluVvRbYi3EacGsuXmTUbDyCd95ylrMYQwh43HNHZhG4GH
kgbejcvyyI3r+Vk/BTmt51cv5jnTTyqRXD2NmfiJ/IRZonAmExMDbzzx4lFSYSJR
2oq9tYRh0DIihdFEpEyINjYAMZMsh2DlN1cgvqNP+5ELDx0L3mxs/yiAbwe6WO7M
GhEP46N0+z3EvfFswRHiHjI91Sly2mlQyJpcaTD6Tp7QTvR+a8bW0IsbkQ9J2wyt
X0akXRtMUWT3O86oSGgfpxo0q+qckXY85vnSwAc0uXo0m+OexSrF4xWsp+LMd50M
BErDFLa66bNK3Yed6ZXAKhY4L4z7bVU6N9VPHPAGUSgan52pmDCafmA3nwubZkew
/Snh6ERzAveSvOCFlwvoZEwpVaVUSspA+zoM/plIV/XWO++mMsQq1+udak6JqhGS
pYu/GdjDUdLt+DTjgYZoJWYgaep5VUjUue2WUZl0OScnn8HmBKQChTLKhdz3bXj3
Zc3YZ9S3rq+WaUPYDC1/lQ9QCp4x4XnoYyv9UnJXFi0pOcko4zVp9vTRX6JxHYPR
3DVpotMBA6OLOVLFZ8ynExVg5KyIHVoSUZG+Qy24WBKHqoA1HCst10cKsKt/O4VW
I+/D0qg7yjnm1CbhbkxFp/kRjHfJbMWDjYo4So6QVi03I72nxNR7mKxzSepMbRp+
wk9Nl+HUA27Rmu1SZja2a/xhHXe51iS1v1FwYTnt3tc1cIF9BJWBjERG6u5/hrLG
3bB2e+3W5CX8IbAFQkyJ3xI6atHiZ9CzLuFFYR3lpBvoek0MuvnXyCtvFZx0OA9j
YqiW1JaeS4onTsZUq5zSHuVVJ494eWIPODfpl2IEAPoNhWs0NtRgOU3OC/zroLIU
6cCuqkYx3062jnA7FD6AoGq2KPtxhRhIAEVmZ4+qQyq6e8xqMFEPkpv1bUxH4vPt
j1HCNNrgB6DI476WZUWisjsww3e9plAebta7kbuzKRLjUp1OFSfQO3IPLHU/6e45
gJwRf1StCVvOVdwfBk1LLQ187/hW38qfTXI19CjgH0kHJApSQza9V0A0MSAV52Od
b0+KShStlamw7tv6FxoJOKxH8eT8hpo3OW5ZEEwd9iVoEIxBVvOMiabo/aFNFFAR
bBlemXg4Gr/HSNLshNpTcKMg6SWjkeZodOUq9YjvgoNPf82f/on49bYjm6WdZQnM
Qfac4p3Y901fOMHQnCX4GsBfCMqb/fp9ykJmR6j49wXJPVBbnuZJfMJWDQ21cItd
1GRt+nu/s5eh1KcxYBiQb11jZturUgOZtRu0ywfS6oL7kYM7EtjwACkHqaSNinis
n7cNJd54eODDfV9xMOrk2Q1SlM1ubXstF951eAPVLv3KmZMbUDKrwBFlGuduDe/w
3OHyiITYslOsivS4V/j7Qe76tsr0I0yPUS+EnxjKZ8jfIHQoXRMzYlE5yn5INKHE
5WfCGXxSYRDtFqfx1/bktbaU1uT8J3HCXLBI4MGnPFHE6M/TU9+9c6rdn4rl9Ie0
iWScqH+T8fhVkFr29n+nZzTUl2WyiLJ73tGyIy2PBk/8gCfjuMY7N7PYpdzwqpO3
dvTTbCAbyf2YMc7ZvoTh0/afpRInZkn6uy3zARuQRGxm1U1njFZ0jLaF5GwURCDF
EcpGmLD5Ob+jJwMS3j5ThtVAHW/71ihKO5O7V8hndOISW9+XPr4KhbMBMpVtuj0H
wsm8/+sdQC1a6ME0YHL63REYCHkiGarxOUiINRQmCvUN5h9u83QxvBX+4DnRnIa4
wzx3HDRwHeP003VITBAqs7qnlULDi7HQ0xpizVPzlidlelSurTSoKWNni899h3vD
VDQrQx7z3hdRBavZeuULCqRAHxvsQieHrPd5WW5t/WUvLWyHpp1m1OW+6MHomYKF
Tz22+xA39dLMP/Jlsc/bXBeC/gXoC6vu/2h3/yYtvRMGen2Rn6mBlhMTBie0diTQ
UiC0g2cP91yxx+F6uNTVnOKNbKlpDdpPUQmT2jlIPe9D/IvZU8wieLQ4BRTP03g2
LhRJO3BHXDEPe8PIB1mDZFfFVLkgPErSGGRLTJpZjlhcQi2rlhx3t1xX1WEDkb8D
oPxmjOhQ+cVXoGr9UPiDlE60JY9JQiQKynGDFDf9+a+mlJQwhjy7juNnkWLzOA1p
hhGhxvMfShob+8iGeh66STMlUwSaOmqDggnjiOgxVq/9Is8fHAytrb3cwPk1eBN3
TQVrqGOXAV8ctL1itVRRJ0FOczCNptAhnWcnxRK/enSLH1orhhEApVyREz0Hq1Sl
tOgo03vjSuyVeuMEUjdGxP5in2LhuwUANTgwJoWWNEVU/rL93MfVJMgiqvmvPwmm
NTPFx57CKLbOHpNpzlHi32r7HuN7LRcK4g8B6aoTiPCCYy3CWo3jhCgE6Hzpx83Y
`protect END_PROTECTED
