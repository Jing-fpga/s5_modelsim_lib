library verilog;
use verilog.vl_types.all;
entity stratixv_lvds_rx is
    generic(
        data_align_rollover: integer := 2;
        enable_dpa      : string  := "false";
        lose_lock_on_one_change: string  := "false";
        reset_fifo_at_first_lock: string  := "true";
        align_to_rising_edge_only: string  := "true";
        use_serial_feedback_input: string  := "off";
        dpa_debug       : string  := "false";
        x_on_bitslip    : string  := "true";
        enable_soft_cdr : string  := "false";
        dpa_clock_output_phase_shift: integer := 0;
        enable_dpa_initial_phase_selection: string  := "false";
        dpa_initial_phase_value: integer := 0;
        enable_dpa_align_to_rising_edge_only: string  := "false";
        net_ppm_variation: integer := 0;
        is_negative_ppm_drift: string  := "false";
        rx_input_path_delay_engineering_bits: integer := 2;
        enable_clock_pin_mode: string  := "false";
        lpm_type        : string  := "stratixv_lvds_rx";
        data_width      : integer := 10;
        dpa_config      : integer := 0
    );
    port(
        clock0          : in     vl_logic;
        datain          : in     vl_logic;
        enable0         : in     vl_logic;
        dpareset        : in     vl_logic;
        dpahold         : in     vl_logic;
        dpaswitch       : in     vl_logic;
        fiforeset       : in     vl_logic;
        bitslip         : in     vl_logic;
        bitslipreset    : in     vl_logic;
        serialfbk       : in     vl_logic;
        devclrn         : in     vl_logic;
        devpor          : in     vl_logic;
        dpaclkin        : in     vl_logic_vector(7 downto 0);
        dataout         : out    vl_logic_vector;
        dpalock         : out    vl_logic;
        bitslipmax      : out    vl_logic;
        serialdataout   : out    vl_logic;
        postdpaserialdataout: out    vl_logic;
        divfwdclk       : out    vl_logic;
        dpaclkout       : out    vl_logic;
        observableout   : out    vl_logic_vector(3 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of data_align_rollover : constant is 1;
    attribute mti_svvh_generic_type of enable_dpa : constant is 1;
    attribute mti_svvh_generic_type of lose_lock_on_one_change : constant is 1;
    attribute mti_svvh_generic_type of reset_fifo_at_first_lock : constant is 1;
    attribute mti_svvh_generic_type of align_to_rising_edge_only : constant is 1;
    attribute mti_svvh_generic_type of use_serial_feedback_input : constant is 1;
    attribute mti_svvh_generic_type of dpa_debug : constant is 1;
    attribute mti_svvh_generic_type of x_on_bitslip : constant is 1;
    attribute mti_svvh_generic_type of enable_soft_cdr : constant is 1;
    attribute mti_svvh_generic_type of dpa_clock_output_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of enable_dpa_initial_phase_selection : constant is 1;
    attribute mti_svvh_generic_type of dpa_initial_phase_value : constant is 1;
    attribute mti_svvh_generic_type of enable_dpa_align_to_rising_edge_only : constant is 1;
    attribute mti_svvh_generic_type of net_ppm_variation : constant is 1;
    attribute mti_svvh_generic_type of is_negative_ppm_drift : constant is 1;
    attribute mti_svvh_generic_type of rx_input_path_delay_engineering_bits : constant is 1;
    attribute mti_svvh_generic_type of enable_clock_pin_mode : constant is 1;
    attribute mti_svvh_generic_type of lpm_type : constant is 1;
    attribute mti_svvh_generic_type of data_width : constant is 1;
    attribute mti_svvh_generic_type of dpa_config : constant is 1;
end stratixv_lvds_rx;
