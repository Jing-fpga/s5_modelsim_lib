`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lz+ET0QyngleHcKtR1VrbL0QWev6iSx++/S0NA1r9dTnv0VDj82g8mAGj5y4Of3/
MZz9rtKqi+ZO/jpi2Uc02Eu+hTmO2pm6aUXuphBEQbOOFc9hiEOBtEMddEFJaHfF
qTiYC6uQBlG0syON2hYZK9dclt9q4QoSzXMHuo9hElK7/nV/OcMN8MBrq4gxuMDW
NcQbTDwPHPVLeQa29EDlkUZzIya2wfl+Ugzn0KZ9AJ3dNR5eObVQ5uHqDKd+2icb
EmygmV364+f0ig4QbcXyDwWsV4Qubf0zk9ywHUBgoJtWm+O278ETKtoh15dPuZaV
6XIeTKUaqvo732WlcStacW1b3L2oRaBP+nc+WhZdPESfBz/JcoIj84CQGOvHBILv
hAYk7qeIo8Rl1kLKafmpRNz2n/yhWfUWF6cshBWlD1M218NkWBvI2bK2Vn0NG2fx
E9L9TGyiSg6En5VIjnHc0R4xkg5LWEAeCvZKLWKArAsEsNncsLxtvbvKGvpL0Exc
E6sWdljMWNQlJHjNsy+6XFD/UG5AJsbt6inyNlTjurBhsEw8jo0VRR+HS/woKNeV
WljhkHo4xGJKJVnZTR4VqvtsXl4lYVxdECwvrSPMxyJhLwuEbfYCA640NogGYr87
y9A82e4bDx8JQSO1T6GLgoShd+ZYxNDHB5szIolxrSigVBPiq4JwtrF5E/JujHPL
ZDGBTkPI/KwfZzQO8L3pYChynYzWKCypov7WihXKNpPKrF2hI9tlUVbWUck3bQJ7
coIyiC3yU/LGDwHe07+ttHyeGPYpeIP7us8udEVJUbqSAPqraakMNn+u3cBAEVnH
nNsh9HJsOe95hm/9VFmMMA==
`protect END_PROTECTED
