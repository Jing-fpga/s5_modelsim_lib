`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w1/31buQNZY8jZisF4u6yKbDZ7m/tTd3/Vtu5EDPyUjdrLL+yXAvM0wbqxJ98vDi
SWjPexdce4lWd/t7PCey9uT23nqdKNGV2e8a8mS9pOoGBRFAv4cH3+9e6VFMORLC
IJo+es49TBr7W8P2tgGfrUPtH6AlpJaESkWcb01IGcGFztVj+mahs8WPri8M6L7X
UhnWE2a7ve6mp4oYbfzPWUESV9qtJV3S2+6DRkOZbQ2jxl+Y1Qz1ZMVbJqmrMR8E
6sYo9M4WBh1gmyV6aOLiIADcY6TD0/Jf5sfq2P7L3QjdjEgREv92wO8ta1V6j8d1
qpndk2Y4qupRCecyd01ZCPuW9KlnV6XFy9xyZWruljTMPjG19KzBJP+DydAS0ehX
1OLkKP/PdydWKAwaCXvQYxPL6Ljn+0bHFd0+0eP7V+nEFWmTW78Zq1BzHRy7chL6
BX+5csGP/FcG0Si1cPr+zqAzi4geDLp5nOHbgL05xkEEIIs8HyeGJbGzRgNVvC1T
Yxpqyv7rOG6HHvltl3ACxRGTeZV2yWEf1U3WEvtJqNFIFOYWK8FuMCo03zRQ0axT
6tpxlLNnUPeeUxoAB1jJZzhmVMde8IPyCVr98s8uMYD0NDLrNmDdD6TRHgc0AEYM
+TlcEsS3BaRxOhJvQsra1MhJh2b8EmPhYZvhIPaGQIu5vGZeQ+CGD7D2wOm8QnS+
N3+kq2Y8Bb6jSymLBaaBJa6deJzNp/w85CRi1ahkVfwCUKcLZy506NMcm+IyKPJj
sKARvVQfb19JD82x17bzTtytlKTp2O+NdfQmzKOsf6D7BKmaD9r/NUozW1qBwJr+
+r4DT/sKFWkmtxOWkTFBMp5Jiz4XDGJOHsNdTAyar3s=
`protect END_PROTECTED
