`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xJNQ0asis8CzjppxIhsFlCz2Vhg8PyjtqNfvOAZNunFuQeWZ2a571XscQlmKq06y
ZqzMa7//2co9dOiIffJ6dMDbAF79SI9H8Aih8qqi5GYXpHqUDEIGgTZ3gVmvNegR
I43Dvu1mDoaA6Zbsns0DF0XQXB+Wy1GGmDiZlA3VjNKfgU1K9+s5v1XG8PdwaQGJ
k5nZedJMSacg8aegkqssGdAHDSBQW/3g7rot75EEurVHsBKedGbFCZBcA2LnqKz8
kOn71ybZ/R53BZz/GUGA2p2Gf+IkvbQlFkopa2iePSiaNeobq72HGejCuQNEtl7K
XyqdyoOjD3YGrpxmDVUWzpODbcQj0FqA09cig3Pfy55o0GWv8QKhI6sMif4ZE5Qs
ANszCiwfYzQfrOwqN1bmdPwwWyZU5tZeWbHKm6qOnDOaLaMYGQWsHEAagjScBoni
p7cOwubyDSBEEEPTtSLiO0+LcU14qWKuZ8kRf3/i4zrgAFGAjhFXGptg7yqR/pZE
qzKAJQoutTXlwJGVxJOV3JXfMa9n/zGm8T0OK7assPdXMT9Rn7j7Pt0SOsQp9Nl3
rBcYz8Xi1AocXXtqo0mJvN8mrzCf5nNAw4fQgAQgXctxxYoRYYCZ8mPp+CgqKn/T
HP73mz9rnCgpA5MTORjYr6HFXQLIQ25nEUA40W62rOFjoJfGUHH9qNLQXSZ9Kr0G
4Du1eAM2SdxM+9PAppzPPg5O0NzRxtFeaOcFU2/R7Z/w8g6uh3slT1mKZDenYQpe
NqVcA9dVVgFwr5TZJI+orJ0w1P44sksI2Zt+GvLI0NRjUcH6VmuOSpBs8EmL4ZyJ
3LaZp81rJKmMkMLsVbxxhKnLiO5DiP8fcpaDWm+p9brppJWaZ0rvts1JL/9OwLwg
mVnsRUQ6FfH8OQUojAI3c7Uts/jF55z9YxHw7wRl5zSZs+vOZOZs+TtxwMyZ3QRm
TDQej3kTQfh4qEF9DJZ85h1TM4XHctC+/Q8nPrJu8aSA9sdKEIsVDvhVF+JydSXL
L51t6Wv2yoPHRXU7HYwUePT+fIqf86fEqlrFzrAxe3PevsN3ogH3msn6vh6UPLA1
tUzm3XFVeLZxp3ycTnYdA6/+ceWjF5TkjYfBxXlMcn85c94edrlih8q7Lf9sbRzz
MEFQDYgkR8lMg192Qf2irNwmMynaJXU3tmXKPU9Kmj5CYkrfyXIzsnMg4aeUCBPc
jdz3vpRW4DkITf2jPBjnsqA15q9IYwGPFuF4LstKtk3XGPk7rZELBVUC1FnGpBaD
h/2YWBj+yus2FRRa9PDgn7nyA7g7+GqtcC0yAHQybJyDCvWXZqAmzow87XWpJkxP
FWCF6qOCr7uGTJ5lDTt2nA51UAyasSoZT7go9+LMRJSzlo4Anv5I1/527r/fXnXe
qbFdz3FPcw66OAPNw1/wTUdkPWejn63D+96soA7llMLW7azyDHtAsuL+bRAsDyEp
PkxOXzrRIMhVguVsZ6KJSu8lSPF8G6tWkgfJIavLg5pb3VL8ZGzWgp5idkZbRDtK
Dun/3ScPTxPNZXArXd26ZVS19ERbdbzFSjjg2DO5lwgtN3sXujt8XYdwfsFVssqE
cA8EoHXM1uUlE05/Bj+SEpOnwG60ywzJFk8DLle0Ndg=
`protect END_PROTECTED
