`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a525srOQkIEs9Vg+lk2gQHu17je/csNBx0h28UEXr/eyvFQRlpVQ6Gze72cKN/Jz
9cYGrzSeCKztAfb2yVSzRbhP4ue+luDuFNlCqVQtbYsgWIRe1GNqAxIDtbsBMPUE
C2ZxMge8CTtiv1SkJKt3oeQfsbsRxAoDbFJzcux7BN6J6sUQu+SfEoAhhZcKvR6t
LQdAVqx1LEjNxQsSFtdnZlg0o4qdO8f585Q3lhi5k7hTbviZp6mx2EhFIgLlSTLG
XeoXtRHlueeJFrUwJ0J34a84qCSk+C5jURTbDpLntk5jW3F4XrSPvcjc1+nkMckH
eLcGh0DGL7pxc1Zd60+RMQ==
`protect END_PROTECTED
