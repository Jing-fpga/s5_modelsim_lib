`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sX8cCY0bqd5D0h6z1GtC44xzk5wq46tZ4hZW0eBP0hK/UCRzWdDNxHCiY9uoGXgw
QujYmpuGHUNdMvsMWzB30zgFKEpKs1IFhvq6Y9V1gz9PQrDhN8IZck4295IgM4A9
y6wF97BlKOAN6XeR6YwX0VMB3jVAvgEb2Fud0tqfErjOEI0lnVs65XRZCdklzKsl
TXwsgBZCt7Px1tboK1qGt7zYvi7UU85HotZIRo+Wj/w13bV/BdTwm4trYD9Qv8I4
e1SLXSiAo/waL/l9nZIWJxw5zvyNW3sQnACuSisLB4lhSwrxxRLiW5ynXN5+e6VZ
xNhiijIyKAYpeEDMZggjD7Ef1XJZ+K4w1zXdTKvoCKEZ9jVcS0a2nvCfbk+hb+KD
5H9yQYm4NHVxuJB9JbQM/j9BEZFeq+Mj9nieucKF5tnhLzUuPpHTnjEKJuuD7mzh
jqpaEzl+cENJFur3DXSy0d7M4Wy1UN/AdI0P6XgeFL0j0jAHUwAQXNkRmS4DDwXt
AZJk6opXktmETAe97rXwEycxoywU68EbwZ084dqeqlfd+cDmiS5iR+v3gsBmakN2
F3VAxm10fXJux8ExwBgjFhTBpBXXWSZtt/Bfs5Rk8itAw91weCsE7YGvXDoUzWBW
d26CUNxseYSG5IqhctCejkW456D0Qm9R4MRW9Y+CY7AA0EaT5UHmyQ0gmETJW48b
xsjVAbT5RrY+K5U1ZvQVJlWGGU+eXV7w0hQZMH6KqVyFPCQ/UIdgXXfwLP4HuTvj
eUWN+Ci2jVd6ST581cmvqP4hMIif2fuO7Iu7EvlpEWYbSYaN1+g/kvOZJxj3qx2k
9DGeq7Y8cZw2jwzTJTg453sWzcSqVgJA91Q8IXUjCsEwBtgmbN9AmM2NhitBOkQu
frN5ag1G37TZLTLUEikbXP7rNh8kcxtMBdD3gj5cu1qmTo/uz/lofZSLqd35hQSU
XencqUZWzpSv8Hq9CIbKZsCwrcjHrwolGz8srTAmeDNhqAAJ2Gd4tnDJiz5oIyij
eDuElwwuI3buIOwhPPcEp6B2FMR8S4jIfBlS11IiHyl/gdaHVF/0G2+ztH7H2Jgc
NHKqIpQchw460JYpislZq3XzOgElwNOKHDsEP2frrz3TDzPSs6K+WkelmDXuj5ea
5Cj9wHJWYwrlkUVPNRMDCX5pYwV/eax8t+f4aTBzDddxpLFrwoVwrmZeYLO5baTz
3lNtW5ehpxOJAkwgyWwmdcwO7YJVdB8BbNrQVeWisEnu2veJNUZPmWc3s/F+6xGN
KMNjAeaZ98guHZoCSGar2iXLOQXDi2MGQWpYh3N/TXwjBiLBd1nVWBEHiVgz6Dvt
L7PnUIX0BIMGRijyHH0B9LAVoLjjN4kRdcBcjag6jwB47Kb/teZIEZpFN1trgLlQ
LOVzsVrn/SD/yOvG+E/s2X5MPmk5imNIk3uXeFoAZ3AMee6tCJiLl9c7rlmPP0PO
dDRkSnL5LJPA5qzxKxWG7BahKWrRLv4rouIN7gnEKq59xLhm0jE6G71RoHfRaxtq
/XrIpb18Rv5VFv5XY5YTxkgfQFgGlj+0eaJvqavow3sUKYIjVAvwumlEQ/soPEsD
LPgUQdp2VKs1jFb+VAT3La6e9Tu70JkCjrxqicfQin18oOE2oAAY95h6anFCOcPq
KK+pA9LRAXqY4dZfs0gtkwJlaCDZ20DvM8i83M+AovN6C87LfOHqYyr9+DOBoJB5
xc1+xia5JrQkYr6Fxt5VobYoQDrC1976P17qFHcHBPeP1SOVApNa6h/W2swPmuFF
QxDqcysVVN9YeQxITEdM/60TSSv6pKVXh4Edj5lMwU7hgUaf4AuAyEvU+XP0YGni
I2Kt6NI9mjEWDEgv7/9QDlP4YPlWJJsk+nyp0t9rGY7QDk5Wegm+4xc+sFTDY4qb
b7mBS/geIDtQtQE9bN+nBd1uYqJbsnnYFD4fpVsLDQmoi36//excXi5A1S7FbDkU
+4mBJssy7RM4nOdzqJWahkdeZGpmPNqoExjKVYXR9/f2n+BxoW5JB34Qb5BQbMaq
vBVTT6MYGdD4U6sfX4Ut57RV0W9hXGA/wn1ztIj3289DtozE3DMDz08FiC3rgD9c
iOhzPQ/wEDUr0OUCfGzN0xO8Yi96CVUBT0pFQvkUdtQxUXfNz7JsljD91DdWwCoy
T/Xmo9Khp5zlx+zkOLoTykSqcGQFEophtRITkKQt1iJ3Wm8ayf8lvM7oLRVc7ZB6
B0yvFOflxAIdhheqAsigREtMtXXVSen3XsZnFKkgxLtKeribZ/+JqTmQsnhWNM0C
6maQe8068GGMreWjIZ4WhqQY1fqTZ/Mc+jbMOg3ZDHhPkrl6vN1uKYIRdqhYGATX
93wNb7ubf6D+8ZDuscR01FCQS8uFTdp0xHrNqaD7PoAxoFrgW7y5/Dv3cXB0uIAs
zgVHr5Q6bYS+tQnaPhitxBsqGA18OrQkNt8M1dNtxhlfCRl6Tn/wCT7O+aHEgsDh
VRKBoUppZdX+gXFb2lXQyG6CxFGEnpLdttDLWLClQWSg2gdqQBh16K2ZSiTjOsGu
y12sOH3H+qAPT7nh195f5k6BiPk0THlvdnYo76iy4Jg37UOL5WNB0+r5Awui53Hn
LJEvmyukgBh3rhPSEvIf/9CnpFIG3GsLIjck/JIt7Uz8RgvXlAcE5JCzSzZyG5l1
muHdn8FXyBpg0dDbDhB198dLilktXONIoF1XPlMz4SJH9Ttjy75p35/U3Th2l020
n86wNtnF6/n/9sAvqmQVIzSLNkdLcIZMFT4Etd9U/kwmH9c6O2TDuX6XoJ4ONPCu
bhFO/VnPxMUKFOibA8JdBSQo0e5vUdIt/nfxOST9aHQ4Ix9cKZ2wqOlrzbQpx96v
J1e592aZv3bAvLbg8xvMwYJsx+s6LZ9DwktRtlMDWjBvEA8Ff/rmFYp3XjhNP34j
ANTY0C8tE1etu57GUx3RyYeGSXfJUa+B1DjT4cVnOjhnkqJnKdRYJTwKX10TQCt/
PiURC6r48KVCl1If0CpCilv8HPnSR/6qXyZkGWXBlRRta8XWd74ePxLeG2k8kbwl
HZPMMEQrS26sXYf0QZUKJCKZQxYBQMcxCE6rogF3nVgO9eW7hG2nH9+httqTlJpV
nhQ6eke5InKqO51UQ//3d8CBPw5XDMmOkyZ7X4X2GgvGeIU/t3FpYr8QAe07BeKS
hJkD5mhPfpImakq5AmYy0zC2vE/X+4KA2lObRG1PRqEYx5myJ8P8YEYMVs4JaeUk
oQF5Ckk0Kxkrh2h+nqA1kuIVvSsOu88oysE1GKyY272LW5xORQjqnNz6vcwq3ftu
cJ1BSMqeNmstlxSYcHGpoZZeWrY1dFk++/bFKaC4FfoH7Riiwba8ExMtO8c6d8GL
i+zgKFUf9IzAjwpBlZmLWtYoTcNbx0kT984nsXx8+O6Hhyq2YkAW4EQSFuVOhhbE
ys97GoAOQTiQx9dV6hp9QI9HSY3og8dKP5zdgVYDnvqhK22R/MK4gFZ4zfUooUzw
DOLLNsjGjll8PK9kiz5358wfGi0/hsQ0jUZwa0n8cT7sEvzlKaBr3TfXW6I7J5xN
xhDqmQrpbRpwixAXBicY0dPQVVUazydCeIQNq8SrSmFlMURGEtb3WDOtmpalbCQ4
zsO4Ip7GECipniRWDd9bnvZUtI6N23qi+3xJZLlUBrTESlJ2bjVsYs7RcW30SluD
`protect END_PROTECTED
