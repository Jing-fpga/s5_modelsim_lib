`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xvH9zUNm6AeMf3kz4Y4Jra9KALtN+uYRk22uOhByorcmdoxip3l6LYTV+zNCkgoE
1rqz2DufdakeHXa25OofMkzcFllaUIZyYs3rPRcqymgKOpWQ4XUAJYbebqdOjga7
xjjbthUnkDuvvgL/bteECr0uisVK3uT4plMG7tbCsQWZI9faGeB5O83KyNjJYzlm
VqBhdSS+UCj5eh9YwB++U8B0Mf43a73b6fuDzDMAkcdTfWbEHMS3FP4nGT5HNrV+
d4PwIDQRGkhDN3mVff/3jgx2omx0fqeoWSGX/afOQXQSwuVcGu+7vvQMKY3X5M8o
boiZU0QmG7KtAPEO5cyxUGsY+Og1kxFLMa8aqN0ZVeM75aEO+pegUWrhw5BhC4YM
N886m0ud64zax5yNgy4kF3NbGIIGlx8qsytBz1FaPndPVM/6zHjPqJ7lZ+KnopPW
uknRowsKpSo/J/9QBPI3Uofy4A3euKV9mjuOpT5lMGDHDcaRb8bYeD5Ni2wc9Lxf
fKy6GmBmADAdi5uOm12dRcpVEhXafmPDxDzfxeIKVK8QA2VAEjxdQiaX3Br30/HP
86mJy/dl+WAcMubNFoqc0ptyo/gNj0T77i25oKfVtQkTWEMT+QG9X/Rmro4KI73y
8fr64dGyToSfcL6lxCTnp72qMS1vWz4D8ctvs0dwYNzYE1l8REFHb2Imz2PBYgYJ
AX7xArLPg8YH6YCjfB6zKXMnCAzaVmGAo527KBzbATk0Al38uICple59iVW+PFuz
pAERwfYPRQPPh6iZRkrP7EyBTQk5oqoCSk0X5vlTQUfq+pjeYvaln+W/X+mstRL0
U1c9kkE9rnZYamTSWr/ufvXDZh10DmuXbx1FUho7TADfTIJNVw4qU3QMw+875hwj
ASfWqn/5eUn0YsbNM6KqoHmH5AfQ1Jr6NVGDAfxukY02dy22E5ssucaeZBXyPZbd
a12TUHjQ3IrLBpRmezVF/VxXPaRmSan1HW1uVs88t8xTtZPdsoEryBHINFiZ6sKd
JvF1OsnNSskUzfEQ6SBgrKePGxFhmVbU3InhAljLj9YZWEDOgg6fRig8HpFMbxUF
QIfZ69KBfj1l6JJlrLV1P0obTQF5QWkAAQmK8FRDM0pDVNvkHgliIkNnUK18Pm6Y
Rzlrf/kT6I8S85fxx2JQCNm0vd4dVYKZzKYTCO32pGXy3U9tqQaC9f1p6M2Pdxi1
fuCezAmpuTHHSGR4es3wSGYLdjiFUuaybjVMJJqHfl58rDJ6bx4Bd9S9XxwMFiIM
ck7+/bMJQvBmSKoQo6MFbZPkACYyoQxQmNYNzVP9igamyK8UbYsO2aGFo7Rf1BFI
85j/DVsTnJR+FQPdabV+RL7O/DXdWkgMcaaC0Ro/A0r/468f/8bVky462OEe2ysp
Kb/T2i8dXvGa7ucDMqxT8VyekaUivyyeH5P3kz9kDSYwI0beBTICmXaUThdRYieb
vmEdOCTo8hZZD6Y4yW4vkw3AAUnE8ynblYslE3lPAny8r7epeA0LDRSoQS7jprCj
YDy4w4zx9PRZa1ELe1G1SrD35MZBhf4IctJeb7meJqBgRHU6D6ThnzPer5F0F8TZ
qbsD66UF3479e9V4qbgJPA8aUSnspND9CjvGRv19dR/EEUnJ+sScPl5uw1aT3M/h
dYEjcQ39DTl0Me+1cwVnzeG7ANOLW9YfI1rL1acaz8cq4IrBbYUYoHmr1WA1//2r
dtaK6vn5VeIirb8S69qeD8vde3Z2tpY7oqmF/Oqw1KVLgY8Kg6Gcxn7z/mYZKQxb
5sW9wpN4SyZjN/KdnmYIaC1rbOiocR/e/vR6/CSsd+oYS7C6Mb+DPp/2Mc2R5TMM
PWZktEAZIXJpvmegOssW12HB2sf6vKn+hPh7m2Lh67B4tJUDZ6SgRo8NvNSir8AM
MSReE2lcHbbb/uX1+JEXG6QBHzLYZuWNFrIKfl1eL4vzOhZ2WKEjHOuIlQ0JuRRi
A/1c1NW8Cq8pMQJ0lrMQc5DaG3YMy66DIedkTnKyZAMqwIqc0rgvTnMbk5I7hlNl
ZuuYCUlD1cWe+rflGI7VoXTP5GHWS7rtWKkVHV5oeqV8xRl8mSZ1V90qnwdyNjjc
D7ivcz8BmeaDlcVwdXHnTeacNAtcDSEzAK1H4KqaIlDi7e0ooONFYeIItwHkwko3
OwLSUHJbIs/VBqbh+hyAicdkz4e4eY4b36ClegcCjZuZvZjHzX8mHqbIZnxJmr0N
OGAPtgusX9au/NG2dBKdO/Hx2NkvenSwshvw4fDsOGwxN1ihYRlE6NTo7j60H5bT
cfZyhDbk2oyZmNNgJ9CWGFkYI6fm7K/2mwQUHWT6qeGx2RRVlu4Ui6tVY8YnkLow
8Fb8A4reoGafZtHA0rRP/5iRFAHEy4ckasbZcpXebuCc0s+AvXXBERae7x7r531V
8ebbNkuVCc/+nqfFmjdk6iE/BhSVJmET2sQaA9rNdPw2TRGYVjVwHBLfwYF/Qetj
r9xASBcX9UNAVcNVvrT9z0ve0LeC03lT55iCJAEhS/GQPux/O87otM5H18Ukfg8v
UvVmU6y7COib/PKnXZhQe7IEE0RFjzTyJNgh/ZC/Ykk09UzhTzCB1zTlpHHaFBtD
TCot2xP6JCwp1+rmO3PB83KCdsNOUekjBkaPdd+eurNmP5ESyy5K7uGVd08/nyfx
iFDREa+zjUVBUZteU7DzDluqy2sckpjCkv4LB2dCssBHy86hDoFXC9G1CWYk1a3T
DM7baqG5Bi9fUMo1KJCfB7IemRzDozcFsUGnvSlQlOOnTQajBGYpXwZGMBdZajIj
vxIVnhkfx0NCS5FKQHd3Bx6yii+wHXm/db/sFnDdMUyV45+ZNycUB0ib9RsrNhxq
g08JjNVfOkUMXPm5MqiOH+6Dga/PMIXT2kCqmYYbBDdQHR6S6XSomI9jDyO9ys7H
WEzhO9TA3UeLoHW7lZjJmibuygVmuT5t1Qg9X3x2aQ9ZBZDRjmD1u2AzcqR8fgAl
Nzx4K3dGqaRrLKXREOxiigxk6q6J5RbaIaYzd8+ZPxoj72HiLPNdqaBsDKDiLdTQ
N0kXWucKUvhJ8udvdqCWxM5FGQSKL3Dret+SCmwWpYbuIemJBdKarcrEh7uKWMiC
7VlRv8xE8Ner3/r2Yzuo3YwnthmBT8wNftScsmd45QDEhd3gGk2gkXaXslVxM2A1
RZpqj8xNpirGUquthMUMruURg1BF1ll0m3EB59U7MaSe0cO83DAlsLAMhhsBiPh8
n2QpHtDTpmk0lxmYapmBTqGnYtKi66ObRmb80Kvym3aXlxpD2Kr0lBQFBRbcENg4
Z7EfbDVOwCKeOnDTem5ohFky69NrLYObt2or7vPGZniF/6bV/LCd6ZQ679NlhUvn
umlTCT65swLOHU5ie+PdknlcZmG7zwo8jJOCz9zGMSxZ+wwHsNuo5ZZpnGrvEiWv
QeyLo/gUWLJ47E4MVfAfs51N5XUcoQ8Z00slXTSR3VftYfg4RcSEmEP6G645AH1P
8h50qoANlmNpVdl5y7Y7MwW1NDsQCVtC41Bdxr4ok03NyRm/sRnSBGljeIURtSwx
B3uFJYRsvo0epqZLJjgSZcgXIhSuxmZcF4qkO5VPcOm63+o6kTTZdd+5oP1tcONl
ADa93ayo7k9Sa6DtQtG94aUfy89fnu3hmjyr/BincpZSY/Wouax0jBirl+2UiXyE
uqs068HAR1XzKeQfFFYXFY8ObtkI0J/6BM80zj7FubfrG3tr8WqyFkPnkWBzWy3g
zjbOWOFfFX52kpToqIfH22+4JJVOBHx1qhJt5fESp/ZE4fb03d6ziLptu8NyesgU
6wTnDicfql0+1NuSX3rFupXWGtfnJ61P3gOYha++xARmsMr/q8Ss+eINsISQTpq2
DNOyeoh6Xy9O996c/s4bp+AKwczsl6YpuhIAzrcEzTdHu5bRFhQQ9JQMrzOJMgOb
/bhmpU/S0UGABiAF8kX6mbuFIa+Fa0lUz/Q+fygxk2UjPDwuCooUT+b+kQtF/0us
yP79DO82Rf9ypJyQe0lb5IM67jqBhKNRBrDOok7WFGtQpeOSLKHV/lipRl/rAC2O
sX6+HSfOq9oSEUABNDKrzpW+CdVn+I3PC1AoR3WA1aKHhlOUG4NAXxVR/OZF9jZZ
i7Wf/pCfGRaxov0AQr4UWHk7CM/Z2jXpfJ/0AiRNe/i1OBQPFClYqmTZo0MkENIf
8YD7ARgeaztBawoJ04B7/iXWH/hs8ZsnKiNqYU28x156qSLcYxga5RjnEZn3LXxP
c2prkeMA+FnxQ6C4o4mJTKKaZWMqSBEeJxqofSoorlkTPhwTWT6TuN/X+QXyUCTJ
ewUMYtZucDcRP/brCR0A4sdH5TaEnJsonav8kMWWUjMrC/xxd69BL8CYn6FOYAVN
HfKc6CdUqZTlZ4O5QO3BD/4UC9xdlYV39EDHRRrwjPms/C+dHD3+/QNSae4+6yDp
y7RcFa6Cobk2oLR+d1r8TOT1vLl4BAYkkRLvrfiVD20jOGj3i3tN4hyg2eTs1JfK
BKrC52Fv0XuDjNjHK6yeZ2kdgUKiYJmoIF50ab79LNBGFmwvPI3sBbF/jF49P/so
hGLaCcZnph7btFDlpyTe5Lnj7t6CJpPGltf0KYpVUh9qhzT2+FWMVF1UF9SXV2QL
rnsYBzeUG53cUnakt4XWYUAwazeXDe92FaTiKW024h+70xIqtrkOUuygSKFAcKAX
FqutHsOBB2oCOXK+HJ90frm7b+1zaJ1acXhLapRcs4tlnbSFKK5WmPHdIDPq2egW
zoxxHTglmJCt3CUzHfCMQgaKJeRy4y/ZpSWkICG/7NjKJbrHC3EbRS2si+16sDFn
nopjwpbmLYhCvrVonmjdf+PZJ063khP+BlCZhQ0/Ab07EguA2rOdgMrZ5erZbIpV
AcmVB3bh0aoah7p3zlJN9mNGwACRIlaGrJOe7MzqrVoMVGfq3jeeSgycCeulpSSg
TMi5JLScNnlBijgRgPhRDH0eO9M1ekipJrpz7r3O9owv5dBZitDXNHkvx/ZZpQUT
bbjXxMMk/HdOn5ogrMfgYfA69bU2//HOnsaRobluYjDrealWJOpfqrZ7q7MkF2GR
TwRLSvkYiSoEkgxqpMyCdrhpfoFPSqDYd9/Q9AT6jH2AQw28wEWf9QhRLWNVWudF
Xqe+HZ2/MwAjPCQqxjyKk1f2ZLZLOPVNGPklSwQ4jgher1u3xHDcwDlZf2n6d81+
abfYtoWNmKu9SSTNs46TD5V479w1Yv4nbc5x2YdWvV9rbr6wrwIsKtuVOQK/gGsH
V7vB58BoRsvNVMc7cQphCXL3NrhSn7PE/Pw2/Yq/wjEDjYtflZAYcXyqjokljkfl
IXJN53oW459FMdZ8a+/7QQH5cS6c0WTjS/uXBzzUD9UA2GcEtyu4PuJn9o46kLbA
Wm1jDn0a5oWcpO0luThFdBqhPfCk9/bODM1rbV1ibTBhwcJUBqzrkllZI9atfMm1
3/JJqXJLB0zgp1O7mblbbjtDNPfC0VdG2h+bcvUwN9U9xFG0XE6Qq9YX/xCSW31m
UE+W6UfwgzPketouSlccma9IXz7tKVMeCCpEN6cMqHyA3x80pgyTueUGlgbvfHhh
yjjLq2Ov7FxH+YEflw1L3af7uYAL3QaDnjD99BjZy17uQlcKQpLheIKiCWtaRBLA
aps7ymGrIyhhILYN6kncaUnYlnBlNIWELXja8732OPLuQm0eSnEIlBnsPb0tD9qA
uKdxeMOcJW40UVh753CTeyL0eR0FXzyqbl20LkneYQVcd+Mat6JrvCfk+DYEFdr5
xTK1AhfAJl+AocotIQbDeb2x0o7kI4KQrG2sKzSz6DTltEoa4wnUOchZxzwmBRpL
bMojfUfEW1Qq2UgieAig0wPhu9c8DrX9ktog4dTK8TwXhajSRqhPc81KjK+QcTGc
PWi0brlpLFmCOrJRnrWTpVbE5NXRjd0Z2Pb2zY66cVLa9Ba/NBF4dO66Ypv3JxOI
N4xi14Qon2jdVdQqcRGHuVHb0HhTObmU0SJhkp/JXVRFzz7wGM/WHuHZ9CWAa8di
vNXBFV8at2mDEyiaKA7vrXGvQspEXKqFXNgKBjGAaoQm/7WKmVok0dBUjh1Nacj3
TPU+cZgVQoc597BJvvgb8qHA6Ed+Pzkrnt73DtuSIS3PdaRyJjbz7/7qdULb9pOI
Xkj9BvKHKDRcV8pJXKJMQnlnB7qCCd4tYCYqsF8tObwbWXd2nuTaq11XBVIv60I8
xsvF3n3uHOD926gediARSkHG9vrtp/NYZtPqEj50Y/Z4hFRc+XOIclKZSXpfiW6k
Mo+aTlopim1l5M6tQ/G5CgnhtkMGQrVgFxbxZ69aZ0ZkhuQFZb8ol6c4fkjq65RN
2cqqb7vEIF9gNFHFwzM3SuFruu4oJqX1PIfHCtQcHUszMeLEwV0pV3j3enZ9equz
6+Q6YsbS4Dml1n86ymTzwPliHeyk+jGUE597mP1TBKpQ7Ez+GaNnoYG4RYKyFOfJ
Ap9bwsqMutt2sebwrQLp2Lb/lZ/2xVRpOrRrKJDLCEhOtMIRc15ATj79b9dZ0mYV
dbNZSWnL139dr2ixfZ8BJgRJyn8siA6JyFX44RJL6V/NdXpUKiA9JrOdlIod4+g8
wqOYnl4iaLSX24eIqF8uhV6Ke/s91ipagEh6yoVF8CitCyEuXmMQsbHsEarptVhu
S+heZD19tNxLaV/JtVj3JQRhvSSySJQqQ/Xxe8QO8DLh0m/+W4JAkzNbAhWjbn8t
1NZfkNTGmItAAdMgtEikOkTFBntqvl6qcRZWSuqk3LMMar5inlj6pxqh8/zFO35h
iPNUXbBKxNYy9E8f7XzEd3PpzvW3Z7++oM5PfTktaqydv687d9G2z5t+Di2e44f7
P9r5sQ6rs5Moic/W0zgQ5GrNL4y6Jhcqu512HQEZzrHOcMC7gohwzS6hQS+orfmy
DA4Hj1W5hynjzOp2plU+ylxC49XbzT5zSYcBILtKL5sHjuPs0tI7wM54ffufJLeU
6maNOAMmBV1EGHWN6vTg/tS1rlLb4GJejlnqfpso2/6SbdbVvVoKelSGw4ZVTFSa
+221ccdaRxm8MKAf575TlonFu3PVRSnq1PpCfsa/ifHZzn8aWLVxCUE5gm1B/s7z
l0I2BAEtlaongYKVmlO7wUSL5FgtYV1NE/eqMp5INCBQW5t3pfylJGEboBKndiM7
upM2SU2tm/fQ8TDQuY+M0s0iD1VT9AqJsdPAg8i0GLgZuHC+SJSo7rHUi9GqrKk2
uH2Ha7xXGvyxOz1dYuzS2yzJG1KR07yWkezbc7LRnGHUKgc5AlmJBqK/kDAr177v
KIuD6BRWkaCsyxvvMZOjTLcTou25ZO4WGsRCMquyRRlFqEkXY2im3r15/Z+f4ZeZ
nES4nSC6CYWpONoUJqRqDeKsftUlAzvzDWqWSkCOJqwxxUcln7WAr4ixc7Sw5iSS
NX9HE5eiwvRxZDRcHwjlsnK1lqbCJaVRVwZKtFHs89IWOA4XY+U605eJxWvHGHpV
tGrXcJez3UpPmTUT2cKYaYYCiJRwEmkw0WUsYanJmgZYCByo6Zw8TzF7ewT7YR8X
+y61X5+jzLrm28gg1JaBa6MhIPB71qT8prJpR5UhMdLLkqtODFCdAFjN+Dpnyadg
yBYVLIPY9MydbbNXrawLRz1MIijm9IvKOOnODRMNVnmjUG0a0lLBI7w4lMmDCoUI
sEK/5DXzTX7kxVfqWs3oBc0ADs53d16DjBV0YRBLSwGGQK634lz6yfTiqQ47Zw2Q
WDbIq+MAG2GZzGbQoUtDq0iu4laM2znqyzUSw/C9K3NIHI4UtxQTLmTZdwndwte/
QAuEiv4olw87TprpsHk0VthxxO4VegLsZqfzHdpXDhGiDf8pkWvxQFBtMeSeG8QU
AGGyo6n1ZIMHfEKoUQ6V3vJ5iu9LvT9aQUndeoI0o5CVciT912Znv26F50nRjm/n
HvYe1/yV1OqFsBxQbxt9ZvWNVmdaUGWWvdlWcEKuoT8v4DYIAS6fKabBCllv4nm1
u1z0n+VzVsUz3cg5Mr8TvJDg7gmjkJ+ZIrvDeKmBV/7yjm/sAE2nUQj5u/BARqx8
SKp7+63U0Zq8QSHxQrP1/ToWn/dSM68mtIO1vHT9v+70VzFa6D6jrh3pehNbmsLs
VgcAiK3FGmtN8Hj8F2Oxwp9vcpsQoLi/wTnK0L133lLbKVaWMUHRkx0WcGGjS+dD
RDRqJ6fuIxvL/VHs789TAjcHhpzsDqVwpIBT+lHO+fge2rYEN+adu1iR6CDHXlJ1
69iEZSAQxx9fMH5IeP9KQgH7iAWXoo7Ii1Mtn6t5y01dj1i7MdtjDnjLxZ2hvoFq
LDjVPfjDlz/w4RdAXE83nolhFTMF8Fa9olrK24rqxYg0ADWqqwMLte9xSbCEluhI
KJPexAWNpkcVOyiv2k12x/SEVb4xCcyhmYS4eVewsnM7GIeJbGkFi/Au08/5ZFM4
wzwm5a9VIDEMFw7rToPtwYtVpNEUvkr9xweTQ6Jc7ZinQyt/TgG9XMQwr6b9FYRY
pfvOCeJYDgDC5/+Pun3dg1fSNL6eghmwxhizxUGe9wdEj9CiJ+Fqc7eeQxri6GM7
v8EGveovAgoyDG8dtxK3XUsSPTx02ECJ4q+XX0R3qFChdVF92RpJ0GVoR+GVXjzM
cRXoSXCU9xV+pMg9tqGazZs2u3zL6Y4F7CZi58SbtbELQoCHgZ7JCpdXs+ykESzE
IxekabXrHd1851GxhIjnsQ+rSNLKetYX/O68xQKLpwkAE15OzZrPIbR7xyNr5t9k
nSnclCi+m63ZlyksCAXO1fZTWv6f26YiAhRaVDd7NyOMjSMhpoMBD/MvdBdgDorU
8xrMDBc6DE2HPc5+e1x7mRLa4qkz42WLKKUvhDPtjjIpaQvHM9T400uZ5A9SewLw
AzzhwpTFTNtiWzWjcsqJLFClotWi0Ejpb2v12Kqa349NwOmGlZCsXtU075yMyhpl
q12E4VSiKy7dhDt/IkJh0X62ZtR2yuBxATP7lLs1XYs4JBq+sVNbXboqMF/i+LKR
rRzf4EBJlypZDR3k/mUs4DC/B/gCCoLxtvG+ssgdK6jqUf0wMZohb63GZk/U+rKn
EmZGcAPdweAw6pwXredpRSyMJF1yrj2Tv4CZwyq2SEYQebZ+/BElHbxE9aPo9i9g
MPQIfrFYaQ2Pb2Gj/7j7uZQlw68yJA9gId5LWBzG7AbkOXOf7pEaEjuFxiX1zXA3
zYR859ylydEi/6GgXh53kfyWE3cucMqIOThhmxUWnZq6PSeL8cFb5fwq/hnvn3g8
VPX7esCPe+5caCA0h5IJUOl6als+3xA8RMjA5lQJtIjvLc8BUn71yMGSinGV3GOG
IneMAsWgRYdop4YDvtZbWxTOM+ikJrlUKrwelu3s1wUU8e4tKXbfQv89Bk0lr8HK
o3znt9CyB5GqO35iJIZp9FA31d7ME6Mo5e7wq/clg+hTVo291YBw4zlNYxJrcT5V
1WTHa1cCbUy2HczrpiOLfw+xniKU42zuuQC0D2pflUBMeN6JzrOAG84HgCMHfhq8
oLCicEnpVdngO5rJwC3hKWADRsQvNn3vUgosUYsGnzhL83j+zPV6jlUzx6qpk+p0
G/pE6Nexkwf8qDt6n8KoH8MnG8DA/27byHRzk/cvncrIkPoUXtXXfby+NhyWk+c0
Wkw8vhRKO539H4TfDChnjq4+d0VzILRZTElnytTKvWnUPTOrQA/pNf2KbYMRP24U
4dp6+KsCMufZ9uTV67cIzcgsrYb03FLXOAfSOVj62mit/HtXuy6DukdmohcJG1At
ULQJyJAOEmvfvoGft575EU/S64uJTl3iW2LOeu9V31WfNtvr8Wbf6jjvMrfzgmXn
QHvX/xljL3F6DG3u8ukz8PNuIo2VLHXaH6TY38hxx/flYouuy4DlAcrJd1sqNsq9
YTFJ+c9G/OD5tdXamW+ATriARMZ1D1KVkjc6ZABgoEYA5CMv12LDVnRSMY5uEtxk
JPLbGPiJK8Cw8Oa4MxYuULBqmm81ygaeJhBOhQq2pAHb8n/+fTwUSnL06LusrrBB
K05ONm0lYjT2V9x7TefA95Kq6rBEPekUO3vgZiHnyfVXgAxE9uEBXsBrAkabhghy
mQ9d6xmzRbPaowbPJRnnHcp6NYeZHssIYR8uoRpBgWg5Z1Tw2iWob5dyJZ6SmOPG
GNKOP3entpEx2rXdGnOEPSFwRgFVr02hph/xoIAxBpJ3fjb2Th9bCSfDMtlAsy8S
7IsG9lCEfqI1kGh4lBUELWvyGcZZQkupp8gv7zoCLLLp+taSHeoTsVTO7VpELvgf
O6wq/grZxw+dsTKABWzNMceBgUdEq0FtvpUbln/Qy/wVBhE6UaiCK5i3J+By6si+
XzadrjEmiaNcaESiLKu2CS035KsKAM0Sn/ny1wWkeawv44pEse7MTEeg8cBIyDY4
lW93ATorAjoBSbD9H8ZJIkv9nZBLig01qRomn+zNSa9zJE7AG2gFSHf8SO0k8s3y
bUiiPsIDU4jevEUP+U56OuAlAMN1np4XQ5ueKqJcwbIKiNXfd3BTE0TiL2JiPkLe
ZaKEAd53O4MgVw4TiJMe/KU3rP1MERzksE/F2qPKzm6xYAdIBAv/oclzR0p5w+r8
xz/3F7YNlRoi/Bpaakf4nIaUvdzlpHqbpPHmsN1c3XDrRodZoHqz0jrYVhl8JiWC
h9G6BzI2p1aGBjTNs/sOaFNU0tLFnRqkM76Feo3Zr0jQqk+jFnLTWlm1QlD0fzVl
ALra3mqVNwVww2WSZGlOS8vB9u8/l4ZiyGNo9JkwMXjQxeJTZ6E9ugEQsZcG4sPR
lw4mdgTHDnwDogQMwPiOdN5DjdUFWz17A8IhvxoAkAWZNom3xTyVmontUpsP+muj
TZbXuWVkxVQXONIepzgO5qjk13Xz9B590IhkeboKLGYU2qjIHksni95cLoj0crEI
KvEuAkwiFtibwbTsN14dPquLrRf+xVZEMIlGLP2pOKjlJnWNdYd1XIjXcCT1DYG1
XOESrpWoWv5kYudYAoN3+cqHJtyd6WkKjc8wn4iMMiQJkUWbb3BNEsvAdqyiXt9x
pPP6dr++UqmkqlIi1wNkuZkvbfBFYQ0ZJdelpolJgRZC001KdCqoEkkB7WupoLly
V16xOgLjohluGQcHmddtU/JdkHPX1EWN8M9XBV0trEpagehEWW1pK8x7Kv9xlD88
z66ScytdU+tv9MZLmjZ9ADy+/21ETvR4RJYofUFiFOnbOXQ+fKPi2VLaLrserEY8
y3srZLnB4W2gxBbo6MVAlh3BKBH/x7X2ipTyuTDClEXhVPcms1ouqpF4qjNE16tm
w+s4XGqmB9XnKmwT4VnuMcVaGgwutBK+nhK5JZTP6jfCTjU8xcJnPowAJ0QQXoCA
ZwVKrlp1BHTYJvstTbnwDMfCPnoK9SfGfg6xv+0eDGXW8F86fMkug8pbaYFfViO6
KpvPd+aZiACYA1kDKR9SeZdJtDY3Qxr59Rqvbw3JaEhqFpLVvtqiqAd1bdNIl485
tnL9xyXM/dFjGNumkxFu4Z+Kj8K5XwDCX9lY0aIyRyil8fREaFvFEg8VJZkd8iXL
chNIC2B7aL6nmc0MANYWRzsAMowe/ycL2DUMXKxPHnJY6fM+gtdhDZuJvc1+z+06
jwD1k1MtdqKzbRfnlW7Pn08Q43z+61oMzPmqM/+qSYNfqM4jKwBp3jqAh+mL5BIk
DwrYDIDHjYMHfSvL86MaNE2y3WbQmxzAL9Jc1pvRTckVRLLA1sd5sFbiAU9ViPyh
9iOlu2D4Ncgvf48Hh41i1y4x7+2Qp0agTglUjrRPW88XGKWSDXk0VATlX7LR4OG6
+wPgrdluOVuOgmtoF94Q0zF4bj7zlCvtzQ558ad7eoBO7p2mN+SS04SAqyVF3Myd
uM3xyzbv+p/kuiyyIvI4UYiBaYnHGZUL/r9X2gsBXHYPnRDZIryBvOJRn8G/YIal
Irgam1QukhHhvFy4o/w8oemeTeNttt/0FFrI+V3PMyZrFtSJwY7m9BCqaHyUUbbC
oUh33UAKEdfrzYKcXtX0Nqhe2PE1//2SaBgCEt0+MD+FQG09VhKartuwtanncVQY
U4eioy0iLhsb/aknckN/hja94Qg3TjbdhFHXa2dSNFFBSGjB5TeWyZVYFuW8DV9W
VOIDJ+2BdjqnfdO5xZxkbC2P1ZMEhLn9PNwpTFN1DrB88JmAro13BVFqOidQOl8E
tZ/y8z6BHMHqjO7h1J+sUlf1GO3WaTono/BJ3kXidKyU+3u6YMFIVsMkfhO88boa
4MBOS08TT6aH74/2PJetHFKgt5gtNDk9lSq27Mh3tz25s56WgG3wDt9smPCHM+Fd
1ss20JJnZ0Wn8wHaPPp17fA87g46TUHCHNRPuGPiGK7L9SqvCnfjostAg3gPik9L
IXK25fV8805SPEcyYu5fcUcxxHWU24B8IAEH0H+DDn8JXQUr0CY6hhRLXdYRBEoy
yVDY3wKDcZ+2Lmg5sJtCyYgcmwe7hl+xxhEpyvS4zKZjHuFlTrqmUoKCC0nHhxOe
rgSI3Tlk6+FramkdzEnoFC0XGqTBBYYcaCQ+YU2urfKWa8Od0R16QiDcXMoPlzRS
dXP4rutxZ/a1x2x5kIpS75glx0A+eWdsn2H4w22CV8oNfkSEsFlFFkLymNnL925b
89h4fCfbZd4d4Kj3273B8jA1cT7F+qWL1H6YPeQTTMDzVs3CbUxBOxTz5H4FRYHN
/CBpAFunPRhNhHfL0YMK7vczS+Jw3+y3WcL9NzRmwPSNt/yUroINJD7k01Zkcfd/
9g9/YpdYfCSpWcyGCv+t5NSBiDrgKLBix77kjwYXrVJstbDuc595+AKGacgFiAB9
/gEd6qdq9ZHUv27BuDP5oeQjCNKIBRNw9w5mqsPOpQ9ePHvojAVwMUeN8BJr8o56
RvuWlXXfzh1pGDcbmU82fk+eYgzTgrRqS/tbrzpSJRoLJeeTTpmOhgTfowpsXL0q
+MkABIGzuMTd++08c4WBNKEsTabcw0d6uAUntm3QAzRdaidcSSPA5J/Hah9TYeuw
uW+RBBPef9lgp91RBAULb9ASchAA24WPQsXZyLueWOZcSacKnVEhoqbKzgU+fF/2
7IUdUnLW8ynmOjVzxP/lzooUCwmvcSxK5fBtlYdEqAmcs1FsZZKM2Ouh4Sc44JU+
5CqiK4/61ohmFDsGuJ/6OjfqN32SbvbCmFKA+zs5Rjez2yAWZNyqCjjCVwJRFOf/
atvL2GCV7vb5iZYBIhVDsDENgiNNpstjob+Tkq/HfRLWQEsBU3pn8VLPyFPNvV9P
XgbeBYNxtV2Y1y1Q31Io35aUG1Ckd2lnGZaeMCbnHTn7xILKxeoBdszhGkGcpyhE
aVpoA9xMP+V+1wuQMdqJ7eqA5EIJv4DXAwQBAyolmrcRBHvFbIXb7Dm5xf0ZUvl8
2vGB+p8zBwGhfvoNdTk5yB0zQ/9lZZK72t9YjukhlbYvIsuo4dLgl1rJeG0gheXX
clflQLLZovKrVoWp+UcXOI2cvyJfMbYDqMxW4RGj1cLmAAF2+eZS2NPVs+58lfSt
v6BNWEwieU4n0ZILH2borymsSZ4oiR2M9SdSVByMKe+kTvtXfpqvtOHpsQDgIk9J
LvyPIymJzBJYKqgufcelM/SFZ3pCSm5jMjKlUeDiiuN8MWzB+25NEdG0FSdMY91j
ILk5aggubd09TPTcHu96s5GXd+Nai7UZhJDNdRy/iNARjZwljl+O1VqUJgvUZtHu
YIo/78m0urBXlqpFLs4uDY540ahXFA2JkyQlZMCA8vtGWrO/3pRenOuHIz8N0VjB
HzRW5aPP4+GG4wkdEpm5WivpcQ7aNfgRWVDcmrLJ17Bq8/+iVrU6uq6Q8LPUoZNQ
F5ZGhgjmFPXvH9dLGsPB0mw6tAJNreRjnS95Ec9KwMhrkJprWAECXMVE90Gyat/f
cA9wwxSl9E1ZXHH8Ce5HKas2e2EafhwQLWeQsfs0tOKU25l0ZvBUsbhmEgva58iv
qPi7nIPC33kLRFSQeTznMfBnZHwq0WDV1TW3Loymjgrr4pRriv6pNsBEuMMOTVzz
PcQxMapssfAUrlOx6g1FXf5satX4jrgzz1Ty/r+by7AKabqVL0OJt+YLc6urv6a+
SOdG5MyhlA5CWHWBA2ektr/X7VJSycYyuMMt8XgpD9s8vwADUUi8uMyFX4zbzHHl
9gHQ3WAyYdGd7XUxb3mkGjDP4nN8GX52IYhdt+qim96lhEQFZKuwWpCwxIV+lhP/
Hm5vYKw3XmNsN/Wh60g1mTP6HtcnML4Nep+AbbsDGmG+hfaR/PqnA9iVJHiJNlFK
cuP6s2cIMMFmngAMpRG94b9ycZeyo7J4gHSLXZZUUaTXYFOJVbyRC9ncC/Zrcc/K
MXMUvc/VRIA4Q3yjZvlAxesqf+A4TNeEbEFXGw8+5UQGew6UgrC7e3qETOoNPaLI
sJDI2fiLBGLeUmMXs5zL6Nqw+ZOtpKOCpmSNmyACoAKVNcUvRtUFgoXp8dKmSK6M
kmGq0mJh3kpHvNYv/V9KTZ4lJEfpzMu49zxZLRdBNJATbDCoaGRqbLdJ8wwfyCSN
S64npaCpbPNGlvlgSORkaZxi40uxS8U5IBIgcBIq1tYj6Ww4+a/sCIfwZe5M0/lX
YTPxJwDtLvngpblgWuZctlrcMETfD0Hf6p1BpSmdNtUhyV7TOCQtTKjgObgeYkrd
xsMcBuwYEHseb9q5D5E9Wz57p+wBXLc4x/RPQ4i847p1GkyfLzsa1NjGeiHYUu7x
SEb/SHXIZyiL0rIsezvx7fFyTQFewy12AMX8Rf/AIBy2zUc5e+lzBYPn4bP/PxSS
EBv4pVN00555kTbuGgljblJnMlR/IAf7EHY2u7izP8wNkgS97n/b4EQn3rrNKnEW
SUlG4SVCJ4zUWSN+xX7+xncjNSDh/MXZcVNZNulQK4oUxAeWfGVboYHudrRdiVE9
EyUhd2pTLkd1QnkA/tI0Petu5R6bAuAeQLPVuwLT78sIk+BsMWKxEdYy5+gVuh77
yKtv//MuxKXSTcf6pNsMO7QlYC+2e+e95XU25N5UWMZ08uCGp5pD0OP4Wpys+Smx
I2AXSpOZx7SVYY5QGfkSV9j0HlOeDVXhnv11kda0nS6fBlvESdnlgkiq41sD7O+t
ZNMYQ4mAp4sN0QPXyCJgkAunFDcrj+IPC4gsLNastsgch5ZX/32ELPcGtGhixIuz
2GWPJ0RTwAOh3Mc5s9D6xObYivlpdjaf9IHqKibLs/cYUieSsQ9uSLmRJw+b7rHW
/ACgO9GdRmxnZYZ8WLUYGWc7cmYdNLkQfLjXFY0bNFn30dGdkX01s8k7n9sNcEIj
g9MLzs7m4dh7pdBdiJ3ddunUMFJ3UPBStwnCVCt95hr2YnWcdNeRyJG3IdDrlOeB
jFNPIDlZBjqmKu+me4pnh2W09oDvwbwLLGtkBuIuHZCEPlGfQLyj6ulN5lLMrYUS
9LRapttliBwHcubjlm+4W2E7tl8IW1qoReXyfXtW7OLR5ADqEo84ov4ikbsmYRq+
xk++d2dyhXxH/mUxYsYZeEkyOih3klQuIXcY8BEOGftkHVz6VaeSRzvn57WaGHPe
0Y788Exrh4hYnHVYAHIcM/fMLd/4rsChIdB919f3dg3w6yzMcS7AyGlsNaj7lqmZ
xyzqeKjRXeKXzmC1QkjioOuSk3KVCk/CQP+dRUqNBFaUQmHdKuVGEx4h5AbCOGVl
zAKZE8zkoU8tL7hsMtAa9OqS11kYr8qEOx8cjq1i2syT5r/Awxck7GeMGgpWBQSz
+A6uP3k+OJO2ZtPPDS8lMUUZj9iCctsauTruhPWLNiaglovEVy9r4Tr28idAB0IJ
o56RBdBA35ETChguxbf5lqeuImRsCPYWf2QP0rwMUVqdycEdGLB69EOKWjh7XHqu
QlHVYu3Zt34iNIjHjay3TpzZbHiz/9kEOXeiBiJyTgB+ZM4GxDMdPBp8uheoim8u
mIhOZn1mb1yaQP0x6DqS1GnsPnQh7ueJJlG8vtjKjgG4VataZFy7gaKVuLjqlAUp
85VyNc0r13LkGWCBY7vev+IbJxVHzhX9Nj2pt5jEBXMwNnoV7SE1viDxzH27PDy6
vW0e01NGlN3Xs+zehx8pV4v7aBCBHKfGvAwDDRNHTWtJXxwuGNTzkoTH4Bfhq/EB
sueuRytWAXMi5hYkd78mcla95WBPQmGqt/P7fTRl1kTjTGqh04orPOSDrnEtYi5U
R79CwL3bRcxM+8/z36X8Nlx2/3DnByHb6aYobWqJqMVkMlqybcQFDTmXZuGCR0Fh
OkHDqvOXAOc9GcvjF9wPv40eW9vT/bq80Bnjdk/UBj3koxZO7/xiGuVWedXBW6Wb
dt4bLE84SbPS/uxNgYfUuvm/qXnAxUozLth1fXjrJtKADh8MO+D3rz07u2DiXBb1
HVoJaPRdZ47OYxFsqYS/365sirlZFhOdzQns45ZuhFIVMWlytD86VZ5iicosmexT
sHMkObTqa60EMc6Vqj8DNTPZB7KlPorc6XHfowSptCK7NK1HsS4+9sohZowrAHMQ
3X3UTwSd2qy0Y4m1nwkzXr5i6ofTP0K2weMkV+Zw0+9JhSQLRV4klFMucecXSLql
dzhQ8GqykffnZ1a1R2S8kUCH6mWbfqbSSnvi27bg1tEZ4iKNpp/Hb9SvVbPTc0EU
/6DNSpMC8MWxiFkZQQ1Tedq5NhSAZRXc+vN+B2XlHAca1XgJ/pDcmpyh6+/FvF9v
PADbSa4batv7Fi16fwylkZHgPgfg29orOmbekUwJ8gYxbJTOreKg5Dh05Ir00dUA
LkzL0G4JpDx1rZp2mAsWfU7QYs8F/Agt4+DIclyZPUQqTBOdcF4rXRpGmUZoSXa1
T6dOLZOjIvWqm8BYCZ3Bqcdug2Df7fN3hW74dOOKFq4EYwQ6UUc2MyjsoiX9ytvR
z0JbH1KPQ9waBTfHepokOZnUDZGSQlPwc8ifDPd8z2/JzzII1exUbR78Cmup4sf5
8RbKgVaCwsYU0VARkdPPc94cJZrt2UWDdqy9VdB8Uegl9tw8hErzXsHYLvN3Zuvw
PFyIvFX0gKPis2s0XN7JaYiz+CWww2Hpdgjq6RZHczwDy9Xyv6Jx2E+C4ZWyU8Jw
ExDPfP7QwPqKkfVFAAxMXWcXjPB2KgYeMbLXS9APA3U28FX+Cp8U6qVr34x1Z01o
cokKSlxeTZ/W3ayhMiLmcQBMgDY/RhcyoEO9N5a1FJDzR8qpqefHvM6vM+ZxBY/U
UH+WNLgFeUWE4+BHTjAlu1AvjrpEShl3j0fas9Dssl9+W78gQf5v2S0cnuQruWUZ
ClcKAGaj5fpWeBkgNBt4HPpkI4jv3uRd4qqJwCqyLXjZoUt4IjFomIiURJ8aehDy
s0952ItxRxCSdS0wRG/Btk2iav6n0P7Sh4V66tms630r6j+IzvqL57MiGR4v1/8+
meW36F/6wBjbM8BYHv2K2JwNpiKQX+fdeGfU6+q4hhVE0TJGig1Q+9FwzgAcYOxY
MzvliplWoebQRFonqwvDatOHHZuhN+YngZ9gVmf+WZfa1uw3nPoDSy5plvbTtnIn
t5uziQL+MZlOPd7wWX1/CspGE4ClwI3u0lkLF0NYb9CUjF3RW6K2fOJgujzLCGrS
EQ+DGMtkjPNTxfFYy7a1jfnAhJ6NN3ZdUDnTdKaVVPTzFR4zQxkyDHzr2fpEZQ5n
OabWibLuyRUrUKVHHUXVVEALMyjhUCQgRilUWVErPJJNPtRS4ACGUEDyV51Sxazo
UDqGM9Fy0zdAVTVuCwThetXi0BdrAYCUToXDPKVf7GZP6lLM2whLMyLIjxtgguIS
QDxbmwmn6ynUqevTwYRA4I5PiSMmsEixKmcZtcXk2khyyaV479l6bLCmN3z/CR2d
oflzu6YteNk+qTZwHq8S9EnuOiIrZqJMWp//m8IO22G0lTQjjw6uIzT7b0t2Kff4
/qqPvzwMMhWNn9fVtKEid/tuzIHTFdU50FXVy3VrH/9GfupHHqEMX1mLeJk60l9S
GIMoVeNF+uRl5fanI1L9wcN3NpwH4lSv4QQHkkbWC65908wl2AR29ZUKvNAA248C
pM8VQlVCasb9Jovnl8Q4DGmzNtWvDb+xeZ/JR1I7gYkCCHHxVb7onMf5AI8hgZyu
cEHZdJZQCehG9K79N0dGAmNfnCpAG3EatjXoIewYCzb9b1zYSGtXv5RxtTYDuIz7
QEOxA7EJpdg1tnmepm5n/qf/0k6d6TxLl0PNhCuV/ngfUK8Ad8z6TjBDNRAceHZr
H7s2SWsNetayjkx3lWbslobrCZbxf+w3PbEvAndh+MmtY7Va2YLG8vp1ov/JL6Pm
EAjS8LDstbGE/VBzd8tWz/l44omwYuN5NHEbnHpUa/0TlacbRtq+qztwcu0nCVZ+
TX2rDc/ETQVveE+VECiLU/5HpBn9LfQuDwm87rMp/BOXCXBwFPQcPrWD290LSHoS
CslpwmUNDqeeWi8J96voWccfaj9MxFHzgfdJUhxj8JbFNXl385Ovk9kfOVeqq9CT
/yqqh7UgLqr9PZVx3DT+falsuLX0PQvjS+elv//39RMaQVK1enUZ0mhV/CHGufl6
MGfTY+O8i9Jo+NOTJIB7kLelSfhd2lisxjz6qcfqdzSOYFqD6U2Ho73puz8j3o4s
m33sDe+k+/67gVjbRI3Kq8nqTLhlh+3kKp0Sf+FKkjt/R0BwCbjREGJhGaI1oa6y
eljUX03eymGJ7rrsNj82QjwQYnlUTtjrwKAZFbmwYRuL2HaDOIPd08hdyCxSEitg
Xo/OV40oGcaRKvED4ES/JerkS8QJAxOOJo7P/HfpqV63J34E1RccviJUBcLRa8XW
9O744VKQw9gbAXU8K9cfrs+FTCjEOAFEp51oJr1uxDRHhkRsz7F/W8mIUvEVXGE5
DBVcuanjIjsDb2be8voQ5q0jI4CRC4jLiTvjLrEi5N6AgxeMmLDuC3RYsv8P5bWb
hGqfkp+Q1zo5Lfqkvdd/G5dlzaoIokp2o3khh7ScRCBK3kAgUBXOQ41B9Ex4icoL
5015NxDUnf7uQOGXXgZ6A54BcF/bYJfbew+H1dRYrqT8fWN+ReztHGvtnd4dqlaU
Jgo+Isgx/sO1rf4wrz+xgoVwiJ0rsISC9zizp+ASIG6Vq4di5jJDq5g9Nx9OzGz5
0HEQtdF9Tg1icTDxHBtwaJX3pkJew3uvBCeAjsA1zlfBmj2yie2Jrgbu3LHplM3Q
p9iGy5Z8OO9VvDAYvnMDTPqD8nVAOfvbR+/un1usfVI47FZYlb1EBU+bO6ajmBx0
kU67XkRhagTez3JyisD7jX247p5t+2ILkWAxXgSWXtPNubULGSRyaOEmKj5ZVFfK
RYbrOqVxVvdDdOi38e0yIGotulTiH8oMi1XfuOJMSerURjmD3x1vyzJFIgTvQ8Df
C7cQ7ZODZVI7WxMpP73DgRlvtIGhSrwls6Immtg1WlIs3UdgU8m3D2EwTPkx1gRr
NmoyObvWFmSP2CrHXacx85317iFmOfigt181QEbl79nMePjOdgZZ4ivdHsy8zHrk
T9sjnFhWSbHJ2O1Rho3LBtHFPzUIrpIrFAuBda0/b1Uvlh6PCdMr9B8vic/jvuLm
UdrouYRqIyqJugeix5ZUjDiyrNrC5jNtPQwOnb3D3qUEKipbZtmZPKD4fyaCH0Pb
EWnXRcobRjrAkHuojvMiYaqxwyoVrzFxMmKtC41HW5caXss56wu13XtoC2M/pmM5
J1ADjMaMlJkORm/DWTAQk1/ebFvfJj+haj8I727rr/UfeHUiFywh1rWXW51y7M9G
R9SOU2bZ3XQXMgPwSnbefywFb7CQPzTvXX+tWs65rRZG47fAWPGvW1rmtAHqnXg+
d+nkuh0Ub1XQAjB/xcVZoz/YItHYiPOyBATpOXg1D8gFsCfLlRSawJKZHiJTrXpO
6SqqxFUbF3stSObXEKbboQ6/wJifuZKiALg6PfcX54iUmqUsf/ji2XtpbleUXYt3
K3BCj3tHYrR+xXt5MzdfInHDsQOeROrXtDK65nN95xsp2hXuHzf7T8Nl+vTcWHyA
I2NyltnxiF+J9V4/czzktjUWXh/hvnrAAABxHs3M4cMxEhc13lRCws/svEO53rIy
9ThJCs++sFX5a20DzByfZd9pLLnY5FCgbTQw0JFVJatjQkmN8XSxxoOYgg+6+tFO
bGAU/j8LCvdBOFpEoup0TWaBXTPmTxjNRnEavP+SgHrFH2kSgn55XnVlEjXb4OXu
Qps6gBHMF+UvXUdmA+jTFar1A0xvo0FTbKBkEvyguDjHW4mts6CSdkDBPJKKuM1U
eWq1zRyJv3SlQy760K1u2U43rVzzPiEsDmF5NR+NGxlSoAUW+9eXYpsC7e4VX4kf
Xmo1BsJQ95/jzSgvGBIZfFGy9rzqgp2R/2cKr8hFQyjwPkGlV4i7D2ENxaTXKEl8
H052lb99QOYc2dPpGS3D6T8uL4ddhDWtALzjao+VaZy9yp2sc/Fcur3vnMszadSa
nBHy0Cg6Duf4kn8iS+O9sjKaNSN1KPnYyNe96y9l4QlOBPdWGeYsUWW7Kk6LI0VX
QNAOSJyhSDCsJROhc2GmGraq3fhMu/T5FqESAPmWXPOvzg0cznJ01vxoRp83L2dw
oDjl0BQRSt4wF3UF7TbEd2n14ctYcqqq5BL9w3VwwKobuKT14gzDxf/bUEBCePcN
dHAf4u9Lk3233xkT+nqh82QJmbaFjexxdfbj5uLG2JOaexi4FsFSooiXf0V05/C8
lxwL3UyMfk8302kqbXgmbZ5IQPKnVjOZFEfKvx16cVPKDUeIXoj0AMjYJ4kgCUKW
czD3iTjWXAALOjx1vCvBYVm/KSG0DyOtxxG3OtHbK50kcOBdvwGBmgoJCZn1f0id
jsdz1XwW4KopR1oq12BtjIDGrIZUGwu0msZ48GA/jBCiajI5zj5qeWrraozQ4E36
2qoR3aGxQEp2EJpb3W4NtGJqLV9gmTxWRWIrodGaKCsmAi3fMcPnvIajuUrK+pxB
hiXjT0qhQ13Hkac/slgDdFm4Yjao6kzlT8XNpg8/yCAOJiy81ZD9XBoyB0JGAXd7
Lsy+pg1IPucppD2RyV3PmAc1sAPZ25p6gyKg8eItrBmkfCa87g0qL8+W/aPcvPE8
YiF/zwRHkoLK5nhREbJ+4H42X9BUrX/8BJgvUSK9udIhoZDDvX/iJFg2rdfI5/U6
HBZ24gZh26Z7Be9No4ccFgZjxR0ZsM+1wlzJsLNFw7u1EKY9ra679Pg1uNU+HBpl
2ahf8YF+52vQfuKDUIdeEzuxyUGDFUpnDxivYhnddhZ+zLbEZ7uAI6gpw2IWKbH4
dOmFsxRISbz6eXfCeMNMrYkpI190ai0n0TFyPEVxI4R+W+biwJphzxcfBaxBcRXK
qbuYNawTYS08Qm89wf81MDFDeHGYYzsBIb+A6xwWCLGMIGIDslcDlMxjnrW2Q7v5
l829G/0ZZBRChnc7QOKUOWoFzcncctN8mvd7Y7bLyk/6B9ErcA9Op8Vd8lyOx8Nl
1TOlFybdhEcqS4cdiKPB0/ASpH9lEchpMg0VVG8WRu6+97YZ3BGSggsDo/DuELMO
5LMTRkX64xBYaK6Y8/iXKChPHETTHogdCAXu5eliT/wb0V0S3bucng5SXwMmQAU7
9LgEU2fSpeaU5vZocjTBdkpba+D3TKbtXtLN9IKTvMpWlCsP5FaWMGH9oJo42c5T
zYdI2S+CBrdHpwL2ZV3OASan0YnwcXQzdgb3xqQk8Sgr+fS9AZBqLb7bs4/r9vZU
0EWO5bhOexrsleX7qFEYYpvDhzf72lNSUaZs1xnpGWgHGQFN3KsXkR1h/YQBwUB+
SX8hooIWOEJC363CE/OFEWtUKhTwkN16VlZ+AaSnAhFonJAnJSUXnSJCiGA7XP9Q
PkpTyCLTLcVoqrHki0vX83Q8LWPh0I+6MQi7dZzM2gi+ffAIquKyUe35/qMCOg97
gl/VKD3V4HdgrCDX7o9gLHtSu+sGvs/w1yLcT8s0mioqiSQJu8iHsq4+IVZPNL6X
c7IZb1GvxnAslDhw0DEU0P+/26xqH5utugp7+SwvcYKD1hEhb+AiypZPUF1Yb3Q5
qz3bq3vmEbOpkvwo7mSxkd4FUKzQEGiP1zPvUGJCUmtphaAbnI3ZtA2F9fPQIdZl
9rWtZNcSrtjzv2vjvB0TavuIGDVOON0eTGQcrJoH6TEWLf1F87PVdS4UANYO94Jp
SftZewkXBtpyB5S15i6EWYWSV6IKsExYIdGNo02PB+nkZQwGUDM5nnhg51gXVbpC
zpw34ak9xAQdrjxktFFChCLv4SoP3DA6cGvTmwlNdb6DPwNEyoe3cFV7GTmiYsnz
B6tWLIIOIUSiH6mtdX4uO2QqWE6+nApHeZTrVRXdz058MYogIdetSAJWmIUTbsFi
3W7eXG14RVB9CURVOyWWJpj2Klsvc0pwL+MkWNq+KCWfwi7QafsMB+8/atLQ7+h/
fTpE0gAFwWoU2TYaJqUGdroeGY+uAWd9Dn+3pHpGkLFn8gdyCt8pjtzLmWQsJ2YZ
mpWa9PlTGU6Rpa+DEYQHjlWZRpS1U2QgEYZ230tkzyBzkeGZWEVgQzQsNf7nExZQ
M80N7DGRywLH4CQXxwXJ6M3gEU/cwdvCJDsS0ykUYwrTI9+ios5pYLwXAka5lA1c
p9xGaNFNKhCxMJxP1EGlptq8DctnOI9TjSl1JbaduArnjnBFp1A7YTNpNLywU3a+
9e+u4uagbhEvk+HCMUMgITYkvNe3a19DiVT0RSAWAkPfdl5CZC6kFq3bgZhN8F0q
gL8ymDm6wajj7wSVCnxPDkGvlvkuFw8x2u/xLvd0kbqGOX45AquM2u3LjfaEDe5u
UKG8TBordvWXwxpX+Gcnot+Ry2RhUtwr5mJhGiGeK/Fd1dFeoD3a81T5n5/P2uEs
HfMhBUJu/hdjdoPi+15ogSIgAtQBehm6DqQ/AOKWqELw+UKVQIdKy/8h8RhEOaOJ
LHLksVVogsW7HBnF15PdGqtfObaUcp6Fkkg0Eb93YVDXPsbbHSgJ8BaI04IzoVDk
E+afc24gJ7tM6d/Ykc35PlpNj8MQQQBLUBZPwiTETZOvS7ALD4XBt7hKx2e+ZTPa
n32y3bY2L6z7uHgetcTCVMiG4058OHKTuEHOIyJspo7hgoJYqnDfOJ+gMpdfuIeF
ZqD/jYWZJ3wn1QAJjzjBhtC55w/gd9CZLQ2OpGT5/MuKwaxJXLjSGub8UiO8s5ki
LVS1esE6WNIdqsGfhAWhoy1uQqI9ESBSh2bJvHO79m7KDON+5USwb7dsFU8mvoRE
qjoHzie3G1oxIIjyntZ0wPzbZ+x76wh+AAvmQ9e/jkkXfP18GFJrrXLDRhYiZMIR
YueGWdJ82IHR2BcDnzL3McR55jWC69UXng6YUk33gg39hfInv4C/XNTIoaoZqGSf
TJ512WgzCbuOVCYCOfnRMSxyf9aPdvCG9KJNx2B04Rnpu+9tB6vz4jAddwXEe2Zp
R64mfwNc+9zxK4OAOgWyeCgJntsiWfIrNHZokuCWMRbb6bob7wm8397e2lZdC6OB
XUhFhvvrxrYtxTnPiy5wJiuqAIsCMt6BzTse4AQF4+WihqIWeXKW7T5PkKaReEHo
uUVEUGf6xXrikznuflxtNBnhaOKznATIJMcWFNeX9jsPsy015sQDaYJf8uoeKdoK
aFeUdKO60oWZHTaweWwKC9/IlPSe7l78YKA7Y4iDwCqHZscipxCq4Ij3ZnEf94D7
qk4JygVO3exI0NGagZ0xlQxUmuP2nshU2lsgQ2FGEvnBnv06eiGbDSgWVODrOR7T
8EUvJk4merly8XVSAvUvioGw4/Gp45Jkw2wZjLdxVDv+RWmVPrfw1y+le41oNYaA
wm0sPZPdicFUY5HQpFYEAIc7H+lYnNwiSq5t5LYQ/9eXjovUCdmjBZBN84HwjX7s
iQmAM3lByzQySYnK7XpNqVKZTSrSrHpMXzaMEFbmMd+VqfkdT8UNqvK6AJijxsZj
gfwJk5roJxVx8PQvM0IkTYU2WhdAcU+HKygpNlnIKS8+7mUGuw/ML17ul7BqeHWl
tXy/baOLqABryaxkc6N+dQq7bWenWxOTucGiyesLSdEu+JodiIN0/LaLM9/OQJBQ
sVCqQ2AkeyRb91V8PEf5kA8/bxWYooRyiII0Jv5j7VdfkzGg6txFWSwY5mzXW3HD
XyKEkR6HXTjLIcqdYZadtCdQs8WRlj75M9/hUJEQeMwUZMqfKOKt7fvC9DKQ0NUh
j4ULXqR5cXgIUKZo76y81gJPnd5Y3jveF9TRvvM3yq1OrZVjb0TKXiIxGMdk21z6
1Gqeql//aXX3d1AkW3sBnTvhtxQ82xXMXiMhG9+9A0itGXqtbLWi4yF7pZictD05
keTLf794UiysbQUqBV2V8IYPABaLQePaXNtSiiiBuN8B/zzCj6pI20YkwmqLOlNm
yNdgZFtAjDCnMCC/wKyUKp19CGvVzHJ/rI46JUT143MdBjrZAqoPBSJGwMtW9U7u
8KDN9i4w7ybbYDMZ1Cn0OSw/9KzuxjBC7IFPZuO4US8TLH0Y02YA8dfsZCqWhxvW
3AlMofS8P97ikYfLfVps0zBNeyLumHbOE2GB02oArhnrdbNQ2AAEgoDFQUBs9WZg
Mkjv8HqLxDRzEniup0e6U55rLUBFDEfq08ht9Lr4UYEtA+E135w0src5gK7BRUo0
fh71dQY+CiJmCzkieFY42TaWnwvTiESVJFSsrxXUffefVA/MIlAIEPrKL8sOu700
2Jt4valSduFJLqoZ4vxKviKCCQder2f+A2O9x5rUA2nUHl+Cs+xbpoRQ+jNmw5rt
koWxFdDj+ucLo7H0by+7vzadwEtMt37hc6AdBSkehl+J6NrPLhc6BbpSl1u3OI9w
08hFdUX92SeyCUcT7HHkgNt/j2zdcF2pHB/ZvnMSrZFulbL3G6EEAOc2qHwF6uaJ
n5T18b+Um5IGkjO4lOBJM1zJinN8iuinm3Lk7hDoc5xmoMsVgo7c05xMHuHf58P+
DLts0DlZUNKbtkMW1vRmBxtWRiEcFbjiJr0W7G5PDTz55H7KKClz/Tw+KmpGD3fr
xSte09vwn33u+YH0eXTBf+ovXE0B+9JWLhdmh+04z6ydJEW70kyYblshXXuc+Xgw
zoVtr6jOIZPp6xvaBZ2USywPJdG0ILsiG5XMtUagT/TWjhrDhPcSgn1drvgu0g+m
woHc22Soq7pjNJ0iRrIPB/nY7R4scAwZO/VSUaj56f59jLNK7bjMBOMKmPS+xXbm
b65t0CIdR6dEaF773cclTBHd3vi7nnfi8JomvkehqWADtDF6Owmn2MyRt0qa31Ri
MGB0WWsknNUs/6D2S60HcEQ8O+InWUNT+CYt+lON5MMkHxo5EDsHxuOWQ6T/tIdf
jEI1yCrE+d5ziso4x9nMk51nvDoyxLxXZ5OsXhgCxA1NDPHJOMiJHaJG8VvSELsS
dvYOARq0IxQat/mfemNaSR7SEe2ENqz3y03J70ySkSg0Vkhh6UuWN0P+y9ZL8HAs
TkCsMrQOUkKbBp6+nw8T9kjLaN7tl/MPigWbhQce9xGHdWPHAAXwqghOLxYMfmrv
sH1xv6xIj6rnZMZ5krjfykhSBt9upjox9cBZ9+aadIj7EXgFfKYxN09Qicjppl2I
1TPeWDnS8ZdzTXg9Ku/gJvB/4ONFTM2jrbV1FNzmuEP9q7XmgM9CWL3do6R4HOED
Rpkci7ZSdSEvL/quo98Q8mYwu4fbh0j/VpjsYa8CFe9LMu8APRf+n1UHSKqH2EYI
xjX1zNYWIXpn+9wnGcnC7vgYi3R08AXW35Y4CnwgFSwrss78FddoQlK6bRVjKs+i
BhcH1Rm0+liN93iFIMZYp3eS5DDhLpDa19M4Fxexa1h5aq72qbKPKJ88WG7tvM1e
b2J4HpLyD58zNUWuWTi15dTO46lWyArdqMxpL9Jr/D5mbM50hGKNeu8x1o3E2Qe0
e17UmYjS88lHizsun5OH6T3nw3snFyXESr8tjtc3JSlWUHoEH+kVDuNtbM1XUSOX
h1zZLPZB39V6v4pztu7Mw82G59fR0AVUujpGSxNOJhDO9wVUQo8IZk+lMBbY2El6
nhNCdjqPGCj4ipLf9CeWDD5IfZ7Rcwx7WKYzUGz4Iv/paEyq5/AtQPz/PGck7XUf
hnwtzepqBCac1Y6D/TDLh6iB4hyansnRTUoD0aZzTB5M3H+mX5BRJV+fA+B2kTRa
JvggI7faf3iBewxigkRonS8W+FO9M4WWHM2U1x7C7vQgzT0ISlzTD/0MMpl0bqo/
9zzWMm5R6dL7/pq43AiIw086ACh90bHLlYQng8HpHN4nGcyvlyYBcdgnubryHM5H
8QHwFkb2XLZCVS6xq1VNRFTIsSYMTNKQPV+Px6jcTWVvQfAAW5vrJsPQrWsYkUv3
KUKYIlDqj3KHaqsvOE2asgbULpnq6bhMoyMhV01TL78hx579Nrql8SQKK0NHpEhr
kbSIVPuVtPUnvlui2ooxQSSxVuIfVrfD46BOUdyaJabZ+lrj+2eSRa5jQCE2yv6P
w4JeYAH0xJathd0NiK7/yyTxpHzfTGAkg3xTF29ja4A2F6koSFgmJD/tEfr7k0Dt
hey0uzC/poJ3MpfvUpxSGqq4rJiLLufVS/gqIIv9BdeCK70w7r80zAho9sViW8U2
UIgqBmNJdpl9MGC44GvzzvfBlFLQzoVEl+9Zy3260XHGhU3EHRkM3U+smZTF7bpm
ebGfkTeHdDKbgsRacjmTHNkFXqukpn2NxzoaLGsctSUI6nGT9ylEN9XnEiY9sfgl
gX7UapJ7y7nQbG2/XOEr4l6EorbRTggAQyPEKfImdvJ72D2xwyJoxb9yb7Ae5oTO
3U1hRt+N0WA4cN7smHH8t8oQOu7pNMdin1Zbkkmc8z6WLkhcXebxQlslIGsExuXW
gJy8imbMpHCwGzKo/VWAdzlHkMHse9MuFbSa4pX1lJHyWI1gAsz6ch4U5czeEIaI
KAJSGdfK9Y4YvM5mQ0dyoP2o5LzoAQJu0MpiUayoIRuXJQgXg2xzK3Ush8VhvKDF
ea682SkIbSFeJrRDZfjKZFiGhB+Gfd/yH6w8kuZS0GvyhfeZSbtroNvhsUbTQJAN
XtStlNQ2x2yG49ZvGLsjjdCDSmANW/KbzPEJu0cTHggeNMKRry6OX3KNoOabPla0
P0qx7uR5pjeQIzR8zLtHEI6R/JLhqd8vquXRaRdY+5FDKDDgAwVNyB1dQ1nNQayR
zeSQF//HsH8A/FnDJqG5xneF3sFnfTIaQ3IX9E1YFGLKMjYFh1lrgKdia7q0rJW5
5bTlihaOZpe9wZv4POvjA5W4yxWgagsqvXRx3RP8KEUUikPvC1QcttTEacYc4RwX
AO51mahjI9fH77Nf8uy/YPugz3F+DOHYPSvr1PaZQVcIAnvPzvOXvMqoSfoL7kB1
8PXQz9Mo0hX/H8WZibFjQrUxHrI/ngJnNCeVXR2euSBX87xWI/jLKa015f1HUOcL
4UIo/Rz9MuGMFfHZlAgb9CUk1ebvM78UPBtHGZCjGXwr3Hotk1LU0RIvru6wVlF9
bDkqs3gEDTfypuqy7hZndVdV4h2d3rSHmy3cH2AjOuyimK16cTE+UumPCQ3BLTyG
yOyqmdqzyVkBoDfm1I/d+Y0jf+CqwSm+2Q8z1altD/KxShXSYIoooHi85pSAwGj5
By+/vpDbmOdg6ewBesIVhIioew4TdoLDYKT+mqSDw7miel4i7vGbo38d4RAW7NDs
2piK6oZV06B4XTStivJUrAnIgPhqrxx9hvtChGg8IOsWGXYU1JIgcZjxCy5y7TbT
yuPPThS8A1x1szt6UxsojOueaD2ImsxY0IapY37Vr2hQbD+t2QDyf7fghal0ei/u
Fryv4gy/WR1DaFbP0Go6gHQg8SOi1MMDVDsmPQioITuqU3QceWatp5K/b3JBhgyQ
NFsVafOITP9tQejbXw9slxLBuePxXoetuGeC7D/F59vAAj7YYWvLCxVSc1hyYx+P
MyI0LUI1nyVt0YVkjkOnY0NfsNOPS0DQ8+iQhvGS8fo4NDahFv6zi3HrSImcgoDs
q7ccazib6ithv6zMT7x8QlmE6hpXDNMHcB/QmPaPvWcBZr/SUlycvKsGFZJm4u5k
P8Xm4XGttNEphr08nOvNgCHf5exJMVyO7wkKAeIvWbx+7tUXwG2dYj/Pr7A6LNi8
6kb9qw6CyM2OM2jBxS+lB6kY6jF/Qhp45NZX2vpHnsbGLtmkdmt+2EQIpSc4UAVU
N6TFmnSrS5XB4pkiZoSl/7JM6S4ipCfsflNneh2Ohub8pAJQZ2iLEJWW2L0H3Xge
WiPEWrL3fs+L1h29+3r+bqj16LQ7z9vfkR/H+/GVkpnPAavUWS7rMypKL297csxo
adLYMdseKeCBSyNCfVq1FDgzUiL9wiXhoaMWMisqMHm/MzJWQovc61fkV768FhZe
hsfCmHNtt3iMx8Fa8tlp7xFJblhNYyVDufqEQaWi8skn4UykYL2itXyWtSIXTXgL
umDVAnI00n0Hmqj/oEXMms+X+XWpjub443f7bNJ8CdV3HbgxgKme5Tcat4AnKKIC
0WS8pomhcIH+Yfvr1c6QGxdn4/nYHuLh3/dUWr3XvWKYG2UXvm2AHgwEB2LRKi8v
Rq+xWIiqxxTU0+mxIawUjdC0Vuuywo/L5QSPJ0Po96dQxR/yq12TGzFvim0pneZy
skrlACVOnQe1EDNT5GI+/qmNV2kI9ovBXiVZ4QhGy4uJok2cfrJ+avWJxyRBV9EF
nhHi5qZJB/+YVCnd8ZJg+iFbSCPDVt2CdXt/XCeOzJYI/rL6+C3IGF2T8CkVkSvb
OaX2XXpy20fI7O5UnFsQehqtY3tP2SoHJucu0WeCqijf0raPBNJE/4JzAysJr9Tw
0WCmIYSkWMeriTcBLUw7SYzZhA3+HNwEy3urihTidZR2KRRS8ibf6AAKJ4D4SVKZ
XgMWg53Bl2hogPsEyPIJivWfab/0XP+Uxb8XAv7nPimBiz1daswj2tnEBo3jOcBd
PQCKAn33qWaDVI9hdE+zgOSbWk5nl7rVi+1RQZB65Rzta67jS+GJKfgLeDzyEQn2
WbL6u2PbkTRvDE2b6rwUGkZxGjOf4Y6z3uMuvqjd3YgmcxCx2XHAQ1kTbehAwZoq
oiMTMNe1x4zLMyxBhe1kl0RC24hdpr+VIoWfpcqrPtPx53XQIBtwz2u2E+dnBTXi
THiOxmySzW1ylVv9GwmnfrH4s3Nqm+iqGfoIqT3937152/loHGhI4rcl5vtxv7Mg
pQtFyFNXMLt0cSX9+WcPq2Jv72z/+BwpESkJQdfmfPLzupw4g4pPJWkiT6pZrF3w
jsZ/yBk1WeLq1QQyQN0bZdLTrhYB8XlBiAVy9RteBctOCm4ojxB2jWnqvCchPgcs
v5/4eAsadN88YUCUjlO+JCXbhL9l9TArG5lafQE40431YdirKvL/4Lr1jkm8pu/6
sjFwMU3iW5GgSTg2iwqfqyuWv1qQvu4sJSIHTOW7O1Xze4V5jIgREinTlWHSPyHr
ADpmEaVQxok9OzsaB9+dVoaZoI8KNJS30BKWD23FKat1ILtmehpVouMiM1MV4SwN
bD8ThXYLFfrPgiDpjbbxOlwAirWN8V4CGzyrOoead72KvpTIRWDQP6feL0d99fqd
LMzImEX44tsJ/pg7q/7ciXN6gBbZIzWtmqjJo3fQV+eWO3SIvZcPUyIeP3LWK9+J
zb5u8owiG5kBMqHW+pzgMxcjy0nijhhUXKj8zPGT/tF8USUGmErEhC4v0SMM/cY0
bPNSdEG8l+8MnMmpu0H3OFlG9TdHnIxbMtweUEOqXeVA4qk/6ZCLtTMaGGn13KMh
oeaCjXDE4Ae0rxHT1X/XN/itswmUmwXUvUXfbm8SgcfpKjUTBbWwMb8slcC4Bo2v
LkQSzzVGaHLlPNE53EewpP2KVW4NNL0Qq9YRuFtqlMmCW01rokodRR8a3ySKn33P
VrTr1pMGFnZpHYym8u29uRsTUiqK2/T6fJ2QY+ePtc44UKnlIgjXg0LeSbp7eTjW
VGs2uNaI8lFwwW7GOzcU+hMsqnsdrL8kulLv3eDuKjf+bOXvrhIogIvvA+A/P8fL
uzT3WalNFv4Wj4vND5NHvHp1+mQiqgjPitesYECaK0MvDix+4eUen4iz3PUxb9Dm
xIAMMi3Rk64W8g2n9QE8701hgkDv0+qJXPaP+XVU1qzsBmeYs97Gv06FH6STgOxD
L3ayr0EQHPD5QDdJ6YXlXHmtu5k81AFQqR1WcH2wQ8UZ8JyqTMV3HG6ABfwd9l7J
OmPB1pfBfx1F1WJ6eHFHNuhMlckvqSklExI2VzW1nO+8Jt72fhUmyVAjZ+SlckwZ
Q66jOcbkQZLyorHxHjtXRmsWwKuGmsfQH4q6AHXsA/694xlNeun2l5EIMnm2ofQd
3eGB8yYw0NqK/f8mSeyKx2WPMeZ9t7GV7jG5OZyzdiXYXjATNhL0+30HLpPyY74g
keCtl71jYREq77Aqq8UM9Uzyyg0rn2fgr/soTL9canbiJhjzaKK9eOGUmQc8FPMj
j5hvn3dWwfoLxmtsLQhLT0vQOSt4Xm+9a5a3Q85RneO4aG23Yo/ivjnctknxBp5e
ImT7Lu6dxsTJwk80BhFnpiy6eVc5R6kvKmH+pNmGSCZEPghPLGnFoiJwosAQq2MG
FcSniwedx5fH8BUcqyee+nxNDjN8fzjfH7meHfcdpYD7PcudD9d4MPK5oBzLmj7c
F56OheDhL4I4Lk8OKpmb6NLB/J4XdWXzHDvCSYS3BLDpq5Q6xP1Gmph+/Mg9Lelu
D7TxWBTqfFlllHPSIRe/RWjHB52OXixDQCvNMmUfZ+b9CO0tKF8R1Wwklonh0Rrs
6TmY4FEjlAJqwwBpPmYcF46DWXP7m57el6UNend9rEYhPymIcbi/zFzeuFnJE76r
1gXdcA4dwYwkjisNC/T9Gb8FbZLJnXgtmBuFY6bXrvWe4itxPzdVAQ02R0DC5C7G
I0HT7sTJpSX0XPZQbxknPo/2NAwgzrqQMSeg1zemjGuXgtWYhmRStsN7o1uNFDZD
TggoLMt1ZDH/vZresOsyAZ0TGZQe+fRQ+yMGWeHC3dLYFcvhlMZI/6zEhho+5bf/
fq+fj7PTiIm+Itfz47fndOrk6V8dBcV4ogfp8DCxz+jslDeriVRzMaKhZDhuF6ag
EsTE3g2kJJp/z+DtPk1Vp+NMk31eWoie1EYsrujYdaV2ERftRn7Is28RsxxOQgWt
Ap74/SkbUd4Pm+n0vMZfCKrGbRbTYOym/9dGDBKQgxU7/t4WPCFHS5lZnhsb+dT5
5r6qDko850ysDtecNwN9YB/MclnJG1hgdWrcumR+mK1JCdvfIDUjRdxSlyi+sj7f
td0LBHvOnu3Fak1K9dpocRAVCoo9V0UTvIGOOKADjiGSJjs4YaO3EZHNJvQPRM6V
rzqGFG0fxv4AtKp7UO7HLgn8q2/MXqyynxwYcYMvKHzLjTOPP/iQxehNq32fSFbZ
kE06YRAEVwN4c3mLk6fyhZGVh1tBVgGBCzQojj+4Q/ODVK3KqZLvKTBoUCnI/DYR
Wb3hv2YRP/zeKByywjtXke/Z6Mns39xVzADN0Oc+tCK1ZQS2qNZE0XojcSjR6rLY
RyriVqfttZFQj3FeKN8/NDhjOdatEmu3Z0AfdZ21LphLzzQyCk0K3zbUHeJiLmrt
MXHujx3Fu4Jnnk9blGPD/I3SjPb3UIsENc3BOA6c1J+6WiAlfr8Iogm5nS6Wlc0s
I80znvVHEicmF9lYOXEWqGhhaCp4gI0p5ef67yFx/QnsfV41dxf2tLj+g+BlQlYC
I0Js5wD7pY/IyQYSZP8NMOX3tc4uyntn5oxHPAJaYUPJndJYqjxcsBxhJg/WwjWz
mYxhPlVZyO9cXvisraJnGWaZuU/Humhtg63hLaFVsIRvOoGlLJZnuZqIb7xRYFGq
OBxuCxP72+NZQ8YnOGF6p/6YyW3fck8e8eL5sNrrpn8l1zVKPY4q+x9f6PgFdxeq
op+82p9d66+HLamtUMhNHWssZIygmvPN84Kk5O1B9Al1A2RPOI3U1dz5aHG30/VU
Uavx8OYCvMHZvjT5oX0NAyVQTOkPVYymc6pc3eIF55EgEGhJEbbdqcL24uumq49h
1YT4Sy9j4z7WrjkayvEEU/4hL+g9xtspIcyqpYMxdFv1843AyeOljtrlPD5eS16g
SSULUY5NrRcAQ4grJWWrTorbNQ8ulrw2n4Tr48HvL0OoIk9koMvSR8X6EKRbBnzP
M7Alfqen8gzPqaWIkQx+D/o6//WmIUlDAPQTVtFQweoWC1Wc065YA1iEGCV5wg5V
lGj/nTlfofypaytxZbOEMvQQAyTivIiBUQAS2XquCSEJIO4NeDxBnJs84o+43dlm
WkoBAykJlXFR1XWXlXIpqATYobnCS/lW9VeyKXQB3E2avOIKg+VfCRm9J4M8s8T9
gJZ/cfPTxZ2hCQ5CbxOzUbDkDaxIVYGXNu1i4DIpmeu+AgLrmY+NnO+NuJwm6eis
6LE7mO/x+Fn/K+tUK9tbteAQdkOnnJMWTW1KsOjDNzlY1pz8zc2uasC7ZM/9c4rE
XGkxihGNsnW6z0GLSB820Q7N4S1gE2jnh5RtzVPThtv2DnkvUOzLQcMwGHAWTtXA
VtgH2TPGvcKtzPTf4LcNUtyep4ybryss7MueYHyXKM0sTvS23ZuppFrLdv9Kn28K
ABXHaTkpmVTf4F8uWjkGf6f1ZJ4VnUc7jBFs39fprDwGiuFvcEVkWKNFCpPQBjs5
63o3/Hi+nYEYx0N/N7ruyzFMzaTQFqdJ2Ue8vQ/YYEcbf9oxfXo1o3d36iUZUSKd
Noi0IV7XL4XDoEUHfp44XTApPKHJx+gxY6I8D5R9PAqDQpvBz1Pd/G5PuIpIu9Wr
Kaz5Kqp9rDZyuPLbRkAwXrAGodJmZAzqGjlVnu6k4mjCzevEOKaYIlV1qwG2oHim
V5bPzsG4CVXMv+5XEIe5rgqnyZ2/yY0VbaOlsRJkwriI0/3wa8s4gxbwDV6jZn3o
UJ7yzUR+twVgIzymEkW2gBHGtlmSisILEFFiRmvTwoOht25bIo97vecKqaGp4nYa
ICG0rOWryk2ymDm56wQa0nls1kZmlsx0aortmr1M5qXnJgp4rE5sPjOOU9NolVq1
0T8GNLDp8d/5q6GQoZ6deLc8XFmW/HVtVZx1S4QFMAO1psWBz503s495/6RaHfJJ
x0piKH6kplJMOhnbXrYhib0xGd1TGSraflNxKjO4lLzwUryRs5yk2aCFroDjGNU4
8u9YwDhOwO49+H9o/0fnNjiSyr0mNzyDZ80YnRbKmotolo6pQfDLenSaTzZjMjSn
Ym+6SmOz35XW2/mpRs+l2ttw5YXrUzGH/TpnGqjiiQaPCGQEUzqrEVfpiNWM5uV9
Pkhpj+qVWIwjzCyolN/WoTs2UHfY9xBvpE0j6Vi9j9dRVIeTUmY5o9CXEAaioFgQ
/H7B1nskZWqCmnXc0eaxmXaFOMsaZljP07nR7haX4pLl8wJwMoaXoKSd+FlJ1gL1
IyfC2xW/oqfK5IGjsJNzT2yVym2Dvxkkp/C8jRGClxU=
`protect END_PROTECTED
