`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gi7MCg//jy3IEGy83QCHX+FNmAMqhdqlj8IiyZzno6t6m9IJuareZOf7ro0ctS+u
R1ve+jZaHrgSpf0whjNoGRUr5AHcmwnlD5xqPyHGQUAFGcsJ8GIsPOTB0B9QKo2x
gEY/kFlD1wkWD6PyhrGneCOFV6Nmxg7iOl3aMPftNG5ZyhCARJkxhfmwJpXefzBH
TVUhYUcXLxf9bGsAYIkHkto/KgWgBYaV4gPOsYwmEQTzp1B9poPQzGOeMEvV45TX
M5rP/K2ug9TSGugZcT1s6+pV3AbqHvhLNG00G85xvb9ZdvLgA1AOnLXnnmSKwyZ1
EgMX8rIfaSLfmjuB8jqfhrWSFVGLTzfZlA0dIZ7ZMutoxR4rAiYltPD8eNr/fpxi
t/cm2ullfhlIoLTXVyL0AtzEl8d5rDdXts96rZNKqPZqQK8bRc/UuEUfQNnN0ce6
IN/rmip9MhTRDw2EBKIYNuRmfPWkNy65mzZ0842FKj4bodLaVJraq8++wPwmLe7V
l0pyY98IfabTEowqsVh1zNedTk+/TBxKz4DgeWMzNXqI0FDPP9SkS48hGOonfFVp
ChzeAyL4cNCir5jLQ1tJ4qk7EULjaFVnp7OO7raB5PivSZbGzUAMTuhzvN7RSdO0
j5tTh2GcNJtH2mVJxTFuoKv4SpRBSb5p54fG11rmOket2lxJFyhX7cCCUagMn3My
dIo3CzgW96IEm5K0Q3RKLpEjZ13WWMAM4vu9Gx49HgRrMH/IvywAZyehDDuKxomf
8pbn8KsXCOz5afghexnyZ9KweMh295DNVKpO2DCdVzg=
`protect END_PROTECTED
