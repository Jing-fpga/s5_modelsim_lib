`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1D4LKYXcK5fEe6hPNO3niz+N7ZLAWV1kgdIuh8rpCWH0oa/hfp5eBOY6mR/ZBeuz
hpOM/OjNF6zDWoXwROExiaPeMdylF6xAW33lf59QkRHoDliMmFBKdmmVkUV6Sj25
E0S1seSDyGJqevAECD7s/9dScOmzYksKAnuCsvMV3aniceQOD70lXIeNEhIy5S7q
5mK+mBUCgkGM0/qvucRsAAMU/FxBStT8jJfuXf/Gms9I+WjaYzYAUBseeaDRzd+j
gOaaGKyVJu+Ys1h7cIWEVlxf3Mhc2lmeDWzz+MWPHfoJFyyQaJx9enVPChFCjdYc
nYeOnW1/RWwnHam5YHpd7fDPk6Kt45Ht6HvOTlQrmkAfROG5biA6vMVQTyi52CTl
Km+e0hUF8lAzZkiFjAn0xeD0sueuVvI7ip1k0EW7M3V/ZYkF3wqq/3oMg72ZxLAb
jw1HDtHEsxWhz1+ll0WbanCNP6PueS55WnMumogMzUtbXr1En7na/OozxvzpUIYW
FeswjYlRNZ2VdSINGKjDzwWetqgOxiFGw8mM9/0ZBKYl2E6RI8a4DCgOO7QHZrlD
32p5FSoA5aEjPD1aqNp6EoWmEvjLGxllmiydzzjRz1cNCSRbaAnYZxBypozSAMri
jZGQE837cPy0QMl+wDk0mzRXm991HyKcvASLUrpyHSFnxpaCILmDgRiElnYlK8Y+
QqfPJAukIUZoxCH8RbqQi9yyaOgiD6l05iAGSgINVjsEgnGrEKV2rwRfz/SIZ/fx
KZn2RB4eHygjTeXLnCPOLptcWAT2ch1777Fk9+a6YJphRwMni4DmtLsSibQH2/iI
G8DRCGJEa5qSqv10l8E5xbfp5pKxGlPd+sBvOil2FQk3tzWjbUis6+e7N9ZQYsh0
y0KPwJ5jwzvJvGzB2RZRl2AnFOakETpm7YIAId8RdhEQ3Z1NWHjNqFSx2EtjUwZo
uJ0HtcOeHe3ZvodAF7TozcY2+gxzy786xWvjGpEWBL5TWjp1JgrYmfFUCdqaFV6D
KIBdIyNmLJtVZVJRq/JEcypm+ByfULBJEpXWwvvuc7BmbmMsw6iUCeCCVVnzkKjl
334qycvVoADs6s7GGlLZvDwDzAFer/p/20FT8hI7C9guk4vB1mhDJS8UzrhZIqq2
ojCwPpl4fNNKptfd7AshK4ihOkgKImbcusjRkEcTy8QZyh2AK0j7u9A+MXL1Vj22
5LlZ3KIj1m1Ste+bd49jKwlOr4zCjGum+VpC/HHiJ7g15Wzb7/+8nSU5+FnjDuoR
eSXctTigjQL/dpl+ql9KQKXSpEeNs88zA94Fw769VpFVamjU7tLYUedU1ZFoY1kB
SFjHYjA+HqNcH0fO4wy+nsz2XIrztn7AJWlfdoVql7v4MfPwV8HExSuZym9JBNf0
7Pb+N+79pXoQfImM2zaDrhWYopg645W8sfBUE5FdlTbF+CWn6dbUhWEznR5HwiVu
3y9X+aF/Mt7VF7zjhZss0DlIvrRWZ5aHDqFqfNm4C53PVWbEiKGGZDqvPGhlt0hu
z6PWz2kaS8dGzHJjR40LvC+ED7pWdpTTamJQd6cENoOM6G3BCZ9yGT8aUe18zc2L
//OBtpKtYK1HgU2JK2qr0WS7sDsLpaNvSxuWqxI3YwHrqc2cbJx8/bpKLzx8Znku
`protect END_PROTECTED
