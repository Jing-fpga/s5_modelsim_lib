`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/mY6wCil+znf1RszDIVMdzNjL+O+px32x4maT1j6WFLFT+vHUR6pmVAXTWf8OnE9
ZyOaJYlfRYfAkzIpH0hCW6ihTlGDoFHmYXi6XA+TjG7rtjFAMGLU/clBidEXnTzJ
8OsVHNCIC3FuTaoK8LUFUwLTFiBV/giNZnjGhiGWpQHknMt8u0M8UJfJNuxi9sBA
PcXb93WkAAPM432TcV2nVLyl92hz/7PeGDB2zvD8+1oKhGfxSMoO6mIcsccx8e5b
qsdTGLt1einDUOGe2jQ706qpqoXZpH/EVq8YfV/d9qEF6OSNhrEC83zlDqpeL60d
S9L6dn5RhsYzqeu81kIzChcVQTZIWOLbh+S8Qn8VWMRnyYrPbKOuIc/eap6lAXtN
+U4+gC1MPaNV7CJJWCw5OIia3VM2mUHQ3BdKJGjEtRZYFMqItGj+iYDo2g8X6GaO
mPt5RC4GyLWn7NTEpIJU1rcvFex1JtMG8lpDHDt78qn0UjqbqufQ/7nv/ywFqZaO
nEpDTTb4uEknvZFQjcfYXNNZlcbPkhjSGlMQFi7vjcjNHVmvpSsXgKehYG/cAHCh
M2x+qHap+s8GcVobFddR3Xpf2qJ6Mmnge3cx8mrQZzMvNbf4tUFOcVpt36f5g6TZ
wQgAWO44dHQfzLXtS32/jRa07uslyvsHeKwAoqEpXf4BNW19UKLkK0xtha6ycGJ5
LCMeWdOV3nINqlH14mi1IbXYMSFFB0NynN9DuLkYnz36qS2Z55IMUz2BM99XI/9U
9cTDBcShV4jp+sahPUiEsnM+t48V+O394rRUSaiBSFv7EuxalePspAx9SCBgIYwL
eyiiDDvajEfaO3aOUKHpjLZAfCCY3iwxEJBlK1MJaWo6stwPHYt8t33En9v2GCVU
Munwayv9dQE+2w7Q+f8maUjBQLjJuh+P5rXthG7aYBll5iNp8dQKLV8sOnBoeF25
t15WADV5DpJYbfk9Oe2yYeGTNdstZMpBttPaVY/zQPHaMJpEHCiRygPeLwIcJ2EW
LNBtCMM/sbfYG9tKam8M/JjHFXddmCtPZimp+z8VpsfdVpYsnfDt5cMeH64ODsWK
BsuFCX5h9jLz66YcTS4kvx4H6HFdnuIcjozxN9BPTibZz6L0QooWbiLNqzOSa2/S
kvFanu2vX3g2GR6sNjGfRrdwMYbbx8b7n8N9IGI/Igf7o/GNCJsB+cdJl632ezti
DGTBLpBdEouxzjzNPr8X8ouqlZ88tWq9Zv/YpzP3qEUpw3xlCh7v2HvwKypeAH5t
NC8oc7UGmnQhDSL5Qa6lce//CEfqaxZdlrfhZJTIDmCj8SDvT8DKhGCclwz9jqYH
cPpUIqYtI50ggW9bWtPBpLUR0Cwaff1h17A7DQFBf5J1vy/tnh1hnHbQPO+KRZL/
KktR//bEIx3PDXlUBx0vo2EHPdFt+tsqgelHKx1hC7O4VF8ubweQTJbymyCgOdgr
pNeHOiDqZQWYL2K2D6jnJw21/XgRL3l2PX/JtOPDL/mN+GC+CKxwDjwVoKWUFnge
/8tECxIIZGKk0I501GH0TdpzruTzNGcX9F53j6TjlgnclTuYYjyHkdoAnYhAdnU+
6xh1lOe23Zpak2czZMxqnNJPE+5etJ59Nb/dNyB4nr55i+JfYjdhO8wyg9KGB/Wb
mmybgyDCdOdLUDhlYmyIoEmTl2cyCU1XLqMAMFrf1WoGPMHMWF20CNfv2/fO3mL0
9RpNCUfeQkRb68mXadI3JeJ8r/meH5FctxNtxWOY7QExaVzdkDdB+4pSMAM/Q2XF
pPcfiAA9mD9wqnQxLegwmgIL3/nt3NxlNr2rhSNVPbJaZAL+qCQGC5eVfd8wPrUo
c0Dw2iSSqd/Vx9CegIusm03hrRbUYlWh3E1+HAbY5EjihYAM8hUwfWfAg89wYTrH
2c2Hmq7Q42kqoMh4LMGSuujdpII2FuP16TN+1WxkwsKCjalP7BZOZT2p+eX0onkA
M/pk3jG7OupatQQ1rNtSEmsiI0PGGOOjYUvOhl1mJxkG2wswqHW94RoMxtePbrkJ
4bRW4GA9gh6h9SMbfNiO+8jWVuY+eFE+MgNnyNIJ0Ip7i8vU8VEGRlAfORaznpLF
E8/Uknblpctb4Ll8QADwwgAYl6Iw9Q1KKGmzz1ymQeM8ZPnQjOAisZvcaADuLzIH
KLJw8uUgztIV/RRl5Nafu6olYdPm6kwKUSbwbyGUgMjgurVyGzZ2iwd04U8g9tRx
/YZ+6urdg7MrgEuSlAdkUBsLE4WEi6kCM7UJXHLI338tvYfFxIhAsKCejBtKVs7U
1cbIzEDrXWETf/s2+5lwkxlKIUuPW0TamAp9sewJ12lgp3J1PHQDBW9gwnsdbW44
vEZa9l53Erx6V3TCK1+9zYGz9pj5X2JR4qQNgmyVPimEa/V3yQWyujsIfZDxc/y5
Qmu3Wsje6BCkyjw0M1IZkQwOx47KrPqy4uNbUca7u8AOKt0mvyKBP8z2r5T5JEPB
0H096DGk+XFW4MA/aUPLaiGRiSY0cM6B4SznZQHFlbGd7p289zJw9qinRhiZ4qyI
xzzYBacnLABosNPkJoWf0NS6y2kFTjmK2qULJc9M0DUvxM8OPk4Nevnhoetnzz5U
Vn+CPIKsSdanJEFJ08thJNmV/tdy5CbIkNKVCt0hdSGG21OoEB52KeiKzORz9q5r
W8y5yogs68hY/hfMeqqZGllMRpXkD2kyG4bC8Qn3V8o3GXpaFKre3zcn3ycuX3fP
cvQhxBIXnLqVdmBemXTI/fP3yRL7QAnsJg6R/4Jf5mkQI+zbpaciZxEofCLYcusM
6QgMQkhVN9aKWu85U74L3inEBNsmHoDRnegr0Yr5e28q1L4BF5fWwUGmw8BTQ+ya
HWZG3YaTdV9CCspW5EFJ9pDg0UzbY5CbNJGF3lCOHXZO+Jqf64gq0AXUmnb836ah
cf1qPiWd9OUnvBb36dK8IjYbIun5OBbMvIMkhYXh4xknHjnfWUYb/gckukVpQJ8x
8L/o6IPZa79ROEfhG5uaENlbaeNscwX42YRlx3qhRw/SY0eTLA1iRB7CQi8gf64R
ArPjBQSKoI3nQ9BUd2dGxgA/8ordFoTLzOp9lRoCJWOQ9ys/omMhpyJ5Y2hk1cec
P4RXJF0N989a0Qz2uNNVJEPtWdVbY1usFS+zFfcBVv05yI/GiHdjxVrnIdk3q3bw
1ZoPzba6xnYer3mwv4ERim+Y1KD/I0VmQ1o+8K50Xb5E4H+fsLMLaFBKR+pfV+kq
gTiZYPnii6BnSq9wUc7Q4XBvLlT13s8d60p6XXockHA+IgXjnD7rYwI1NcWGtWSU
5bWblyMC8GhxOFGIXh5aSd5Kpq7cmLVAN1Q6ocvNiV4u2zQqQN52gLtB0TcLNSv9
fekCtFxvXVvUPmPHRsHDGpf2X5Ek/nA04i0Wn3cHvJjGOSEz0HPs74PXUYnzNHl8
8MPF/r0fdRhyZcqm3GvYuF61TfMNikhOzOkpj/bHMsAMq2Yi5+RMnexfVIE6NGd9
Z71JRwE0knia74hIMIgvK5EWDZVGjVK1raK73yz2JhMPCB2k09/ojfC27m6h8NpQ
piEw3lOJ56DsLJvaXS6HmI+zEUr+SNszN5JXA/AZvrvgzYfYgIEnRJHKwPXu6KT5
qNMKRhIKNkBiReu38lhKJA6vzMRy2k1K43iFHYspdupCQIHksawkNEt+FvWovdq2
bXSvOs6EDpPep5R0vwDgbfIEVVEvESWNwl124qDGk2jvh2TNqAd0eyWkAbbzPCTg
YsOfwl3I+Stnr6Kx6PZbTxlL7EvIuU/qvLQOj7Ft8QFXl23Ib1yORHxiV8Wpos0K
OGXz6bz/JPUT2nYQUuXU4dW3AU4NlxDdudsPX1ueKIIB4FNno+dj4XuNt35IZBhH
IJCVDHsvUJXUQXfcwaIX5yyU49hZBD1T+afyC1e1S8xgm6h7GoVL6CxioCYbv8+E
TtunGcP+gwEG3DZ8qDC6zz9Oi8V67PzhsIpZ3I0H8wxws4LefyXBcqKzIbexSyEA
hjv+OCyRQTeCj2jEF3Gp9lq9+do7WADc48kURFTiU5ClrbBmTT+eiMmC7+qXeX91
raKQHq7REQHVrN+Xys2Sdnx+vzVLXhmMslcU1hB6Cl48MBsUAvubEYEvX647xPZe
pXsIP9ur9sgUkNY+KdM05Ls8CzfQnexoT4xvIbjxKS4cSKoLb86ZNwqGruhCdLOs
7OVgahM4UxYM7FHGpkS/3o2kK/sZ4/YFefGoX3r+aVnt6aDYwERILcqlUcUV2VqX
ncpi42Bm/qWRgwMgKRRw/X8/J4zTYezaAwzjpmDy4vHbpbDkx5ugfL/MtpD7sI2S
t8nUfneES6/dXr6WgbAGcPdsmQw2wdifaREkmot0PQDBm4GDycW/wRi7x2lJedIn
8p94xzlasv6UI6jLP6LeFOa/XZ/DwoFoUGDxp9/gjlrcTrBcezfWv1ZJKjOazIRt
9iUXi/oWSMIeQpub8lSuE1Ra2MSeGk69IXzsnGjJBLIepETMc0A/Q3s6t8WxoafM
KcrfG7ld0s6VarnFgnk+VRtkVzUy+QfpIl7ZM3l9509KEjgQCRzmhGlw0QxIEFIa
qmvUYfbcDsPf5FR9CmHgAkUJoXRxQJ/gPLWV0qPeIBk/4YlfQbNYOkNUdj92keEN
Z3gY1bUBxpFl3m4BLMx6SZQQ9r5ffofoWWSBuG1xraDAUEiPA0/N3Mv7GOr89hF4
+aUefQrS2hgBmCRDEeKkVHzHkFaEtT4Q5bTktXVaIf+zJl8T+ipJ/yijzxfPKzPK
ScNfjjkd1HyShKdq+GTlVLko3AocsZDsYKmVWSzq7aKcYZSNElvcg2WqJ3Mawc4o
QSgQhwflcLYdxyTsI/ndCAH3zkEyTqNQFwN37GjY/Br00Q/tHMWK9OyxCRqf8ogW
3QN67GHQte4Y15QXOb083mgB4WSEk0+QCTThgLEV6GPlwELe3YJohwdta2+0NZ0M
jkC0A9yZxIvmZ5+oa5RT6QhgWrjsAHB38KEX09f8YkWmbtiymg/Y73spKBUFoc1j
rKLJoXimqzdripH4iLDuZPFO9m2IKLK7Gm5S2z/a4AkfzspZ0cEwrQ13vYv8yXax
7oH5w4BojhPcREcQA5f6T077C54ODlywBVvo/vyQlodbHmD/E5TkRxkVDs/9XFwO
8+k1QqMYDa2JTBtAhKrpoeQPCEFtU7NjFwivRoaQss0IiOENoLJzo2s5pzBm6w/8
I/KsUsL2jSet1XVRcBt+IyAUTEfESEYJz3JU/GWMINxEILxL226bi+tzwBX+wlo/
IGThwDBr3mSEJe7ImkhaKZUGvagJ3e/Wi7AOBS6tq9K1/k3mKQHTn1pGv++fZugo
hi6ULW+5l8CTJQo5ou+3ChQmvrAgT1R3BzLBpU47YJI4QtrFp0LaX9wJ1zwvstB8
6HWKeJohxPsINf1MH0LA7Zmm0DoRWqfZRLSdtv1Pg2rTTwJK/xXbI6YXCv3uqZEC
vTaBAIT4MXtylIEdxbW8tucGivdw/ZBeEVEJ/t1Ffh2FySLENbPfgSNOxbLcVtNv
sebdsR/UwghRNg6yifGWHVY8C92dt3rCStarXe2cfpTTpaExIyai4D1ILOtTUKGS
PMntVvbvETqGootm9ORE6BJfh32hDPl4NVJ+d0bzEw6cwwRpU2XCLv04BM6FAYiw
ewY02qdoL0CtcRNwg6vOxYXv6NK+YsU0qLGohPDIdiLPck/IvBk5HEcTd7oqX34A
P0iDP6dCKdteu5PV8Qc6gqL9La2aIvEK3Ao9rSi6lcPDA1pKryn9HFRZ2RIlq6j2
mxdxchT2afnCgr4+aBe+k/AUIRMDwIgTHjZhkTkPl2sCTzCuB7WDiuYoL+05fc5P
C1jlKEQl53wl1T+PNGQrQ8tEsXtuI2pOc1C8okaTdBw6Di5ilVH5bJ8SceTplKJF
utvO+drbzcfY++iVNxwXxT3lUs+UfDdGS4FhIRhD5+GpPjvu9oXHpiM4zgbyuD/h
zyt9t3kRHvGBP23lLpJuTPg/nFm6kAcBEqnfpufJozTjgnx6/BDhKO3jcNXMJLdc
EOluPQTgoPlTssq2OvSb5i8b98BdE/fHrXWffvxCS1XX/ZInYt6CtXAWzpob0OuT
kFBNXLtNqVVuLqv0rFl/vXagr+K+h9wxjhMf/1d78ykTPrPZjttQwViyacuPiEry
oFqfQPgi0oMNvTboBVaFMdg5iSeycHbuVfuqTTGIa+qJE7AAZbG0CrgJs+zW7N7X
t6Ra4aleTvcHp+zB62y8Mn3K6FkW3h1GBaFa+DYHZkd+epKU0+cZ5/vwSWYFsElZ
4fRkEnp2N7m3dsTNKeXN+yoZ18GUYMWDGyTeu7oXx0F34TB6+9pFJ3mROQjirsDE
9zI4OSenmQdlkO8osd+HXri8s6I0EHSWOqUA+YVlUAAFD9JvWVlIMc66iXbgSBkD
NdKG7oaYJMdVzoS0lj+wQB+fYt0fzZJgJquJtPobjSrXA+YOK2MhnMiOHZukcRaF
uMR2ItOebugaa3MLo5IW0bTX6Gou+HziMkjN9s6bVqWj3/Q6hFAFdeqLFLiyxFvm
RDTnlpD5wxxiFltgUDyflyL3oBc6vmJPXXkjdzlE5Eo+QZp1QL772m8PSvvTCgOW
RJVdlKPmH1Dx8AaHp21oOr2vlqnxtj1r6Kbx7pQdeClxejZvXYJxG2slhiqj6ug9
2tY6wtAsRNF4gW/5rY4m6X7fJsvvb7iichCFCNDDtKTCULJ1gNL8xWjoja3Xop4c
3OPGmcsNELpz7YgJvV7doMvsfnLppsjHyvkkUIlEjQziZy4gqdV+jNbk9adHShri
LC8t3/eXObsq97TmmXgMmGptIsLlQeZjoLrZL+bl4JqTkX9OsbDU2NcMteY0C/7/
TL3cq5o54CX1GtnKSlA9hKQJ/KboTjsVEMknq5bgSeeXXKXdmNFD9ijp2RRKtO4q
HLhsHnHMScLC1rRfW7gxuOTgiqqF/zaLmRm0s8SPAOmCrHhJ5U63mu3oQ7Y4JOdJ
nZSo8gNGvWXGKgw1zIlh0IU868N3tIPB07MA2Z/9Cfx9UXPqFkhUW/NCI5OSu1Ne
x3TY6QCJxOvvnRNx2csQG0zjB4i6UKwGzSuSFfoYe3+MOCqbanp4TgCZun5GCTWx
IrlpMVPVpZG4rExB2AJQpQpMyzMUk7ZxlLKStCy7X/8gVIeSn4x85wZSITVQldea
o5S3sqm6msnmjJA9UCBuzM6j/ogxDQwtUAorC5rPl3/IHXTplKtScOc4wPBudaDB
QyNZdBWquY9V/KTKD23ddVKv5lg+13hTCERPlRLNlzjwq8t8uExrYyHg8AvXowDV
HZZTM2daNo/TStzeH9nqbeF2FbUe9TwQZ4iTjOcdkJhFJtRO2oWakdByGGGvadMB
rxbKzLf0twQXoihEZHNrriPuv27MosZOGqahQxc8Sv9TEUj5/oMLxGyqFkCxJdTZ
w4C0ax6LqjNHTmvnoSiq0h7enXg/hr07W/dH+p+zaYNq1KtFDogOM+r6TFs+YVGV
O5hZUwFGtBNB6xYbjeIgJl7+kvLxeI3OC/Ozs0wazoqygjMu/fAVQwMllKOAKkAR
zAIwvCNtuBa4d6YUzc0kUxDhG4Pc9UWRqs4tl+pbNuBQerEGGIli73RGOrA+vEuJ
7V+Do9z2HtlVFPRA6ajfo4wSBdo5sxmn7j/E0SfPlloZwa9OhNK3DMKY7RWlAmtD
OvOJM0f43c+LWBGpx94+e/rJslpVrUhSlhkZ5jwuQBJAWmoY7HcHL3hPSgaBFjgJ
2kKW3NgjrI/sIbIvKk2n0Y8sIujplIVyUwZvw1flrTV94+HEsg+YruCbPiW2ta56
xb1PwOpYgj8+BUbNPNGb6NmoOGrLwcTfp9aW04/QZeuGRpkbO9jwdqvrE6UO+DGt
LV0Eq7v6MEYkR2ausrW2cFeHonLhiktWwLoo1mUT8jSFJ97ez/JlQuhs2/th/3I8
rziCLLKSVhusqh06VgvfmlEU9ibkrZL978FsK7/AAgeO0epuKFjKMIBFSdZwm5eG
UTdJGmaKP7h/OMO94D71Viazj8BQOL6eu8utuJAiQspvqa1oFK5Mp+tPw0EbW1//
qrzIhSm0MUwj8cYJseoZPGjcFwp3spZ5f/8IHBB1ZlSAAAQb3vP2JujZz2L856Rs
LYtFHPJc+cplx8kKiXZ7kDjT10Z7OBxOd993XcaNwAdo05zj6bLB42XVSN7bofvS
El1qsEAQuOTbqjI76PI3P9GUSS7N66/8Hb8MTqNd9TOecUVAcuqbIOBewyp/JRes
rZAVN8Zyg75vRkDC95yB5/geBW4nAoKe6KtCyNFl7OZM20c74D9gdIN7AdDeUYRQ
0W3DdJ9/h9GvxwIpY7Pj9OkbnT66l3XJ557cDW+8emY5xkXWqivwIMjc72U7jvaj
C/Go7Osp61ABdK13MdLuPUwa8/cg9jQzxFNIaeBjJekaDwcbVUu8BIK368Yu3oB/
GvNClvtEu7hoMDkPq9RXbhBknreq7CUxCKMyvovZCBguljs9YI0IgWQKRR8gkSCT
EZsntWk25Zizz4MAbey3uIQXpERWeHC1+uHCpowbPy9beeQANkuvvCYLmo96YAiY
+zOQ5teBv14d8Yqi8tkuQVLoeWJapSWxyaYMmsvhRMP4UXA6RToeHcLwg09KUBBu
S3V6+l1BKQJdyvK7UYa9SRtNbuBbFMK35PKqQ59wrgBJ/38SzIiE5kFrM7U9jJoe
2/MNx7d2t77ZSLZRX2T4VHMnQZNPfQVC4gjDyw3hH66gVRbBUVIAI5pr5+oMJokU
0qp6+fyxu30ebHh9uEE6GT2/TvvHM9Kh0rOYgcEOnIxO4XiXdxSf8TWa3qXysIYa
7ramZrunC5HGZG95QEY9+PnB8UslW3gejAa+lMelJMvbkKdOMt3Lj/blmUYr69AS
WBQ7nhNW0sqxk/dakdq+bX+1Jpvsfx5yir9V9/Cg2mVWmiQlnDxIDNq9idRLYKnZ
L8kAYFewFQE3daXEMca1+1eiKILuzlIfbCzZhoyTf6A8ugrB5ZxhxFcbp4vrYOyD
efhb+9r26eCbkHLiquNolCZViQj6Vq8U444BWAD7TwJIHFZNNVE5RsuBkeggwKFX
tGJH2uQWJgJakBtZfVnyDaemG78RduX1zfFQrvyFzbOgmTFJnecz4VNsA87nOXfk
Bo7xG/MJXItT2iN3QbsAIq4p5w72lAsgtZ7CtLysLZZh/fEIlCY65vaHQUv4YsqL
IbmCuuMiYgAZXb0Di9CWuzw1w8tQ30hIqHMeRdip6ZAQkIO6C6A5wgm4gDA82FYl
SDuJORIOX3jS9UhzVrrJayUGi7g5mhAiFE5Rvs589mXBhlC04iVUeAEBW4dCmo46
OsolWYJxyYWJwqtYwbNJIllIuaBUFwJsxeWTgOXHpU1slWxImaJ3U0nKzftNuFun
Vf5P2p0BWMy++q5AfeHqozsKGvFn6bNk5+LTdKMgmPFWjdgWhB0fhYuZ5QxfNTYD
Vn3UIm+PE8/5YQQLleEl1rZPuhpbZV/v1cobDQtwGngyrL1RPXeFstqM0QEnwAqY
shPr/Cite/qU+Go7NbKpKhPdtxq/qAqZi8B5FXQoo/YBnhOP5XMbqlAWu4m+4712
95NBNx2bZW9+YF6d77fanG7VDuzSxUmCEzq2Pa0COviUFY3Xkns2IgZF+eQcfljW
rK+YfANbH+LpJtEYwrzE1Ca2Hr0d2k5Tfdmx5AJLqd6Tc9wK7UPW23E9rAtGj6OY
b22dlS9HuHSRBgdil5pW0k+wgQU3IzBh+PjbUhSpTfiOpEvk4GtZlhJtfjVYotLi
yCWFAO7vaCczQmMqj7pliOtOQvnDP4VIdj2CNw1+Ef5Bin0MZqvShEl9DVfX2Lkq
izaQiBp+uGlIRPqoOm+S2i4Jl3lTVnBPq+ZRFZd9dRPTPbTtWJSTW0CD3k6MCz+s
zqibu1OpU/BLHyjJHSUDiNSakccml4XE1ig6fuYLdamWYDxahtwQ95an8mkdwG+M
lCsO4I0dbnSv8rgNzOfycgehwrDOonN8gsA0nUDmdPT054VbX18+Ojs+sNI5Wcyn
Fedy6CGmkjCoQTkneNP/qAVvqMbEVCcXehlp9wYtbuKMpD+PrtlU5gLJ5Mpebfch
6OL5vXJNAZHWRGlc7ftuOmogGC1BaVh4WTABvvvWdPjdl7d7XGVVdhkHtZ7k24CP
xSYMv7ivUbmg+Qi9dA3Sc07G23KZ78Yi5KOoa9ZwHDJoYBm56Ac/6LQvJCbusiWM
xNdD2CANu31/K1NIcxbj7ru3vRBojiQsOGzU+SId81/c3iZBKdiPsAkBbOiwMXpH
P3Uv1+VKQ7Kv8ufcYCm2C2ocZlXI3IZXY5XSsOTeJ06v/4qclx6HqwkPmyKxHVi/
NQCGr1s2gIJ/gkoNqORfr6rTQyE4390+ouvkoMceyWNvmLeF+c6Bj1MfST4PoFzC
Zxn7LO6GO5hUEHAQqCE87nlLevmQltbWLKkz1cILj9gj28ttEtDT82li7Ih5c2ub
NsN6JRC/sjaO7tGy2seDpy/OxoOX2KypgMO0VyPrtzrwMIcy2aSzJd6L5yu5B9Ut
q7Wm6QpG9lIqVjx2kPyHOkbmms2hgB4s3t5rKvwpxY9oXlu7b02jM+zVyzpUgRI8
ygeHzToCghIq5qg4dzGzI9pF8frdINzQ+f2DtPHNl1o/xJtsT6VrTwupMu0jre68
52BALORtueMlWOGhPNFiFgBS/Ffbcan+5fnnDDDez6shHLwhk5RfRlL4ljnxeStA
7Eic79xJazFEteQKYWKIoQu6kp30JDcYUnGwGj2bopC3dVl+ljZDwDyp3OHnrqzI
kF9qf9hsM/sZEmlsIYOzpbmGNONWb2+PkE5PaA+K5Lt5m9B5xEcTOjE1e1DJS0ep
fCqznXb8xzhRxEa2RnYNvZYbO2T0Ectn1qgwpXUgDyKJAFedMvShaQOjkLq82k+r
kIfjB5N3bynMdoiOaVizgSQ6TxeJ1ygLol5Yuw+FFz2RrQSLy8GCnkNHiOpc0igA
h5SXtVNk4ffvEn8VnFQEbtigwVDu2MbV7sff8qaSWJ/64WVc46jYjZ7ZMNkJ8Pep
agh3K0/eAQZ5MhzQM73LjSgF2emBPE/PQgqczgg9IkboCAolUIYVyS5T/ebEMw9f
3ITO/Y7SxoTeXGBCumkZbjblN4Oy01+L4lC+Yw2g43l6OFW5orkG4fEqZZtkfnHP
dYWq5G5bA2qO/YRdHE9CnVRMSJIL0m0v5S5mteyFA4Z2ZTvq/ltEBykgZJVB4nzO
FH5w6C2Wgl+Mxnm8OK3VETUMA33gX7OZ3iIoyi/Nyuvhhbv9Pq89id5kJpX3K1fm
uVIwFDUl7lmaPkOhn+SzhhEA+/f8TGT7+5hTxxfAlwM7k8k6oLsPxmkwlyoauDMu
bk+duC9pD4s9hPFn9YjTnXLf6ZalNUcnAcg1vraCJp4psYRPlpccXRVnZHR1X+A9
Y3gg24ugizaGQ6vWOE8joh1WFfiIG64xTq/vsIKNA3po0V9arbsFKu6m/JEvGPQf
r3X89JnstWTItyhqgdRD3kpWzQkKpubUNfxaCDJ32Cr+rkIcwZu3ZiXXIdwsLBEe
5maBcmPEOQyxPNxc5on2Z+USR6fU2oE691DlC/wYnPxfVC4+qryyZrBChEABaREW
UmPImPeb/kS/eRxEQJVvjQHCIDzgYxEDxxM2ijuJxydtKbruzsQUOlKozf0b0wWF
2uw4vpfBFprXE0lzZky13SosC6+M6i2cfdx4qrpzAHxJ0Dr8sqa6/dJ3PE0iI0KL
QRzKGFlEiMP86NYBPlclVmOQvVJyrARE+xov4/QvYMaWC4Ozi2cvGQvSV/GZu8TH
/x4/a0COwXAApqcIcetoxO9DHBFdZiIkS4iHL3EODRnRYhEgF+8ZLcjeH9vJf6kl
viyBGpRGdG4osvzCFcSfWc7PeAny/Eij/yH5nwMfPayWzclxS/tmmDo4sAF/QXhT
+nDsNJPQ+OfgZnXd5hxDC7dJEPlZaX4vfkztM2AQqdmVugmzRodpLdLm2Sy5lqcO
/Ft+VIbvxrFakNz2Tx/mUUGf6o5edJaVW6IwV1rs9A27Sqtr0AeqBP/2Af1GM9N/
S8WevYiauMGozfZY6bOBZ09zadCAqxu3jKSK86XphQ6uanE2sPFfi6ltIkmZH8RI
xx2Jc+WAa1jX2jMvG0Cg2Ax2S/DhvPfJLLCBR995XDmxXzQ+MJMWSO0pBhFvKI+9
TLdvOFSP413QU0DWhku3oOxGu8ror0NCgH13Bgp+Al35z3v6GAfFNPWzaeuKcdst
64lMZlv5Vcha2+tKVKUfQlRHgnDCvGCo7N7aoYdN3Oc/al0XPZ27Zf/GdV/CHzrc
Z3eVcsmavKkOn+/FKuSHqpA7T20K9INsudtkBWFahNLpiCxUGzDzY+iasKiZ4LGp
hPbNIyb/461RxSU3j5oIx97n/y6ryOUmLxca4pVVLCEiwIVAw2bjCV2yUDqf/drE
1otvQr7Drm7OoWYRGpzxSuGD7I6XTtSVBUqQa27THN0oq4ehufwwH3zRIIANxalc
37dyczs/GVZR9oYUknvzF9Q+Nm8bG/5Az3EN/8+zOhBwgtSTx2wF7bIY422PNCcM
3uqo22CNxzcJbI8j1W7gPSxo2Fhk7DKOXWJw9Ns/ETCYPuZkjvWRzmcnxb7JuEI5
VqnzbQyE79l5hLYSJqBbp9wlYobwsJfMsS6PUMEeg5IWE3uBgTmZXFA9AV2OOJ6S
e3XcbzaZrKeqc1AEa3VM8lR892O9Y4M3jwJWJw7jqRpTpR5VBxasQdb3MabmQCce
ITc31NhlSCXwLd7kFo9BiIT8pOqIg/ji23B3vZqT/iyselyFwFPRFSEZL9Yzbs2H
2Qd5yJmvyeXI/XYYAmmMQpHRFWl2khDsOmM8vxJoh8K1iz5XrPVKnuyhOHam0qKz
FS91H/dazW0G9JVNCvU6K6BlqZesUoiGlZ0/0y5yFbWxdMsZo/pSbWtZp0HOgyJV
+xxbQ6zbE9DM/3nt92fSAEvMwvqun91+XYChmnJwgabJ+M+lxmeyB98RI67pDLGl
wsGWfTRyp8iBnJc2OR8zNKU75dlSHGBoRv/Yx67OSXZhs+fVXUUpJtv4iMMJ2t6T
IOkOOTvxOWK5MWAZcJMqGNLzYYO3zq9LRLIaN3ef5JHOnUVYCTwqR2SQo6dVtDFR
+kicheH54qyMZ981L71GXkuqLvSgqOp82smePeqLZoSIrYh9FuOubbzZvPv4s6qV
PuKxQLdVS1TdVJfwuh7nJO8ZqFnFg+CI/9tOYTNq9p96GTxogHg0z2dAOeoDz82/
sbifna0UA7K0ZZIme5ZAesfbSQhnfof56oLTiUYCXEomo5y5RLUlt2ovx51aH71A
U/Z9dFlZF3nSbSTZVVweAzlxCvVGtoja3jXkYHKsP5vM6Cdx6mmF4jIjmiJY1mOz
gLYCYznaguFlu/6eHFPL2smgaUFA2YldCC221WlEVsImt94Smp0o/r3o2KL41q1K
Wpp7O+L0fTVplB5VD9o4DYTv7y4FrA+eAMnCcGQu+JI4FQW/94e1+qYZcqnPHbUB
XVhlad71qZDBc9bKbK28iCpFiXato+Ttj+ZD2WAdvgpIyR5FPSmkDs8lEFPU8xkg
dgVGqCf/BWHlrzQi6jXfR+FXKfknEoXVn/H1S/ASztwrbfDYpsrb0kc6tUhqjPny
ZvH0aNUolkNoTSls+aRNsMak7em7gnUsugjBUO7YGgtWHTsrRobvVWoCPKPKfNxv
/1a/1r1g1wYy8tvTtKUYn3bnVFwI1ZFLjPY5vXS5vwyjY+fs3o1y1DnU0W99UcSb
978YU6C67w0sSIud5el/rrjkYQ82nXDa71leAXruIkrBI9xFEI9n7Kc/sqYkjKx2
LIYp/pA9NydA+zcK8gA3QEeTkA1S+q3PO1ZTIj5aJzvi89f+m58a53+dQo8X55Iv
atvJAXmFtiQRMaUrSQLDLmSfuLZYwfw7qXmzIZHb73VtMhrxL9Uula7myDUdWzmv
GPhGxXq+Vllvau7Mwri/gQsMk4mYAM2/NHpDDeCw+GF3DJMmYhqfsTXL4YODspMX
tsNCbpSffSrLaqDfj6yJp4oD8fAWBUrMiy7db9qUR+b8QSS8T0WxuN7Y75ErTQxc
e842pSPszkdx5neWuBCh4U/AdmoUH+ZAbadYpkk7uiP6qS1WbwTlNHoDTXiq9VpH
D4jMitC5mggAiWiVd7zH6psQubF+RH5rlMXvZADBZm2G63O2kbEH0jN0paG7kp4p
pLM2WV0OLEnfCsHVZDZWPhzz4G8gz11026NHUfEDuB0jOCeHV3Ka72avB1Efgn/o
9jy7J/hPo8eYwm1oQTNDI9KekSHpFYpyvd5NSuCIiINODhpONafMN9+89A4OSJhl
pXusYTacFY0wv54eoFeFOpm8bzoap+l8x2AA3kad0+5n2jS+G2cVqbsHVCvTxroK
3rNptxeYCbmobx3n13uoRdu4I2v9r2hMfHhzAfuyxNl3tsC7ZXsXvJ8OsnptIo04
DUPRRCp1vBJK0rQzfpBQJHRvezBxVDjXx62+16qUjIgjjtpC6RM+47dsGfZs5mXi
i9/BDcLU0WIecUk2b0CNgG0r7tVJ3LfyEFQPz1+1yy7Pws21jss88LlUWBq5qkhq
fiKqwDFTll0EYs3Mt/7Zdfo9hd6jsOYLxwxNYyPYnpf2aXkoX1liAmNNka1BWUFZ
gI+v79uWMrQ96ndIBZ19dygd1KYMT+9KKX/zRFVbJxkOZ8S08/j4mdyWXXp4vn6Z
HhvBhrzXYOSQyNJNcv08cz2mGbR5UzhiL6ihb8FYcRVpph768bc/MZl7tycxlw5n
/fLxIWrCLJnMejSQIyg9SZXUuU9HbTZFnwojCZFIwsfVlpIIdmNg882WHozRVuxX
TMc2MWN8C8D34RJoJRLhgKiznx+AJZ+1RGQ7Ke3uHsETm2hVEX3RffSrJ1O9/Mz8
WXe2Q5RC7tyB0LUdrhselLLiSBa9W9zMFPJBjfbgeARY2Rm8dDlhQ8/bTKrIG/tQ
ATy0IDkIm6pvPQw8+Xxyu2hZqt+Q/H8aQ24hsjwBTm2eUL9F2jJ4ep3zCoUo59Xl
XGkYp27MFZmiQe71U8177/khRmvmvjYsC1mzzu9lxhPZRLBzUlLAYKz/cJu7ZNjH
db4I+2Mi/mBv7P2m2SZynKPLBlIdoS9nDqGAxh4Nx+Hj5cCzvC/4mWlWaBWuuA9S
3KqWWBOzyS8+euWIOJ/nIgEfpObMsNLmtDZgoZQy+1gypJb1HwJRd0WFtsnBr9m+
3YGfh1MrnrO6mYx4gGZr9TGCY86zxVdW+p9kFVgj1nprFi9lJ5WGrSmIDuzk58Eq
7hBVlzCAOSsdO6XHhw0TcmMB/YkonUcpLPAumuh8UIESAZN7X/C1bLTKfjcLevC1
eCgbAmAjh5wiLlJAN98M+167MxSrdqRssdFUIkcZ+Y0KFNt2Md01Clt5lx6NZze5
BID4WwsiOdKrhHia83cRe0aqm6KB9v295h51NQBXqpuvlgNdlWPfRYSStFVnK1Yr
Tq16N5+PwvNB0hqZ9EoZXcWbweM9tmND+v2maR7S3aSzEMZZ+7csrUorQb5jF9wd
7aFz6X7z3KWgV5sy8WKHCV3zD5wSVjUJaB8mlm1ALmR3yKEIj5TLYLOqm3F7WJb9
Ld3h9cBjsnuCjWujb6wPwDZw56dmx2JWfDw6u788+HFj21NAuI0GlZUwz5hI3lNl
QIuVLtSshw55mgVQvtrcu4ZyzwCgMQjJ3TbOYhIP1K4Lte1Q+k8d9TTD0g76iaSQ
y/CeYY8ekBld92nHLxvNR1YmS98b9xaIFBCQG4boqK2vgJ5vPjk+W1pyH2Xzbo7p
O9Xyg3+xmqxQHIh8KEZXwcT7npzSvIpxX2NeUOU/sg5lYIKRyl4BlRUQdCD+qQty
Ow0tpKBjspSDsaUwEyavYhz7M3NggTrKOxuNxbKIUzhtKx/rqgKCYi0pKa5F5H/U
DLF27wHcrcFN7okb0WGdo6FdxkzxBt2D+IdUXr7gNjuZzjNyGEm2rCjaYs0ZsFzD
2oopR1GbeFY/l6+Hm0KOr6vBKdjF1FHHZPIghu0H+ihIdZdWbDSjamJqkaklHaaI
tfdVylS7pRmKaDNfNOKMRLoDsA5YiPXg6X6i20I1PW++SzlRBUDyHkRnQJMLtTu3
TQHlDIpwN98t0qkfPRJgxgx1dRopMp/DKv/sueyUlGOf+aJWJqHlSCr6Td9oXZEX
4w0AsaubIjmYkQ4c6rkbvHtmz0ZqCYLrXV7ZyRKRlq4f5PSs3H8+KxcSPBr6J+nI
XrklxeUrEL+zHHU2QEHR4TMv3VGiu0tl/zXKQorwMzmbG/D8wtO/kNGSpN9naW40
Fgu9FMJekjj3RlPGihaxsO/mL2XA0aZBdUDM6ivafYDE5zjo+mT7AnZcmNUQwNSL
QNyyT/vkYI/o/zXiXESHQB01xSJLLRflfOg9Lj6Zzt8Filt/VbxO+6o/y9tIdCi5
2njY97LHxWS2C+wTot0Z/vNUH6KiMMMTJXmsAiDs2Ia4YJ1W3MQ3A9SgfCagejn5
j8ADJsxMOwyVrFPzjKZGXyh8ghgLD7C3BDBua0UEg49C3Pg1JRENjhlSdWOksd0r
Ra1TRcZr33fuN+h0RufYBFcg8u5l6c+2+JAf64W8P30OMteKnqjm4Qj9aKewqaeI
RKw2/vMqb94bM2i5V0+gSzPCgWdhIDUTxxPZlHbPzvPjixYGMOpRlyqOXTTWO+tp
4DkdZtxuEU4ggD2JsyCSp/GhZ11YjXn1rxlepyEvl2L7PUX6kVGdafFqt2a0c2dF
07y0/pQW6BnXxrjsPE+bhIxo2ii4ry7hu0yrPtlsfQfgnkVkOozfC4mY+NR3IlTS
UWSxJjMNVC7jdZ4k1UIUOKQxHkzdbsOkFkEragxZPewvG1b4Nkj2BJnDFKyh6zVJ
O4zVTaHJs34sl7jyo+NNMGdGP+TJCYoI3xG+BkI4VzC+Z7lJP4kdfMMAfHs7BcW5
3WgE/ChImbsZUHD5Ag0gd6ipOfolULVwEDhMj5MMCCFNEnXpwme+iCpJaDy75vC4
bqkVioFUPEkDevqxhKY5MFnK9huKBZvLnAexwVpPjqVNYDUV2b1HTyVv9zG1eHmW
lmp1jsH5Lg7VmERU/H2laey7AGILPPmy62sqW5nWXq4HUGSL9cIjIWM4fF8Ept1A
DqUt/5iNiPvTOB8XbvoRhqvR//Cje9vqTjVVqgF06PULkcvXSebWM6g5ODBeVh4k
p5LtJL2QYLKMa+xu0z1bfDuAhSvPGi9q3lMfynPFi+yQvypypVfS6p0beZ8m3d8o
lGZhtbqmESg+spiT8XkETKhLFaUgccarHOkSmAXjglAdthI3PXf80DNZwJLaXa/o
taVDEqaqPPj/XKNUjg+YzLzFmHE4sjXYRcE0MfNm7I7qoKgeTMa9BsKo0tH7oIYf
485zCP7bYgk9kXU53YD+MCDKgtx9746s1Imx4M9B8q6F8Waa0BrcidJ2Mqfudy/B
4BiJI2ZiZsMWl9wGyoL+S24K856KgC7wDmXWr0chWGteu0Hc8HfFp5m8sZ2s6x5Q
A9sevfotLXWYSJ/+UU9phr/Xbr+dfcUHWTRLDLMX0fMG68B2vK2U7r4R4DqocgN8
cFh86J0F07U22Fy/JJLr5mjihp9nU2G0dovH2PjxmLCMeO0HJBXh0JzsT49ipHJV
L5sOqAAr7fzC5PVWfctRpoAEDM1LkjO1CW0j40W0x67Bvp9Nwn6gMEMl05SRqvED
fn2ksdQcLD2gcixa+aCz8unOJ2CU2k9Gs6bMYvg/zwodq9AFOXbCUzZbKVQHNPsV
qtCQ57prYjaK6ubkp7QtMaRmgFUuDb8D7nt9ovsDaG+IR5Eyi4grQFD5jKbdgO2+
2d5E+Fqbw36cAt/aZMiywlTuhIM1D4l7OkhtKdl1tl8wTugKLjQ6yNAnQSsoPF9X
y8yDj8iSbwUg6wLXwY4W7bBkGuwtAkpLyn5WeMQMSBh1k+fBp4qSm+cbIdLkkBTy
K0xcySrgvBT30P0lWvgDDNIyQS4f3NOtNjsJiWYv3ADUW9tINP8IidWW17T4nlcg
i+sD0dceRfPuH8GYohh/2CtZ3a8vId3rV5XC0tIc19tDEz5EbpIa+2W/xIWzB8um
K7gQSz6dEPc763SbJ+0GpwPVglC/x+UUmXZtChGmIk+lN+PIgqs33Pzc/SxYYz9O
Ap0wBNw6cQmdV/OeYQLKdtU7RBKN/eqSD6h6fn/OCizI0zjp+kCUd4ZbL+nUUxFQ
dFVgwNbRCRgs0l7SUQtwVJT6lNWcncQ+tWmcoxW+E9hZKfxpw9OJVfM8KoqBGFU5
K/DmFUio1y3ToOvauqZBt1EEd0RLQaliu1BXviBFprtwQDEOtG3E0CU8+iMZAXo1
HsOYBmrsdG5D06Z8FXu7bbrCdJ8BEwmWx8MtnSOV6nB2kJACwC9KuEhR0d1urWNg
zpybl0+mu7wdKXzp0n2ev16tSVJxNdS4wtGfBvYLG1pU1lDyQrJFSYutujT8Cxsc
p2gzM4Zz7pCqofmQQYS5U0qAW4vknkbHkijDWiq5Q3yWv99ook1df1MERbaVK6yv
1gOkoFksS35aGm0npe8xpYMmdhNLW2HMF3xgQls6ujbFlgu5QSPS4lVWCbk/ZP2V
EuL8y6CyA3CuvT5GfADHS+XD35u9Gew/czf1TBnRcGxl2Qer99fsF+GH5J24tcF5
8lAlXdANuBb9QztNBXXxjqwSqcGWwCihst9uyz3HYdJd2Z5+pWJRlPjKD7alopdb
D6ibJSTCzdDuTwz8sIQCQptJaMyjQgf4g97QluRMgXYUbLz4ZApp+mh0seHTUETJ
drSI1KvMiyyPA4q7EHzwK2Wiin5EQxJ89qQvkRXM8u6r9HujFNPIc3EjLmppVVzi
pRvmSoRGVJ23uZwpIfBtDvsDdS0lH3/yLV/QGJfPmfMuNWRzgLHSo9Vs+cRKAPbR
BM57Tellzaa41NIKo9kgqDN+j/h7VcQD2uVxPxjeVosgwXjfGd4ftHHyFUqMWqcH
hRXnozIZcezhpE+qCOl6ivcTDijNEbubmAAx87yKmKG+A70avtgVkr3NOlm1Rao6
hARZWhzUu+iEtYdJQ0YbNohkPAkBZREZmbq1A3J6Ib7jy+tJuEmX7X1iGQgMVzKI
nBWB0+cSdGO4BR0aCYDWcuPM9s+k0RPkeRaVhrSrPDj2P/M5heP6NkOUfD91pfFq
1lYFqlS3kB0NU+1CBu+QNNaRhiPlfJnSMIzGoaRf7dQbI/gbRbIvCVlvEMm4eMS9
xIbwKvtKwPw32uwUiZJzkRzajuYrgaeCIeslyEP6OXzQ3+tgPEevbe+uPmwnr+bA
P4h88ghAbB6UnZNwVHCATUpJurS5z68l5pkS+KJg71LlFnwtVM+NURmDs1AcHJ6Z
GpOtzHGcVdy4l2T2xvCVLDQ6J+fIyEJdrWhh98wCqzbnHn8auGIKWioLejMbPluH
19ggKeEz5EoHSEAK2y1XXoh8SgIwNyze52ZSauRtzrmxdhf3SAFaWM9i3cAP98+U
+5WI48rUMEJy3YXyqZSNtJL5uuQaXNVnX3C0hmu1KcDgEDD0Z3XuhqR+1tf9K/GF
MFEZHMO8qjmAeXxp/21eC/h6C2sLcjJxbjlfYVVB328gFP08eblnvy1bAroqDGPM
1PQRS51Tk4SlEFcctgPHb34EhsMWgpqUGGuoPnwOfvp+rKEYBeadBhiTZfwAyhoz
IuXqYCD0HTjAD6yS+U8lZmJkeCyF9bZrCK+z2w8CQcA2MoghznWX3+oHL5BIy95m
ROshRvr3Cn+d+QMXXyPbRCv5r8pzd4oI/vuvNl3t4I24dH7yrO9WFDl+rD/h6BQ7
v2N4hN/Lrx2pELO8r4aN9dXD4YEqFvi8OyvwwOgtHK+fp9C0gzzcyu99Wa0zrCbA
asVqU+/R3CLQOw1F+fTSKt1tdEW1dMdVOObtmOx4ZAbUejTX1xoAmD1GXuVFuS/c
U0zaV+w3whBfmvWj1YD4r2m4X8A8n5WcjYTUDCtRLXPHoTK0fHWenp75Xlxb9CHc
kYPXZGyJoAQ/Me7gKGkHmkydLn/HYXwW7OGnmmPeXDCuGFExNNacNLn3iHmThfQw
f1aY03L1uwDLPU2GZNfy523O4qbj+k3JmeRosfMPJdfdYMxfgzyuFCgHimiuHewb
9KzDzH1ZiSdmOsiN2nR/JzMVlSpFm5S3e6zmPoeVyI0ri+ya60wxJ6chYV1OH7sb
Utb0UMxVhtehyLhvRfnVIYnLPfp1cKoHfb6AGyjKsrk7OuvRxo7VQAIXvFwZMPzq
QZyaNBn5BTLI7g6CdYufzXHuNmVsypxkbQlvZUOSuXr2tVx5gSFluWgDYn7i8X2O
mf1H51zPrCJart/4MvI7BfhjSbKdgX0Km0ZPYnBsAfWXjLFav4Ek7kBwsPKbJ+Lt
exAyXDZYQ83mOyLqPnAomO5UxJsd54aF64OYzxEsjUo0SKF2jd6elG7cXE9XMa1+
LG8RIFfesCXgyfIk30XhgDUtlIq3/rtLEHvgNQOqZTIBNS7uaNlihq8qC5eF1aOJ
t3jdlXNaHE/ACWaiEx3WO/zCyiS1KVjbPHIESFpxrRlM9wZpqRds5yBj7HLjtpAz
IxZGC7prmeIVL1zVRe16MRKk+X/+k6PYzADN38HKllu9SDkIqDB6UHVqBKXP5uX5
UKULKcuPttchkYIhzYoV8AE2xMFdnDW+4AGHPJTuEmu8OboNo4zpg/zLVM58Kuw6
fLlM//D9XM/FFxzGe4fFopSqrMLqXTmfDlGXpTqrb4ZlNX81rtVJYtpDFQOcfnwV
32hXG+jty6ioO/Bj7VCQej+ihmVurHXXpQ1grTpgMgvBFw5baPjHRN7wyPALoUko
gjmBsanieoOEMvpFIbAgjF6Ev9vJ+Jh0P5QQLz+colQha7jDyS1paB0Jmw8WfB8z
w6j71neg2qu7CI7+xLPZJxGcb6eN29q4UWfL8oeAGoxuZ6UXYEaqIGkhW1tTObEi
NotU6DkLNF2wmJFH+JdejEkVXyAymV53ruBM7oC8Ys9M4adi/n5iRBmre9i+D60s
04sKrHakuTgfS7B2DygC8wzdG7fqFI6mUCFa9x5USbY81rRqxo0Q+NDE0Wn9l6l2
zTVciinSj6lkLZnMOufHIaJLSAQov+6NF07WO6KGsCITBTf0EfM8JxA0Hv62Z4tZ
YQgk/KQ2XrQYRvPH429+cL87s44hqYOMKtRfhk+vtY8wmZIvYvTcAxjN4xcBNb5M
l1EUQ8JNRv9E/W24XuGOJJBCjRB/hArcobgsdiDnJ1DLN4nsKw5oURd+5ThEkAfm
48/s+C2gcfgvfRLLgYNeI5/Xx8NjA9yBOvJ/saEUzMpkk/XfwG0A7yaKJQoN0q/U
YoswSB/B3+6NT8HvHLQc8s3pWW+85Fr5aGwfiiwxDI1eqPyC3V0dL5o4OWzqOtVT
v9pYwsTZsHG6V33wTPNUbgIZEqvoOMB5BO/06IkILK2Oj6mo7qkI9jBIJaYlDGjf
BfBK6EZyoTg5tWhw6Z5AhuaNiuYWfEbYtsUe0lZmCkWsGPuphFGiF8+/nOZBgKoo
DwWVmGYJ00e/VMgfxU10FViCZaqLwitWkxGDCxJxF4d28WUD8ZBxSQ/CIy0/0/6A
zC0+U75Ygpcjyfze0qNw4xiW4ugXtqjQLQ6sg11WIUGxHv0K6Wpnp06tt+4mhh0m
DbE+URDDX4ubdhOZjSBtLBnLHVNo0BSze9Yh5aWd5VLp80T9F5+3PVPd/w4ESxsD
9XxSZhZaVx7r7uiE7gN/VvbTXYqZQMVmE0HqyrbFaJ3VCZ9YEXiM/afKp9rOF0Yz
`protect END_PROTECTED
