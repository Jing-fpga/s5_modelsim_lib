`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sBsKCT1xvhjaA2wAOh8IKO0QSZjVLf/G7yk5qp3YU5SrJ77sTLPd1+5FmjgwKBme
hD9mC2xGHa0HfCK9QKKxH1T4PdMa8nwYrVVv+Z6+LDAhViNqev9GqEdno22Nam+H
8DW4HGR8KTEQhItWFN4neLzg2q6aqXaPhH9HrkiGwrSgUTynfmn/CWGWLS3bzW6Y
o+d5q1vYm4P6JQu7eQwRwgfl92m0oihs2tKAbyCiUpi5cExYJsS5TuAazjJV+pjW
EwecrxU9Af+c8HJyklxT3a+pyhC1IodlN+KfB5QaNzQTLjcP/yP+ham3QZnNrmho
31zX5ddW4nX0ED39dTtnhaEhwa0ndTR9KzZcC61TMQRCazkDDLsm8IR9CdkVNi92
Z0mFF30etNvlHqgnjdV8w3tKN+b2Wu0no3wy+Cfq61R8KkrM695gL082Zg8Y85Ur
/xhoPkwjVoPAZgEfddrjxrolKyHlDmIkKuutPEbQUG4GjUGo0UCIpT4Mzs0sJT6g
xG/gpvRKb/Dr15Cm0pTbj4Hh3ZmYyEBq7zA/qnm5dqAlOxE1xET4uSCg5U1KRCh8
42DKuG1hYtA2paePHYH8BJogKbPWMFDAz6eLh64QlovwoPGs5QWGqO/ZfNauHLfO
EO70p5HAZFf0Z5yL05JomA==
`protect END_PROTECTED
