`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YiAlxDDGtLHH416reQXU+YDDqgRHlw6Mb1mSFhx2Jjad/p4SjdtQVpfMvDykxQKN
2t3YlYGqVjX068o86ixureDnICidruRdwrjMRv80KQ6RrrEgIw4rDKj+CneoVh5I
C0PLk9Jb+dl980g+31qqf6A1Wi2ee6CdNCDIS+EnNRtSuGvVYq3h6Q2G6kpBZlbO
PGGzsTt9YWMztl6o9ZsPE7dZGKkQKcnwIOuu2I8v2WEgv9rqwZxal3YyXqHf0Omr
OiIPyFOqcSGvNolTmKcKbCAzdBY1BlJzwZjufN5N1bXthjvKftgwg1zD46qn0RZo
emywZCTDvcpCAlQhBQUBiyxxk1+nmR4Z7+QL/A7NZZgQqvvsdjq0AiZccDoDBeyD
ccl/VPgx1KcatukskCIn+2SOeNFIsk67akKA7bEg2bftifquQKiX0wdH2CXI7ocQ
vVwUf0Sj5xIxzD03zJTYXoUauXO0UTUFkUmeOLwo/jJZ/R2lAsSIqUmi0W1QCGHX
9MJiD2svbdw7sQgH2ccVLywQx1TbHL5B0LJfvCF3oYBfWb61Yz5+liU3AYF9Vdf2
ABu7nfn3ZSZHOllczbhBXG/wHMPXuy9xfXtM+yCRZGR76n0w9lUTm7zaTwVhoWQl
IUwaH1xSD+oQtBorXvtGOoZiGDPTiTcidjeB5M1uIPFC8yyP30miX44MF1UEEESf
Jk4IAT5WyW/wDFCFmpTKVrc+m0P2KFn1wXMUjjH5WuFiVcKsGNXuW6ULMCPjn4gu
nlC+mbGdaBv6pjjpqlmOUOUD+a08vN0t+9fRCWbLVAl8oC17rmz2LV+vRazMFNY2
5f8OneExsdfVRHLQVMSstVBtGnxT+HxvjcRUFD90EFGjBv1GoHp5tjQ/zzBOopsN
SbIqEztz4GDMu5u4Z67JoA==
`protect END_PROTECTED
