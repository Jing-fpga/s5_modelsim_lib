`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sfy0sq0CXoS8qdXdLyYaCDxjgg3L0vnS5jw2W4rXrrC+8akWTXewj+FETFTDSgPR
m33pfx9ZpsvSE6or5Qq6eztrKOuKH2wrpr7xsbCKpAVwvT2clIp3FgE80pXcE7aj
gBcsmrcPk18Z8kLoUo2xYjmPTY4E6JOjgkptQqB0LdIsKtZ+7aDTwbCzGONlGZaZ
NM5xDd/exXkwHY3yx+g2K86a9SmQxfuCoNvAbAfTf/tSe9K2Pt7ltY6pJXRaxPhc
KKYdOxmBv/dZnrkoKIaa5Ewwzg/0fF5B7weYMHLqgLb6z3ECrlKPwOfBnH94/dRw
aoYyLv0MYBE7Vi/KF4WbRL22NUPiNIl3phaI8Gi7hBK8Xsbbl8TUT8/vK6WAP05j
+TZ6kCGjFLEPzIrugueMMkz1Ksqch0VQTr3qVLAHyLGLYuegMCGjpFPHysXoiac2
3H8ijcX5wi/X2vefGAfvUE9onaV4OC975yt5AXo7pDur872Vx7ce5RANszPubtB+
ZA1h4z2VrBRrJzlkQ/jc861acT9rLmuT9N+JCqQGdveuUc79cyjoQ3zxKC6Hmrun
WzuS2ZQWqNA4E7V5JAmAvFdkeXEEUnrdIm+Su4pkftE=
`protect END_PROTECTED
