`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bj2JNP8U8VTrz5KRl5WenC+SxHUZ+nmBvptd1tI8xMTxQaOm/XW64yo/0WC6VvcT
NLUUqVK5cuakg9n7mAT4I7IUUUqWf4OiICzRLE1xNByx6Z/e8rNITux2ZeXN4b4y
DXLMQlk4V+deXI4gkfdhCRJwj2LWUF6Ofmq9ExQWs9SiDbHpKBmiVRfKPuURGsEQ
lWAwO0uswOyl0wnEBFeC/RruPyZsdusjYC/48MqgxEreLF8Kw50p2+WbfeXu53c2
cUuBbZATV2psPZDuSUa7lgDqfCAVwhnTXE+X+X6DtB0hSCJqVgF5nV9tJ42dG6PL
zAFAfXq584FKc3bygSE3PJmy4Vgcp6wz4VERZHU+o4TtSFm7z4Y//0AuTGusMgOZ
jEyBAS7kSUUkESTfXokqCmlRJSMgx1qQIyeB4ecOvrPiJlYCKBTGG/dbuzHDDW+T
fE9TgToupdfYYzpdEBjJslbN9wt5SoHdtgXNuYd6XKW1g7oAvEhyvaXQynvWYLJI
lO3E3+Gais6ag+pUaNYvZn3eXbmdIFnC2rzh+vpnRqp+EVPPQ28PbOtoBUIQZWbK
KXTskhzrCIgHFIYYlYQygYdy6snImsMcnCQuBrm/obDZm83V/AvfkhMC5DRDmpnZ
oFhepnZHzBlYHihWwL4MCzm1EvNBWgDF9gC1D5F79o8Lipn1XmTXY96UwBaakNA/
ZTqyMjXRcG0PkQ5Nvp7DWDJl7OWzqcfPvUCIyrE7vfRORFOgr0h8WqPekbnmOqb+
5K9UjelRUa7wSYdOdOC4Og7l0jNnoqCYdtYxuVif574ryBtuMnBMciYhLRmGEmgL
3xO7nT8JhLUHvkJ0Gi+bywCc1JZ7mNXzeoZ4b+hzaqiKcmivdRUZm+kzJznygeYS
m4i7RgjboPPtdXbfmRdI7rkxgn0wO5XRqXyJj+ooJhR+Aahh3+cgDFN3mckUk3qD
k8eL7u1kYpQiU9tqEWjR2YY00DvYpx/Ncp423EI+/JcYy/gfU0X4tq/SE/0B+vir
by0noESSDdR1nVDFZ2cMO0ihWV2Wjr8ZKNtpd8yt/OLKPsU3dydFoqOITdGKjiVL
xavZm8e95c5iATF4H+W+l+kSP/KUtVjg8T6AYG3BvDjo6KHA1UDQ6GRabZPQbjrL
SdM1NunyGqwrp89nmjwn1KTsZhpIG7Xs8LZRD8GDKXJQjRXKX+chAv/0otAZ0oz0
PdJozGhM9+teXPzOmGGdvZKvEZgeF+vFZGMg90Qs5M6xKbnBzIa88NlCDW0aUhde
C37JlhBhuPTblt7NKdaDMZ6x3RblEiGIEE9bwtHl+Oc07AyzymJVzGU/tyGSjDhK
tglwiycN6z+4eBLm/nLmjG+i/75H3Z9f3GsQmsOQefi7AeFq9uLHyJiSamrL1x4c
7VFHpULiHJAm4EgDupw+7ud0A3JbzC0sPWoStEZfk+Hh6NDKmg/e0KYCsDCPAV7x
XpX9jV6eQKgKseB+k8KwsgX83ym6dE1sh10eRJyjTgeIWrL8aCdCVcW9HMIEt2xA
g+VSCCmK3wNpNawC2syLYKfsxoaVGvcHnzxr6Wt0HUHrOC1HV2gkh10ElPPhwgDH
m6CBsJhoUEhtQncgsb/w1y5GrYQd6BSKP8fTpYt6H2LADJo59bi9+zlSdTsVCd+x
TNPfCUPw/q8SEB9XqA4zZSVCDC5yVGHEAnc38ntfoq/2BsESzwXkyJnYUPRBKggp
WY7R2QgCW/HKQmU831JVQET7/s7/zkxB4yr3W/OKwMdtffcXb82cRb+jEYZy6QHK
bQMuSSmFNPX018tZJ0bOOgXVUZYARLecCzn8m6FJ0p0MlDzieT1YMzrtTUhFh7jq
DIKWc3as8AvCT+/yFJg+AqEdf3fZz6hBArq3CJ5wSbMw06Xw4gbqBS4uQHcaUDgB
sb/MjK5weE3j8O5fQLkwEKeZZGMKa2lF1nyNLSa3b0hs7yV/vAyH1koNkFT/UGns
yUWJi+qgO0pZLeepu7NbMdCbuP9QC1CdY646wm1VVddJh3/2yfm4LqZCstdhDUzI
NgkdZ9UBDkHP6RIbYobFFA==
`protect END_PROTECTED
