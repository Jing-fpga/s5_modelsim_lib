`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
io28Sw+/jIa5I4d/gWYwg2h2NS0Ksw6F6g1tAccAHXvYESqL02pPThTaunGsQR4k
94VaaGw/da/d2ZCSJI0qDoQ5R8NTEr9zdTrvZjDQ7hEN1HK9pZiozvchWPKAxpnH
M+DDVwXqKCvJUrEvhIuWJD8x3UIOtpUSSFZuNe0AfUi+VDZs+1Ukpbp8eDPFZscJ
CfnhMghXE2CMw6Gt7fRvGunzjXxMlrrBU8lT0Rnitbz6D2zLlU2W2Lte5mcCA/hA
h0PsLPlFZGgXlYm8liWk16Y3XQU7se0tz5Mj4SJ2uuPFwd7oNskAHdFTLMq3fSxi
TuL3E1TiTeZMw2h5bdcWtbXw2B1H/nERZLAH1uN0Ge+wzJih9UHJWm2/jxwt6D4c
i7kyiQByUQI5mlcQb0qq3SVWVlbvAeOHdkQ9xuEajusY/qYZ71tQAXqDgIIDsypQ
5n09ToQ6KckHtvvCaKBBJ6X4O0pwi3hEh7noajsvyUKXrvAAnJWl6aET5tF34aBN
38i7uam+Rva/n46kkn9hTDZTRoAozp1PR4sVfdYM0gfX1g56Krq/3T4OHOAONR+H
ms147lA0G1HRmfOh7ekanP+uP3klLBf/5r3NjVzS5judda8ltpfkGaHK4QHgCuBQ
Vz4ABEVmo2LZLe8dy7MbodoLM8y2l06fcmDgi5va2VWGhzCVk6TmC2BI/HsqLTbe
hrHoQmOicm/rLL8vhOjGGf4J9c70/syo8n1feL1oVEdR7N7lnPDMvk21A8/hHpqP
oxYV5dspsxmW99F2onQeLJIhbt4o23DsWXjscVjPO0Q=
`protect END_PROTECTED
