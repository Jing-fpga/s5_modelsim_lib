`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NVZNAyHUQWSJK56NS9wrFHUzHWwHQoB/ZVeVffwxh8WZVVMtzptA0DMfgWqd6N30
D45YDKTpbrzOCN/IDw9viY+3lE/SMAUEyzG9RzU/nepCtnaj8OY43HxeisAvCoLL
y/RFWxkN1TplslKcukTDV8s0sjTECpT/XEYCVB+muzcx4C4RwdubxSAVc76SzNAm
lPtdf/wRrPrChrnCr2H5PK5+MpO6ZvzyghYysEt4aCYhfym43IQ9AyZtzp0dC0+5
SASBs0SgkMZnAdHZMczpaXPijvprY11Yu17cgFEgQbi1Jt2iYskM+ubbgFFdyZ1G
BqwZcjdYxYN82vkF9ItEotM+iu1/+71LzD5/xZ34+SbQs8hMAK89hDe5OkQUjIps
kVt+lJ/s4mNzufIEoSbR23TD2NtxVDkM0Du+qOMcD4SmWqqyjnKxIWk/jBVd8ZaC
VDzGxoIJAcU6XKGoMni7ZHxF13fbST/OKXOGHoyLMnCEbcAtLVHVPOQpr+n7sIa0
wXL8C+HeTFa6sVJqfADC5TCsyB4+o42Glg8ZuZ6LdT9eLKsHQy0772LEi9cR7iU9
QV3HFcFrXZlO/vfjc2FQl1kPrUA3rmNA6FCVJ0WjMG1jR6TeJW3pBXRPy4+CoDev
4d86KCDDMEhNI/Dvj/5cH+7u00HCZ1B6ywyzxUvjYBKeTrDCI4cPF+wZyooTW9dg
18sHK07kEuHax2fnIpBQb2amHIOEVyHi4mqJ2dy93pc4ijKadl+R2dm2PPl5F3XJ
q61Ln+YG2pADs6SqZrEb/7vYkYCB5BhE3h4TN7ofb+4jrxdaE8w6AI50snHSOJH9
HHRa3DxXJiHxC/51WGMHf3HOha/K1kSKBrkXGtYDr7n+2x/2Sc2yLvsrYW6pji6O
MpEMindxmm3ZISOFUEfdUfHKLpFrP7ZVSU1F5fLXe/JYwonztbzMOeEJ7kdyHjae
WaOu4fqwLGv79PpeKJ9qNEGtcWHcE+iyPi+t9I9zwsiTjqhhlzFAI3A2Ia4Sqomd
OP1yXVQOjeFw3btnc+9QfUZYtjR6mPkoVGss0NOslHK+4MyKSR6aYWrK/6EtZ09x
4Vg6Yufjj63fa6dbByFqJVw837eXxB9dsbRfNDg651tW1Sm6Aq6MHiqXSBXP8HZR
otSuxsKlmqzhaD5rt/CBHrioWjwwQ8gnc33I8NGB2bp+08FJuUK7iGgE1umMD7k/
DZ8og2OcdHtBXjCBqERxvWfZTyUkLn3RdWz6BPs1SeUWM0lLZbBQYlBcDrVpSUPg
3BJKfbWHgbJNXrTSZRjXEOCaOftghSGU3hX9I69iWmHIf6QcCg1y6etDqiqQH7uX
cUfB/4VLBpdSOiGg1SaYjkKDdeKt8ISqoRv5yEK7r+nIkLo+o3PIopxyWxpt83TM
WFS4bWD2TxpMcdySR49jDtonQ19pezub4oVn2197lP/V9+zv6OKJehaI2+Wh2VTa
h9+wzSq6BERIBgYpfjLzLLTGf3D6ljTmFfG7Kox9SZ34CpG161XRIqatTryA5Ray
KnmqBFFXzM2BduqWD17HuoZaZW35dZ9/Sh9uMg8MaPtocUv/hBiOnle3cMzcYWnd
WQzxYGHMnjcAwdtoPn/VAPLAYa3gnECCcCoPCWQmvbkO9TCoVLk99mTAQCl4lRbi
+r0tYmYipFYxaUBnss2Vg3LRjxupbJkr0wFSHWXunlPLIDnedUU0O3V8o0mBaht2
iK+iIWaLIqZ+XSAB+LfD5V1Qb6nSzhGuy9cyqsZhP9siv/DUrwfFra6X17r5C9ca
Q48dQko5EkBMH/I5gf2NA/a4FyFm4LdE3leI8uo17fpkrLm/56yyd0qDeGcl7YEy
bcManPrpf+SzVJDuIjOIFCaMSLQ5qvxygdqGhPEXrLH1qHCZ9AddBaNHNsPPo4DG
`protect END_PROTECTED
