`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pfH1MwNRQX4zRe/gGGLtQdGUFC1MYP9efzVkqrMhmDB4e/UW/5g9SXpbFrKFUNRB
SX7xs9JZhtZbEtOUDTPKd3UZK+9bO/2dhayuiPrdh9Pd2/BhwPzKpcTLn4QArMpw
F4IUMRZ19efB0bgsMBScbS+Pe62H1FtgwtJXQuw3blFg4WN+sVaCmnlZHUxlSCIZ
sgC+zqZzbJQduOkB9t/FrPBT54NgwMkY7M7gCkAwMknu3wC1LgyfG+l0uh3xBnyZ
8RbxTOxO5vahf7i9IH8/MtOS9K2Xt/Rng6IDB9vjhS0Wsk1EOECe+2OutN2v1tFN
oyngoYDABhEBiWynHHaINkxHLIYu0jx4t1H3135M7Sh9o1A5pJWUVRmBilAZODR5
zlomQJP34r660+zn7K+4bYxL5rUnGREzeWmMOO+QKZWLBcODnnPtEAe7Q+WXeAkI
fwuHMBZd9sD/wwSVVVQiZkSs4puA5n4QmaGMeACDxACsEpLPpGHHBLz0K+LKs8bW
jvh1CvuCRHBay9M1GDYfERf96ZCBi3Y/2Twnb+DWDfONgs1AFs4MxLFOMe/IH+ay
ZxRMr3rg0DzuyYbg9R3mMMT8oWmxik/GbCHyDpVhpAxDC/3golOJMuYl8toewHIk
9A5hImIBYX7dCVxyZdhOrpjp2CTlReX6hWQ8myUqTp+/NHZu/L7v+st6L2ICqYId
B1OagL8YutqHUwBdd0H3gZWE8xzbce9+mDX4HpKX1gcfIZO2319LqV8xgQPgfJhL
XVp/rLH5TEcfNKxtMlqUDqjsQvcNTGVqMGwQ2SVZUkJPTNF1aEdNCn5PFHkv1nix
iC4PBXhVqzQb0edWmEFjkX9bL8PLANxJw/ie4NdFfKtLfyfkWI9bgneGfdtpgKAd
bE2oi3TxDegK9cgGFP35frq7c9AIHIISMe7qAR88CWnX+bZP5ifA/76pxPlueS/u
5MsTAG/HhhEQQwPUhgXyqFH2UQL6ba6cCRpk8Yc2xESmPr1ok8f+R1wV1P06OWA9
P9hWk6YF7TZ+iPBfhSHh0yLeg+kP20su+yr2j1+ckIVHsVbF0eRF2BbODMPeIbCE
oEPbbGkGDV9TWHWIMg8JYb4rG6q74x5jmgfYCw4Bnzapc6VcFcKAEYyHoAl7w25z
+QMDSc3VS7i9US17Hpalm61OOI72XoBBksDkTaOC6VTEdMFclh+4cM+JBENKhJPs
gfC7h8tstaQR/WvrBD/FqJ1ynY/LFdmMYr04Ff7QXN5xfMpCDgWO318/AQ5J8sQL
ku0nT7jewRKJiNELKLVrV7OWEesrXuNbClm1192BGZTVzyf42i2TDsJXvhV6E1oo
JEvoFtj0L7Z2oC8ByEHrut/xQLO4HYopEG9ooC01OO6BgknvPddviQdZ375GqURY
DEmacTJVf4lUik7+bLQKILOrEpSSfpbpdM6Se7fa+V6iMCQ5kVCExc5TsBbLur6p
8rVcHTUagT1bFqJ+HFgoIOWdFqVYxutCZ7ir84WeveWrsCAYbwWCXNp2KTAG3vSa
17on4bjPTu6W4iq/2JxsJ0QP+mWoEBf8ypDUs5dwKHDjBGj7LwjEDfDjPCY4yBHg
n1d0hlf3lo2r/l9OtEWKyAYoTuLjKNcFvw2PtjQy/Uc4Jyjx/wEWC8WeoJKc5UGF
f0uaK5R4L2cgcsdxhX/DtwZyUfyjUW1iz3nhlwKDZBrtSPaVwbm/G9zJMXUNbI6n
egEFbt7vc7E9CgB9emx5rYQ74VRBDNtlMwWP4pSxJQoU3042mGyybE+BCPJCr6lM
RU515NB1efPnpvSZJI2cZxFAKAGLJC+/cCsxoUrxdhCH71Mm2ZijMGo6n+bFAtJt
+gUH19hY/lDXLmquV1vRon6t3YQaODyDUSMDllD8R360bWNLQedQlAhR8PyNCi3O
CDNfrwQhoH3YjmgmiCAXW4XvsNhQdIcCoOCL2y910HbJHSqTlndEE9R7TCX74N6J
KCCWMeXC/HecrREPgPeaOq43IWKvcXVaa0/JIeeLna/fC+GxEeznr9z4MeCo/tn3
y4viDBjmWjJnHJrW7jZLQmMQ/XHCQ5thELNeBcuS1Vo0TCQ/CPWM/wKLcpWuogjV
HHXCACSm6k7rkn/fYsWl4VOn385f+8fnPBd3mekuZ4Y=
`protect END_PROTECTED
