`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jk2cixFQuoQS7BO8sqMMYum6cmFebS5QnkUCBv5CCoOyw7miiSdmjOceaf2Lm5Mu
RdQGIQZORWvBIZXTSlxY8TG+xCV8dcKgDGECusGAkh6NXng/R1fMsffIf6kj0pEY
9yv37HeGbcLKZFR3XOAQsFSkWEKvUH4J0A8r7ruHWeUeorFOPpKKscVrCmw3L4w9
ivOeX9v/QZRQFXQc3f80FcInNeJZxh0fmCn2y0GzE5zfrAQsbxyfyJ/WkozRyb4Z
3TvIhrY+3M0zIlSeXFZkfHpEWKbo+tnPjdFZzygCG2TAlzIQZKdd/9PfqsRCmdIQ
nVFtNGYMvBiztcGd1uQhizlel16pf1BlUPOiPGWuZAD7XkxS+LNXWyrC7k5ZVGnw
J2OInkUluciGGUKjjwwMhPsk1oAVMG2eFlfKTRAhCcI7mXOpEkWJ+NBg2P/sdtmQ
MnZQWCD40Nz1iyDQLX+FmPnYBVvH6/Y5VUFF2vEzKBm414wPSZ/FFrCNzo4blboG
L5muzfNkt50Lm1TfLRp9nWh4uMYC6OtekndZlqP1FYt1bWWSLkgxGkg1QMjcmHdU
E9ng41d1McBX2FtYpXS5H6YYeIvNxK1/tNj/rlYJtWtbjKcGGg5KcJSIPNxZiLIP
p9Zny/fjSYyOLD9TNgvfyaIPqHfY1yAB55GCHLXBB+8RsIkLqjzbDgAlYHtWqvI0
kaffBb6tvxfBBwNyYstrxvnZ/vG/Js1syf4TtdoW8wsmJlQBIPYa+SLvUKy8lq/i
JkKFBZIS1JiTl8mv7p53xEDs0PStYoDKqT5xyON9qSL5l9voRP+egWELbOJtp0Z2
+Ju7vJtJpBTkxn3j5jr5qUTuH3nZEWiABcdmI6/IBRYjG8jvnHSZ1cs2zljJxA+V
mxCY/AA1w4TW3QA9ZC52jA0CN9RcB5kH88z6CkS4P640X+pWKIxvsBfuXkuagwMo
`protect END_PROTECTED
