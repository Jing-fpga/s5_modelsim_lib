library verilog;
use verilog.vl_types.all;
entity szmkt_tb_sv_unit is
end szmkt_tb_sv_unit;
