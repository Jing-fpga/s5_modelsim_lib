`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
byFDKqY6GsPQ1tpjKlnHDmhDdYlVVkkKiYYfOs/gWCKOf+LJ4DbM7XnNYdxPqe4X
jBoXrjknwukqMMEHbZpsfzAQ1dt2w4OBt+6xORcOqLdbc9tDARr7LU5v9fmQ+5qy
tAr5utCZC98u6F55rcS7Ks6xbR3tlN38bqEo10rJwf0Q3smnIu/IK7oI+pomcD0U
a9MuLQyKUjdb4Wu1aXXgsH3o5yBobk20uAkwVB7IrSnhsMJbL8tQkSnXTSkn3cM6
NiCR8IwYYo+Je07wl/DwZJOap7Tr0hseijV/FrCEZHtYISiTVehdhPbZTWgZM5DM
EFd7AoWO5MT/BiB6mxv8pNq/qKu1gU4FOizaKT207ZS12bkEOU6/WiHO6dP5E48v
6sUESx8K8LS+qGWCvQI1mumGXmXT+iAVc8pxKdRTPNLUkvzQLfCOOuWUfdSjxVjC
xziGfGUEA+WyVvQNxnS6PPuWeEFKmHEbRdxKgVbj4CalXua1BaZAw6sjvFGdHu3g
VHadYy5LHe3vgm0hZwU8+xhmFkXALBlJZxIGrADmCGmpIlFxeieF5otplVjeIs5x
oxVV0r1GvGpyDIbj/TB87MdVusd0NjxxO3He6x7X1ULOhVRuxKPaD3gtZ90ac7zg
VIiTJdk9ycBRCxVVOPSXmkZwa7mKlI272a2HUdbymQUiONZNdtX8fNLEQjDkLXmL
9i93YBSlIRJ3DpVVpFSBppj0P22RSvN4hK0+mhJWoX2FH7cqlA0gw0OZo/jz/62X
UhbLMFO2kNkvoULxr8B6RzmveXKCu6kLCn0exA7evgIsFyATwPmF24qF3xfKdxmc
P75miA7rNrCD0/DtYrfEJyWybwzg/IkPONQiHpeu+QDBW3YJAQQzVGyCdvk1Ikke
/wsLkKezgnVttoGi2+caH16P/vad6H5IxVJpMKiwZ+dMWo4ehJUatYrm08rE/A4r
3mtQygmNEjbRr+wvxblSNhkgKt4HSHbd/vaIq60Y4O2Ft8Td4dqmHTdo+2ycHB4N
jiBNoIA/VtpDH3vcQb57xatbSFSLxxmNVTxjj802Fp5YPDAFvAzNM0xhLaXs04kq
Y/3fGzkXHaWhzLr5XrgHbdE06L58ncQXbRNcbbwul7wUtucICnpSOjWVNegEQ8BS
mrSRT1HjnXAOj/PX5aEfIsQMvaDhzyKXnfDh/RZPKPbqQDIc9wNXCwXLYWR+RpYg
+Ob8vB6Hb4wHwVeuakAgHlsHrqWirR7V/Gw0BC+iIFVPbtXFgpaLYzJRs4n2Ktlp
6pHHfhBvw42aJSXVgdPx5NoPY2oSIi8kpcPMTq2RHQj8P+M3yTlUW+No0GvR8Qdk
mn/rAmlPEdQGbXlnevQzqg==
`protect END_PROTECTED
