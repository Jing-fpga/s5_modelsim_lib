`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5/Vl6MfpAZqRWamZAggQMeuXZGx/AedDubP9ky1oyt3pfc5ttS484QKkYj+hQi1U
VCg1tXpi//KMKB9J2yFEwckEtHMmN92kLjf6XVzSXqr65jZTSZqknEFfGPdloTq1
7QZ37riSDQIaDT4xnBbriuBLMqA82g/AqU51H42yGJvv2tMZaFG569CApPm2Nyut
0N9nhCUAfnkLKgtIcnjN5ioF7FM9G8cTBwFTl/j6NPNu26yjI157eNXul65X3SYg
c9l+X5erlVVu3wX7m1UuquhEgAkcbJbL7BHNKrYS0cv8UtVJR5qrYgUrCJbJCv1k
fh6bZEQawPUMiTFvkrGQNNf03nICLyHDVzs+SJ88absRCAS8TBFlkhhzodqRMuWM
F5Z/C/cPeTgI8YYP085c5IGFfYqpzkjhGTzDby0glFAtR8raNE/1ZPThHm+EZo0N
XtnfS/JRnKmTV2/JkE9y/U8WWei3r+P9GDNlQROlAdPmOz8/aHQ7PFnDtCvBPtJw
z/wi67N/FH76vsOvhbSqBuoctzWOLYFb1111f4GkhBK1yrxsPeNuX71aFWIhT4Jj
vO1QSudGCbvPOYrxhW3fPnrQ/VhsxQA34Eav0qTWAfFP/kV0yKWI9+zJ8uyXTM+w
I0uJM0CWaAVQGUhUiqvO/7cjitOFKyvH+3b/ptw5ebh0Bz4MkUbCpzV0HQnXEoNL
eGs91q4vaVqoXpzD8+H4Zm4sXBZAfmtl2Mo4ZkjqsH4H2AFr1p0Q7F1CBBam4Pz2
oG8IOoi8cmix4QH8jYMMPgDxV0kNAutb4hVyYi0LIGyBL0W/bEz772qnAsiJv3uc
r/z/rIEGfP2KVOJrU2WC4jQMxHuYsG/ellNkSlQNdgsw2kW0viUmnZuqLdLEHP80
qqA/06xFk7vRpEM03ApU7jKW5K36WvjYVEbTtF3J3PR7H0d1Hnba3f3HYzuSZyXT
HExMZKFbZWlNKLFlllYERbrTxFKLThk4nvo7EALAgnPAfw3NxVH+ifYld6RJ22O7
fk22Km7i0wnxq+sraU50YT/1pPx//3wHVyJRA0oZkkX3oSD3Sm5g32cbciTARpsX
i9uLnfue2g/x5GRm/ZSAlLWYp51RISCj8qfULy2jFKMlwugyYRFtLQFnT3eEV3VZ
X2LQkvdFkECFZhr8IcfkEQhwMTslfgmnoAeXowmMt04wyG2jrc8L4wldEkcbgdXG
axzceJSFknFpxP5/QrT42CynFCkMfhY5T8RXkYVFKEIMJG5wKOkScTKXW9/n5YKv
5SbuKR06wTCiIDEF3UxENtosLrfq29o4TWZhB48Zy0xEI0IRU5XZPUJKuuEPLxTI
BHuaUHYinKaRAwiyvNsMmg==
`protect END_PROTECTED
