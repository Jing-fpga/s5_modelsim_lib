`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5M5NpR+0a+LXUdPauJIp11Q6/gsVwjVOIgzOoVkZ68+MSydipqRw1RuR5KzWESJ3
td499bTUUmXOEgUhl0jEHFSHq76gbKhnLyQ3UOPPQnvkn4I6Es/2fReZOohH2ez4
PPta9+QVjqDLxXYggDPHs85JEVMd5d6jyukf9o39t7qnerY09RsA5CQpXnwijw4u
KH+U9GTw6jlWSs9oy9hKt2pWX5BJma0DkzMuovncG+xB+mQght4CSN6pBww5maIe
aUlKu/GuRQZk5gMd89taOJ8RK2S/NNhjsd90XbiltIsIQRewqoY18tmYbYi1EACe
iPp0+Xy6WNVSdtu4WTeniMHq/BSlk24+qoMpRm3LS76tmMFK/o9M2PFzXNcjb0jp
wJzGuFAcBgjf8+gTHthoLQegtUtPxDLNznRDsgrVjEoW6+tv25S8VBvRiQcpRrJ7
7nO8Kyoe/2O2ukUOfy8d0DU4p6r/Gan6aR1PG9BSJ6T9SjBiartXhN9V/98lhFjN
8utdzOu2Aq4a/0kXhTgWgBJxqNjTFanxzQiWND7Kjw4RCeWi1mVVqMCSIz3CYkrg
PCRmK6NDGUEylR2ApZHWt1EdsuXmnVzeHRbNJX5n5cWDmDQGS7O3B7LKgd///VkS
pKW0TSEZjTaZzeWlG/r1iJZLS9ugp4iIV3bslGm+bMTVHZ6IrirC/o07l/IKGpyT
ETYxZ4lNPP6Nzcb/opr+tFxz5Z60ysHXDlDeqd1MVuL9An4ocoSBysZIB6CczFEE
tUGolviewFwRuH0E9BeNs5VbPo/eCwAAwuif5knw743lSrGpNwXNqsLfjDpUb81Q
WvP2UGjuKeKzxEuBiH44GetMS3/xiIscAB7Me8If+UvLurIO0iMC5xZgAvbE5AmL
6AvLGs8LuvlPbCsf90GQ41CPc8wnnsU6NmiKoqCRqtX6xmBVEn2jbcM0G++L7AYq
pcjPQEFqy11Q6YQbkLgUCchseJwODKk6ivnQ1mkOQwIakcz84IIOKRz6HgjT8FXp
vA6PGU9A92xMcZFxv0wxVfVMeuOdeeoC6nfCZSNO3W0Y+6b8U9oCMrW6hpKIBINJ
1MNT1DkWQsWNKTbcQnnfAdl1gVB96Uk8fvla94I2MU0NnbNTFDyJEpjBh6zrAtO6
xsyhKrGhIjST8Fci4/bbxQQSyHxO+XnX45+K0PYOdzy8yzpnV77qYkALkp6Eq6eH
2SZSDn7C/ac9QUns4kxY/taA7ZFMsWyDjaq8QGrWC2JGRSufu/V84uBg0bVDUptw
opCzu01kMZqyNsu0oaVQgcD/JHXz4SAzobvFx+idaVCIGeK3MZnIqLL1dabOXUTk
AIYKbY9KaIj6om0aGrZ/MoDAESv3OWNw1hu4FesNYEv6rvyhlkNLI6OrXdkg5aK+
zdZMHZ5fN5E+w/mGxypSp2eJUgcXqsN18+8Wub3rIsG0tEG0v1WBgNQNYypAiJTd
cqsadcMAVLPlsaZxdKkIGUwsCX63oAJNMJvv0iXOe3brMvhxhUyWcdmLQVX6PtPa
`protect END_PROTECTED
