`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kH0ItIHolZ8oS6vNHaVuVPsoTYBldJp3e20taD1o9N0U9UF15Lo4aq07/KFSJmhB
9+zMBqbxbAVryFoHoaat4s3ewddE0cLaWxepRD5U/vfiq0T26ooFMc+xq8p+Io2+
Qs6OZ9qTc6UqRXg1YcttY+0hqajKK9CwSIvPZmxZMengfvBWsh9Zaz/uV6JRDfm8
TfCp5TSA8iUezcE457OafbCZ9O7IVsXioW6pNZmYMffv9EFtFvDfQKtaRrTLq0Rq
tLaxwxpCc/6wU5xx2auvyr5a/Z5OAzrwBmXFXLeCx7QrpaONqXv8wWPcwh6B5wbR
uyQhr8OyQYlQxbpuz+gP8XQHsj3Ml5q1Gwxqv3kkwqIat3WJOslKn41dsn9qhDLn
71r8Hb0WvlrXY1cbxgHpRqiIAFuI/0yuuhDmca2S+n/J1cAxTZltVWTTdM006onN
DZdXRAYU4N7NkO3vum+Pr04ppSXXFscJvmsHmf5Xposm7eo739Fdtko2fb0xpZVL
zu19Lf5UFBPsdrSaR91DajNv42xuM0yWt/DjDNBvM2D9zFd7HYQTd8Zt1B/SC7dt
oX/jpGbuzsNUQCJtgkaolmkdsUyVEmOF0JohNHz9x0iFsCJzXo5ipBJuDPUiewuv
9+fgrXJX0WsecwKm4tC0GkeqMT/+jKizhoVZQ7767xoTDxLcDsNl8gDrLSFwi09o
/VTJ17UqePHEthJHzgstSnyhNssAUHpJFKFREQmUcyQwyfe/x8/ovaMeACkA+KQp
VJlJTBx+Z6sCho7tbHshQtn2LYU1YknIgk3whzE1JBLGuka+qE1Ghey3Nbru6hTQ
iYKx3T+uP4Fl0UpakCbr3249/PoCY4Fkt415p/4jzCDwOINOjzewEapFQCauzWuI
`protect END_PROTECTED
