`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qjDa7n8ty7RiJJCJxxGc2HKZ1u9Qd0qCWddOvolMbzJr3pNhWIuxWqKTHcmQnG9z
RR3SSYAgUtz8/UKvlQCAxorVVrvI8dLTd3qV/PQkiiJxKJxIts9fedsh0v4gwNAc
6GFSiZ59tt4hvUd15R+nKxY97XvyxsPitD+E/VWs8ycA5RLDKn7gRCKkfO6MdmB/
HahS8QdeVDmoYOoWULABmE84O+pM6Wcw8y9i81p7m0OxPJjO8XoTl5lx/8IW3QY9
UcrqHE8TTDX/vc3uEgzggLTkkkYKRKwxrZhUaqOqK8lJxShW1fCN2zhLnxtNBbbn
i/DvveBU7ja9lCR2MuL7ScitoXPTmeqqHiRY2V6icZdKQPCsAgLUMb1SZeM0sjBj
wqjSfvDjU7OO4JtkgwDIn1B7Z9CvA2BPL9DlJZTUcVgeuXbnUoJGDqo4x3zXZSIv
bHKLk+nWYfzPhcu/7k7dWZlXbQ5OtgfMXNqmpBbCn2/IezGEAlGsW45ih8K/hyTK
j6+500KphVvZQ30Kf8GOIHi7xH21OuLNkUtnvVxUpaJz6BqFXuwzhcFv4bh1VOt4
FTTL3IwOeUZZ4Oubd3FtVQ4Y3nTsyZelereo5LGJAYMNQygyT4+TLAKPta4GWcAs
2dhgkXrQyzns26orrKg04wenQVqWP2AVwqc/97R64Dz8t05nuDZFBJbwoIyKqqtd
Yi+HErASQy2Jk6ySmdOIC4Whdqcez1U4rofb96bnPShsH037N9JmK2+JQwoyxeG2
WmoFLpn0I9B6pX30TlrIfKdLKBylNclmeEdijjrMMWl/wMdUyNdrGBMCnGjS1m2i
w0wXGsBX2wHCpiwYCmPHYnsq5cju4OYwP+F/3FX+xsKNPvSzSKsFzkGBSQ6QeHfq
M/4Kt3TJlLX6CwqarJiW5821H9bu/pjuYbhSe5tCZrQ7sNKgGjPr4srinBEcym6Z
iOAOHHo08D2M+sGH73TVTGJTLt1fXakbjYN/Wp+vsZD9VBT2pkRtrTfvP+EvYhh6
eAYKDBHAE70fcJ1Vy1RWJ6yR2FCZbrbcJemKQp7djMHg8+Q+algR+wjD6wG8OOXV
L0+GZaMukp8MFcFzdNkxzLdNN/D5lmsJlFAe/owP+bArba0g2Ayj+plWKoN5kbku
06IaXKryv8kYb4d7+3s5HhTvLiAkSmO2GBz+wDxd5BUwDs8sK+EouwRuj0/xvpvv
NpRBO6GZbCkWp0zZiXJdZ52/LCyvq2XfUUSnnhc1fSqF6M4BJtH5iciHlVynZxDO
nHHUUrWxoAVHuT3B2r/rT5Cd7mj/5A0WGTkRnv2pUO8CcwK9RpKoi1J3qIym6gBG
irEtjgGRsOHyysf23FwhI75y449tqGXGRD6QwhSMC4E3Btr4aoTjUU/NW0GCjpje
gk/qzlQVH4rjyVi/jc+agTrr4TLPWCddh4ZN6he2eC6TSqzhRq4Ap4LiIvT5RdzA
ravA53oPkGVb6RsEMpViCcodMyQ0b8ppvVyqUxky5nVNqXyB87DPpjrCcpRj7taN
5+aPPh4sYiokxZUNOMrI/cSKY8WUbmIFYHwXPAbq8tWVX+OPg4uit/6pZ0FyBbFp
lGrJ4ZtEI4xED95owDtJn+FBWbx+F+Pb5ir8pA2sV+NcAIGPl7tL93WQTFDRxpg3
WPBCiR+siNHXwgWqacPb2/vFVwjzHskuYAsV8SXfE3KZywX8kW+lKJkCVxGPbTp4
PMScOZ/QWv9xZgiuGYpMvngqrlugwB1xeNEv8uWWae+cnw3Jrk1leQji/+/jZ8G/
vgk8gTFSYXahlBE9bYqTfFQDVN4VlVAp/DqV2LZgQJX4AZx60ksKjObh+bq21RPf
kIFyv+3BUyeLI5nKJTqS44m1Awjg9LX5TvBSLcdi1qFrZ4WXOFK9MJP+OPzZD7uZ
XAp0WcPT4qKyHwmLMKLpOA==
`protect END_PROTECTED
