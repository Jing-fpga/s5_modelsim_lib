`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
42xY+R4SYU8UAvz0vbCFzw2jE2Hl+qY44/RMzrnhzzxLUvWvzIcZQcaq7tVawREd
rxKTpCdx0ZqxIsdcHeclMj5vph03Qb54XXNTmWTACIsrl96lsw6qCqpOwsH0xSZ9
N32d93MbfyxmwOlWk8XL1rwIjaoE/lDIMXp0YVNWV0Lw4EeXfmUWMpiPFBde/e+q
lT1oM1cLLb+PNQLLBfMd1TpdHkDJuSqthpo6cb1TDv82fy6mDWqOwf6wUyl2eERd
cba3HA52n76rVrF0/mMAxZ1uRj3wANF2IhWePEG2a1MoUAchNe6/gA7rLwHBN/YZ
Ari7X1pYQ71PVluw3bkrybTbGvxxCZ00Jmjz4tzPuOpnIb+zAb+MC2Ejm+pPtY09
YF3FKOovPOnC39vGUVcn8Mjq2f5RLjNwObmkoPh8cnZNxPztBX2JNy9/HVqczFPX
FY6rA28xoqzjG8FKxTLZEwPfy3nLwE2gyHKuRQsR17YW6iQLd0tezxwcTg9O3pvg
LWFWjUfubvGUtFJHn/nD34+DlEvZRw8cEsvC9xPMIEwU4keAJsicgP5JBkbfna/p
A2YJFdI3yU8wOIkYYAIw1w==
`protect END_PROTECTED
