library verilog;
use verilog.vl_types.all;
entity stratixiv_hssi_tx_pcs is
    generic(
        lpm_type        : string  := "stratixiv_hssi_tx_pcs";
        allow_polarity_inversion: string  := "false";
        auto_spd_self_switch_enable: string  := "false";
        bitslip_enable  : string  := "false";
        channel_bonding : string  := "none";
        channel_number  : integer := 0;
        channel_width   : integer := 8;
        core_clock_0ppm : string  := "false";
        datapath_low_latency_mode: string  := "false";
        datapath_protocol: string  := "basic";
        disable_ph_low_latency_mode: string  := "false";
        disparity_mode  : string  := "none";
        dprio_config_mode: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        elec_idle_delay : integer := 6;
        enable_bit_reversal: string  := "false";
        enable_idle_selection: string  := "false";
        enable_phfifo_bypass: string  := "false";
        enable_reverse_parallel_loopback: string  := "false";
        enable_self_test_mode: string  := "false";
        enable_symbol_swap: string  := "false";
        enc_8b_10b_compatibility_mode: string  := "true";
        enc_8b_10b_mode : string  := "none";
        force_echar     : string  := "false";
        force_kchar     : string  := "false";
        hip_enable      : string  := "false";
        iqp_bypass      : string  := "false";
        iqp_ph_fifo_xn_select: integer := 9999;
        logical_channel_address: integer := 0;
        ph_fifo_reg_mode: string  := "false";
        ph_fifo_reset_enable: string  := "false";
        ph_fifo_user_ctrl_enable: string  := "false";
        ph_fifo_xn_mapping0: string  := "none";
        ph_fifo_xn_mapping1: string  := "none";
        ph_fifo_xn_mapping2: string  := "none";
        ph_fifo_xn_select: integer := 9999;
        pipe_auto_speed_nego_enable: string  := "false";
        pipe_freq_scale_mode: string  := "data width";
        pipe_voltage_swing_control: string  := "false";
        prbs_all_one_detect: string  := "false";
        prbs_cid_pattern: string  := "false";
        prbs_cid_pattern_length: integer := 0;
        protocol_hint   : string  := "basic";
        refclk_select   : string  := "local";
        reset_clock_output_during_digital_reset: string  := "false";
        self_test_mode  : string  := "incremental";
        use_double_data_mode: string  := "false";
        use_serializer_double_data_mode: string  := "false";
        wr_clk_mux_select: string  := "core_clk";
        use_top_quad_as_mater: string  := "true";
        dprio_width     : integer := 150;
        migrated_from_prev_family: string  := "false";
        mph_fifo_xn_mapping: vl_notype;
        MPHFIFO_INDEX   : vl_notype;
        MIQP_PHFIFO_INDEX: vl_notype;
        DPRIO_CHANNEL_INTERFACE_BIT: integer := 4
    );
    port(
        bitslipboundaryselect: in     vl_logic_vector(4 downto 0);
        coreclk         : in     vl_logic;
        ctrlenable      : in     vl_logic_vector(3 downto 0);
        datain          : in     vl_logic_vector(39 downto 0);
        datainfull      : in     vl_logic_vector(43 downto 0);
        detectrxloop    : in     vl_logic;
        digitalreset    : in     vl_logic;
        dispval         : in     vl_logic_vector(3 downto 0);
        dpriodisable    : in     vl_logic;
        dprioin         : in     vl_logic_vector(149 downto 0);
        elecidleinfersel: in     vl_logic_vector(2 downto 0);
        enrevparallellpbk: in     vl_logic;
        forcedisp       : in     vl_logic_vector(3 downto 0);
        forcedispcompliance: in     vl_logic;
        forceelecidle   : in     vl_logic;
        freezptr        : in     vl_logic;
        hipdatain       : in     vl_logic_vector(9 downto 0);
        hipdetectrxloop : in     vl_logic;
        hipelecidleinfersel: in     vl_logic_vector(2 downto 0);
        hipforceelecidle: in     vl_logic;
        hippowerdn      : in     vl_logic_vector(1 downto 0);
        hiptxdeemph     : in     vl_logic;
        hiptxmargin     : in     vl_logic_vector(2 downto 0);
        invpol          : in     vl_logic;
        iqpphfifoxnbytesel: in     vl_logic_vector(1 downto 0);
        iqpphfifoxnrdclk: in     vl_logic_vector(1 downto 0);
        iqpphfifoxnrdenable: in     vl_logic_vector(1 downto 0);
        iqpphfifoxnwrenable: in     vl_logic_vector(1 downto 0);
        localrefclk     : in     vl_logic;
        phfifobyteserdisable: in     vl_logic;
        phfifoptrsreset : in     vl_logic;
        phfiforddisable : in     vl_logic;
        phfiforeset     : in     vl_logic;
        phfifowrenable  : in     vl_logic;
        phfifox4bytesel : in     vl_logic;
        phfifox4rdclk   : in     vl_logic;
        phfifox4rdenable: in     vl_logic;
        phfifox4wrenable: in     vl_logic;
        phfifoxnbottombytesel: in     vl_logic;
        phfifoxnbottomrdclk: in     vl_logic;
        phfifoxnbottomrdenable: in     vl_logic;
        phfifoxnbottomwrenable: in     vl_logic;
        phfifoxnbytesel : in     vl_logic_vector(2 downto 0);
        phfifoxnptrsreset: in     vl_logic_vector(2 downto 0);
        phfifoxnrdclk   : in     vl_logic_vector(2 downto 0);
        phfifoxnrdenable: in     vl_logic_vector(2 downto 0);
        phfifoxntopbytesel: in     vl_logic;
        phfifoxntoprdclk: in     vl_logic;
        phfifoxntoprdenable: in     vl_logic;
        phfifoxntopwrenable: in     vl_logic;
        phfifoxnwrenable: in     vl_logic_vector(2 downto 0);
        pipestatetransdone: in     vl_logic;
        pipetxdeemph    : in     vl_logic;
        pipetxmargin    : in     vl_logic_vector(2 downto 0);
        pipetxswing     : in     vl_logic;
        powerdn         : in     vl_logic_vector(1 downto 0);
        prbscidenable   : in     vl_logic;
        quadreset       : in     vl_logic;
        rateswitch      : in     vl_logic;
        rateswitchisdone: in     vl_logic;
        rateswitchxndone: in     vl_logic;
        refclk          : in     vl_logic;
        revparallelfdbk : in     vl_logic_vector(19 downto 0);
        xgmctrl         : in     vl_logic;
        xgmdatain       : in     vl_logic_vector(7 downto 0);
        clkout          : out    vl_logic;
        coreclkout      : out    vl_logic;
        dataout         : out    vl_logic_vector(19 downto 0);
        dprioout        : out    vl_logic_vector(149 downto 0);
        forceelecidleout: out    vl_logic;
        grayelecidleinferselout: out    vl_logic_vector(2 downto 0);
        hiptxclkout     : out    vl_logic;
        iqpphfifobyteselout: out    vl_logic;
        iqpphfifordclkout: out    vl_logic;
        iqpphfifordenableout: out    vl_logic;
        iqpphfifowrenableout: out    vl_logic;
        parallelfdbkout : out    vl_logic_vector(19 downto 0);
        phfifobyteselout: out    vl_logic;
        phfifooverflow  : out    vl_logic;
        phfifordclkout  : out    vl_logic;
        phfiforddisableout: out    vl_logic;
        phfifordenableout: out    vl_logic;
        phfiforesetout  : out    vl_logic;
        phfifounderflow : out    vl_logic;
        phfifowrenableout: out    vl_logic;
        pipeenrevparallellpbkout: out    vl_logic;
        pipepowerdownout: out    vl_logic_vector(1 downto 0);
        pipepowerstateout: out    vl_logic_vector(3 downto 0);
        rateswitchout   : out    vl_logic;
        rdenablesync    : out    vl_logic;
        txdetectrx      : out    vl_logic;
        xgmctrlenable   : out    vl_logic;
        xgmdataout      : out    vl_logic_vector(7 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of lpm_type : constant is 1;
    attribute mti_svvh_generic_type of allow_polarity_inversion : constant is 1;
    attribute mti_svvh_generic_type of auto_spd_self_switch_enable : constant is 1;
    attribute mti_svvh_generic_type of bitslip_enable : constant is 1;
    attribute mti_svvh_generic_type of channel_bonding : constant is 1;
    attribute mti_svvh_generic_type of channel_number : constant is 1;
    attribute mti_svvh_generic_type of channel_width : constant is 1;
    attribute mti_svvh_generic_type of core_clock_0ppm : constant is 1;
    attribute mti_svvh_generic_type of datapath_low_latency_mode : constant is 1;
    attribute mti_svvh_generic_type of datapath_protocol : constant is 1;
    attribute mti_svvh_generic_type of disable_ph_low_latency_mode : constant is 1;
    attribute mti_svvh_generic_type of disparity_mode : constant is 1;
    attribute mti_svvh_generic_type of dprio_config_mode : constant is 1;
    attribute mti_svvh_generic_type of elec_idle_delay : constant is 1;
    attribute mti_svvh_generic_type of enable_bit_reversal : constant is 1;
    attribute mti_svvh_generic_type of enable_idle_selection : constant is 1;
    attribute mti_svvh_generic_type of enable_phfifo_bypass : constant is 1;
    attribute mti_svvh_generic_type of enable_reverse_parallel_loopback : constant is 1;
    attribute mti_svvh_generic_type of enable_self_test_mode : constant is 1;
    attribute mti_svvh_generic_type of enable_symbol_swap : constant is 1;
    attribute mti_svvh_generic_type of enc_8b_10b_compatibility_mode : constant is 1;
    attribute mti_svvh_generic_type of enc_8b_10b_mode : constant is 1;
    attribute mti_svvh_generic_type of force_echar : constant is 1;
    attribute mti_svvh_generic_type of force_kchar : constant is 1;
    attribute mti_svvh_generic_type of hip_enable : constant is 1;
    attribute mti_svvh_generic_type of iqp_bypass : constant is 1;
    attribute mti_svvh_generic_type of iqp_ph_fifo_xn_select : constant is 1;
    attribute mti_svvh_generic_type of logical_channel_address : constant is 1;
    attribute mti_svvh_generic_type of ph_fifo_reg_mode : constant is 1;
    attribute mti_svvh_generic_type of ph_fifo_reset_enable : constant is 1;
    attribute mti_svvh_generic_type of ph_fifo_user_ctrl_enable : constant is 1;
    attribute mti_svvh_generic_type of ph_fifo_xn_mapping0 : constant is 1;
    attribute mti_svvh_generic_type of ph_fifo_xn_mapping1 : constant is 1;
    attribute mti_svvh_generic_type of ph_fifo_xn_mapping2 : constant is 1;
    attribute mti_svvh_generic_type of ph_fifo_xn_select : constant is 1;
    attribute mti_svvh_generic_type of pipe_auto_speed_nego_enable : constant is 1;
    attribute mti_svvh_generic_type of pipe_freq_scale_mode : constant is 1;
    attribute mti_svvh_generic_type of pipe_voltage_swing_control : constant is 1;
    attribute mti_svvh_generic_type of prbs_all_one_detect : constant is 1;
    attribute mti_svvh_generic_type of prbs_cid_pattern : constant is 1;
    attribute mti_svvh_generic_type of prbs_cid_pattern_length : constant is 1;
    attribute mti_svvh_generic_type of protocol_hint : constant is 1;
    attribute mti_svvh_generic_type of refclk_select : constant is 1;
    attribute mti_svvh_generic_type of reset_clock_output_during_digital_reset : constant is 1;
    attribute mti_svvh_generic_type of self_test_mode : constant is 1;
    attribute mti_svvh_generic_type of use_double_data_mode : constant is 1;
    attribute mti_svvh_generic_type of use_serializer_double_data_mode : constant is 1;
    attribute mti_svvh_generic_type of wr_clk_mux_select : constant is 1;
    attribute mti_svvh_generic_type of use_top_quad_as_mater : constant is 1;
    attribute mti_svvh_generic_type of dprio_width : constant is 1;
    attribute mti_svvh_generic_type of migrated_from_prev_family : constant is 1;
    attribute mti_svvh_generic_type of mph_fifo_xn_mapping : constant is 3;
    attribute mti_svvh_generic_type of MPHFIFO_INDEX : constant is 3;
    attribute mti_svvh_generic_type of MIQP_PHFIFO_INDEX : constant is 3;
    attribute mti_svvh_generic_type of DPRIO_CHANNEL_INTERFACE_BIT : constant is 1;
end stratixiv_hssi_tx_pcs;
