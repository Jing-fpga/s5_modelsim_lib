`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p8ii4JxUXZQ2IEn1PdwLivTl4o0N5UsKMkdYO4R0fe5WA5NPzvVPZImLvDajIsEx
mJ3k1DAuw5XBkl/k//Q4TK8u//3R78NLJGRjlKLSBulA3LNlJOuKFxc1F0CRiBCs
xY3EjEa6OnT/Rs195ZAkZAHXstGvfB49Qq6Nh/0VOUPnnm1tD2jY6IEWIZCCFBmx
Lq9tVkkKzfNx4UEbg6Vt8nHI3oVvtV7np3CHJrJ4eVs9qgkar6mbw3zNIDzWLdlT
J7oiIu7dfDcZcJP+5xjMQBBfSSLpfdsyUF47BeaJ/J0XXsfS3a5tJaM6e2KGsDyY
06KURjdIr8HFDId/2zQEDJp0coHLg0ykr1r0AuQIME2kGekC4heJK9AtkCE4bFRb
FuRKa9u5OeHhNtOI6OVv8BX7DKCRYulYHOffL/eIzzLBtWhfpMgLIOBVh5D4Uuty
6JMJctW+aqisZJJjJJ9kj9UiW80phEKOwTmgqIWfnIm8p16LTD6pmGiXuHBZ71gX
vCKTO7mZgR0nxavIhA0eNU8LgD+iQY5aG6UUnhlklIg3MKCGKL4lYNdwzjV2DifV
jISSvxaHIVzWyql8Bs9KgoU3bOmhBAHv0DzEQl7+Yg2/pmox0PifNhtpq12Q+c3D
1c62kWJ0TLjtW8thuzSi0Q9IKqCiNiz2nyl0TYosP5nMEuGIvCf5X5fs5RR1Ufjd
zWMgz6eGY3B6wvqzcI4XjkY4BWeZ1A+zshK7nvIzoejnM6N0Ndt5xakKsERCr3S1
p7cfvhd6wNkqBLHUoR4/QuyE6wyeA/LlGNogPszc2F0nzm8AoO6ROZ7bV7FpayVb
Au6Ev5DSxeb/7cFxeN8xBLRoaGIsUd5t9nT8J4dpe1CcAfk6gd9GLtH9NfmsOXko
2+yHGO3Xw0rgUlNnst32OqzlORgLhhf588QhOK4lEH722cD1pM90YXkrzjhXTUg8
v5RVDL0wTkEMQHoIRi4lSACjEgM5yESCFAcSs/Nm1FqAGN4V5UP/IOb5N1RIuEg8
PkbeGqgQf/8s412N9lVgUUWj8RVZ+prua+InTXylJR7ivd3NwlfJHDpvK+v+NAGi
bN2RqLwCa4Nsut6ZS8OQD0SJOOljHxeDlYuiI6sYb8GW06Qzb6KhShbohGX3fsKX
G0aHXyjwnRyKYTKkK0FEkeHVdTnW6SlrK/Gw1X5aybqQyLlLFqgTX816uzOQCaum
m83k1fHMsixXwK062oBVBvqya93uAjkab3OE33a5eEXkD9+UnjFyCGYVT+Wnf0xz
lnyrx3eTxav8sPtRueBllWcfHs++cNLCqL5/8o5Prpj4LDSfQbjzdUs6ag3ciLXo
0w8vGTxoHKXy8Prfad7d0IY/Uv3bMWjOpVx4YOgvO6Gyb+UIL0JU/nP/Ri7uCNWg
KYjwH6CJhfTa0M1HUMikHHnuHFjNgp4R5qhdSI7Hh5YHE41dbp66NiUxfJ+pZdj6
Ey73XGPxokOqBHnyH3bUJfZvZvBozCZ88mUR1GMlk1ESYCzEBsYYNKab7y2Trr7D
xcRoDQJ5cz3zUYnxPJYk51HHzzUUYkBc5l23j5aFD1nY7dD325O3A7W/GckhDzTI
VQHWHr0lAT8Dw9234FnXa0aC2wROBX6v3dsNUYEKx1ywNUI2zv/dO4ESUdou+zKz
CAEJ7q0l/J102o7H2sq+IqrwvI2YcOnM216/W4vboOc8PqQM4J9e6R5pR4YpqZRM
itGzpsFlxTWOWTLWd3MGtntSV35nQUOTwz+/tYfNWcN4l4Ips0ttWTTlgFwEUFEG
L30uW8PGHyX6OOt+aMzyTE99lSd+NLNM3biyTCv4lD3Y96OT2EaJ9LTR8NCIe8nU
buhp2VPsbPoFynsUGpJOJsr1ie3WaAEUt9PIfwhTlCgd+c9fxHQm8Z6AYZ682k3k
Yv4qGpJuVl9nE8u/FuRgEw==
`protect END_PROTECTED
