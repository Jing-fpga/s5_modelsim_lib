`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1aG0MjxPmD2mTuMCGvl6lwJJni9dyJSUG4IsMqOVNjVH3P45jSRUHTZRMTHpKePr
VomokZ/rGEWMj5wtJj+kvEK+wvvTJ5zhldDQfNpJPSeQY5o44H5v+r46rg1WHiF6
gN1jnoDUU4tAlN0xY9x48qGDUa84fjqzk6bJeEg3EKpsOVMtOWlNKoyKQmGR0nBP
sr1cZNrEYKxCCUeaZRlnMCWW0lQ7eXj4yemunIwit2Hgi2cDwuuePSXUM6jJ0U6A
U7OzoZEOiUv8SyXHVCjZER+pARNNP3vI63yQFNjezEU+lSSHE+BmtgivAj1r6v4r
lTtk1vfMRaebOUYweTzH+MyblAnGyfrxsbbOxD4/fzA=
`protect END_PROTECTED
