`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PguEFi6vcbznhFy4Dy6V0cde62zLR3yMYih/k8qApQNpf3WYeiZHsBg5MWmgc7TP
1L/Psepb+Z02W4/j985GYM159qsFgyoJ1MxZCl7hV4ouG2HdyHR6t8/wgwiRNvpQ
hu1bKKA6TBvfLpIzbFRO3Ayg30guq6VjwlD5ahR5azS3p1J6Y7gBBgubD1EZpE89
1UfOPaf5sFDOFP8YLqhdRmcadClEXRn9kQlEjCrq+y7F++r9v5uVT7N+xyriY93S
sceqx3egkD8O2l4v73y08ABCTD6DHGcRX2mFWsSZoCGGGYnU9IbqyUVjcgFx3b86
CY/4VdYrP4NomjkhSvMXcINVbSkPhVPpIAXIQ8et86GGR5CmB5EXHaiUS+4N3ur5
BzMAg+sf/7+l6Cde1QUgimBGy4vm544eXd3pmbfrFxE48qblka2B/kcpWUef6Cjb
MMSCJe/g06iiNbLsFbgsxX0CU7A57V+MfgemJ53xB7XkDRZDmeRN/YWzNwkLgIZa
bJWpHdmDHFQRtq62DVEfH+RnmRM024EGDlOIJZi8CjVEA8b0kXtyuYIoeGmcoGG5
EHly3oNfVIdrSZ/pERhJvKw+a2ZyKxso2Jd0S9PwTREA7t4qibPN8M7c0UBi8lOU
3Vw7RSSJKcioM+vevVsaJDS9G4tCMIMnlyHZ8XP6Qsb83UsGE0aM3h3lrPjQ2Mp9
OjggrfWzW4TKO0yU3pS59wbftJPEwpEJqy18DXxwHUpFzhJpKY9/Oi6MUi1ujK+E
O66DZAMFhFlQnAG43lXAO7jBgUFETXgfxZZa/rirpsWINjY51gHIDZv5YFUd7CxM
pKMj//rTT3kYKfcrM9CU4W0vc0LrP99N6TjX+J+dlZT7lOSQs7zToI1OgXaBxCdw
A0btvNYXIGuG+msZdMt+im/eP/znkWTfqrYuoOHCepjf9TFJWfu+4tXdkupTF3lV
U5EiDEJlPkeDThVvHaYJOHcBh5MtxFyS/IX88EZLSZQbpJy9++Pgvho0c6cDYugX
GcesAna9/cOL9NoKxCenh8SSuOFCIh3QBReRoK5HeUisrF432PQZS17v5Cjh4e/p
FnAdqyZXS9yrg+38VNybuZu7KKtAkd8xDLY9k2sNtFxcstQ+QREKPZ2Uw9sjiiiE
BJnQM3DvSUG4vRDFooah0g==
`protect END_PROTECTED
