`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ch/j/vjQmcYZi7HN8fbyLbz+CJWlYC5UBjo/DcMZIcDHB4+Z00B1Ca5HkJsb4PII
bni0ZbpzRbZ8M6fsd2Xr/KofNBhmRk5eQIFPu+9AOCQeAhlrgDBWk9Zs7+N9TbeB
QXOIczpcwokYQRKIvXe6bt35tSWzQzpAALUO+R5sPEpmu9h1h+R7B3SbLhBmTDRl
bxkBmOcvAdN2CvmcmOMjD9Qd/LexQRNLGSMA3SDRPgqvahbweWxWUao1tLPSqsoT
VDvxtiS0TLbSr/K1YiqxTpZMcCzZGrysMfGNIDtROvBJ/jWdrKLnNGSbeNxlTbdI
txEjjifiApp68hc4WzXoZHUE5S4wLNe34DPZdTcQnU00+TJg7N1sk+Pa0+38GhPE
zEjcdsWthsw3GAowenl+wGV5yzsgphMDJF5jv1gzQxY=
`protect END_PROTECTED
