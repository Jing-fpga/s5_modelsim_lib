`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DY0QzQ1Vnj5w9v5V6kCfggD9nEyvc1zReuRJOJC558/MddRllhtT/R6Hm2gfE8kT
RA/ehzpefgJd2jKRoG7J5Hy78lNujbRnB3vmmt5PxSXreS562TV+yk+SChzS2807
APUJNihZEXz2v9avczGVAAJQ6zI/Sl21UuN4q3uc97/+oL1zvYmV+47dGQuPaVFU
K5R7+j5myyv/nO/2j8cijkpBnvJIKxjHnWkAepfHvU8FrkFmylkbqLTMrbsWpAbE
M6uW+vBexWaie9XrDFQQPBMk7ji2M9g0i7mH8l14pvBnuAs8qnzA2Sd00XHqKVgh
WZMwFiOVdc+zeYdLpuOcm3wW1tau88Ptw/gSKdD7+rGJ/at+TtiDYQLAlqQI6sGW
nFVUlc8QcdbvxvDkycaOr349QIdz6kanIpgmzFHsZRuqwhy7gD7VlpxOUbr90AK8
0CHFwIlolKQdlYmptTmo4AU3x4dXiYxXPx/dVdlVjZk4o034CB6Po5/QzDfF42wY
vsaXbUxWMCn0psg760MHhaIWlCfY6Q0h53ccpHPeAWvdRRwzs6v6cBypew6yYVq7
f7AsXP/yW/RJ8VODTxHyZnvNV21QC7OPU4Al7PQ3nevkJQa7OLVnrMTqfoPMuPsj
d1yyF0dfJMEZE/hhok5oU8FRpMeiipVBHVS1L2lZ1kd0qmu2z0vBYIGL7LHoCZIV
AgDzB3WjPgAAKfW6dTWmiEeaIPeNpH3cqZPCAs6fCSkj9miIxjAXMbrZnueYnJ36
lqRVVWj2FQGBpt9m4gar+Y71VEO8bWt+pfFWw7yGatkCT5IRSoo2GNsaTAwDve4Y
jhYZ3pZHYmveWjXhATYVsY5lMVBkpL+4OXCF8Wkf5bl6q1bogDkP24TgJ/j/xp02
BpZwTKeuoreTFmUVxJM5+UV0fyzhUfqhoHTbExoQU7oaJ227CLl/hi38kOo2ZwW7
qRd/jt6DXOKFL3//t4KUxQprEqUW0lbm9MjHTkoRYsEYHa5hwZxvRLxBt5UuIVv1
SCGtWM77HvKw2YANNoZrkFyRiloizX5k8a9qBuRLtSpkoizDVpldGXGL5Ra6XEAC
U/auJDt72d+1sTzB6bjo1ivJ0X7VrnzQVrPQTiZ4cW+aQzm0lVwiLbzk0AWFfxmp
PJ6Zto0+kGNxDvMhkbL1b0dISHiZ4tuW/cv2eY1rilHwpgJ+eHLq1FhAk2LwbtLW
rhAfIvyzn2pde6f2FIfFJJa+caboeno508+BMMcRvdGoUg0/ostKN6cHlQU88pAs
5K2EH4D91q5yi1Q1x05u1nug/x7NOr1yzXPty7T6vyp21STXMWmm2O1qoEm82t/j
6A/OU4NvhG0qNsKa+wKDP0xssshusq7qauSQRez0LaKKcBnjlXzi/OgD/ABCpCF9
8fYMTWg0Kth0EO5QZK4EvqaUtOHkAN2YfV6qxYbJ37ah1w+jDY6Hip4mJeaz22wC
1wh3ZbQvLLqG725t5ieWf/69emoacv/whMW4z9vahWVTW+eh//RC0Srd5jILbv9z
+TbWbUV1sQ21P1B4mE3RlCICJTZh6626ZJciT1FxyIQ7+Muxb6Ps3IfAu3O9ADTZ
qOtmzkuON9AGtSibytUNOcBbKcRQ7N0i2eJs5hxbKpl41tSQerLYHsdGz6ISPP6t
efJsWFnBXi8SxTTujJK9eIUtFmqW05uh72y2Vn8B3qChohWXuRioYKB240ICrThI
5HnfgA0hMSiqLU8rMWom3m7iHCY9/MBc7NS+8n/jp0SWb8P2FDXROhhv3/gMgOWt
JTKR8XCPZ62kfMXc8DV/FQjlzrmJ1gxz5ht9z+mUjHvgJ3EN7DxZXUiZRXfdXq1P
Nq7Xwc8xRvxS1JJtM7fzi7DZZ5iVogaTeJZZL9THJ/IoFazDofuJJF1CVByc0qip
ajnfL7nN14lDVzdMzFgOCafExT2JzRhatayO47fo4M63OwndzN81rHrYEMKAIUO9
Rl+pm9p37yy4rj8RQRT3qtAEVg+WS9zlWZQu8PCjoThpwKSdZjnYhI02Cz68H+UR
E7SoDL24Nn5dU/QPncHfkrS/NZULKDtItytUsCQ6Yb2JJh6/M1NIb41sjkRkXvvo
a+Np4egnqSz3Q9YTdWBnBQgKjRkMgmfUlhxNXGwzzF7CAe6IDxmRYS45lq51TFXm
1Gu8eH3iwSFJg32BgPCUAgDx2EFRghJDB4p2SSqbuQWTtKQ3NE/dS5t1O9lQaPtS
iUSBZTqmCfJTQx2iJ7fTnoEzT8rWWFAhg6UAI2PeWxRFYQGpZrWPIR9MzzlUm2+2
66nwJ7SWBQfGD0b/Gja+G3pdr1wneKtYsjlp7q8nV2wVfESJTyoDk5zrObkZPQW7
TUerykNHwNqkpxdETrvEXA1UDm5G1QsRA0Mzi6k3SW19gX3FktmcFgbb6LrKQfNH
4NvtiRCr9LXvGI8mDaKAyc2TZz8pLaTehFp0IPgInzH0JKyLy48fUufFVpmvtABs
UtwJ+pAtx598cIv7PMG8+GjpvQqg3NuUAHVVLRM2qjxhFBXmKdbyRAoqoE7uy4aC
QXX5h/efrjbSepbucgusEgRtVpYpCG8hUusHpMJLsgVJaySuLTpx+xIoXE64fbpG
HYaGGy52rzegrC2bc7m7C+Dgd+etLQjz4/1kORJKH1bwscNmJ2APlhushAW9IOzw
0ZKvGTe+Wduyc2UltDwvE4LwjOQEld+RhYvVJ56IVYslUPIk8OHBHkmme3p21ZVw
PrWD/Re1BkSZZQrXzPGKmxAIh8+Ulnk00wOssdHPyB9O8ip4rendIYtqZNex+q/4
1EGx5B9MtQ9BYy3ob8PTwkFTFJdmP58V1Zh69RCYVD+a34sQnZ8IO5L7zGsW9UuG
zDRi3Nxhx8Go7Q37mUReyKjOFgHsSrlXgPcXZC6XF/YFX7aB7A2492bnDJxTpxm0
82nX5HbXAmZprCYMFsr2Uu/9qcv+Z6u90/+pvB/z5tIFHDvxlM9gH13syY4zCoCw
qBc/xQJ0iGfgTyC9MZjtpMMfgGb822bcV8cbHEvoy/r/RQ69rSEqFl1olgEQl/iO
MyPwAj6LJFYZ5Kc3vTdef8SSwQrhLw/Qx0SvMtq5uvs5SogJMatqfq+4MP9VdpS5
TfxySFS9BP/VyPIhUZj+d75w04UYGfZUOGcDikDH7SFyxgJX/D1EI+g3HJeqU8mK
uy+wcK+mFPIGk2jDXpClqmBChl/FHAz9e+tYdb+DDKE3DWxa7xA6lsyCN8DssJ3e
hVtrQMwL8r8w13jitf8sbmGBUBoYuFTobHISgQhEYAlUB89fJXqfGv0+ULuw+w+q
7BaLQWotOPpUnaSbNrGnNL8QM8kZC8bqBtJVBp2R7XjKY0ro4gnD9ug2Nuev84pc
4pjO40nUneX8vUUDoqjsvI5cwD0UwbUMvxi0Dkd809VX8xHRjbrCLjF4uZwUxiem
azxX7uXNNH4okck8BUVQYACK+3bVJQ3T1Kl9T/qxcVUhEJLKIGKQiO2jLzkwcR8x
eN2G24CVj25u0+G6A5q/9jbqj1HTPtzjBn70IuD1A6LzKRKABA4plKjR3De1z497
xFfOhyfPnervqIiKKo8Zyxj5az16MDdlKCU1UIg5ve7EEnl2tJUUiXPo/d4T4BiW
POh/HtvJojT1Zsocoz9j9cMr3p3iSbyjTCCxxD1b8pJcGRYrJbYjuQHYySrZPeMV
m7Z90CMOJG3S/+9XXvr69TrdXGFFbGhRSmCHh4kHT+XJC2DVRFDnrlkKk9kWw9KZ
dj0HHFpQEssgvE+9DEuKnXHNx98TDQ8QkeR7Ip2GhD58ZjpRenrgs4KOlFBahR9S
7ju+EQtyR+n5njX1wyQnvJ6DwVSknAzpwgkMu2RIdBRY+K2RiV8qsfkoNBXmH+bk
aBcyoydsZ3p9kdY59MeiqnQ3pNQgV1mw+PcZv/06DjRp6PqI+E3DCCLFEfOGuVqD
zRBsifBfc4RJWdmML+CbdnLEauQTxFCSXg3jxKtdbk9pXDVIuIM37oFABUSCjxDE
WN+FjJ4zKxCAP4n9rPwq4p3s/STiyzKEKDRezQ5Z5T1NgUCoj5ezZgrBfD4p4JlN
Iuy0nZGMnXZJKqnetmNaz5lEMYEjbrYqxVHzPsrRVVP7Sql6pjiT7qVrX95F7glH
7b13/JO7FCRuLLtO6/l9x4c0g3PBuqFWIYNIQ9XrJaJwW/9l3HjKcbINOOFwYuoZ
p5Ed1Imh3QjxM8lbYiJmugbzQHrfWJPxJJS/bBn0egl+9d0gA5OeuiLe7oLztJba
/Gi49Zus4kCsevDq5KHRH+vNw3SRfOJEdXN+pfVDgtdw3B923rZJt4obEH0LcvBy
1KizMNzuz9wbfyKrvQLQmdtnv+59G7G/paVSfh5rirEGPJCHdKzYboiJhvoKCvSe
Ncee+9JnNmNoqW/TsFupf3BfduZLaJThrRqSBm8GGbbgHoJqpgFq4pf92Q82iGNS
OBR5hh4rzD3xlPKk1fX7HcboZsK6hF2m1dbDopICAC7mG4DEF4GdPMc3o+g1w84N
kVax39x9Ttl1qjrQzE8zJkt5v93i8SJaR/ue+rjY0KeVNZISNzJQK2GVJcRUMm6o
EtN/5qigmhR7er8zz2lGtfKvbZ6vvXV//jQ+XHuIxWcGvjonO/+dbeu6hxXJtcRw
OoHN8apil/wBMTVy2OGSVPWXCzKkkZPF2b/x3TLlNmWf40gpDUvT3hB94IZ5rYn3
wKZ4MJ3VE0lRlTjmPmvhA5nUtEVTDnSWV2FdQnqrTmp27ljxW0RIAdDT/WK+Fy6y
rkSXfS439a0ROs4VpgUJwbCiafhpdq2pF7nCy5CH/oEr3tNH6byGJz2geYuDYAtX
SoSt+37hBaFUeAANqDk2GqGd8irFafvWmf5++a4xYNYE35ZfvVz3d0M4LSPyhNiY
OOZJ13rp66B/YxD0NstJD0hURBRP26um8E+N3+eN1eG84Pt3PxNbo8GxFQ3eGmll
qShqZ4UrhFPoJvvlCGL4K/e1yXj0IynQoTqBF41lRAowREhA8cBaug/AXt/E7K5b
WcSMVsiKYQpeDBMQzrBxsG/mI26R2lqzKbXxUGqk64umhXf7fpVel/1TfWUwOzHe
R4gl0a9JRoTzdO6HsAdweNWlEY8OERYffd2sXUScCF5uVelhzn+4ZxmatREyNynp
nprUgcPkNwxdBZvzj0rZfiTGuJwYFMC14oOS4VwyVtwtT+vYui0ZQ88gLEMscRxp
b0DxrOL8RMI9M7qlLCLoGl5/y17Rq/ZdtriGZUhGQp57KE1IZzWAFCS299VuoZtM
jWtQfoJh1TK6Slh1Tt26LLA8QtXzD9EmwTQCC7sm4V7hXYyIt4rj+J9fvzSp/kGU
RkJ75Epmj3k5TcE6juBCmn4X6jGYC89EJa3a6T79nDJksES1RkPEXubo52I/pTMB
NbgRb0RqKsWWpsy4iul8uXA4qQinN81TZ7N6a6SguVkIlpXxG1GfpyhqCwfD1NsQ
jVYAZwG1lXpQ3RJJj3rhcHFKBFi5SGUJ4lP20XEwSANG+fnG26+LMJonmx++J9xf
c7ITqaQyVqICUVLSk3SFbAGAr+UMQ+GxKbOk1xdv7fHstzHIgeMoLooEnMOJuGO/
NuZGD4M5aMGe2R6L8gzkxsVjrB+vD3140ZlLjLGu4WNJd9gVVM9dCmkQLwfjS/oH
tqUe7ep6AKNLbeTnBrwj91vM3I5Tn33CNiHrItU0lvfJVYk2yJWXRBle83Zr6/ZZ
xf5Q+Q4YlzW8tcu1mN5+GGKBosDROtcGPHFRu3+pbM1IHo/UMwWDSjShw3LKB6dj
y19zb0U7t0jwrm+NMhxd8LL9N+77+ex4Z3qjWvv5NgHxWudazJrQHk0ZLVTHiaUv
q+YPG4FRZWTv/Qt94Y+FqKRoiDE3P3nr44sfSN358QsL+x8eIn6VyXUzRVg0hceA
ZHcRCH4AR+8cYpluDFegsZpdcTEGXXa2ZGfHBAU/4RrLQwdXonWHUNJwyp+lUcc4
6yh41vfGBPuiX9bdSbSlcGMggolWfLYwH8oQf2+cZMwfLD5dvwGN27JQN/F5K7MM
6a86DxulGziXmDpbEl+UApFNu+vWoJ7Rqg6Bx/d4wc9bVWEC2HbWxc1k2pGgssTa
CHJqXM1yUREufpREc5KJwpBusrL2MhkKG/bBGQxXM9Bv5JYm8Cr7BRFcpbXv7Ea4
kGMbQ1TQxIhuLMzLnvUpDe+B6PMQNqQuz7QIJjB6GqdQkrDiEiOWfbaaIY8h4tWJ
nu2dtld5lIWTxlV8XrIm6GdYmHAfBmFNRPfL0KXNnNNmiJqFrD9mQZGoq913eOP9
FZUklARd7D5eZt1gL6MEp1bKtkoXYyALQ3oUI5Xrl/koagI4+9glKx8RrmjthAj+
im2ITdAz6USTPfZPeiADUi75EVSj3PbB3VQP/YJaIYTnD1pAipRzixkFDz7HTwH+
0EkwF01/+DqSLoN5etnM3Bu2hEV8NL+/LES/vUgLEcZv835ghvJUvLn2JT1HYBXS
jkvwzjWQ9qw45aMiaKHrGtLjQfrT54MHJckwBPUGJkMLNt2APgXarD6Y/o+v8AQu
1HdJzxF0vyjaUGTHQ+k3Jzr3bTTpBIB7VrWteU2gagJoGUEIBlu51RE81iS69WRp
7KfbxvkZfFEEYIX8l3XTQyEpgMi9e9Vcg2jxSO9NGYr8EsOtJSqXSV8VBxn3y1FA
PVWZXntGCEsS4WIljQegJLqMTw6bCRbR37ocgVch+IHXn1YnLbh0lvwzjvNn11u6
JgnBxtc15IJzWBFU6bIYQlwZJ9q84dUrjD6GRADZcWFLE0n3ehVn5uzQm3aJJFFC
8iEuvLJGMvXzjxEagLMGkSUyNABbV6mhYmoZyFGxl0hR13l7a8N/crq98AOrx2q+
X/a5DqQgRp6RTPdqq2Pp5geSII1FD4k37SUmrLUEb4d8d2YaSRcce/jaTvkiWDdo
ot/HyQu4E1wQozwAcynvdkvUlXP/NvhW3aEeqQOx0wXJ3KVw5A3xmF2hN4JAFuvQ
pbyHST4gw1c4cMUx1ZSisSl2BOPKKOjJOIU1pyWngvUWiuAjwNw/z+c/jcyAuwMl
2Hv6ntf30rrST6nIJOEhkqW3kbZp6mA9p/aDjmURzbRN8l6n619RdBExbbulXTOl
/nVRtZR2lXSia8SLxbkBHA+q3+U4Omk6XFnf3fyKoPYnYBJJjoKh+fRt0H9o+2p9
6Vwrh1ATjkAduc8ED2U6I1/ShhT0I6Qxqmjfn0/SM7yz3g7P9dFcrRKelvv1JaXL
1TGew6fFsTF5oyyqmiV4RfZ71lFOqQ8EdqKu6dS+50en2iEAaCr3tuIO869rSTY1
znkNHSIbsPMiizGC1Yedm63gCNQjyD5Ghm4aPYYU6OvX0T2K4207WDwEQporCdzJ
m6NVwrIzbCwXC7iVH2ziKhcG3+o4iPNVYkkr57JF13Pwuru2WOzfFIqLLU9LA7CC
wSEZ8MT0GnfhmBHNnnJNRaRZIbEN2G1AIbvfNNNZjCVoa7BqU1Xk+CzGJlBy3k/p
zP7VeoglTajKcyh088I6FHI9+O0R4jNQiMgZUDnK5sRyTAnsSqPmPrsV/Q4dM+op
Bt/esa1sd8HTGQUNP+uA34Ssa+QmlysfXRjoCW7viZ82Ls3WcZu+v4+vDfHG4mD+
9J2sFJWTKl021PwfaXkOYFYFrk+fENriXdh44jh1LSErcRbHZPg+AYG28bQ0Igpa
vleW/ExKA5M9c9v8I1jqrZCyTcw1W+5jkNRZ5+MZPZxl51SVxjNXYh2MKK6EkBIL
8nwd/FOYEp7YTM/PqvTI9cYlM53t1B9fSpUVCB198oFt818sX0wHZbkcQAEhLpTA
96GLwtem7OAVo5WfdwgI/kn6TXLkPEse23VqVl9Kn+F9038HY0Lc/x08wOc2POmH
pp1kZWp3Iodf106Tp6pl+y1NszI1pdEi0xDPsP3+v8mYWQl2mf5myx8Vft6UYZhV
7YdrXH/eehRntamlqcqL+pGgbodUxOhhkjErXnFeSCQI4S8L4Q5jhBeM9J43Q6Pc
XcgPtIT196OJgF63MjjMqoQePXYd6/nHH5nn0pQpDTCMue6ZljXWvr5lGDqPW++8
z6jVlyJORd45D5uJAmtpWEvOrHXPAO1nMOdPpWCLHtFN0XrDp1MaaK/05ofBspWl
5EKs8qUNQPAlcddIU+Gy1CWhPKqGg9J+cfPnd0dyr1jDEJ8W0lGZqqfFW9G8M7Ri
SSlfDjjWY/dtCP1fl50GjELmV4EOeliRPGdI0byKiG3RfJCi/Qswzl8i+YOzZSez
rr7CJM/TcV6dODHn3qX4c700wL/QEMcrARGghHJ+/dt9w+8f0XNBgo9Od1ef1n6q
u/ofTsto4pfR2SrIfEMCbLpxznemeZ9+azYRhm+M5C82lr4vUBIsFQjnMYLcDJ9n
kSwBVa4ogdReuQoqA6t4awN1Qmz/M1En8TYmbNT4+BMfTwBpWTMVE7wnpFrx89uQ
KapDee0jL0P0eQBarTb0EegFZj0hSxrfY48nWx9n6ckULaSGELbdAbQQ7YIjOmA8
VkYbzF//xoFppHSxsUsUNlQSrt8Dv8I9Lh/y3Npf/tsiHeGHXPXmBoEG+R0mD3wb
tInUA/Fcz+mfNdUwCXWVMxw+34e1/NMUUpXFxxMV4GJdBEiyLabVms9KCHsOp16L
/eWh72uyVKTtvITWcZuQVL9wklnkcJuz2F9bwHWcuc3+YxeHtneg5VwjWhautynn
nxCVHFID1QSWA6qLQQYlTTjRNaiQpBCBrwekvW9GaRRvvC6YgA6X0TjNAsjkeibj
xTtUHnkKT7LnKRAv0ng9s3hEPU1cejd5RCB9Lop+RzhA6UgUsonxYi4I+u9rIPWe
QRrZQTdm4XXdDFej+d9c6gE+9SxnGocIFJnsmBmwzr2NCSaOCeecO4rNpD6vfuIF
N/wwCXqmMze2tHy3sq1/1kOeuXHXMxHFORvtHvbNnWgn4Rov/Bmj9bdsjuqizcU4
nfi+NuYcKqeN/RPP0+hmeohd6mC4g+YigKshA7kKegTJ8+71v4pWnMTEfalvSF5l
nJHzaENH0InlL2Bq9n7qLTyBrdZW+RwczroReUyf6i7YUMLy9FNYAKxmgiN7l1DJ
MhWW6xin4xcjYJvEnf9ZawfXE/mCj7STjLfaKzj2mBdhACUA8aFzKlXsMvdDbnVQ
ZIMTx+4254uf+bTMliTZtu9s0F7CIO1/lONnWmXPGA+JfjY1vx3w1ZI04wtUCCVZ
xF3eP+RgrjAJbBgdfqMNYF32I+pTAyg/xP8E50LBb6rI3P24QrS4NYxMst38G1ob
Vs/ReK0mbcKv1kPtYklAGqH0aUuZ6HltPe2/H+O/xmptWIX8/vhdUIPPi6DOtqxJ
OYLLO5iNQAQ8ugJ+s04xtZlmFNSlyCs8G0l8gTgD8cdEUd7FA8K2Vx1dft9TerKR
Eme5H2J6JlAaxSqFc1cLlm2a8rHJZBCQKoQggvP3UGQvACc4SHef/ePvmwX0C+vH
uckAJa+yuNhai/4Swzc1kB1GlcVh0w81uz+ZxN04Q8SyWgSnL4yK5Snocm0RLTvP
SAkaNxb88h+mX+nANnLTIUbFuDf+0VW4P0IleUDaY0zXzjW+UhnB7P9QP7T8pVfQ
2dfHPARCJNoghzNeG2wLXeV7vwQ5HfnhVUShaZvtOw0=
`protect END_PROTECTED
