`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y8ttCY0U5B/8mPtgTPLUofQalc72q3qoWgu1zowjc89hZdrdQZrelb36u08pYgtS
oy3bXA0ax8ATm0aW1cgK9aPbDfn6EHQAr6kW323VUhq2mJLr349AeGgFtUrqXE1D
+pJJFGJBBqGAKZ9FgPeivoV3bX53Uy4Y547A+3INru9s8456M3K0V8mrPn+TIfjX
Bi8nfHeZPBdbASuNO+mnG/TtWOtis6mvcQDFWfvnhYq9qbnkQ0jOYCyA/508eboI
Ur1yyCXmmMmeAeaNUzW6MtAfuQtsWgVXffoOcmVr5Ga/zluGB4P5QTfLq9HKKvrt
iTjypLjWKDIDwaMuqi0BUiqECfBvEqudblXU4hjap16Cpb7JP0fe/pb945Jt036V
YuvPvD4lUors8g9cKktakQxhBsIoXBgOFuUA8pAHV1agU1tpumhf65n2ppknJmsW
+WCrHg0XyRBLEZk7vn5SJ2lXcS0Mk9brjw8tyEwiSvpZ5epmhzgoxtvtI+YRin3M
umwRByWVE+5HuMalGwNmGEWH9Hektv3wswKuNBc4mt4FkXbwfCSUQBLGmKBz2jI3
aFwt73xSSQ2A9D3VA8vs4nS9fq69lu8pm+HE5yIHRXVuQB0ONAOa38lX1CypKkXG
bvD69SYr8KuUwFuAfy4Vm1HPdXJxIn2pz7zL2n+Bwj69shvzFXaNaXSuhZFkhvcd
Oh8WA2qBKtRMuKC+yxDSENKK5nvbGJ3O6FmlbJMa0IZn5iC48tTKcBfN74sudZs0
ayP8hn0JUCNZuOvkaThkMoshcUQNLe+lx857QZHuNhxESUQxlzKbSOBedfeaSaON
jtny/L18PmNdkNbkGyCobVDwlBJrD2yTI6x5m6MPEeVYDcJWju1UszwAgid3u7C2
L6q30YZUJNmjr+U0iM2nKxgs+Hpy48xGxIPRGOm+hya4XxQUWJ2ZvJssL1vo0Rmb
o+bf+q9RH0IJvmXtxTYFfjqfekN8DjIX6SmBNOPccQs4M8cHMEOJ4XqbNWWtIuov
Fur7MuAGUXPRE6YG0jeja3bAFiiIsyvNNhirW+6NgHa/e30RHyucKgGSUE0cMLbY
XCM1YyutbRCdXfXNO+Eyr7qdyRadK1eoQmEcH3RdO7aKDwmNCfGo3hDvCVfdTzxL
bMCaG+aX0TJ0Qxg0hdsfa4jz7it8bHfwL3P2ZL9aD3SvtZhRVIWZLg9K0POFaDv8
Kdqoh8o0iJ/dq8x/lrB0Y4yBnp7MOmTiblLwzYaNjCYT1TZUmsW4D9TIfADE9E3w
5V+aQGWioGgBjEd8iOTbXHhOaw3y8heepVuYVVYl+CqlpCOrJWjMTo5zHBwIxltp
ZbX9yP/sp3YIpmyRNYszqkkJVVoGymrvKxj16pDLU3HO1lLuonjixedG9RuIDj4w
me3aG7PRs0GfY3ZhW44Cmblia09VdfKAuEFUrESTN3EcE4mXhO0JfJ1djELz/d6d
kf+jM3WHygHvEkJqtQelSYvebuUO84p3CmIGpAqG/crRxvjn5LX4beSYD7bM9oXw
iKM5zXRdgLzPffGCnb4KgSx0VFvvJ19S4a48b9lvtS0D97cRgs/+thcKHpXGrKV3
ZSbCbb9oJAnft1Qvw8mspuNsfqMrLwEOj1FXx0v0lscW+qx9DFGDhPP/DIr+Mkxy
bxRIIRTCyR+w/rqX2xTvUGW+jKpNYEUi8HyavbN6BETza6orDJlaI0Rg5C/oLBxD
k93173qwL5xyxkLHweoRi3vumairqBMsUXU/WLSbMfSwmjyxYDpCSllI49nPw/HK
rhFQV1zxb5rxANsD17obJcc5snALwpTG3I0n1nsKGon0qoSLnSH+E/NR20dwk4cD
Qv9VMtcQfxDUZEykIgdXsiiOft99Jw03MAvSo9dgPmUw0hbLPUJNTDoZZUtDhYAk
RZBq5EVtXJtaO7poq5/TUiZWDlb0eroLFex6iqumUa3FSd8JHlfngCviorfHTfzT
jxj2S6n/vEGWATdw+jNmnYNaC2vuMABO+ZF29tv3W4AjAhcW0e+YxOhKw7lild8a
24mxOfbRVKLg2oRp4Y/BDVt6i2udc31Z5Tu7ICLa4bQ48lAAqLV88Tq0RqyDytT4
z43XDN84hdKDFZzf8pPBSxx4DvMvHBkx0P68hvc2tnLimw1JEeTqhrOh48g3UI8a
+EqYxqD36phMVIij4MXV2X8U5cMiUI3ExUzc1E65PCOzHkkEItassWXiHwGpr+eO
pDqpORVLBijPLPY7QiTYafz7sfllJT/2as9Z6qVPA13UodflKy4UTUgDCupztLvu
uoHbEkBamY7yjWfll5M9U24M0Paimv8k6MBheHjnqUB0WZB/YpqKF4YuG/WPie6H
8Iw5Ws9DGuykM6WShSkf90h+NiT46MtfLL3RIc246tC4MtI2Kf0Q7dn0vSyj0D5e
7G7B9C9sG/X41RCoP+xmfFyXv6tj3tOBLvOwIYROMIg7WNJTgcKLljWilm+cMBNF
bacviJVYQnwF5qxolovt7BQRvdDvfIezh01/wlzpNt47TSQiCPIOcTZDueBI6mx0
YpIkIGBB0JwPaH1BEuWwXp5AFdtXa7X1//axuPu9xB2AF1Gb7eUmVFtmu0bPo4Dm
DWW0i9tzGIm8wmuxSeOkWNFAGrwylROD9X68AnynLdRJdpTIzlCYVYrdRa8qk4Fb
NXPjfuyodfK9Wa9Trpfgf0dWh7HbMRwO9vukmyn+0l0lYMtANtMrF8A5FYrB0Vnk
ZXPjhBW3EMeQe6vbZ9D1i0GE6fqY0e9mqZYQU6DcLuxKtBsQr16ILwjhch9kKpeH
L3cwDBHorAHyqsJvXSUgpUWFGftwadDQCEfrA/XdkoWqlH1jBlSOUy0d2LR4XJr1
uvkXUWUJ79fesVaGt9VzFU3jcNCgPpkj2Ip7XkWCavDBBxBxkg2omLvdQnF8xx4V
PCzztz7L5aLvbsBuzmBnAvAqm0VXhSkeSQziTwEb4Cd1qKlpb/13zMeimesBiEQ4
Nr+NPGTmyJZOMly7d9FGqYNzj/OCtFeuAyZRnxJwU9YPaRtN+LJxZB/gvzW/Opxq
mg0r9CkjOyz1FzWn+OLoOjX9V5VaVRdRWn8TlPfq+FmU4mlvuITTxoW3ERTNP3+0
2/t9UROR35AaYne9Z/1xaLxkNgJ3gXfyNqseyT29QnJCkbJBXpNmUIp7XItdlsI2
LAwoLhjvfkphwHoJRfmV7RhtS3q/hDxe9Hn+QMVnVPFL3U4Q5AwVXditFga/Pecj
igDAVm3d3yQKZzJpcnFW8oaCyF/4MkSyD+JINh2fiVCtE2bZ5GBXA1XvXx8cAXq+
9aTMriJHAkU+62TPhRiORACjeXIiESegMLlkZkJEqawCBbAyINSh3UHKXkvB8Yqp
ubhT4qJJV0VCeZ5zfwQALlklk33qUMhHJp/raYPkl59nhajXYhazHoTxIYH7I7YJ
rxlgth7W89oKdPH9l36RE1lZrZ80NpRC7SBoy6KR5jPbkLa9iKnUhAnB2m5+PrOI
3Y59XGO4buWddc/h057W1hBtM5Y2DGAQ3TkK5K4gCjxPzKR+qi4XdpkU1dQgQaaX
mGti8qhEC0WAcVTn2kuhZZO2rEiGiOZZHj9A2ubf3LwzjnvfLQnTPFzWRnx7GKAL
FTb6eAnnKQi3kc18VKR3V3COV1aCI2S6h8TZzgNTZC0Vv5LihA16RjNvhpWBghDf
N93cUhru7zf5s1Nh6cD+yJx9Ctil2uiLrsBktssccE+wZ2ZzjWNLLCyirWNo+k5C
GYQjO+OFoiGIt31QLm7XYpKoikTCDjJwCEKO/x9/+m657Sh57ds0IwSxvoSyv03P
dsOJuFJZg/u+nYBONoCkySWqJgdTGbujjI22ARbAc2sfvrb4qttjZnZhIWSG8sLq
IuUMwsucOqo6taqOm3o9Gef8HLwCuKSx2KQxlqk11sAVDHqbYzJIFZmas4N4ZL7Q
gRRimqWtg05EWZTGZLV/HPYM3+hF9TSCKcH1/OquRP/tjeyjv46STAowKQOXcABq
QDkXkO8lqo8bX45Ef1lCFxLPL2C89LEAWm2JhwU7VJOrAxJfbgacfaFelXAoGzgc
OEgBNbEM66XozUstSiiXkSPGReTBBB7OxijMRYRFt9/kSNnLiJf8wgZ1q8uJG5/b
SZUFR2nb4VI8a/eJsnWNjrTfAM/1wmKkGcD+8ZTNOowb24wVMWvGVLky1hbZTYyb
nxGDvs44a6deUDgSyZ161tjj7r5YxeceahJ+IjIZzCU7dj5bbYEva59dLyn+iL3g
RGXjA3JDH8bipip3Qu8OVbT9hyrUbCHEAQ9p6CzSbxQLgZBk6yjUantikTlVnOYC
a2wdwt8XYVXwL44AxU9C/rLn5GWcSi3XPXaAkRVNLFFclqOBKYlogF0k4qR4fT42
m11xWKcieY8QhqlMniKmNg9Oi4BFYvALcWhTfkwLyVOBaIABQyDsPL9XcWjRk7X4
GoBWIknEDijR9MxGkVpbtPmwBjflAekuay87y+j9jv+HZv5/6O/+UpSrXIKawV5M
x6OzHk4sK0sb4NGZ/4xLYI4c4Cb1ECVhCCNRwSvpM6Oq+vAAGlsej0V8RhG09FRy
4zC/cNNPqdSVG+heV2bYWwSFxIqf7uEdyBVgUh5q0xQ=
`protect END_PROTECTED
