`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kvkC6GaT6riMoGzdA93NWtChKDx1u7rFsIqBNbTNzRBu2wa1/ixhxvOhitS5Q6xz
l8383kjtV1Srq3Pqqk4NF+nDg2sshUU7yHNheOPPR7HEXFxC34GMzaYVLCKM7W1M
u3qJkBrO2UUScIGriBZfKPVrrBBbVgVmOWif0Mm0nhnAw9eqjzOFYAZSTNYkvZnr
SlBNNkK0G8dl+PNhVFq/RLF2e6xbx0mKYaYgmNuB1MieqPc5ytofimvEW+PtiBAh
4syU6+BFf+jJKRD6C+s46dTpwKw/Qy5ymz2UZ3A/45Tudqg2SbmtMxC8/9iH1Vll
2wwO3NDrwU/jp/MzrWnYsfGOS9/EJTPPPhVjrkVtv7xfUghoSqWoswTBxubQIuFA
vA7qztBSUSomRc2krjDhAXNu8Ay49JnvwGQ2DE8xFSQ9xnJzrZ3gJLT4zLBZ12S1
KBLrX0WKo13rBE4R0s/CNVkiNukuDGYpTzIAtEZ6n6WOj1nFaLUSNpMe7em6QEbO
PgDhEzpoz+baB6rIXgttxwLTUnw08lPuI2KG54KbFAyRmzLKGLJ73t964Xa5StBE
a5ZVcnvviYFeTYkCeOk1NfXpNuq1n9gaGFkIjcl2Qz0YUcz7SriTUNuObGvAf6Kl
elYoK/5vHGxxpYV62WDmtw==
`protect END_PROTECTED
