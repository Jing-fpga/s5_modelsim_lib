`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z8Lww45uOQcsx+jz8JSJBxYDpyyoe6OLWTjTujqhRdrgei0b+CC9xVt72MAduF2p
h5qgCfl558LN8Iz8sLFIx1Dt0xQe/HW2gIV5GQ6rZjOWK8/Zyq0nSbUYR351jAiQ
O2IgZKsb9P3YezUpIwXVsk6jyuvyTpDxlXhLhn9IkKjb9Ja8ifcEBFVX0t3FBxQs
dPlAa/62W7kxhR1CAzFawPjQ52DRJqD4YF5tdg5OhbzjEhAcxUkJ8RwDq78n/SHb
Xco2gloKGLF0/V6xcjy8XIlgKDfvoMhMK6DWZhbBdbb+lcuuCMQSM2GotnBt2RQH
HvEBkeeUNNSlC7JeLo2ADuJOwaprcrC+O8siKHtH6CjwSwDH9c0n1z2u9haolgOd
cM3yRfeax/Cb/w2K5IL402l5l9JzGW+elCO6jB3aqsa1j4gxQB63VGkUhqhU55Sk
wCPkQSdW/QrAXn0xpLj1RBiUu7lnJMWsZH5g8aNMzGWcZO+SINZLWLca8hppAh4f
UvWulyhd+PNW04aeigO0ay+0y0whuj0SY5RK0E5bqvtiaSZyRjupsZ4oTiM/ptg2
C1lLUlFf3Y9PLZpDrNdodeJnsVg7Y7taxcvZuiCyyF6PbxZHYg5hKRbBluAQNsBp
mB0+dAvtu722xFH3F54WHQF9aI+yZ1A2GvYht3fEBmVGHwg3N3YVvTnQYPv3U4SE
Z/20HPNjLc3SL/3iw7BE7yKZslvWNcvuOugd9Mu4mA6F0HBbmkmLoNTgADSXeWUb
0V2E5sER2JRDFCDeVhx3hoR0xQhv1wsUCDW+KOk8gufWx24q5GAsuUgMMZQj33y9
VxjJ8+s7J80qal42H/hbwuwiMBL8w3/UM4QfJD8Lq4uUIEMqezZue2qpx+Tf92Mk
IBFAUParDVIrmbspaxDqkxMgmm+n4RgHwnZZNWjU/cT8dLzJzOBlseNrcq7dyTOW
p/cgrL2fJu2hTd+OZ7q9v3lLbteTsmwI6MizPSzjzwGpLihT/AOoB6aL4XvRUvAS
2L2I+LE+H81CWjaS3lzrnllZ3FN3ZUOxtjZ0J+nktfI0LLKy3ULGtwWgA561+bPe
jyH4vmg4k9/UXspT8eoVA2dUWzshg54zTb+vp51o0ZpumyjnyyMAcsWMzj7mcR/N
/8Us81QQzIvYD/c8/TneZtyDgNpDyZWxCH/Aygdo+S51IL6I+sWPUZE9dTvnJ11j
q3GQ2ot21c7lYQcCS9sF//PyxO5L+z6R61YuUj5thyqaw3DS3h/75QPckGZH/84a
YbURchE1iYBG4PWlBPrEzevmOxoB+PXgZxCRpka0pbDyjdcj89Spd1SrkubJj1UD
e1ZD87t6vv3LsSpkAqDOCHGPCPqe5v5n9g3Abg0yaczGfeqgFbITBsoWwC0b/RI4
BNW7aaOhpJYT+BV4+wcPKjvsag9X5h6TXtN6C6kvvvylQIRTY4lvaYtb6XlKYsP7
35SMiQqVIiy104XwFhOrPRjAmPAV/qYB7/NyuMzzCndkkyxuqNWNc3DIk09fSRCO
KTVN3+uEy09ndN6Y08KbjhcNIv18m5VTqwHZSqyRvy0NClX4+z0NRkRoJLllfnRj
wXy9jMxWNv8N54kc01zzkjpmj76gce9+3aihBlK3FIAK/IIv94FsaKBLTtw5IZST
XR6B6iqf1Uref4bneUB3GFGcG3KnNfmCNPizmxcUzoDolioOPNf3kr8nv+ZD1bbN
8jqqK/9CN1voJM7m6E8Qohpcq/Vv/6HzZolUSfeanoAuVgpR7uFoY2/A9hoWOg7e
SEnOGpyDuIYQuOWzy9NwI6/+BvfrcvpTrG/CEOUwB6Y=
`protect END_PROTECTED
