`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oiab+GP3xCXHPACiYznmCgoaNfRmEtDscCJbmQqgOYJfEb9hDEa2GkYupi62Cbc7
HmTEox2F16uARTRk0bAOWLNl9QU8ucuY7MAJFUISu2t7g7uaKjQt/FnU2UkIhf0e
8xWG3Ck9z/zK+ZJ077r5eG0aqLCK27D3ExmH5Q+YyiDlf/sXlsFVRXS5K5PuIM4g
rppjWbIwkDBkkzXLJhAbklXcNTVyx5YhbRKOVFASux0c7AjBg6PF68wRK9JJrlZu
TQNe42sqnho/pHvDjVhYXqwAb5DWuWvsi9C6tJyvuGnvYZCiy2lFWgzKfzVAsuRP
hWeKjt3ehxrK+1QySd1II0MTgMHDw1r7sXMU/at1qPb2M0AVr9slnoynJOO1nahV
yj7KACn/x9CojWcq2b9WXDAIHW6IjvcKf+up+hSQucqcCqF4WwdKWf1NChAq3GBV
qzUXPMeBppyH42tCfdou4V47kX6m1kbUG+dUb8XzjkeKdrGTe1extDd3SmVLyScm
L5OFDaWM10tRoVhHaxplHB+SAx2tIj+OPrkJxGHtGiCTNPKsWkyPlL2lSNUnbuqU
FDR26Lb3nG/8zwE0sDZivMOig6urM+GeJJ2BIDtAYgoiHd1TFwrt0rUS7irIDh8L
i9HVYenK2cBiygxlCD+v4Wt59aCYE2Mpvd/U66QVdZDPxw/q3aaBb5ElpY7z5GT2
hmJ6t2CR7TJxALwlnNUA2HEXHm58umsfvKuPOkfb81Xf8SMEALAN9gkO7kx4hAfc
Bq8Q5s8y40x5mnN/cplJH7acSNjWhk+k0sW2go+5jGhSP90eaps+SISAXVX3Hfq5
BNWR77vodUfv1v4MApMr9KoXG2888bZ4JWs9S0oL3hxTmUstORHcZAvf9HUcsulG
POH7X3/PFlpJ6P7rh077LtEi7yX4zgVWNtaXnCTP2kuwXTAC0LL3w8s5XO9NVe3z
JNDm6s8hSaM2Tj7Ik/qHhu9n1f+Q71pkA0EesQ53QPRqpQWJIRAR11SLCeKALYpA
MKaWmvR1zl0AkVq+gQY7DF2sILB8hcZR0fTEDVWQE5yFfhso5XeRW8gHIRE4KzTH
7S02c2tdfuPKBT1mAdJ4QisBD2g7wf4xQsyNhYAF91KBBjcYNq6nJr5T4QTg9dUo
r50JkAV89Vauyg0EL2B7/qTd93N3Ct0z55rN5yEzplvjvooeBEwipNl+eJs4QsW2
F/OCCvTK3wcr7/jZRLPBg9/8KT2mI8daGz6NNVE8lhekQWFgho/ZzfijVXOJKVdc
1V7QuAyiapsy+lv1TXxa4ghxN5GUg8hqN9NXRRhtMrkt5ZaVNe3sQKPo6t61qh2N
yPRV8CRGldzKc49xLEwfJIA8gYUPs4cjdJ0aJEEnhaF0xk/PjR33MkzAQ7zSZiaF
cloQ7M+AZ9CjOqoKO+0F/kO/s02u1+qNrNdBDlAozq5yX6Q4fCqvz7wWWhFqCDCF
HxL7yL5swzKWThpZK1u1iWjA+2x0eJlZLwFtO5pr7LQFpmlMkQiSyEjGSh2ce6IU
0lL5Z6azR3u3wXdbWOfBdqJwEeWNXvlOUyDIbsMKKi11Lk6Sj9skxhHms985arKy
2oS6sx/QCHcvMJsLHjJgMrciB09lxZdFpVds7oH6FOeAtWwznFafkXhCJOtecyoX
wzk5wiimXvhwMribXF29vGGi1m+LBXq3ue4EPK07IpEWVK9C6w+DRfT0MnBCyLOV
wkvrMJWFTCZBuEYLOwIO+GN2FeYju614E/peZKPF95b5WSkaQJyQG7HOP2yRuXP4
8M7uBU9wjRfRudOFJKzENyPP/BCR0BPvaiPyrYlIQMEV6GVvNoGELi9Y5PpIpa0C
v+usTdLenmaKANprhiREC07QmT6ZAz/QNWf7hvp37FYu26S0zzh/2gy6YYmF3sIe
j5JPKFt8Aw7pkZytBkt6Xg35l7vqgGA0sDmIHzvJrxzCo91GKxdGw/8nvmopewpX
NJqxEcPF/pmPGgLowwIBERjywN0COpjXFhMHcgvwq5WmyFjwCppaskPJCnV6jrKS
`protect END_PROTECTED
