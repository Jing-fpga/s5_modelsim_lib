`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TaQyEqiP2RRMkLe3Zu+/ypL1oe56b1k2D5yWl3pPi99lwQPoiLwmRJoKC/VJjChR
rltbqkkwUUIl7YbYYVZZX0C76MMk4mX4zXLMuHcidUbN42Mfi9lyLirHWbtkE2WO
/G/55WW9xzjmh83VIueuzK6ajnMqxjTO9I/+YXtQ6rhrYTP/8/0XzHGLgPLHUA06
BeCcqji7eoASRcoRI6vwO5YyDHHIcS5dD2utzqyqwl1i/cx6c4VPoMioXNI83cqD
csdQkFkU05dnAOZiwcPwJQawJreVW0NKtLLXLnGZhJMOFoyJMOVikJktcHEev4X+
uRg/luxekbTJyC/bw7xBQmj+DIw12mhHRfDUmFQWI7TsExj1oeL4dMr6d0rk6HTw
XXEdcfhNL5sFLG+7sjDhWC0B3Yq5HTx7knAq8yMnvEcc1YzWadnEJOyQhkcH1UvR
KVgBkvy/jtmd3DATo100BADRikYJdLK0RzAqS1vL8+b7+rnV+QQM4XKXhXXWpFUu
QJL3bpaQ4NzljVBazm8/gyBiuaK5JXeYRdXl92G0Nf2ZgU1fjwwwyov3LOnIdo2y
lNFJi6GPCh+pWCiI48fKFaVzrgLS4SWz3ObAOdN8rVTZZvGe+sndPOPzTifaeb0k
OIgOyMhTUQ2zHYlv0Yt1XDwnqLi3O6Ki5qn7Nx139g//s71qjF0dBgXqACjeZMNI
mKRNfY3EtGIwwB+PuyKlACjMzwBje3kxi+V5sb7vW6YMNVXaQ/Q8c6QkytTL0mYh
jMiv8KzPcc8X+F49vOYyCEaQzqt/IOSrpkM4T/Yy6rUNlMGIyPQZZ1srnzGofJ3B
DFmsWJfzaJJF75bPcu1XxBOIIMqlYLVLb1TPseJzLe3JoqKVs+yTqsW4CXDqBnqX
LlO+EcrlMlguVBN31gd4wIsl8fNk9e1L8I9aTLN2tWbTBOhMybj6NWk6Gc2bpSZL
LZN9CRRC5/WoNjXnVIMv9OZYFUp4Wk484AygC4BM8ehsmbCyl5GTxxIIO9oYfPh4
bhCvoJVzFKPlCyBsh0GUDRR/RTJymdBnm4EdVLVM+4YJ4GRJiBj3dcQCt1pxCL1a
u2j4EDjuF33mq9Sodt0glu8ZSQqfhhQThTdtgQcwU526utJf3KveMnzpAj4xPk4Q
5s8BvyL66qGmQ4ipcHhD/TWcp7aXXJ3pzk/SzcSJ28a2K3Pbqmfh6Yl0TYlqYKHK
tKU14G/6NjPJItW25V/qPQ==
`protect END_PROTECTED
