`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V9DIZ8Il2d7PqqvhiEWrwUUEnzXI9pSfKKXvyR6oys6nC0msAq/lx9Y2o/yCYQsY
9mjJ4skDNe3H75Z+y5w/BYVbFGEUyJCSrO5JiuLboRGt85hY7JVVl2RxHgnf7M2j
Vl84WRFPJZXGmzLIMfWiwZRVA27Xk2UAAWt4MgFG+xQHNLVNxwk5N22UrlxkJ0Ls
Xtg//hgm0KPyMSJij8uA5rp8HzCmxWkPi5v+Dtrutyyicl3e58h006rnvgkyeaVc
1X3JPWYSnIYKnH1wsLbbEZvy/iiC5Scfp0hoAsgmXiGFPpOdC0qL6pLTOTelHYf2
H2XmVdanypZDvO2khE+fc5LItI110rjeHzFPkpH3Fap9VzyMsYufRHLnWSD5VoYj
CvMNssbP6gFJZ7wTfhZ/oxQ1WWztt6KI1T9y2HYR7aGrz+MWTj/jFVbLCT0JS2Kj
n6DLQ5T4yPMoCT0gJfcvxspTJzefU1NKfe6wc3bwRlooGz/II3cSs3drhbWcjnpK
PL5/D3Au/3NeoEEa4TAUdbYlFlo0waq1wwipeI09AgbKPWCFSNW/hCpNi1Zs3J1H
u18zYI1a1tej0jctdeKuJIJNCLkAZ2ZsTsyZ7PJkEyV9ChBt7GNJ/LFnvNtdQSkw
df8E8R1cZdY6mLxZOWknEEdjTkYQ+Xp0YG9oiiMaJVOojAv8fIB1SLov5f+cp5x9
OfYx0lZBEGzz7IVOYAS7wI5jBrOpobncbt9PrWp/mdv/DPUsk8MLJ4FQKjl7eEqI
mhdkZ47e6sZsFKRx70dRKrs2MDTYNaL7MWywZQhHZm2RJui7saB/h7flTbXoFA4m
YXHu8GwFk7X3R135qX4NucbnM/tiNQgDlEn6iXlHOyJdlXNZHjtzIw3ViSR7efsu
sVvZLmeBH8RoWEo6vNWJ6e4P/EcOCJiosfXXB3G+9CwZHf+PkDiqvVHJr6r8hlZW
xjzQN1IyuuH9kZZypQl3d2TQKN7VUBLpo96Qn/mug6aa7GmlOdGAvCiDYLdHFXqQ
PjV5+qD/pGtTH5ib+50PL7IB6DSVgPQsB67l2TEFK0TMYimuOsOIDoKZMz477uK1
pYWRX12RfX9SNJRVinUSEtKM6NRcHfytU26mpBTVrZHtzc4uJmW5/qhiE1+bWm0V
dcnik1qazTaynNeTG0GnM+fliuLzzUt9sTtnXXJW9y8lQqixflcvcyCgNQjWSl64
I36U0JjPv59nzm03xnSb72MTSnKvarYNT7nh7CzMDI++T4Imc+/4mkzjtrDUIM8i
lIc8yCdbzs8PNzikvHCNdaElEDfy49bKOvGh4xFKXrUqHTtkbH/hXh083LuAHrj2
OCz8x6DR4zhKU7ISZKDeFQLeK5KXZb53sa8YScHiIk4iV8fM1preRUOFjKRPsVe7
1INB4GPyy/tXUXhX9tLsMLXj6tcQ5nK62vLerttKZAJWYhLlWRIMyctQZDmv+7aj
czj6wKm2GCI+IZFZZt59TnUE4i/MR/xR8dLvUryRCk2podCNb2G3yJBBe0FRALWg
XL4uR+TcPBdnK1pbZ6b7+sa5Y55POPk7jp0QAwdJGM8F9kJ0EC0btTH97F9NvJJ/
sDaSFfXT0cXo38SUaha29okFmJkOvf2KsYJcLqfmfFpL8xQYkZQ7UHGC1FXzCAPU
fIu1AaKeYNsjouKvON1WdhSNM0tZaEy8ejYxDatuXPSg6P2DTwnctwkL2mrVF0zq
3slEMIErMoeZWoKD0T0TdulkCnD3JY9Dl8GeeljGemixJlsNzuQ2SG2YW/sKBdwf
iqTy/Tfnn8gvwfqyC7xeKARc1km/dibjlINA+afotFYJu4L/HxXADYbUg1fCzgw7
ymuu3S0byZZzfFmUyiqIbPc6QmBcByDCC7CraCSZrOjSozL4QoNbg5fIiIvHxydr
ewu19HvLjawnKCvRIiHlYAryCdH3GvSB6mrT8gVmcsSJoR6YIappIrMQl2jocBBM
tMAcszwIbyyrL08QTOfyIXCOdPgnUFXSxJe3eMTj0yFuJIst4JsdYpSiN2VUtrzV
X/XB855L3Svr/ulXd1cWBP8dar7Eo9S4stEujUVMrswo6aLuFZk41gTPVbuTbVnD
KC/m2MLf/uIXFdVNJnEYbkwjgICRQRwPR4xzceFkAa9iCETM9fMzjW5HZsMKkO15
85ps+jgppLcY5HNnoqTADPKiryYmVYiiUsS0yRs/icesFHkcRgUkJr7Ytt0QbExz
zEKfyCNiufcQX6QDUUsQ2h2dMu3l2spT8omTr0JrK+3idr7NUWwMwb1u0pUW1bBa
y/uvCSNEtnRPuE04NfKiw3kb3Vy3yC7txxQJJUETa0Vl8/7/BwLyiwWzbzOSjA56
I6Uu/Q+ekii9RdyIS79m7c32K6sAov3l5g0MMBz4Xn6NvIy5/BVA61mFTLNImFh4
Da6ILmEKBjo/fC3WrN6Fyqgn4BsWRt5W1y6h0elzCSWanirSJxMpMWNrsnjcEDk1
sgvXU6hIUq4U9xEb8eZ/Tf1vi1VM3Ugp7WKsyzYLeR+lFcvwknVxH/atkTa6hhNe
lhmOB+cG9aXqBLwmnns32MRNTwSg5mTmQU8WUnlR5XdXlau1nxXhrXVmy69Xj/f+
ifl3bGlHPvrtWLskDOzackh5TgagkxhVfqT2FP9hBBxtvP37VkI/lAUZXph3TH7r
5m+9K1pJpuY3octgWG+ZnWJqkjaYWf5CQw6IZew/jx2ImgB5AcVA4BpToJHX8NMr
iHaokQ+IJ1lwW0pTIMtvbLR3k81hBz0zKs4E3Szyvy0KQi2kk4Nty5XBND/ScnbU
SHPpVuBeqkyIx3tCC7Y5pozWpSyBf/Yk941299XsZ6u6hhSNSl0LamZP7xnFc7Pp
q69bVxUNd8XOz1IF6eC7xE6sMlMQDLA4BxmF7QWE23RK3+CfyK6rr9kgJCW2Oodv
R+E+JtPoBa/Bg5ijAVkcdqGAGaCDbKImtMNFR6PZMt3luFmoyhbsy8EF6PT6IIbt
ldKD2PwGxibxvNYOcHbzuRYGMsjqztEgZjcUnmgRi2DrOW5YxU8UAfVCTgFhuBB7
pwIXsDll5tlu8McDWsrYQIsd6DZVyPQULGnJEHR1oFBVBTM+9fL7IAqe2rZsDdz6
5qZ21tHvG4mt0AszAtq8HK0jHKEQDwcLgpFBytIN7HkhRhJmyLaPtYSmBF6hdBYg
9khCstGBLEx7cVa7UQAJQxNK8dURV6c9lUT+PEJ1eDUbMQ+pa7o5fOViIttbEWz8
wyt9iule1lXuf2u/wCDj5xQSQfDTepoyrhehXOuL4zr01SHn6WKhkEHuStMXALUj
oqlMhtCpx0EAGo+O/89wgbMm5/yQdxvWaGxTjuxztVQjQ3gEiDKkLBBa0B++P24T
gHcbP41qRNngWxo0wMZHxUnNSQFeajLLLMNVnMF1Z2YGWZXfaM+JbSVSVwkxEios
n01NY8IYSos9YcRkmdUGtU35QhFkzYj9EZGlXqofUiKjRh1lqaAlNEpCFFWC4dGI
oPXquIk6KdTV7oXtaMg6h6ht9vap1E25NHbAJATPng5C6OpTlP6mItJZFw3sc3ZJ
bpihNLxFmaZ+n7m/vmJ+ocbB/goQsH3aq3MUMSv+rPOXMG5i9NHsURf/xqn46E8b
VzZ0+hsPBWRtkvbjt/7mK/1GVInnplOlogzv+U06W+duSSpu7l5+Kg4sAK3A6bsr
qwxk3yLS2m39w4Pr33XsuLYbOOyW3Vvf693N5sso3mzDOpLfiq55eZ7QGfff53IL
6QX72X2tg5WjmpGIT86a4s4tuQyEY+lku7+4JApQbZGn/SVVZU/6bGbRCf09RcTi
o+A3hsjaBdEl0yFJukjWPs7ey25wZBgldMoOyDOpIrnwV34/OxSdUV7Mney59oa7
FPjBIo3gLUJlFn7R4Yc4CckDXkbRkvunhvvMQfbikkwBsAq8luRT8bhixqqB/ITC
mCHf3oSXMtPw2n/jTCl5bKMuxCkc7eDOaUsHzDriLUZoGtmpfc5xaOzIJDuFsU9k
OkoAbidGBLkUYKgG0RCSI2G3EVKf0NMjBPHK7lYAM8I1r80EpFJuoggocHbEg2TM
MXvIUdSjLq6L5BHL8moa+F0RrItVF3/c3lTcehb67Mu1nRsaLjb7EXicLM7+3THx
JQ2yry1/Gwbox8CPXJsJFvIqtJg1b4EeXKhwRK+z0YEFd4iuq9AqaBo8X2deuuP2
Ml6buDG3k74gpcgBfQg6dNVKkAxsFH/Og6IZsxS8IzdmFljXFRq5mn63L0+Z0Tzx
crj9JQ5MpshyrINq4weY2WvPsQ7RIbI9w6xU6xdkPI7l8m1JDqjTiFlJsQOBH3oo
iN6pL+ufv061xq2L05LzKQyy4eB6vsJdfCxQDklnS1/4s+9DABCnq39BKdKTPvwZ
/lLKH9h2/d5f4M2nxTw3JTE0cgVpcCF4Qwrg30+yAN/BjZuYvVlnckQUT8vWBjFQ
mT3TiZsqXqXfygT/GQdNDmb37BKE8x9oVV3tmBQCe/t3qeh6gCEkI1IG0gDIirCk
nkFKXhAtsmLmiR60fi+DOvQRdRoZ4yebj8zSMHgZ6S4+4zmUtDuFV0I/n3uT2C7X
C2+TL0icN+GIP8whWLeMAh4Q/ch95MDIIxRkH5gI6HUbUukrM3sadw1jbBGymSaw
Bvi08psltYAclATjJeMyFR/8WHs4/vo5hW8SGqi3iS6AdP6alBktUwBe6oz4OcF+
nrKjLtbe1Q+ffYM69tcRWllavtg/AHChYWuTOjiKGcFvh10qKbmLtJP5CTI2EWHI
baH24mwmRqZv6dlonvHc+RdEVLakQmdrBwqYc0PYGluHzN989X9W7eaajTM0Q5fD
vQJlPTvjRrKYrcGP3ZvaRFYHtF1Bg2hi9C1bevQiCmWYSnv47Hz3dWuhV7bM9Og4
Af5UNejWBQCWJ1j0xjPpW5qzncy3g2V4b1RpZfSaVM3FsjsuPwRTR69LtxeWNRu2
ghwB2LaPL6VvHAmiPH8JtScd0kfTY4oqcACMLreA9AFy+ic3kaJkt08p2H8Zucua
rX00qKe88VndiY9f0ydBQbGvaOz334AGUYbiTwuMXvYdDa2JnfgftqIflLiLqVE4
DvIuZuqEDaiHqfqhxehsIDalzBTNCLhIzStOdQ7mOeznfKBFtPcHypXeQU86+1Tp
xOMrtM4NwwKJTFPwREmUOUpIQpvtT8ZKnY2aLZFct48XTJVluyZu9v4Xf60t5+f9
iwWaKLFuj1/roxFXoNDOmxtL/qTrLvubFG3BPyo0KUNo/iIgnlSBNzleIsak0Be3
IphoH8BdBB3zxDFxHmrTx+L9LCsD4QQS5xry+hnirMtUquPu2Vs8XNHw1uVrC8hV
HbLzMJo6XNK69m2pg4YR1LvzcyQKexKy1NVAfKve62t4DirWhifnSOqOKFBr4krD
E3apeU3tJTC3KoVkg2JTled8Qg5NIlvVC3/fmtYwdSziRryYtO4XvBZ3/JHtgh6j
zvmJM3nZ/xiah/L6JneNQ1q6zwX6D79xLA2dULSbDYwQBBGyUZvmAHLEvHq3+FL8
z4dZNTx+6NoN9BA2slrfJe2l64jzuk4OTPnsR7ub2SMZy77uPMqZdgBjlpugDqO/
17WRh4sgVQ2AMi9arOxf79bisQNo65yRqVvw9UJOW1fwBKQTDs4FSQsxElKhKYxT
Ha+k4D8Yl8z+dgVD+Zr5A6DMoi3wgAzH8OWuENmYHCHgv50oIgPxJEUqeUktGkNZ
tvhzCqUjUhDCeqt0947lDNog2T0ywFb0bHjRMg715+MaHgrfzoGfx/CSCelW0gKZ
W2MI3dNjTOOUdSju+zmqq11ASCS5ziEmO+9EoA9f8Ix104jwn8t+p44FNPRH651D
/kKHyd23sbomQQ1F4oA8wsK4d0spGWSCAaQYIUtr8PWxI6VXsBk3ajGl/XmM8cHl
f5A4AU6lxeShGOxIMk86y0xB3M/Rq9PSv552972f3/lsH2VD9EVGI6urEDRMmpeP
LOrGOWxpVzAlMn38cAMD2AF1QEc0tLJwhQB0mnR7Ls4+ICC5eUWCDJJVIO4gcRDB
cV6hB702U9RsbMJ8jfuHeA03wLtYz2yRP5oArvOqEYtIazCljfLTX4j2eS/0K2IT
bAa4BBx0b1luCd3U7ZNPpF69btZ0no0p1FvnnhKTTVV8yjrZS4Re+Zv7TFz62eJx
wfj5t9xRNSbonhceK5fpu+GKG4w3Cxl7HbmoNgg2XB1cB7agcE5Wb6vXKFcuAkd8
M7Qsdtm2qqkUDuoSF2KWGTA0VgBPvi4cbSoWB/vfyTqCxmvfk5BWfqFkxh3meA5G
yYEHUtmxI+fK8qYesZMwvdFagGUQzvHuvgTGCsq++LwY9yu2w3kZWlmkrCsHQ/s9
WH+gWKzZflxI4nGxPUf6T8gTdG46l7vwPmg/Sv1EALXlpU397c9JMlbbblsQcT1v
tUwHmhwViXIl9zIzlDENT4GZGj6E9Y+JpX2IloDyLVXquLvRugdJKUYvQGPAEQP2
W+m7Wj+zuis4E/mgAtEIUv5ZO0+/HBqyfCZGaAqowD3CxS4WOFoerSMiBQFLphsA
LsCADGrIDmLEVFDn+o6oRxJQXFnk42WqdnlhIz05myEcPjfFHU4/KEgSsmNhmbMs
7GlgcRgaIlaUaKmOJ4uK+woWhWJdyIDDveS95DQ5wI2zvI+aRg2zFNnRgM0QdV/p
9SiNKN2OPQzLOUAgLMUWfl4kcXS6oC+720RMpNvWfbnOhrbBMZiEk5WhpX9o8nFQ
vcr1fthp7GvOdYATphPfsaUg6QE/IRkbbWfv9r/TneSGP+jx+ana0v7Xs47GDQEu
vKnjWDvhE1zzDy1Glrq2bVDHvQudKOZqa8S+r4ri9tpr/Zq6+FS+75ATlVPaMZhH
wcBkGI3pxNFv92Qvnv7aUeCKaVwNTgLvrXKKcpEzxZVne4KEChWacUBQzJbtCoYV
1/+5er4R3P2ukLYPnL1bC8Xon/8T5p+UcEuIjJexaLbAK9rtcCDNZlnl1QnoYbtg
hqt/c9d47Qq+z6UzcN6sCAzKfouCHkm7buBx0QzkonF2jHiVsH5ZhQeMCjBsfDoh
BOkAlXYsrgQNy1KIWtIR+dO8wAeI5XROW7TOqPZ6WMRuqt8GAE5Ro8w4cjvITJD5
iV5roIC5QfIGyv2Uq3ZTvjuYwbQGoaVjJZq2fcRawwJwGkWH4/v6GfnPHgpiI5Pi
JAHJ+Wl9D9U49uerFRFiGxqTmDailete/G0cJT66TNHi7EhNcniPViQ88hxyaQ7Z
gPKcCrdqLKZr7ezIdGw4B7JkRvAnagwIJgSZxB2ACHB1M7EZp3EcwAe/o5ty/ZjN
eykN/vfLx3AMZ6DUOXj1PRZMznASzDURAiQ8kVX8qGF+0hghWpmhg6CBrq7+tnNZ
XQiODvHlxXLpWs1zXs+bfoyyzCSuEAyPacLOVFkulb7zhnZfa0zTvM7OsnLmpJwh
hZfdZrRNPSubgutcln6WYMMCaNIkTC27Gunlm4jGwFfi/Hld/eTOVBrQV//WvNYo
4qWMDX0rk3c+LTYzGMDoLVaYCjHpPJ6TPYz1rqBgRGmoHr7kzcEZZInHiXgPzfwb
/pbsb2fqcfh3LZf6l81xOX2eHexSPaMgZQfsaRvYX6TR/1MKlgDvWRSRZkdN4KDa
7dbe2VR/I9aeCrFjmndB0F12uPWsDqiOLpmrwRvx8UcNyXsZ9LE/UK8droztnRgs
lG0SWCFoUuzVnsf49DPqJvr8Xf8ryd4ywKC+jO0SVoP90PYAH0/SggLbbkqx6I60
lva1GhwUr1ZpghIUVlVBGh3FiqM6QcOPLlGj4PQeIE5RP0r8ZV1LFJ51XOPm0NL/
O+0SFMAN8DpygIwH8x9bOgZmDOTs9AJehHyQNDiVUJyOphaOAcF+z/QMDjVvvz19
mR82wZl7DjXMfhD618w2ZlwRnINfT16H9W898Ss/WEu/2d394oji5+o2Wjj6Okyg
iO8i0cy27BA/mOH4LAFZMRcmydoPJuZ41TQq+WCf/PIg1GsTSKIZedGVZDBZs39C
J+l1gEFY+r1vbCW0jOTc+7R646symgPUX8kif1wL7OW0njjn9IJuZhBwrGQoZ8Hu
z4IpniY5JsIauVVhR5M9eq+URBamjVfLBBNnyMTFJayEDv4MFqxPkf6nHvfFNsyV
DDfImzVFPZ8CRq9C9y+zu/MxnUE5rfiHG/4Q5l9E+T8v1Qc8DC6U4Z6anL+q0Ciy
ED5lPAazfru3BdwwyDelrWUR7C62Nbgzqg8Thl/CyFiTsfmIa4dQ9AFn+SN92uF2
1ORVcRMbwqv3FnH5V0shV/a09dhMndaaycQ6Qnealfb5dN+vi+HzpqNBi325lYxR
0gPpVPZxzPWgCQkjotAV8bGBRxhepqB5MrZjZ+CvK0cBer5LewejtcezftXO18C3
N4aeyB3axcbBjkKyHRDKZzRrDc0Y1dZ93fPoihTRkjX43h25yQwKe6nRA23ictL5
iFYCupoYI+Xm8f6Sie8S7XP1GciyQIBREXgH0r74EpAhFr028lDaOWwQjjrP7ac5
iAqxJnIDBR6YIZhTS0+Q2rog6yB96m7znTjaCfV5TrNqH8cG7ZWbKxfKRtpx4CtK
y1+UFkgKy8UjOBzlABiXvsWHcN6KT4RVoHQJtuwq2C0clds9Wb3W5jE319ZDv2xj
s8AGur4beNSHLQm9rMulJY572UJ5sIeNMG8QXg+C2VfzQl6AIDdv2mOpso5TsJnd
Cli22fQP2jvzTNOPNZ6cpdtHLLUPiIrOwMol260J/SW86D7EX6k21dJHLXsOqQvS
I6PG8KyyV+yA7ysDRj/YgZUAwGrO5WY/LGycasRF/LGkJ8eZHb9rd4uuF+Jxg7jh
fDEN/jUeMWzmfdsQDEqC9KLEBQK26gycs13QicJ2xPIQnej201DBW19bMIc+7WbV
PROO+OhoB2MxGhhYi1rFHPbKd9sV7u+YNWhO8fhEHPXtNGdPV2w80E1YqirCuEPB
mZfRyQUC+QjH8EQ2dBnjj9dBbwVl5+vqV1528oCPaWgVRfGXd6u0xFtY/Cnx7Qb4
xQ8PIWQrCBEZ0tfYQ6VM5Kkx2gktC7ZcHeYA/QV86Nq7NG7t3VHlxoPqLi/LK66i
cxgAPT48MlYZOdr+KTiFJ6s1obT4aGKMYBfJ5E480tcCbTJrisFrPJEkjWUjH+LM
VKdMa9kOYo8eX0AiOnHSfl1vSnkCN6TDmUE4jZjIBSc630tQCNtfJXx0pxkh4MoY
JHwnSlHVD5QyFp1eAUjettB7DoH19jxFJMyW1LDEa7kUURFCAMFpOdjNOFf6AdBq
hC+STvMj9vGlIh6kIcBPMXY/3KI3MMWzwNo+EvNuS9nr2eaNStXuue+/ntAq2liG
AUj6o/aHUZuMri5/eQIo/I8wTj+kmH+60esoMGozge3ED95ZhqFWy+C4ECV5oN+3
SrNn+kjj1rdTIz87g1YL0HUB3bQn41nQFmFHhoPBEWhEeWMtTPMFUIqSJ3+4T7f0
7aQQsz2K50DG0O1iE5EUVgJq3sMHojIyQ0TTT+pQYeDUoYfpjEqIOnivsdqgJIBg
NpFBQoFisJrLl4aD3/FtWgAc9aB3qh5hCh3EpIOSkq7CiVhsMkNnDcN8Cw6fRcbo
vvCJuApH2knM5UfiP2HTw/e47btXQ1zBklYYusufTuzP7B5o7IdtBpsyGVe/TYzr
OroWOB6YLDKIAoWbWdf72gHMpN0iR2IaxqxBpj5+v07dARWF2XrMLTbiqWejKvBH
U338hAG7s+U8m1d+VlzpO4pVwUQTixlW45nRzb9VUwmwG2a5cthnOvSZcULaJWOp
dKE3CzlxG5IcWui1MFiE1xlliKF+qyX2cAQWpgFuqPC85i/923+l+KWcvF5XMYhk
WXj3cP/uPLswrX1U0C5MPYpW7HD2Ji3N/EVOE77pa2Woa6fmyHqkkAxTHniYJ0yS
92CD/1D21apA8bU6JndGYrPWVSK0Yty8jZmxMrsDtg3IkXr1UXHYtr1zIK7UoJL/
8gC/Eh3By+JXazIV2BpHpVA+PGP4gRv/NjzN0cnxDBEIKaxWp+GMKb9XY+WcX4n+
9zNDjWQUMrIZlRjhqT6jqMqPpq1Y9Ao7RGoGseqAVhzdpV4/mugGOGWVRxh+KWap
+rO+16UkH/UX0uNwa2+7af6yLEZoIQD5BvppfUy6ueLySfBxxF6L3ZaL5htlAi4V
5O7qV3nPSYEwOt46EGpLMuQU3a/AxsqusfMe3TKnd/dtwAJV9JwLMzRjF6JeKx/T
wyrKzYyy3gyaq66Y+ddb+8dJ/bvYPFKpVAXX/0msUoERiTkIlAvEnr6nf87hSavB
/nXHgnNt6dFQDXVbmYmS5Nwp+BWtRVD+fjBKaK30sCT250RhK07yWzn/r+4BAmP4
ZJFgsClTcw8bl8/6c0fPWBmU+fY/yaTOvKYHGDm9hnzApZPYi8s5dRhb2hbZz8Fr
WWQGDeZ3EFAQCvWBn5MFOOtclK26Ccp9qVvJWn/wNZj0zndRFeou4bkG5xc+dS9D
Grx94WjQkobj9wbxUUDTQUP7OtIQ+T+CoE9Xo+tRFpme9lP3ANmewdSCXpnQ83zN
UU99ME5gWyGokcnTciLMHMtcyTD9z4HTeH3+kn0KOg3L77YysPx46nE77SX5cHkD
SH+E2o2GKRTkjjI/UY1bdeLYgJfKmjkuQ9m9Mpp/mw2PnmREJJ6XDUqDtGyE4Hpl
TUFSj0na4CUkqT5gK+c0JR/1U4dYBm3sjUfuM6xiNeW5c5BC+YNIdmJOPKRoHMWK
aRPdZgfvr44APpf/8JHEOMSsPPkNeMQ7tXNj9AVvCA2qVzRfijIkwo+F9OrcodK5
xlGVvfdDVLD04ziKKEhP7eKfzYw7JhGk+Ve1Vq9gEczWSEYFLa2JAZHu6cFZ+oKC
ZQqoGX44Ei19HAb0Ts5TGKt1hlBGJA1sCqJgsqugcO6Thy6JQLNqDoKSaRzI4pyq
yFuEaHnZCPtZ0yakZe3LCPl2mIzZ3l8AA+DmkijB2Ol0tSv3qIn2CJUXH0huG5ZC
3Fgo5lu2/CoI8ZwVmSJ70FEu4052qda5PfXVa3v0Kc1A8wdtZm+gYcUZqSuZHL5F
XkG9HqLR3eDPfA4jj9WEMiCA02koBGAJVlsjS4vkF3aTG7JAQJwjJcj5nQ3cGRbV
clNVykgBGOj+PnMV3s/D34SI+b6E+rwEwR/pZTyrRrJrSGjOngEazXbH/R2i4St1
Jkl0L2lt9Arxst0nOMemc2Hc+cmvtd8wC6oihAdjjPaofY92JZnkv5rIdu9FPwM+
/jhzfmY8Z/mxn1fCl2zjmhykXXBeRrCEvosjGTygQndeHBfJ4B/mX/ICWaD9Iyrx
ntOSdeFXnyQaRQ1nsFFzWDt+Fv/u5VxQTXsBWREnlHynO421+XBaWmBwli1r7QM2
CVXWyHE+sii/Kem6uHUgffK47tlvPPj8+OjUnyiaEJBo1AWcORp2xEi8CQxk0+Q4
OkP987dZAcX1dRSqWtzWkRbB3bn38L5DgwmzvnK4NupCeawFYimUPNbh66G9tcYE
H69KTs0xpCY1N80lHz1KYLKSX924XW96jir9ZfpsV6Q2W3xLROyo9BNF3SfiA2vh
SSkqTnzPuSRoUvtFLlnfosLlcUlcadEnCz9dsJNEYvVc5i3aLyjfq4T6T9OGpSLy
LJTbiOcyZQ9tqvn4fq3n5II5F7xsE4wzFKf+OKo6ig7HIfUxsrbNd7UL4MVAm9di
Cpvw5iRMrG7wiqlgvdeHPO3cxRFipc/KIrkXxG5UiEdcPQ1hfyOotOQabyWez5m6
pW3kXiw864nC13HuJ6yQn83FB9GNu/xvl8CVq+cmFOA=
`protect END_PROTECTED
