`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jrk3JbAqslfyuDK6WLbyF+VYD3Ku7uTD8vemE+ltW0zcftQAh6vMSHuOEDgqC/FJ
3YEYg9Fiwcar6OnFLVJ6T0dfq5OKf03yopET+gZ9MOXey3fYMhJLHYXrOlmrYZwT
Qwk4UJNAVAi8YFO309hUwG1gr1JihwvJnhOWXOeUrkLJTkcaC2JtelOSan0Mr5Me
P3I+3GP3ekcsZrRENpibG5IpMhdPkyMee+eL54IU+em1RV0VeVR/8ZAFMbEfk8Tf
b2drs9uisOTGlw9KWO+Cr9DR9Z3J/75fTPRpjkvYsRCpbW+OxbyqqY7b7OEubBcT
TNjEo9hn9gzT/W+5Va9gMHuzmBjTqdanDpDt2ScJ160zLS4TeALsShhyS/PjTW6X
hkEbEbQrKCHIOuliGRJiXLi4z0Xyh0lV2G6vQ3i/ubkNgSzecwnMgrJKv5h7SRIl
symozut05xI4yZEXM/qNqFsDIqUYtmSjqbZDcw/4w2nzL9g5dquCngKOosYAgcxp
GH5cK7OgqBp7hwuUDsLM66I5PbtnOEqDlQM/7/kKDS3CgoSuxuhlSrAlAAiltq2U
bZMbGdvOWAIbYq/6LXIoh0RT0McxtLFZKZ5GqruXLcRxqOexA9EFqC7YexmScQuw
ha68uTKuN4l5TH2P4OikoNmGS6OuA8zAj9XFZb2DysTbHPSYpzxEJfsbuHeZfbjr
ulCOS6kuHJ7a0stopX1a5+NXeWOFVFFCHwTSpQKR+QwbivCxrV+zcRjeCeTmzJDc
rFCBRM7Fy5ePlaD8ywCB4EABHIZgrD/AeDMwXq4jj74xhRvgiNFCJvDhYfdc5idq
v0q4LmBySedBaJ4/6cWK5hY08PZ2PnEH0tRYYmOjmvNfzWtpGPQ4Nuqs8ynQ3Dnw
J7EcUpcoC6GooH0q8rFLmgP8c61i9vx5QXWeaJByTHDefoF/q+/HkzL82UX/qa0t
DGwXliS5pOqa2evua+ErkCs8MdpgMxpOCRNXCY4WCTgIMRv9iKE08jL2T0munnBX
28WwHld6111HFF6JPBhsfiWxMBZZFkQ+CMELB9wBqOgwIAyM844Igfeo+Ivx6Qn8
aEyJvNBEAZO1vgQru7ESZIJA7PSx3JBKqQ6EVx37UYBtcds+p/bBemEBGiKrgRlj
J7ESDRqk5FTUkBRvm2IGhB+CCRh0S3RYHUjbZ7nz7P19iE8Sz+dGqJ4tOx39VO4k
fqnUuB3fxVzL8J0b9LYRMv4aFZzhERKszlDPo5ug0AflAOfsOR+NamsFFL/Zi1y2
E5VqKLGNjUj+m6LqM3BWfWIqAjDv+RAkhxj5zKqR9gqc5/fFBfj4Gv1c2d0RQ8U/
sQU+g/GE8i1sZUW2scQgpeoul8JEoXnytm+v/gtcmpTfpFWIZ1FQ8HS8Xf+YUvPb
hSQ7opfBhiXwxEAOYjC59I9VPvEZMDpAZ+MuHl9aNcDYsllxJqfB6y4bkJVTPosr
Rkqf3t7PID2pQTCf6Ktysq12rIHBWA9TGatImuuhQjtN8wmuBqunQBZKggP/deHD
xh6rKcRK8DGB3bfEUbOBDF8CYbmljIn+W6Pxho8EXGxaa/0dZdMQrcrDOtTetY5j
b1RE5Lu1HAJJCeL62+ZIv7uEbLa6qIhAcK83CFBPDnfvD5OaKAiTb7tWQIJVYxlU
QS4ji4DNFEqoralLGaMl5bOMGHWejCx38s2jxpPB7bxwamVAj3Ps3sLiNhEOh3pK
4uwEo2MKHQNz2IIeBBnP5Qwq5l8i4HtEh/mjgYTHImTAc12x8GAJfP+iFgNdFgN8
oA1Fua5WWVRMW0icE8pecFi3P/v0S57+j5pukFQK5uGbtmYXuPvlgr51DXUJAwro
lTuvVoEz7ZH3z6tY8/6zuffRdcdQmMGHSsgZm6X9Dn1WHzbmySmCQXyg5iJ8ICV4
WmsS5y3TuUxHDH8l17svlrrHS0CiDUmPfGORaG69/G/lJXQgQslxwiEH94Ij9bqy
XN2hwHtsD3hjgZNZoAwTvk1Wyxv21HbPob/6lnTAw7v+psdZzU8vieYwThjXbFIK
9E+PsnePQsuxt9MERtVpMG0SXqE4I/36wDP6hC7v1jf9tPRoJ2xy6kJk3I7OEIer
UppJQIAsziulHnJVUIN/GWy927R4XvAZUJd9ZW7UDcoUHWnkdY8u7XG1FDUPtjXe
j+VEu6H5eb4GRmt+M9VjV/2hjKzHrm6ozIim5+nH3CDcL8Zivjqm4HqfJ64e+dbh
NULl9XTM3Mf6BBOjNNdMxP5Jysa1lIOJqXOfTlntXMeZp1ms308hAO1cSfsjwvea
fUYaiFyNEpHO6xt1FESKynDOW1Xix8FpKoyoHhwCFAIftjZYxLAgwEckBpEm9tGY
Tw050iNUrA6S6CzGl73+HMC0y/Gjgr8aHF5d5pHramRS6bsYb650PNT1h76RiRKR
gGGUkRDc4tT3eF0rz65+6wlj9LNoSzsfk+aVNxZ3EWnMB+fW55eyvSiaiB1rsDpk
ZcGeahiSXMt/eiBztszU5fpJ4wTztazHqPuTWxQJr8056HZplYTPdpFGvN08A1In
luNVePSTu63v9zCykJglAYyXdrnxF+TG0+z1XkXiANHVJrZ25/Lmxnps0bZELQsG
K0faGKZrYs2pn38azpe+EIY5Muq2iqPnZMXrml2VpJdKnfuqWEU/xG4bnlqIb6xX
nxVPd/Q0qKy3xuAtfksX4iezoY21SpMv/qsdi9iKVXtb895riBMhIqCN6L3PupKs
fH6buNnSdrcaVgUTXuN/IAn4pTufMouvIeb85sZYTHF7GGpOVfHI2aDWWMUgWMF9
3aGYcC9bxD+cEjioQ8tdVBXi3Eczq6P2ZiKEHqIiYIyxKgYThMplXpRs+iGIl8lG
hwpyM3WLL0jk7X20B3D//8LtEXd+whdgtNE8arFg7n8Y4VpcVVrPrlOwRD0ah5qk
TeCd902X118IVAPSPz5YJt/F+8FUvUvN5mSzZPo1tA7dCkYje1HlPFhP7xChN8U5
pr6hlRbqBAHdoAnsOlkmsSf228ytmxjlb81PiMVNe+Ab3NwtnAfykknav9snDtA0
sOt0D9vKYn9DP8zb+sXWIBZbVBYrcmh79YeiRutrxeyRo716RNn7KjaohD1/03RR
ms+X8l+6dGBbMs3M89J4XriGJoMXwJl2yVpx7D0w1zHxdDTUgPEwKQP7orJJz8hW
TdO5KFHDeQzmqIuq2aAQzZCtlVNDDwTVVo63XLu5SxKhIn3Zj13IMEBDmLJtn91A
ZbBmCB+BW5eP2yO2M+q821611/4GNqxUcI5m0N64q+VteshUzOVK6uN0FevYoUpr
kgshhKXLcJ1W61uHK0pnY+3KHBozDEO+sdA4K3ppJaQpAvDgABo7iDT77X6YRPZc
vtJj7NqSae45Z7kr0+x+RxR2jA+n8tlqfoRu6ia1rkqP13XnqZvocLU6klUIc7sR
AhtWqmtsfqQbvA7sViwihfNSM/MobDQM/c+VVQIPL57iiELPoH+XjRWSmqeGAE8w
aRl1klTJ1+CuUynMX97pJ7PthBkd7+4/3fGe4aHDYfZQHUzHKhcWxntwiQ8EccZG
1M7GPfpJ0bLHoxU+XB/5Lzy22c+Den7kzf5KQXEwmavc740eV3zbfkzwPFtmgBZ0
PAQ9t0I411COe5yRtk9Wp0xvjRRCDM0P6IgkY8Z4Ze6YfM1vLYrww7GRL03Rs5z4
A5zcz3NzDY+z1mt+RjNTdypfGr9LV9TgvJRvfsmM7a0by5oCoHaUdMraJbceYt1E
0khZuv45y2qDTYtfU7y4uHeiyeLZAtOAa1SK5NgW6W6YrSV0QU5Nc+SxpNbS1eWr
tFDCDnuUmiSiGHXjeot5gpnZwBQJF3lJj6mLl+9ggtQn5hTDig58FY9N82HKB3NJ
29/RFHRn2dPq0erKYF2dpwJ7tMBNFqNJctPTrJngeL5FRrpYyYAEDIjPTkbu4l5R
rPhAtVS8iz0YsCeUdIlVrjbnM3Bkp+sE3at/8ymQgSxinXiyuY0NiGVu8HKN3yCI
tgk8WTgbALjah89xuKd5badQZjxFVEPgxwvUbv0N/7lH3R8xVbhP4PkhP0bGx+as
KTDbXD0y6ZOTtmAaD5Hr0KomVROoPW6sh83aUnbpi+DT2UqpMMignVY5qLCL4hHQ
Qix0YkRAn2S+ByTZn9KabFjRY6KMx+nyqxdF+bW8Iutifi76ds+WVSYmGQkaivu4
nbymeMuzbKVKoLtaHbJ2/RczI2GFSW7oY0mei4qg7fcG8vdA722LBTtQWDR8MPnJ
Pm4VfOdFB4RlU8JTSOGvFxbkayEEJ681DjV0QSndjBk5vz9HFNLsq2DPrQeVj1BJ
gH8dSUpnpqvOItnTQgk1kbwoJCk0KARGkq9CUyoiS0V7l0Ba8KVPgLONEx609Qxm
DoRL65FfchLTuGEAZdGl+aTm5e8AEJFf9mCkmjydlD6c/WcPS9igfrhd5yhT5/NG
eD42+xBPFZlC/dsTieQWerrOL5L3Lui69JixYKGiW11CVZvrN54SUmhGfy2bMx94
HkTZs+hk1E/0QUWPhTr5Jbt9F0Bh7pXB+Jyzoy/ESNJixJBfEfifxnCYseCjcAIt
BRS6Lb221QRrgU2/9IGNm8qa1nFaObohBtowbgE040dOp1ZPk605AOEjR3JSO7Vc
hwBxF8s72ZF2PEmnVFpJavx1MqEWmcM9JIxQn433kp6s6H4WmB9gj7HrWiOTjK3W
ZRooP9f1SPsF1gGTbdLKTqeNsWfTUJvMfDQDCPIaYr72R8yRbrmlqRLEkyYh5Xd7
3CwPTlu3KS6squv9yn2T+kVlvDLduNIgwbZwdreNptuotIcL8Lgvjdf0hlkPCICK
PzAT5cF6HiRxBMLNBi2pfrcayiRiLj9GSxoTov9qPIYHt0A8Hkc7qfygj5nthy/J
`protect END_PROTECTED
