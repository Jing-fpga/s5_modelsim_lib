`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
adty25bpowqMvqPvG87yrGoQ5m286syUjJo8n1U/plNbILkzWq83nBn9VvShrtHj
e8nj1ahJGAnQMxnOBU/aMD+K7eWqAbOT+84PQiTE5OJrARcb9Rqpfu2J+okObCGi
k667C/MFUCwYTlfmHva9v0KeInhIPAUV0q48LzNXvEcuX3Pe6D6z7AYZ/SDtTCYw
x6fU/0n7PY+FJAvr7h7X9iLepZ6tHO18OkJFx300t2eiswHDxO81epgQVAeaEGNq
qMhtHyaxthHYcolVtzOm446WiQRx6dGqlVJClOIWusfKTMa4y0ZIoE//xvbC/Kxf
k7T80p5/vpc5LrNAPG0Ltb8Pov4zMqzXepQS4t9rBsxLgmEa8r9sZaRWtnapWqYe
e4wzpjAC3/ill47HQSTvInb8fJsMGXAkjLQbtlVludJjcr6SUvHWA84o9WEBKF1v
Ss06Xzb5Yx+N+8DnLajt21rM/yixk2t7cZlhetQDqFPADoaGq8Y8WN9omvNa2AkO
QJaFugsNLFWzQNMWHN55WZHmEOOIhAQAyFNlXnAf7dt8/Rqwl2NZCxmC5L0bxRGD
RmGmkAxt8SEzPS/pfYm25ajQzgaytQ4TSFVxM6ZlMmGpwmOGCkHKff47VO15o5ve
yq3ijt7YdgDtu6FG5ZadfE61hU/Q3lqcNNUi8G2wFucP6jryzlMVGlstOsd+fjX3
WAUJRJc7Seu0bE9JLRsVfEF9ENrwcNuu5wW1uMxRWkZ4IoFY3HxuEmPkrLe03NMu
QPiW4j2jvTGOOiuofWvoWJxlblTHrV8thLhL2WNZvyOOu7xLJes7j/9OayuOgi/9
wAExI8O8Gx5PyIdYERVRWGzsyDqnlM1RLhnrxCAOoJ7ev8wHiyhUe6hIYuyLzUZO
JRHNN4K8mVOBLXHiOUGX8AZTKJzQHuWu7L2VrsETnksGXL76w+YbranD0X9UQvaz
rkgD4woSCJaL5P2cRKwMT77htEfBEiIV3OPhBuJzbMo8gi1qwReW9H4PkmkqLamw
a9ocIE1qAscKj/moKy+kcl1SII22+zGQIukDmhS+4NVsw5yTOrUvAcO3wk5YEx22
nj383knsSxbRgy1nTS+DucHWyrjOqominRYyUFm/2N/bvoApOqvRlUJYSl4Mj5Vb
2hyUOWxhAFtmaTQP5ZbigF8oEVKs6U7DJwvZacvhdqKKMfmLLAQYmctBRZjWgFr7
zk2dwIhD5IyCXNoKBNBsp596kmC9ELPl7OWMPif2OlxidtWqHMgPPGyYBJido20H
EWpGzjLYd0u+yKU+BTo1hVIu2opsQgL8AudLlk96zAp+7tQLvsbBrGMAXTcwbzn9
8buZPohvCVx59Uk1+qSLwI0bhD0J/ZbnHWaV9eDakLAl5k9tjhHmf2vJnHH+MUfU
ZvvKx61PTqG+rk0KW/i+ddSHWr6PP8L5Jgsy+r6NY2xbKxypC4+4yvA8vH6X4ru3
OQuE/cjdHFSNwrzg8V0ppL3UNkvVkPypg2mYZtcY2vtsUpY1mh9/F1gVkfWSC4Bn
Dp0imR5CF9+dfCRTMA9DxIXq68fuGfJ12znnmBSKojciCxJAylkI5DAYP5HoHPic
7EGUyjUa//oh4bok68H745wO32qslSHMxTLjHXtiQP4rPqj1wW5Id4XhiORuK7q5
7gFkKQt+bfhqGSILrmc88WpArDrKOM8OsDoY9KMPYDntFyCDimDUt9ttKMDEcwm4
O50AW2sk0cE99sZJAm+3xhTj86XR/tKjmmanGM0WkCAENa49/Nb6va4Anwyks84K
2Z5yjYrNOF7grI6PxL8QdCLLfsLKX6+WfOBpnATPuvAcJgIwmL45szTbcP7AvXmY
HoxsGbAC3Y3wxL6341Fumzsh9TqbCvH3+MFtft5qL9/1ixlikHmJpqcpZC6N/bk+
B0gkS07nKJMiT8JUoZ2SUZakLtCWoee5hx50o2PugQnGwCT9khXHGBNwSBo1cn3k
wPaS1G7sAYhzL4YVSj6etQxYHVE/Ig6EVsDiomGF2ma+ZnoO8Zq1rSkGoOgY7ODd
XQmz9SqxXpVIoBh2bI/4xLxk45+9MFFjUFcbB74FIZC2SOTamV07JIl8S0uYe1DL
jnJ4YMAsVPbW+VONBRsxfYevKdB3tDV79txxvTezJOgpDfr//HV4ouspEjqDgTKP
n5IKTi65A3Zrngkf8SFG7buf4wH78A4QY7st+YxNmQ3oGZs2noutarxsn1cphFOO
SFhEI00YqZXeQtb7xlCEYCV781a/aEmB3wLABx3CejVc8AgVeFNS7qA82OVX/2jv
BKYTUEtKpCLuU1wjkGgQjXILH1LsalK8icfEGJ/ldfxgGhj3utTdb02Xsi6QZT7/
lT2mknqdS1PnVYR4IX8dXuK5WexKuRKdudaBk7h5bqEKPtBdi/GH+aaGyvy3kY9M
mDiwHaXvuTRQsssHcXE5NO6xuLDtO6VpA8FC7tNELwe9UKmVOA6t9z2r18Cas0sG
NYp/Skqw/KJHsdCZOlgCk9Z+imxedDIu6ds1Z1CB0Pe8FpWSFxCpKyBjnvnXt2zk
TcH8D8KZX4L5y0ct/+/Q8iF6XFgvUYUHS8MlA7tsgXRcqa1lXd5eQtDhUio1/L0K
20M5Ww7gavjoZbU2cj5g0W0HR9DBa+y2Bgz6igHG4j1fnRBQqpKR3khIBjdmwifV
prYp7PKf3F+vHZQN8wKfX2/qLPurhD7i6H0IbyPX2ZQWe7/W+U85xNGNN3cIbVj+
4ME6kV+X6iTUJuQd4HlmXjW7QfyBAayOkMCHkTeroVnc1TmKmUNqUbboUqe7oRVj
xgnrUVHaeL7V5tvXfJU1aP887IV7RrHyHs3qnHuTVQjrSBjGSiuwx/23S9nERmZ8
EGCjWGtPcWrOYFj/7BOlUhW6Br1Td6CJXZfbG/W+c9o2jPCs6BT7JaDxejpRUc7U
MxkdOeqIUnpdV0dAkriLwi/jd0bUeJa2N/7d+V7vZALzq+Tyrbu5JvluMcL89DQA
5xqFurBQ/iRFZgr+a/iGcFo4b28bYnT78eE35YBg4impdZmuTB1cnqsbdmmO0OJU
dzzh8FV8EtJHgO2dP9A2EbIs+4yAbDG7nB7FQon1kHT/SQk2pLmk40vhHMawAM/U
RcB+cnU0n6XUe0/mKB1gtpCAD2TBQCTwaAt9BYL0DfIgW7t9bMsudfgI98DxCXgM
xfxVnWF2DHj6AdrHQ+YlKroAzLJ/iC5UFeL0tSoOtxi6Mwwnyx3Bhp/R1VH/7Xfo
GT4g6Rz9tsIt5wm0kgdUHTEXNtVoD8W7GR6Ygg5zAjBJ7Emmql4hRHXbsTzTQTRw
3i8mEEa/htdsS2QF5l3MRqXg/tHS8/O59+UQj1qaZDRoTdOgWiV90mBDtx8IMis5
TtJ+0BHInl8naa+YU2532pzrygXugWg92+Dg+68ZpyLOmWZM5A4d1e4IY29yReAI
/swihcYYqHQPHHOeTdg5+Lp78UKsCll91aG0P7e01L6wdei2j4ZHjw4M88FvuWbg
KV5/DmrMFz3jh7rPSXWRqI34u5Ic4OeRnajErTPIeG7fmR2hmPiLmcy9cNvf9Y+p
qH8FI9DXKuVQXh1gM0iJat3lUSX6diYjQ+kaDpBeX3QfAS3vw4gIVQCGejC7K0nJ
ITiKQU+Bky2fhKTkf7VZTCJlvfwjxO9DBDbBZ8vYUFUjw2JhEWVjMTXCaKyKbSnS
zL744TgzqSDRLI3Sh/0RW8WfZ2c9TWjT9nCJGmageuIYJTAGoDPAB94pNZtjA5aQ
YZaB3UpdIiJYjBOnseF0/DFzqXcvnmQMcZPn8+GdDhMeaF/sef8iU9CaChJVMNYE
M08zZTKKtWUIGOe5MVf5hPlN4LrF+YpAPLrG3MXAkSTMdUxJBN6aYyg6H2//zBmz
eS2vMufsnLKS0nf7eywg2Q3CfUL2ql96B/8I77wDvMBtM6OVzebbdrA9aKLNHQsP
F39RK6idL2NwVHV/C6DOr/DJnqWZW9gJkcWqXMwh1jOh5LENa4GHKXSBiFBzgNVs
kP+0uyTFYiVUUrVLRI7pb5aqlUO0QVfplxZyJT3rUasfd67T2ndQ6dx66bb8Z7om
Xs1CXmJXR0k++o89eB17FkWxGtB1fjHg5DXXdlmQYUqzM1ypsS3g9j3r53KPplDm
FpCILAXGLQSaDGZgMKjsdcKMbYcjWqk9nMYGRcFOfAQm1d7wtm6IP7vHfgI0DewB
7+ZBnM7+eS7pXWPbiTsnzC+l2oAey9P4a7E0/DHWVQ32JX6bGdEqNgpaE4oYzJuP
iHiG1oR5vQ4MV+iv64WyL8+Sch2YRrwBfrIAJzlPFIbUMLUz9T17kTQroC8+l3q9
U7yBO1G7R86jLU5hFfBwRQ3cjzK0iKx0xAJzeXKeyBMnwhKEXUlqYocKd2huvY7O
mzY17Je7Y1tzX+rrI9AGqsndVj4Gy2wBVU40XEr/a/W0sZmUltBBryEVU7wpeiFV
8puUJkZBhQfJwGEThVlHHxqJVZhNcBT+mJdcLG37GrcZtdjNmkDk7ifUNy0a5RFz
Ssm+kPR7OvVRIq1Ovxe44+dygtCt/8CPxhg2wLWMfXgV5Dm3wchWudJ6eHvQaG44
InPOZxmvMKa3X3t/4BF64/I1Ec/9j5/saxqLOz0IikK12umdNEWUfbnir2hdqOds
VirSEQwHQfHmZ20ZdY0pm0BZpyn3xhQyqJrnNR3PRNoEuaxsleAkJNRR7CL7yYE3
XiobQFwO1MnHxv4V39RLv870cUtWzh32mfT04auiVizSC96uDlQL/dI1kiYuy4Zj
syb0YlpfXeecaIph9/G3AqjYZ8thhW9xMETsRhTR7BO7/lr5ntRDPwu9catCeMCX
W8yhNUiNo5mBvfbBG8/WU+ngryfqBcDu597e4utLzCqueFO2RfRwzFgLO+S3+nlA
Gbz6IWlcrZHAIme0b1cNFJ8xXVgY986FL+HC+S5SnRgpaBvDA49vymPU54Xv25C/
fPh5EdcQMHuY+JOCPPp8Ydu/HMNTiv9/DbJQ2BPFXQJZUPQ4HLkYFI4IkMhsCiZU
kuzzrlL1mqFYpJ8qqYrIE3NHTldeiCPUMn3oOJ4MyFzloA4xChmOG9xGmwxx7Om5
bSeuh0WwGuPqcKga4OZ6vxCQagH/rcdLQXW7KjBjDYRoga3+tXY2+ITQKBOidf6i
qNkcvWNPNLFG/Ucw2bST4COxpWWYxU1nOac6kFmApBfRVq9b3EVKtz2XwVPOptmJ
WBeTRBuZlRKBotyBuNNlf7EXYRlejryDMfb2P/zzBg8be1wfroRLrSxqiASO0Ljo
kG+UE+nXysSd3lopFZOtGNlLncNpH+mv1E8TsYtV2WbDUr3ZwF4Wd8fHqTD6Y8CL
aUPSa3tx/uwvyme4AZdW9ia6zE0XKfz2OQatYugqSy4eUcBrdC07u1cO3SsCgDLo
CWDHWa8y5GXmp4DukSaDnrGI6hQ85cMq2Lmw5XJL1c+5gnrY+Wp0o1Ux4ZDXUf8y
Z1zYK5tB112oxEKH3aSU4t3GxjIh1NX+umjD39j8xzL1C47OiM6Df3uUvSqVRgLO
JZUHGH/cKKVmMxZ+IC+ZiYWpW9Qq+bXGmOgwDqUQlllUlcJhbGTzTjcL78rRK/Hu
oUBHaCVZteg3n6/8X/GxZStJXnrMY9WRmu7l/2yqRaJZmQtvadi++yZZekJmcjUL
s6LxN6PMWrizPDPyrXl/sgSiGYuSssK+EHvHhesOuOeiAqX1LiKJ8vJ1Yt+RVJ2x
2GGSjAweJLyEOJRNy45EBLJ0sZxAiPTR7W//k68VIG3laiUg7CtkxWY6WHZX9Qyx
oXxp5HEAY+FQYRvjqzzbBkUSU9fVt3bob43h0BrUMBJvtwwcKK2iNYpJVsANUmmP
kt/KMltBnvWOXetLXq/FHlmagf614EZ/QqxJ/x0g26eusr3dAKFQN/AYvSc7mN6v
RyojGVy+AGGLzms4uBg6tpLAXENYcyI/d/Wcq9YEebZoS8PGmPh5kVU43DxSR/uK
5LMQkZI8hlpPluy3Wm9oWZ0aW3RO2whPY3kn8rWLWCOZGRBA2DooRQim4vqwT1S6
KT2qrVnT45o6VOtXbtjeRwkBubuwVex003HN5Z42hSxPqFGD9IfH09oJ/uyv/0YH
zuMtT7RL0QHqGKwl40Y91+Fz9ZPW5q5lFtn3CKF8cLD7PWlp95ggbnMpH73j3eo4
nLs3VFUi+3kC59zi9WkEuSzQUDSuIURhIFwkqtWq6GTqI/JDJd+HmeGsYk4PElRB
KwTUHd07dq5UKeUnyY4PtosXU1mnDlKs5cpZB2wsQ1VFkawUSNoBHMQ0KCH5k9wK
CFW1G0+7a1ooMvOI5L0I9lUgVzOTo8ZoJzuFAhri4GcclKnTNaTY/8fJlGlqfe7s
zMgqgTuvl7VShGyYjNHCNQL35AtvIf+F6VkD1VhE0PCaswf5dJrHifAVskhFpoEq
R/2fu0OHs6qryPIcqg58oHTpACs4eIX24QuZUIplHiH9V9ivAAM7WLvwobZiPK1d
lJgKnhXSao5Vtwdc93fPSfPnlByFSfUlPaxzL3+DWAF5dT2xfU7BpjXGNirs/iua
7BHT5DfbSNHrdQ0dQjjaDNhgse9VV66DM6mEU77kGri8rAUcDI67kdr3Gw4BOcSQ
/itkRfpNEWpOxiJnU5cyhZmGl6227/nHAuD6+QOyiZFM5AyENbx6duNuJgrW78Ee
dQm67AEWRzWr7PMobWIar+S2qVFwuk0iLfrzJn+oZmZaYQ17Q7DiMeczNOu4DLvd
dkl6yPKiONrJsXdo8Q6O175IvhyZy5s/0Zey0y/X34r8QJNHKp3M7a14M94kRVXC
vdMeVzUZaUEQPJ/UaPnfwuQJxWL/e3uf4Rw6BQd/eOW7wCyzN4l+wBMbgbJcUlea
3+IIh58ScO1/WlLmXTgocmEhw6FQt+/LbBHoUtCLrzyDFH9rKTJ+qx7hGGjs2rty
ClFhNJsF2GdbbGRNigjMma6yOu/wllyLy2haSORaTcbmQQ63ju+V4ho+lzoUbLfR
V+nFjLF8CWDjMdMU3N3JKWTIenGWOaxwlnquo9EH3vI1/5LvmPXo32MkIsMW3+Xi
YwWRF6qRW4A9leIrszsKLmpd8cliV1Q1DK7IxLNNWpvfeG1TLaQvBLNJZ4TejDne
EaBMn2JsqBymle/I2Lsg4tTKZLtZb4t297y279IGB3nRpa/spW/ihOPSSaw7eK0q
It7b2pNvkddN4NYYaIfeJ/2xcnTHS/KoYdcuaGgCk5iULsKSi4FY0cYAy1Xd8zAB
45I7dHK1+hfpUFic42YfwqrMfggdrzFkx8Q0yWLo0Uwu8+nz0XhH9HGGUfKFF9O2
Gk3pTnbooNvRXvkveQ9MDa0AyRCZaAMW3bw9KG33w1aGpnLMi0Y2MgjyTa23CdAY
Oip2AHVhY2bQAa5mjQxvnD6LLwQfwK0+kiLCUpa1iWCXu9pCgnPKfQeEd44o3EyG
uQ+NsjyQMBsnU4xbmz4xl3me9LX1HKuNYbzoRwvrR4noLDtJkUjV/p8+EA30knKt
F0dXIDCa+EMp4ZkyyCzuRVET8HTaYePphNnzpD5K/0Hnlq6AKgTKGqKLgX+zfKS4
xN+66M7oCHbLuhYLXoI0jUZFuzdz5MvGMWXyD1RWzX49PPtP8eEDlAwrxo0rcn1M
F0SddaRu6Fhf+uUHvkaqjPvNwy/ClqlUDMQaKVzsR26hDSJGq8VMrnR0vwxgSX/9
XnhbbSwVpoSGNmiZaTB+VQ3AZ92TyO7xy1tfRgdpFVVmvDlMfTrWvtVj9UCNgVmB
yaYmx37eRv4sm3mcsw7hbAqCsQwahqzZcHwKLcTlZDaYTDFSiQ2NCWejCU3ZiKwu
jSwynOHeGZNiTd7+ZJ6Bw59Vkw+9lsED+IWKzh+WMm47TjPH5QnSiQdWW2p1efpN
AbWkml6xnICL16Iy1uKl/7RBcZtDIWdO5APG9MqJAPdUp9VJ1YGEoBbBqGMdUgQ6
hNsDqz/RnUJRqoBzM97SOMJPHENYSz4hAfbgq6lEhR9fAWymAvwL8h2oXjs1f9x/
g6kHlCi9vrC3OF1vmCX5jq24pDUATc1iXL9PrIWThYsr1GruyV+pbI4ZkD2r+8FF
zHQs8xgK/WLyGbRmDBdni/UGcYTm1UQRfsTHyhclxiBYORY6/zpXeOUVhK2Xk2Gn
ig1YFCCfNqFfD2hmTyeWKd7I1rBwSnTXvinv7Xe3jxTonoENm3mKUG6LYUK/bEos
tfkeBE78gLDJIjxvq3h6XBQMpzTlB3ztBjmVMKzFoJXKAOVoZ5a/Y07YG7xG/SiB
QnxE6piHpnRXT8sBhjOc5m0RbIs9BP6T07cBqvW+7i/TEKQfPXMNp+D7Hi/OS/jx
3jMD13vcXRjAMCITTrUDmfcSJW2HJ8306rT/zwEYnlJ8IBhu7/7Ph1T+o7N6XYla
2NhiZnB03eUjD40k+o0JZBwoThVokLPcVKycHR41fjlr1dGANtunwJV0o5Ilf6tE
Cu+toT1M9qXJH24z9lzdSrZd51tt5NLQBd4uvtaGF4UTI5OW2GBcR7ke5hKU6x3o
NeowAjxFwAmrWFORGXKaGS58TT9COdIO3QPRtgZ+MbQ4ttfQXY9T3B5LmujeeTzE
rZdGia2t1GnSTnEmfM1sEYMsS42fMlGerG9G3ai/7zNuUQaCGdEpRkza73cT1K+2
An9TyvvIo7BFhrm/brF4Unh/sM+5XxJ99x/qNkIP25RIEK5y9r2ZQZyLocm7sGWw
rtJhdIlWCnDLuGJjv/HgjeL/YfYsbl+MRAsePZJItyVlZLLGIEawBVJ7+RbPpRQx
k90fsN53I3KVnZVpzx+vkZPdYsWHQtppwIEOnDYBGAho9oJpq1DYgbja3ZdBH1Fi
dlGY409NtXF9bYKb4F4MP+rGexx8XDMCf+8eLC94CrHRpyeH7H2mWsBwj6xWGWUc
usgk2D//oXLjv+hAbG+5nH0pA+oX6Ig553H+acNWaFHpUhKznIrpy7KhTzuO9U4v
6aNeoDC22wApU03sws9E5AnIWH2pUggatJJGnSOR3LAEi+pXZ/OFHW4LOigE+5eC
J2NjnVs9wTD49xLIJP0xfvA+t46wIqJ7UFIU7Mi7z2ytXfSuPLsWwMAGZ4BKeeu/
fnnGkWiMuXOJ/9VwOfJHsE6wITpvsuIeyKc5AnbDw5/DW5TW364/9N4IprFapaH9
YGi7c37XH3aBQotYokfWGxgglmNV/8Dn37Mt7LKGNQZ5nasL4DWct00PuNXMo9ZV
T2s1rhg5uY7SCuvP4YDXIyF5pj4VV/HRY+JRBVfhCM4On2LM6UWiT+pRSEPEJM2G
qpsGWwcuUqn0c/eDz30PGpVi++Am7/PlURM51yNslnIJFb4rPtJOv5xqO4SqPx2g
9ZLmaHYaf5/x3bZCGgwpRXh4SGLHWdCA1pLqFPIzODl/9GIpiP0cJ5pQOJZGUxp5
+xUv+qa5d9AylysHdRHbXvU4zWHENJslzzv4NUd2l0f9Xy6yvMM4wr4Tg/M78blF
IpGAvYIhCgrnPFh8JE8mHtG7KR+FI4NRcQMN+B46bB66IZz4NngzmoQi0m42FTyd
cdXBVJ9bzdDHGgLjPzegbJ+4/+nl6N0ZYDlbjevO1TPFnMsZgECx7wIjFbRpf1BC
iuhRb++j4mzGPvpHCtFnItImcO46vNkSURj6XvFR1kbNx3hTbRku1umRo4y1uGs2
mWq0bRQx4Vifuz3tQV2QmovnocWzeByGW2ItCJdiybalk76B4zJUso/BYTlXgrzF
hODQ4A9kIECnXdpP0JVkT2DiqJGLM70h9AV8f2bRrcuJtsRxwh+a3PJGPcoaq2lM
J4zHoPmvfFoUNkVNFgFKoixtn2pI8RFTuxLNBcBVDuHXIO/adcOb14zJShHzMz7D
9M4i93LPvHYpJV6yZkNb8AzIMtmCTyJXIB/CV+iy4wM8HvsazCEEfAleadTmAZQX
2k1q53FiUq6ccT0d7iOV3IDj2VAOkJt+Kn8HaaT0yW1XU4wQHnvUswyKUB5fF5DF
gtjlj73AcTmD9zJRSYaP0qPZMhyIC3yLIfxalXuePpdqkxyhLP5KLG01wF+DEreC
RclAs0UdQiiQgw8GjI0dcWyRiKrYLOBCkMktXJs29N3DFyq/3oNpcHw/5nIa0DyK
FF0q9QQ1PCkP3S5RyKiGFpvMt1utBsuZgQ/l4COF3bI6lkzzq0XQUmMdxpb5FCqp
KiyQpPOs8yo8a9b1WbeAF1C0jZzud6mdax+MrnmkE3lj1NGSfaz310K5I2xkqH29
nSKa6EzcQYxLHh2n1eYIYiDhF9V0jALLm6Ly6rudH7Io8Yu/HNMHNfpeEothvN9C
jqRSqsgAuC0UgFhvNkr41j537FEWC1c55yNjODCt6p7JxbkhWRYec3UgYVfxyamh
66iFHZ3Q3GLcLl+2dYExuI/FIih0UE4u4miAvqy2Q8aA77ePN9Q/wzL3cPgvqgMw
X3qrGbSZZDsQuvMxj8kNoME/m5ROmz1Voyamo0gzI/9Wq6DBYgZ3yhMhlEzgWArF
Ff7qear3As1icVhSB3pUp8kRPLWdV+KaNvU/AWEk5bMyzJpP3Noosr2lwouKWEzl
58VGsEyaZUDgH5ARYb6mmPLQB+9ulNOmxw51Fk1JhHEN/Fhmpen+ZDIhwcdAEYQU
8HWjOJZSkVzPLE6PHafrhXfMUTNbjHu/eZJ+al+BMd+CEgX38dkruV8HZgIR4Lvj
JUIZDbgQDuFTervU3Z/x+/IjzXbUexwUausj1JbipIUOWSQZ398qcHesZj3XtlG6
2nQtLgRRa3/LOTql1QtiHPrv8Vnxr/3gNCb6OWIuUa+EaRPHRPQVQyiowDs3CJ5A
9xRPQq5iL5b0bPSjyixgGQSyHN/Hpi/BXrQHKN4WQDUMZPBpQnZZfVU3wZv8UZ70
JtX23N8gLSD2t2O+3raz/RUXKKWQ7lsOlCNQWcdtbjuFuur9MXbhOxI2AUZV1Xd5
3/ek9niB74GiStAj8J7s/mD+uqjt+7psXLnJrMckAmNbiVe0bxxbE0Sl92yjjH9L
j0pAMMZpfLOEizqtN6k4xmddXsheYIIJEAXpfm9Qlv8Nc/tUUBvVEDLOkjAldIoP
qoVFUi3v23PsXADiw2FNNaGPT6Rzq+znCAaXwsSgA8wz6tXIt5wvaDudb881GjgV
fSnqqBSBAytx1BVhfcKMFbFPULhL+ewJPCO4s1153Ody1gAxZApXWEc3UunFi0OR
w/AYwEs02fyfQZiWFxXHuIMBRcEfkpIqYK1iHJd7YXyfKmhcdxmd1S1Z/NRZddaY
TP7O3pcPBo8RC0M1VhJ9RvY0Oyi4q6k6sHppnzyhucQxQ3mjroQIuWMETftACnGy
IeCJQXgVrVwlVhbFGbgFWSZBpOKl66/+1h2Ssg+3KiuGdqpLMEzyuc9SdCmCS7dN
HR73F88mlypU5PddXZux/ierNUGxWwpbYfAhNBpQ4byVqRqqpS9WRJn1zzlM1RFY
xducdjQbmiXZKsweDWQzNBo9/jPZnfYecyxnFpxLiTkNfY9T6OYlnfX4T2b373Wb
b6biP25gMMnUFuxjr9WiODC1LtIzzlZ6tWLRgqVvgXZhqPuI628aj03XIojWwbxP
001NjPAwVsh3us9l7fr6itEBB5/4wPAnOW7WygiBjElZCG0FgdUDK2dqL5KEaUEi
SSCIX4j1U/dpvb+FQOEBLZTlW7biuqip048e63CCwLs4yd2O/PY1SZNvUhdbO9AN
DBGSqf73gkGgXvAaUQt88iS4n673BcautBC3gxNQ0C8kugJVFrG1fRu8uLmszzbL
92CGSk0KvSquiWIubBSBmuciNW+gDb/lUbZNRTl0oJ2YC4FgM08McR5eoOacTxvl
Wey+D3VdjR5wBa9KwCsomQBntmRe0E9crm17cgpYuHCEyvx/moNlG1LmvJewniMd
kNwLW6dghYUnCgMlpxrVEZvO38jV1MyDt1yrrS8wB0z8Ye8vMzHlVcvXOuiABcpZ
4hXxxDii43nv9sxPKwJqRQsKA0TKR34YJ800RJgcN3nSm2V7Nbx5cEfnycAQcgSa
/j/rPpS/K/gnGWbh1rnX5QYpo2uqyrxrRQ0jrbgdUCneWqibUpkcDzLqsgaJ1eVr
3zowyaanaMB8bbzYjiyfFRFCLlcdpl5twCuK6D6cj1kgNk39d77t5o1ijxjnDuHU
p4JGrr6TNhOE3hT+EJghRfvPZuI25anCWAnQS3dfDDxECyKkcu0aWcD83g02aCj2
u4Bu0IAKht2u/o78iAKLNECqUySM9CjJz4X3EPBYes6h/mT+mRisemAvJx6s2ULG
s99cLf6zFUJxo0A7196gzhW1AkIOnxoscda3ms4KtOeLQHMnFg+2hD5FtkcvGVRS
VuXaP57c1fXzgini+GT7gTTdI9FTE0dStEcZc3MYdgVFD2d9rmG8Eo+zMOeMxIHB
jAIR6Rjz2f0Am9pZY104B8HMzWCkqvTnytwgeMvgrW4QvUksZ3eq8ukmJwXv0OS4
goDT1wP1mUktbe+Kq9Ac7LAtAWd7y8mvjofjYnvyPCLgzrQ0RPhRvTEN/Bj4WXOB
hOPE6Ql3NqznVosyRXcOcDRKKO0rhn7KyGsUum7F8FSWUCJ/Yxf+nb8flh16+fCn
JDeKLk2Y3Tllxj7ieG7MrqXQMbV7r9pQFCyXRzS3LBfg2hMRRjGEZ5LkdouXS0XG
lvuRKvilQtL42Vi1fcVQKn78Zl44j12iaIsGGuJOmenQw3d0TpmiKOZU6B5CyJAr
pspfgZcjZ4itusTZhktc6euxtYNU9cgEtxG2DbyVWHKy9ei4kaDMRxfkrLQwtV0U
hS4Qib5CHqKF/jkqHVRa3LkkpdhKEB/m/garp0ki3gg31ZyYH8A2kG8ISKsNxB79
cDLDY5oGkVOemEFGe20VnmxVXJSb3RBCdJMnPGMUSrylOIrG7RwGn+mblZFJefBo
IVDQ3leGGf6FaMwF5FeffTdXgHdXKuyzfd7GG4bBkr842nHBwLPIDT7MPxsvEpXC
GmHNlH0BNQgXkJCS36rsOQGBXxHtJ4oyXp3pk+/iXjbfhMjA2ITcmWVfO6WESVOR
7xGFOo2+3ZgmPnv2irpgaAG4ynVYXDjt5rdFgC2if2FqjXs1OVWhFgHBA+MdDILH
/OiqzjQ7iEHlDIIXtZQfiXq0L3r/1kuyQJkj5HbVb0NYQKN3mCSaRJYyzpyy/QM7
9Ga4ny1yQh6Wwb9nOfG7xNoKS4/VFcOfos7b+rDlB1XgVCYB17eAIrw1Xv9Y2RxU
`protect END_PROTECTED
