`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9hiHaEsg1sKFeO/ih/LT3XEFyUDyewCBcasc+AfJ30ENKH1jRUEDODsipXi4XEfk
rKSeIl8/2ZAwIeiUO4b9b9a0YoUbBS+BUOcMwzkZ5DRT/UUYLV2YYHoA66sGUNzO
c9BLhfWmOCYken7/RbWXJ6pVIgnr6L4oO6BkWAMkkU5c+j3dJ2Lmlh0/whouaLKU
KcuPELBTH3em8qnq1dNDOwfXcUXfRaYJvGNGZkdL6P5O7rqif4vsXeYgKvX6ViQf
XT3D6++AeLLp6RcTTYW7iqQ5EFlrM/AS1DqN9IZzIDwnufx0FTDc7k95cfpntrVo
UncLOn+nx5sPpPmwanHM1mE4tTvXuYPDycLQF+/N08BPtWekTmp7mMipblrvNpJL
QOneR7xjjnF8gdX489GpoJ5AYy6DpUD4A64XF3kSU59xGeZCPwqBsrqaipNnGKRK
Uig4LwefqdGS7t2C9DJObGROnWGZYuvtqeaf5nKmyHpCRFKI4b0hS8WG+EAwf1fO
yZ47P4o3B+5vKeWKrdURfwsCJEHYfKu1r+oMB0yGtzVDQgMkK0gGoHOOBeuchQ6F
HabjqhThimY8sdWmUVAeH7LsrMm0TLcaq+pF6ZN5DbHtWRPXzB8lzf3jhna8Kltb
mqx84usK6FnNwcyMyikNUvTz/OL9y65HfZKok8E25lBqT5dyyu9o3ddbJmJbVOY7
c1Z7rxhMAVlfSfQp6QXnJfBNc26LjlMWHKg6wTTniHPYzLV9HG/zul56SQ1ZmZun
n2QfRbhGKy7lBYME/Cgzze1WhfEvi+IuBklR9bDT9a3T1MruMyQK1fSWtOY0cmuG
vnJpeqtq20+lTeT7n6WaCetIuodn9UnuNrLk6b1yQKLXRXXmHHcxB3CFe/O5+AY5
ipaQE5LU7vbrnmnI9OtGHCQrxZl58sqATj7aJJRSpPh2N/JjCoB/frLjPbnBA4uO
jIeTdyI8eXc34Epd9qYXzZNPSnRJDjl5l6xY2+c85BNFAnadHOElqN8Aa3JzvRBI
LS0pgs+TV4IcyxEEsNdixSXsaEVrnpQoWmxNLDNw+OWC/xYcE7iNjnZLpCO8q4TL
pW0iTFklEzZ90SbarQTjJzAdohywrq4lRFCtN3wsBT8L3BxLrmjmo9KAgIg2LdUh
TNHLsJKE108Mrm45IKj6oICUVZPkM+2bizJkjpqk44w=
`protect END_PROTECTED
