`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zVaZAH/np8vwF1GywVjKNT9BcUgB2Eyfu2kf8bMTxCZIkX4tmQ3+ceKqPQNfY40Z
SJGo4rJflnePg+9bDSq0m4Zar9SZEdD1T+xEonJK2ypFQ1uL+8swAVh/6KauMGve
j3ev8KVE02nKqBOYkCpZFz2/+cxXgeC3ezcxUoElGPF7dZREK9xu7jbs/GNrmZXk
xGhTd8MZN8U26qgIYy3m/VLHklm6+1zg9dzoDEJAG4ffMqpwIFu5w8RgkNqo/j8m
TO2FZuQIgC83K6uLgMRBpV53yhJ0rY4gDDVqlN6yBxPH4MvII62spdXoZVoKvsoQ
onKFc5ecQut5w4lmELkRWaYwNYccMqWWUFuEr5paDamQvPCYzm3Zss9HBm2DeVn9
ZmWkl4zUewqaPiuUh7L2VpEnvTPp+bulsvlBhdizhJtiAB4Lt0KJPBz/B8ocfmvm
VGt0Y60HFlnmG8kWxUKGjLxMB6hs7S3edwNWpq+6vT9OAdtUh45cbUxx4OTrXro6
MGs4sipw0iJmgYXNJnjl45yZxf7sp4YT+plEsSzoB0PogifdqimGsFJDVL/Cfu5o
wVscopxjkP5bSIVy6K+573tvSMX15vr1FzZMBeNeoK9+YxjXHUoCWBO3KwC3QpOP
varqx+QbEKxr7H0v2szIe0FGGFra3A3kMktM5T/Ri0a+Bq4fZoSCxYQrJ2dcC3XF
BV/MeF/Cl911CLx7R5h+xIuacxGpUmFtfsHSMSpujmCKJioZ2u5VZnlvYWhYWUXV
o0QhkjB1qfGOVUMiILhTveU3dLXLJFwHzjPKdsidFl8RdvvNY/inxTbWyk/tzFpL
0kJL/Q7MkKRe1j+iD0h39P1AjyJLiqsbIau86O0XmOXHJr6xjCRlqNYMJafJk5/C
rsRPK9hstoAzEUxT+wYV7A==
`protect END_PROTECTED
