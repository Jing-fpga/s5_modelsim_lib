`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iMcIdOTCYuKDbx036JwKLQMpdgvbVjKjIVVgzM0Xjq08BV0Jbw2o3/zFoFjMY2xM
PBymEGDWn48DGD0jJ7sDTyhAz8wyR23AtliTSkXFmQv0TYEFihc9qa11Ts5s5KSY
4w8Vh9toYw5+idcWdbFZtBDY1iKd2EFnjHJNNqo3/J/58EoriQ2EjKqGqou+HU6d
8/Q3Q8qTafXkL77606CCYiWWXmluqfD3vQ6v3gpGaxLyyJLyAInvqEAocJmikcqD
ME9VCUiatQP9RHxSYum6dlpwDJ3Rv3RxEsbBBJGXb/pvzpHe16Ey+XKHW5Aw3OER
LNU+TsM701F8Ihjy8P0kT3T0n1kI+yoRiU7Y85FkJagfHgM5FBXbr7+5apmo6ygp
z7+o6kuyqa5caWYRNR8H3/66EdnDFYffkcPujXcl+GwU/Zy+AiGaMGk/46EEJzGM
wpJzCXPzWSgzFeEh7AOiDTjHb4mZt9+wxS0FrFS3Wp0bpQuJjX3i8yH1mucv56ru
TgGMwxCC8YFf25Vza6xBSrmMZah8W9kSNVdcz2p46bKbcII+miRZ/0k8O1b7FJrd
W41GguQDmhuknyWDK/UPKpgwK6glm9A2iwny5uuQBLwKKcEoG27Spaz9O5k4EcX2
qYtkOyXNtFQQZgA5jTyj0p8ieE87bS9quTxkY05bo8B5hiTbalCLPAlpN/lDhUih
jrqw6qxGJSUT+QBG+YyjEyLbekJ5HhL8JvprSmfIDPPzprLqKsXnUAascnccDNoH
l/jQeAHhpJiLhq9o2OoXfhJopvJjx1B/fJlcyQE6t0AXFgtho2iBo29YPbkfivyo
0voXrjvVMD3PBHKpNEpk1Ou+BjP7x/UYKdXxPS5loh1rsrXtGwOPeJGBQTuBHaBc
1uS+notag/f+uan18qA4CxOj/ct9eFwSt9s1X8k9Ig0xS16qC2rESsMLsG1iu6m9
DUKfZgMFCPI+SO7oi7ilgfP0FRjUvZWhSdbbSqh6qnQfRdGIvaoNbLkC0s6Lkuos
1HgFxH/h4fucIdedK5gdzo69mLyKcW/KQ+LCu23AjXUxqIYJnBRhCIasr+EKETwG
buH8dgYvXKub3IeKHwcXZCi1UsN08Gw22n152sfv5Pk/G+HRuYX5nZuVQUkswfmR
VJVqmqkBSA351eDcN3nvo+CPFUqthqcBg9+C6kH1ngcsaXvCQV9HGWOo5PV8xkv0
Lkx6cWhh3CMxPo+47sQvNFnLjgzzXEB7E307fhtmZ6znWqVwPi5qsV1GjixWFiWJ
+z86F38igUz2T+VhNU18WJDAWoALytUaaE2cpFC8E0gl6S0lk1SKuC1+5Kv1pskL
TWgVkA6elsvviHNQua+VzON7XvYb3TOTX4U3RW628X8SU8wKdlATjvZcWZ2/bxEH
rAc3SUDgoBgqTRyDRVFORyjBvoMlaKzMpX8ZkK/+GQbEHZQuNDBONI22WsJDxYiQ
EwGuXuDLKzbnm6CIpjSBVC5JVdgvH+noXIa3AiqwpXKSqF8uOU8AGv0lGDI3TtEp
CATX9gQe4dB6u3Pfy+d6JRTNMQdAXwmZMEaqiWtTHRqNJo4SyfOYXh16Vc22ajy/
7a08LJXgROE2cT5+x2MXlVo0RmRSu3RV7kVNbYEgY6Qdhz2KvOkD6lDvR7geKW+U
Ajr1D5RJ2j206VUZdr/u32fvLAJVLZIc1I0VD/obuUlkiRRDSemlwdspFCPMNdoO
bSpXTB+LL0+trFhHU5MtM4zTjR9/GQU3VRr2S6x93wD+7N/H6YL57ly1IQCyk3MP
7A/ApoTTBZ5/3n6oFGlVRUYzES2dSMtWM4NGK7nwq2I/W8itddUgQgCMZeUNCVIn
UMtOfKB70rlLDf0AO3BByQ==
`protect END_PROTECTED
