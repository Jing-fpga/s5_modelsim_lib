`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HyfciJ8Pv116Gnd/k584T27CKFajaAtyKUBlt61JI1kidy05ygVp3Rgtc1Hs6X5I
PB3gArCvWbyqFN5FEgkvdWE96ZwTvxOW3yXyugBCpm88zwoeXwunt7vMAPSM0hLD
eZK07sWnOfyC4LP+AId/a0RCG3S3vHl6nQgjvlIYZppUPnGr3rdRKPUoRbPlrQMr
RYi4/yMqQHTcOsk35zo6VUJcoGYJ8mtQ/KK0mXBUYVGoPYPbYZeYMfDqwlyEb6u2
CYuFi4tR73nhZUUYCsYqjXvHBhDUvhjYAxTkuBMC+QNJYtreeoeMH9NadlMmw0C5
ahihG7b4Jzz5rZdM8SS54MIgbnw4jmrNfbAQImmY40fAp9V3Ewe4mAfAk+6IntZV
eNOhvwj1pDI9wxA4yb0aMEA1k7B+fyRxa/gc8aZdkcOK17JFjGlKIZ9FNx8iENMp
43B1CFOweyXmM0ty+tMRDoCx1tpz7QpesQ8riJZbcvzY5UhVQitkhD/7YWK2Wo5K
zO2nwsme2WE8Z87j713n1WCqAhp4x7jZjoAHoPSPDfXc0XNYgeYBBdq1qrTekGPz
oF+J9APRXl6Jq8orHbjvopDn7FrkGjgvly1AV4mNOgPv4gkK+8ncX7+r96IDmq7S
j8jzxbaROhAtCKwCi/bphW2Q4Hs0EUzyugNbt/SQGrhZYANFtql29MTFsltGYRN1
jcWCRm/04WqT2gCQYrRNsOjgUTEY0cpUWK2FicZoh44ENaNYVzTavOiSVdRb06FR
0Oy8yyX+bgS+RONkL4OJ641L0nbmDotT/p5xHtiaqkmOTgfs3/HVa+KohGhsZ7L6
gYK2reC0gtZ4z0qDhqEOHNGMRbfSxF9vsQDRNX+9Pt1fF0gFcNSROwLnSA4aSsa0
CW3M6pzGvQ0Vy1xHJc8qUNvLnfuOrVAxYfNmngtMR7Gq9R3r9qfTGYoQOUBOr1h7
BkYLICeXMMcpF5Kyozi7krnMMg8W59WOhs0XWc4OCt6c96tq7XT8g2Xy/nIHOlLq
DoISTBJS+Vpwirdh47nRwAOQohJnmlGCWwoROzICmxANC4kaYGzhBkbbgAsqem0X
4s3vFrzV4xatl9N4p7Zu6wy7mxQKfyBuokZXZxIW5jqQQDdON3HkjhmnDii4tpyO
x5JfjLWr6WXj0Ca/drOogGgkiYvfZSHPN+nF/hF5bNximrs4lDC321qEN5H5zOK9
rSe4N7RwmDjd0tErTtOONWvKv63fZN1rfjDNvHYpGBLP8sZKfZ4WJ69+gsOhoyrp
TevTBVF2jx21gjHADMBvGXbjxRem+Ca8ylsja6sHL4/plazS0hv8fPUStr4aTavN
vK27q2NExmVtmWX4iTP4JvHnKuZcDSjSp+9OcCkqgJ6N55Q9hLkflnYgOFjjHsYD
FOtL1zw4ExDcH4VMIAR7JyhN88WC/8YY2mFjeGk2M/D6rs3rxsIx3uKmWRDL4jnk
cCcMIglZWbLDduNA8ILBScja5dBmeyMav/2caeT0uEl+8fcj8bYhbeqF7WONjNO+
NTPEmj4Ra4NkmO4nev+gC34lXY5qA29DAeN7zzAEci9Mualad/UNdam6uZCORA+j
nJCOJwAv/dvdBRZywgrieFAzIAnDQkiA5rOd3qGk1XXZOCUYMTtCQhbVhL7EmjQ+
wPcno7IEVlmHAilsJOQhRuIzUIlasIOlpe+AtE1yk4UvF8mpEKWAXsmJuYkCZEiV
2tnhNKTfBM6TplxMr7OO4q3mAxKW0ZB8R76ShNuu9x8Jc2T4nHRQRQREdnHOYemN
hOg0Cqx7Sja/afDWDEEqR8GwiUckXjogFUTHidN4d/sKBLATDJuttZwP/itpS7oj
D53eMl2sDcgW3948Y9IMcCE2gMAGV9GQ9KJ94XbccWdpcsN/pB1iwOqbmZ5b3JOf
4wsuH6mbZoO1FJ1iqlmpBfFmQ3tiSPwRfaQkTV2/SShzetqOVQ98iXCTuCec0OkX
41cKEJDaQ5Jt25+7+Pv31vvDP7WDHybmrRvTjgBDUMGvHl2bbP71cysKt6d4SDGy
RHd4+b48HGPWxzfUkfgy/Qa244XfyqBSPKQWKnEaq3LgRZlXYLYKB/pwAx+PIZWv
D5Fs/2vM6S5HvWDbT4qzI+0w9zO9e7fWz41x+iaKuCfH9jHxM8PhOrG+Ie8CrRlM
4DwNucAZvIX7nkDehhRuEuk2perZXqH+xCc2KLC7RNyiPk2Iru2qi0B+eAhWrmX8
4aldRjjHv2dA0xB3cdgAOdYZENmMHhMbVKZXyOdJMcVI9Foeeuyi4aBMcVI6XQWh
juodAD/Za436kXHYjgBjhmBmIPm9XO58GkKUdQMoICLG2jzsdEY/Y6ghjra8kiV5
Js/0cG1H+rmuHwvhcRn2brxRFy/JS674BfMqm9zrpir8i/7NlvCE6cJIZh/EzfTs
Qi8dz5KiZG/bvP0q9rr/Y6NpHvKwGNnzvd8v9Y8FwNL6xn61QTD2ZN98ClG1j5EJ
+Do2vEIwd7ji6mA/NdYumto6iO7pLQ6fg9zl5CgohXYQ+M+8NPEKqZOJQW2XfUEI
uub/QV8kvqi/4L+zQVHYwdcL+W6JkrmGh3BbYcbTwXKrWHrSDD61PZR1E/c9Ykho
f6PX+cIMtsYbPQ22dIu8J5fK+JZ3G5gKyA5SlX8UG9TodEwNjdinfZwrBrteiVfz
PO5FDj9Kp+8N1aJLXzEUdhL1/YGkoFntdVU56aL3X/SjzNWdjXW2yBVcPb6BRP3l
L5YY7v61dp+WnltMECoqv/jcXEd7GfouCQyGGGoQ42wdKr1hBwGNo/GAZQ9Wc8zb
Zu6RXReL3jFc/BAIoQcgNeFKyuy/6ScoY+pXaBXN61wj8J+v3sBegbn06vYV5+Jw
qJno5WixRYbTxtPXM5xR+UBFHn0Z/bdw3/EjACLIC3zmkCsd0wgMRID8SjY+EKaX
VHB1bdBOMwjze3Bqep1I6qx2QG7/s4cV2SxNAZbLc8vSb/5uoLCC5vX8gSX1JUjO
DkKDAVZt7uvJ9o8oWpebJsWKCyLGIquS9Li+AkDQUI9CI4oiCVVFsmYq1UAABzyJ
wHWfBzM06queckfNO3hjXP1v9yuqrSV8Cmwq3bk8f2zYq8P/8b4m+RT3urgZ1FKo
pO2q4dybDK0tHXs1bbNk+QLlKLnVSpbNxva0HERCCeGlrkrrbaPbCx8utKP8WVoL
uIXyHQoJBql0SE/O1yxY11PuCDOXHfvydl1VnF60zTBp2NFll153yhzfwsYJPv6w
+CsxNRV9a3n+KS6RKVdULv523luHWPTEN7bc2qXk+J3lkQ0kUnslvh4IyypjjlFn
HZ6R10DX4Xr77wiTaDI7dwlJwkteUAEZAe5alObbpCTl2uiVFvc+LS/L0o/6Nkck
BDaGed2lTMdX+3TlE7p5YattVqIQzZJcmp5EvzBpNrdkrBeAkXdKRBeegAxT6fmF
Yx/rMdIJIYewa00YNB7V4u1OvgrS9VRp/HGFhz/ZfUHf8HRBAlqGWCcDjwNQaZIS
w/d8iBQBc+RdT9NfX59Ove5Kvq8wQHJPuDAvRHFlpqzV+yXOSh8udKBPErHaUrir
iuPAbt8Of2DjkDGItAkFBanNmPtz0oxU8tN1Ua7U6ZUgDxv8sUY7F/7EfpjWo2hI
oN45oPRHyHc6Dq/ZQI0T8fLrG/ytdE1Hf21SZXUq79RUIFE/BILleGk+GuEU5Yln
TbYi/8GzDUbXlqBMXb9D4EqdqPoZFP0iCtMj0cYQ1EM6vESKLfG9PBtvTAJkitmg
7xz8e/tPNxTrZWF69+zNEl78OziM8ks9oGBVEwOQGbsVddbcHDOTeiMAbmiMK0Yu
bQ1o62CCLGo/BioegCMavCKaw5mSO/VBRqeQSD9+nab7IUiOKEdJ9JimDhfGC4Ay
XkvqdBH8IlL484X1f8BrRvPc+QsbMJEPcZGbXqr3iHlCTg38Q9vUndkUfCo3cC8V
9eHd5m45Q7UKaTI4Rxtyam8YXtL/QxAVv2iupC+ZjASkZiymWwK82AQ0RELjnm9S
54SWQdaRrNSCfQ5bEvZciE/m5233qX51BNudxAOTzY40meHQ3c9AInxp5h3qMo22
6ATqj1rcC6NLscH1yoyGCIATl9WIer/vyZf6qx3+9jVjTZv1EStGX4YzpfQB7+Hz
DnbH/gbZjrXd1bPUk72FRS8MiBmFdnzNsURtM4LrS5WL2nutudHOdSDE+yJzb0SI
+aSH9q4ceASLLFa69JGTfZDmsOWvjDhUjqSlwR6HDjXIFmMlTX1l6F8SLphGRUNk
lf2p+wui4AyX7obc4T/jTmKpHWWiLB6RlYZD6Swr+bus5TCB/4+2yLBAitr8gxjA
wk1qqfqY38gSh7Xg6BDCBaDfvwelaLvECoVPd/2QAQv7vRF7Eeu+wGbihB+cDKkC
un9K2hs9bispOi7bTNGnomiMaa9JDI2N/VhhnzOKT8s=
`protect END_PROTECTED
