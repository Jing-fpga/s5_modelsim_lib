`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KcKD78n92nud6GCmg1FxfDhVJRKiBx+9KbrIbWqor5vxd6kfMBqOv8WfLtWgtatq
cJnduALB907xj5vjvsyGMEoOEx7bndEMyOkFBz73uoW0psyz3yZeHKxrcdqKIwrq
PBlHKqDT3nlJxb3ow8rGVTTDV2qMifKoWMH9e6BiO1MmSb3+JadeE5Bx50W+26ZR
/tLYDNFnEw4/0/MtExaii+o0fpI8L9ZPPUObs+oobp82Ghl36SwAK7b4OIPCrdWz
w7BU/bGXGZusNf07dNmh+d0RNR4DiBESr+J5dLyjh6nXzqWS+5BNzK9jB1N9bazA
SIFWA+vpoOGd7fXZwNDYSiwQeRclmiYVP7tQTOM6S0HLkUAYQAWP4hIi5lQIMiM8
6VAlQUQ42jJhQLz3ULz1afZRAHWW0jMJ7kPGfGrsTmRRDUDu4TIcPbKYLqeElKiO
ji956BGsBV4nGGoZs44BWMbgJvkaktxrGcn455HYJYNy1p2PgaZZFkwcSTOuC3R7
4hASNgJyjGqgylAqSch8RH0wPSE30qBxGbcHpiRvaiDEK7UqtOpZE7DMh0zIQ0uI
fim3v34bs/ManKWjhO8p8LX3+p4HJqP1ZsLRWjVjm6Wrob+QIcd9Knw/XCObPXin
m6xCzxgpx1u6O3WJz9KZMFkTjx3JaBogRcLEhCY2S3n/kCbdRtBnvCD1XPA0F11Q
jez7afx366ZuLmS2pzA31/QN8YG/FUFukUF4szq+raP9fXsok+NtlBIhZ4DOrc5A
G/GMCzmz3mZveJTz2JoR/cKfRS0FId42/d6EcMgi3TlU4GPXDw/QnBIwC3a+o1Pi
TjHyXoKPpHLOserDFqUm9lJuhzf/JnQJ5dq96OthLEmIJQaTUDDjLjpWs/8vPhUo
MVx7LvbTepE+kuSjqA6RBt1vvAhW99QZlMYkx/h87D/PnNapUnbeAXQE/eMa77c0
pxb7ZK8r1pwB/ROmVMd6ZUlm6DUcxCElbZXYmrWU6nHs+XLKr7f62vIspiksaktA
3Tzr4m92TtZ99nZneCU7E1y6b0azIUExdgH0Glgw7Qyv8pUxR/gWk9DY0qUzrOs4
JG23U3lPV2ABY1F8zhuemilt5VyRa74hjXx4XSK9RJXmGBQrF37/54813TfJaA0l
JTKDt0tfrnHFRostslsMRlpAKpyOObVwg6uU3IDpECrzBftzXWAFxo4oiZR9VwXu
`protect END_PROTECTED
