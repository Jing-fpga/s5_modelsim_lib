`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DM9D3Y0CxdXNHTx3363odmAOgvR0mdI4fYJcuEoBuMHOtt11jcL7ouxWtQQXENgI
TTA80Z0IJIHoVd0gOT9Mc2ktsnAvmETSLTpo3FVO++u3IvE2PtCCwCnqyplKu2wh
tB9hd5vhYiiAWzKyX/NYNCX5eWzur2ivd/2XsQePc5urMLnxyFIkGwNEmVbLe5r5
tj/m0OcR4Bw3EQkzUyoN6V9ylSx1KiGGobccOLyFAjfgR1Y9A7s6hc/z+a4VNc89
OHFyXyJB9Fi6OLJlKzyth8j9c9b8u4ekjdLKmQH9QXwH3tPx7nwiGXWcoL3s/Nob
dtWSnT71q1+eOrL6HU/vKZL1X9WItyNSXHeEyQG3IEOPcC8KgDzovjCOE/zRzltD
yCYo4wGSHzpxaAce4RavSWFGviuxIDqV4eibXEY8mUdRrHO7eRNHb0YK+hzW+udS
0npTRpeFzy0cXSe0uQqRWcgrV+2ryI0UUEqprOnTGoEWB3YUpyEmQkwJUDGTnF+W
mbAeI9lBGLGeavRb7WQlAxbVH6vXFIn+ayZ1Iwdf5i5AnPXkiuFOts2xo6wVlJvW
/0/ppmguEfM8Oo0nPydWmyx/jXOTsTcIFrPICl9UQgbGuOBUQaxbx14cFHEPiLx4
ASASILFmAwRCGfWJw4JPyy4R9N3y0bsG2zL3CKdc1N0bwQhFGUzIJ3RxlVZ8NFGk
jkocahp++OipUPjQod4LZA7dqWK7AokNzd2vEiSbmNC5ZFZ2ZGKONtw7JA9+DhzY
LKM8QiK27LlLnikweczz6V6CxvmwJtfACHxlTgxFwH0aEczJ+jE88qk/v2fTzVuE
zrG0PraeRe2jpCbWt3q7xVEhFG2SSdjxy+hrzr5xBO1BtYoQuJFOQES52vVQcg94
GxlTWFy+NCXoB2Kt1UDfA/SDimzIvBrv2Log93G4lBI1ko/Fb87yUHKyX+Y9t91U
RxRU7lIQImVpbf8tWK1U6PFPeVYo+He1gVe1PZc3cKZm9LcU4f4Vgi4n3lUkFozJ
Fsa1GpByszn7Av7AVHmnUw==
`protect END_PROTECTED
