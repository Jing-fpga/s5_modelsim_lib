`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fn/B5N6mE5aLrGPDSbFTaBJJuH6PQ4W8kYGEGfsmaAcmMiQFl2WzR0rXnvLdSt/L
NyOhMR351HS2YsvnyT/UQfnlTJuFHEA4qxOEhFzsdRbPdWfxIaC2C0SoIj3jl1Ui
El4vUE/5p5MLlRWxOb56mWlUGUHRuWOPdEVpOaCYX6+J4iMZ7wGQVbMNdu9RcUcC
IN+dfsnwnwkP/cT0ODJvjtOdd9ylTY0qVu7PkuYX/zjY3YqMt5p9Pc/SdM96xMia
DWZ3YRPEr8SvxOs6dz0ZpoFS4hwT8/nOE4Ohflregr8bdsLDsoqgzZYODGttORRV
770se/e65EBkazZfEaHGHR/DokCs45hPf3ilB9+oZloYW7f7Rc8QZ2tFDclkwsMK
44++HqAXAsKuw4cM6k0ptIJUCnLYiGiMK5piu1jkfXUzXJqiUJD6w0VxVgoHIQt5
5C2JREQWqkhDQagY9l/o36uJMWUznumMmQJNgTAaF0DIM5mLll5EqVH5ft4IBsUl
207uQ008trSObCC60M0onEsk4876PcdQiiMVKpctdZ/xKUkfZE4dF7Nav3dctIQd
7OIcqWyIKYarpa8xHiUxggaBF1oq7/REGf4upSGOHp7A/yA1erj117+WGmIQVcYa
X15U5rEXNt6jacwja16g1NAbhU1DqqXWxxlStCXg/Bpps7AmQEkplw6SriXHf1bs
VhA8VJUuqxAG1EmZ7neL99Oop5Bg7mPQcLSEl90OS1xMuxx/vcygt0vaY4DRuEcW
mXt+UwOSySsb6BhG6UYpSkBKaWRYhONV4m4+Rs1p8LiEBTwmbHwxCJ5FxM/X2Yod
QTYz2kzBK7eEkixyKLCZIPC1Rx9J6jOtraaeBsDCOQToYsszH0dX8KyQJEIZVH5s
zUZ8dmuAyt9VSZWR4JDTmFNwSmzdm9JpW+//eftxI9u4HlKZjViZtYM4ENLuFAwQ
Bt7Qa5+mBDu4NUmzpzMHb6IW3Ug7pKHqF/jmVO7fyvv6lIZvVIb3THpOZUZGpto+
WG5+KLzZ776u1c2kE8Kofiqf9Mvz+StcYzMvrS79q+4=
`protect END_PROTECTED
