`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eLtHtISm7RhTpKe9SKSJDNSbWPT7TRcyY7nDtgOydtojtbzJnYmJ7Ak6uqfzRaGI
4Gjh2KIVerCYzbpWHNp/dbsI2f8Ps7tiPwVIHkNr8Q7spKG2xxgFsyy+NWt8T7dx
afSrUGc83ptYdHLL7Pu8/hrnrQVr/ZyHrg8OV0eoROnOZx9CbWDtP1KdHt8aHOLo
9iF4dJIJbychYsO7EPwnICghyEXfcrgeOH8DBNFww+3Zgy7oKAMfj4VhZFHJvZTd
ZOmRgG/5gfhxvCmPrd8UA8l/cx4/M4iZ+Fv/2yp5qvoNTGCYPgh6GzsyZC3/cZSo
zQ9S+A9MMZHd8VY+MYp+Irs8hE8p5BdK+leVOh9OJmZWOTGMhAyJB1SDr5DlK97W
EvRpmVvOPR0v8cEV5e6MeGbLQdhWEwFqZkSxwrNdG8sV+IKPiOFYa389AO+hA+6E
VCDwYmc1f6hnVFpP9iVKOezEofepvMSGUV4hUdHdqCuaT9e1H5FfoDHY/tpKpePs
FFuyjFPqVRVsfmcdHsH2YjTO+YyWhftkOeoL0Y+aqqpA91pWAEWREyA7hsq6LlL7
aVcOjOZ6E+7xzuA3eEBlwcnp4//woRyiSNIz6K/1jTzq6/F+W09Vc0k+r8eZIhin
XZArRrvePFf5G/zkub9KBJ9wbvCAvW++VSrCDSunJgVf01SP7WYPKaw8tlo3onHe
KS83BmyKzdC0jlxr0tiZ1nDjUMfV/rWrtuXbs1ldXkzTYTRFTeFmsctOvAjSMpwg
`protect END_PROTECTED
