`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c8xmQHcxsxaLCUhL13Z2l2kYNlYzu4/2ymDOclo6BPsNzb75G1GwDdW9h+RDRClL
9h9pTg+ifPqSQfB3JX5G5vW8DqJJhJ1f3Z2KvcWhQOCTJaXkuuTjtZe/aVrHY8Uy
+Q+cFNLlF+1BfoKl8ug7iWPrrK2RJBf50a9MoRsrD5d+MOO7E8Eq3MwPQyZrAfTr
/HJ82Tbzal9HTtXMxV5pHjoZNM1YVXbQBqEulUpv1zLGGoW1gujK823lRVNLMDfe
jTQAtu1KZ2k3laLmICfDYN6J5zoKTMqZwnj82Jyh5PClXzeIOWhVeOB1Bq50i0t5
qDmCP5kI9tcVt91KOPXFrjnJnNjgv4r1x4v3CPRX2Dmbn1gBIJlF8tekyYL3Qm79
ZaZQL4MSmulOLgCqO5Tfx9xFXPB0JldIhPf63pdwczHqzu6Trzxf6BLWjw3R+1en
pft7LegZznZ+OtDuW1RDINBqhbNsrgQ2QrfDGVgceBf4BZ9Tl4a3pYWRvLvXn5X/
LphG29N+ZM7noW/KsJ0T0iuhkTbT3+ISPoAZkI4y3KFVhbW2iBS44Cpn96pUjS1t
/2BngCjVtGRkkM+phf+MjrIgV7lxZWHws608h55E++EFz7mbXgf/MV7hBl1yZKMs
OnecrVIyyUSJ794YUP2IUv2RCXNzCAbmpNgHs7FQ3/O7Rv84eW+ZSSr4F7EB/d9v
5UXFsbG9HnlGREHVyTVIjuxVlQHmR9gbaq+RcW3mnLzFEz84/Vy0CbVE0XU138w8
jVHiVZAuSFWtKoFs5PA2wE97bTuXBE700of9Od+0zPhBWpIYH/VDCxhWm8vBor18
fIPYYmk3v6hKJsFM1nEp1whWTJgcfsYRhn25YpGUBVTCQfGxiC2njwfULEcdGpVr
JYx0zsinKvu8pL+FQbOEoyjprosZ49yWZ+gJ6hIcXeNOcG464nK/NuwaC7+BM/G2
d6lszhuDX0VT+SMy6MaXHjSAWAN1UzbwCcbhg6hILTycEvcJJigcYUbPnx0HGAHS
6UF8UMrayeX2mThJNhsNuCPYuDb1VgZJFkMyWJK0UZpAULP2g5bzvJN3CYX5WtQg
UtRW08APqYjpGIDEQSTcjq1fttzQ2LMAlmKJRbPbfJCYPNOiSyjWRxGCYq6Jq6uw
kom4iuXE73hxlMGvdU0gRqDjFWup9Z7bRBMfkj8kyJjewDpy353gWJjeg5WVGTmI
fmG3dqByDx9UniyUZ8HrmSDXJCMne4gELQsFiknEXh97ra31/Ww230Qg9tL+FwXm
zgCGTRVFgtG+gxI5UIJP0kxPfveb0mbi7DdynrIRrachnXoRwWC93QF9JO7IhSgj
zOqRxmqigJ64LqCOAIfwXOf34Md6/DbZE+lrRwZ0UVLb8WYzbli3EXPh5cbkhiCC
x9RjWabBH5OaDflEWK02vBpoopAJjLgzQ4Y44+VgbA9y3V4ozsFgo+iw58ZAzENG
GJjns1lQyTjCZzdSajGznxTxAVZMWWSuPknJplZELtVXurZq4VrwnPxXBqF2FL5Z
YBdrHlDiTykiC1gP1TU6xNS/ENdKK/4n8dls/HYSLwev+MLiGDtHb189dQIFFqVk
5vELbYQyIQz3NZedM/zDksm348NiOGOqI6qX91imWEgOpessAJmka7Ugv7AUun5j
cadxjJHfZ/UY87ecW0SdvwORJEW7dcCLiuW/mQXPjcqTisaDDD/l+JKASjcgXguI
Ew/aeuIiKsIFs4kg0mGiqoueLLm3aCg4OsQ6ZIufOfST+m3BU9X1B2N0L+6Mrr2m
ub0Nl231sAoWTVDKqrNc5yTVs2Iud0FvTsHKYtgG3dDoyMFuqQm3juW307R9A7g4
trWFKKpNrV4uB68tK1bhHbcqrQfNIWuq29+JbdFbIYMfkszueTZOalig+HISdDwV
HcpnsqieQZhQewdyoL5b61tMbfCD13laPisJJFWdqUab3AEAIWV8QhMiNRhFHJoy
HFRCd5Gzxk7xNqSX5uR+0ryhbgdO+L+lURJbk9kmhzF+O668Ooze14YBl9uiEG6P
2oNoYQqHItFFZCyAW6Wzktfk+OtfuAKViVZE2eJKD2v2DaNpx6zUJ5Xy1GaxBBRU
m5QR9ONcVqQeE0UWK5AfYFPOZAtFERmD8Eccvo0VHFkKSAn6Ysezes2lMa7uLlc3
Lnv2TvkHckyAeED/e3h2AHf9ghSiZdwhuH51gyZPI/MOApbUaqIOO3ian+UpKM6y
NBp14fmTpftSgNrlUbnWuVWpP8EC1rSG/xmFyaVJvlgl/hMpY7tWZUa7dq+mRV9j
wWDLIGUyJiWLW2Cz+/r7pRMm6X9zYK+qGucIvNjzpsL8fn/d6vd7kLJMtpJxJzz9
cs/gT6DInkppg7MBC292OLL1lWo2hvZ4UomUHlsROOoqdPdA3Cczsy6DBJlcXEvR
PT1gi7vVzOuSF10ThWhWduQjq+g0wPswkBenx/oA6SxPss96Hp8Ub8JtcJI1lXEy
cVBT6taqVAnCJmZ9kFueps0kJZCP/gKXWJ9fqpnSBJ8IOoCWrtYr02SwRFwi7Jd3
xYWZpCvTNuftA28nuqQVWI5l3e+FJzDe0YYmAb1d6UGUEgwfuuWYG/tqo43kz8VQ
nD4NQXYXlFvvPpZJtCWPwSlIJYlS/ftFYAukORlpHBzXCFsG5pDIoLwCqwMU3ihY
/kKd/PGG1PQac4PplBrJbkb+VW1qaRBndiRJwL1jsiRd/omKALzXpVnQMS2s/vyH
NW1jrQBQpBElQWNssHUI8kFPfxzzQa4xQ7I3kKmH4Cymw6+GaattJREjJPAELOuW
AaPfJ40OtDCQqLtSUz1+3bgWOo31s5i3AtcSw6uIDo6+uF71OedQRPzRb6hqttvN
6c0qEJrwZg+OkhtlUePOMWQ8GxnLKJFevcxQdQq1pPVmN5CMDHoKBg2q6rBWtQF9
HKKuOxH5gbopvItbmQqFgk1EklvA5Yc7L2QoUTA118hvffuOfMl6CtLLeZ5wAkje
gLZ4hhHwOfalHFsBx2EiSASDxHG4hlvfNO5jEkor0knbmnviLfvU6Y4FVAnIC8g+
8KLZI7rh07PBybXNdI0pNbecq8L+udnoqn66lmsaB8aZ4ePD2TAZyBkvrj0LzjN/
BoEeaniy40MWlOvZitfWoPXRSnCtXRUkdJXLenL65hgVpveB9OxmoJ06rITmlDH0
SL1k717HdM0W73vRvDx2lB7g/zO6r0qxKWkYejRmWU3dtg2Y3NzfZZAkzG/WKUxK
FpWjjoM14sxVblFmspgOfvbpQeNePLbThyhKaXB6CPI=
`protect END_PROTECTED
