`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ki8PewB3FqFRzZyJQMK5S33OqDVwfrOVPeQQg4lwtMCHe55C1umA2FhRyf49GLQr
oTcHiDIMhj+vorAPB4UwC077f6Gkk+F/yJOQW62E/6RafPtvSiXo9JH5IuQfLiNm
XVDRwb/OoJkDe/Sgo/si500wwj8fl2qfBeD438bEkr43AQdVo/6j/0R9fQbmSUUA
dIB5oLW2FzxVu8H4KNDERiKuXjC/UAx3EkqlqD/WF4TtJ0bssVeR5ABeMPaVvAKt
dsHE/1oV7SzVqXWlegmN/ibrxWNJbAimeFs5IqxvuAQGS2fNH7MtGZl/2DoA5xuP
1NBPkYJpwHNOE+9dVUu7WpYaDBg0rOeLb+Bt5ezwICVLbenXYreskbmQZ1Dhi864
VBTIlyiSOWOM3cvH1Cmsfw9hFGX30RPcILDuHE4h4Q21ITSvpGgYWn38AEArbinc
MhzKSGM/8Vzszivzxo3isgFTxThUG+N52HruCpc99isy078a+Fs2nah1m6f307Dd
Y0wJ7x7Yoo9pCdgZNqHCXVjXnSffk4FgAAAl7idDCjkZ3cbY18MbYW6Ya5PnCYzW
hOv0VNluobyeNJMagL4hiZk4CeldK+pBlTHQ8XPC6c0jiPsJUR1+NgIL8eGeWv/K
yFE6dhSr+0hX9HoExflibY9Ez5l9kwEtLEC8xt+RWxyz4hSdTVmZiGCrntOu7dW2
vgXg/xW/OUFDLFz+Spe47JPkzm+chZZH0BCINSHanGtixwFoNhyIah9C+SSC6EHY
4610RoiW2ZyD1l6cHoyj4RiMkHDOm4Xp64ItE6zshkOLqkU7VZcsTnnIz2M0s3vH
f2qj3MmiAyaZtwa0h6FJthvlJXEWPQ4i22Ql8I+UXTDB2tQOODP1YM5LJnqC6rjC
tEw9WKtu4JE/lH+yDXpwVH8aePCvF2nNEh+G00hLP2kTLugfoGyUL8a+9wrznzoB
88VPdw5z15K6Bir/7ZkRne3p1yChihlE7I2aDnBCphsRb2uIaRTb3qyPlsah5asF
iWwj/z0T22mZi1HMCn6Gmuk40HgPE+mrRkYJQEaRQYnuYi4+D7rrO1i3XznHhByS
ihjTJyHB1MTG7gzHIs491ANEqmPvpK9YpFPvb4GkfdWNupd6R86CNtGiU5vnpB34
gpyr2fmMSCJ0cTUoizWE6UW+QTNbX1R9gsmC+E3ROXi+YDt2tPdWgLSG4CNJaCeA
pwN9/cyuo5gyxvOhguUta9eCkZCksoL7Sp7Cq8TTndTN8bzvJXGOmb1D7yKvIFyh
A7+knUcAKzHEG/TfkFV7mHINd43dVyeXF77LBKq+VAlx5vtzRsBwOZ480rzJwnb8
N5OxFonIAO0cRz4i/NicEBMWc2k4zG3Ad0iKUnrwWFqvGxscUBrTAXGQIqOWUcsF
T0J+dAQMXsAzFpNYfnpZzGtuVQYskumlM0FQhHtphiMqy7CBe1h9YX3HdBjejAtp
RHD6Xg66S+HVwEObnzYuRkOlFxCEP6QYh0T5LwjngnVi2qPwCgNO+FDuiSXxBaF0
WMJVOt0fOnvfw2ijaprBxkb+swAdJ1/xZeLYYOeUCc6reiwrLE/HIhR7avQI4GW1
1jIKvGsgQFIieYKBbGgE2ImXixEnXx/6a7ynYgcP8j0=
`protect END_PROTECTED
