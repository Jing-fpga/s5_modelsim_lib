library verilog;
use verilog.vl_types.all;
entity stratixv_hssi_pma_rx_buf is
    generic(
        sd_threshold    : integer := 0;
        vcm_sel         : string  := "vtt_0p70v";
        vcm_current_add : string  := "vcm_current_default";
        qpi_enable      : string  := "false";
        rx_sel_bias_source: string  := "bias_vcmdrv";
        bypass_eqz_stages_234: string  := "all_stages_enabled";
        cdr_clock_enable: string  := "true";
        term_sel        : string  := "int_100ohm";
        sd_on           : integer := 16;
        avmm_group_channel_index: integer := 0;
        rx_dc_gain      : integer := 0;
        diagnostic_loopback: string  := "diag_lpbk_off";
        user_base_address: integer := 0;
        offset_cal_pd   : string  := "eqz1_en";
        channel_number  : integer := 0;
        vccela_supply_voltage: string  := "vccela_1p0v";
        pdb_sd          : string  := "false";
        use_default_base_address: string  := "true";
        pmos_gain_peak  : string  := "eqzp_en_peaking";
        sd_off          : integer := 0;
        input_vcm_sel   : string  := "high_vcm";
        ct_equalizer_setting: integer := 1;
        enable_rx_gainctrl_pciemode: string  := "false";
        eq_bw_sel       : string  := "bw_full_12p5";
        cdrclk_to_cgb   : string  := "cdrclk_2cgb_dis";
        serial_loopback : string  := "lpbkp_dis";
        dfe_pi_bw       : string  := "bw_10ghz";
        silicon_rev     : string  := "reve";
        adce_rgen_bw    : string  := "low_bw";
        adce_hsf_hfbw   : string  := "full_bw";
        monitor_bw_sel  : string  := "bw_1gbps_less";
        adce_rambit_en  : string  := "adce_ram_disable";
        mode_adce       : string  := "power_down";
        pcie            : string  := "pcie_disable";
        adce_rst        : string  := "adce_rst";
        dfe_ibias       : string  := "dfe_ibias_from_bandgap";
        dfe_adapt       : string  := "adpat_from_adce";
        adapt_sequence  : string  := "v_d_c_b_a";
        lfclk           : string  := "lf_clk_divby8";
        hfclk           : string  := "hf_bypass";
        hsf_hx          : string  := "hsf_2ma";
        dc_bw           : string  := "bw_6p6mhz";
        lpf_bw          : string  := "bw_205mhz";
        lpf_gain        : string  := "gain_3db";
        hpf_bw          : string  := "bw_500mhz";
        rect_adj        : string  := "amp_full_leaker_full";
        rgen_mode       : string  := "high_freq_mode";
        rgen_vod_max    : string  := "rgen_max_vod_125mv";
        rgen_vod_int    : string  := "rgen_vod_int_125mv";
        rgen_vod_min    : string  := "rgen_min_vod_125mv";
        max_eqa         : string  := "max_eqa_125mv";
        max_eqb         : string  := "max_eqb_125mv";
        max_eqc         : string  := "max_eqc_125mv";
        max_eqd         : string  := "max_eqd_125mv";
        max_eqv         : string  := "max_eqv_125mv";
        min_eqctrl      : string  := "min_eqctrl_0";
        lock_lf_ovd     : string  := "lock_lf_norm";
        lf_offset_step  : string  := "lfos_step1";
        hf_offset_step  : string  := "hfos_step1";
        lf_offset       : string  := "lf_minus_2mv";
        hf_offset       : string  := "hf_0mv";
        macro_hfclk_divide: string  := "hf_macro_bypass";
        macro_lfclk_divide: string  := "lf_macro_bypass";
        hfclk_duration_value: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        hfclk_duration  : string  := "hfclk_duration_val";
        hfclk_edge_lock_value: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        hfclk_edge_lock : string  := "hfclk_edge_lock_val";
        hfclk_lock_for_adapt_done_value: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hfclk_lock_for_adapt_done: string  := "hfclk_lock_for_adapt_done_val";
        lfclk_duration_value: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        lfclk_duration  : string  := "lfclk_duration_val";
        lfclk_edge_lock_value: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        lfclk_edge_lock : string  := "lfclk_edge_lock_val";
        lfclk_lock_for_adapt_done_value: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        lfclk_lock_for_adapt_done: string  := "lfclk_lock_for_adapt_done_val";
        adce_atb        : string  := "atb_lst0";
        adce_reserved   : string  := "reserved_default";
        bias_rgen_enable: string  := "ibias_from_ibp150u";
        level_1t        : string  := "off_1t";
        level_2t        : string  := "off_2t";
        level_3t        : string  := "off_3t";
        level_4t        : string  := "off_4t";
        level_5t        : string  := "off_5t";
        phase_steps_sel_dfe: string  := "step1";
        vco_phase_sel   : string  := "clk0";
        clk_source_sel  : string  := "vco_clk";
        polarity_2t     : string  := "negative_2t";
        polarity_3t     : string  := "negative_3t";
        polarity_4t     : string  := "negative_4t";
        polarity_5t     : string  := "negative_5t";
        offset_ev_level : string  := "ev_left_level0";
        offset_od_level : string  := "od_left_level0";
        offset_evh_level: string  := "evh_left_level0";
        offset_evl_level: string  := "evl_left_level0";
        offset_odh_level: string  := "odh_left_level0";
        offset_odl_level: string  := "odl_left_level0";
        offset_testmux  : string  := "testmux_off";
        adapt_en        : string  := "adapt_disable";
        adapt_bypass    : string  := "adapt_bypass_off";
        speed_mode      : string  := "high_freq";
        vref            : string  := "vref_level4";
        atb             : string  := "atb_off";
        pcnt1_bsel      : string  := "pcnt1_200";
        pcnt2_bsel      : string  := "pcnt2_200";
        pcnt3_bsel      : string  := "pcnt3_200";
        pcnt4_bsel      : string  := "pcnt4_200";
        pcnt5_bsel      : string  := "pcnt5_200";
        adapt_mode      : string  := "adapt_3tap";
        adapt_vcm_op_en : string  := "vcm_opamp_enable";
        adapt_hold_en   : string  := "adapt_hold_disable";
        adapt_limit_en  : string  := "adapt_limit_disable";
        pdb_odi         : string  := "power_down_eye";
        vert_threshold  : string  := "vert_0mv";
        v_vert_threshold_scaling: string  := "scale_plus_0p8";
        phase_steps_sel_odi: string  := "step20";
        bit_error_check_enable: string  := "bit_err_chk_enable";
        out_to_nxt_ch   : string  := "out_2_nxt_ch_off";
        select_1d_eye   : string  := "sel_2d_eye";
        rx_manual_mode  : string  := "eq_manual_1";
        select_testbus  : string  := "select_testbus_a";
        clk_sel         : string  := "refclk_or_cal_clk";
        reverse_loopback: string  := "reverse_lpbk_cdr";
        to_jitter_enable: string  := "no_jitter_enable";
        to_scale_jitter : string  := "jitter_setting_000";
        cal_eye_pdb     : string  := "eye_monitor_off";
        cal_dfe_pdb     : string  := "dfe_monitor_off";
        cal_offset_mode : string  := "mode_independent";
        cal_set_timer   : string  := "timer_fast";
        cal_limit_sa_cap: string  := "full_cap";
        cal_oneshot     : string  := "oneshot_off";
        rx_dprio_sel    : string  := "rx_dprio_sel";
        bbpd_dprio_sel  : string  := "bbpd_dprio_sel";
        eye_dprio_sel   : string  := "eye_dprio_sel";
        dfe_dprio_sel   : string  := "dfe_dprio_sel";
        offset_cal_pd_top: string  := "offset_enable";
        offset_att_en   : string  := "enable_12g_cal";
        cal_status_sel  : string  := "status_reg1";
        cal_limit_bbpd_sa_cal: string  := "enable_4phase";
        rx_det_pdb      : string  := "power_down";
        counter_0       : string  := "setting_0";
        counter_1       : string  := "setting_0";
        counter_2       : string  := "setting_0";
        counter_3       : string  := "setting_0";
        pcie_qpi_sel    : string  := "pcie_mode";
        rx_manual_mode_test: string  := "eq_d2a_test_disable"
    );
    port(
        adaptcapture    : in     vl_logic_vector(0 downto 0);
        adaptdone       : out    vl_logic_vector(0 downto 0);
        adcestandby     : in     vl_logic_vector(0 downto 0);
        avmmaddress     : in     vl_logic_vector(10 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        blockselect     : out    vl_logic_vector(0 downto 0);
        ck0sigdet       : in     vl_logic_vector(0 downto 0);
        datain          : in     vl_logic_vector(0 downto 0);
        dataout         : out    vl_logic_vector(0 downto 0);
        eyemonitor      : in     vl_logic_vector(4 downto 0);
        hardoccaldone   : out    vl_logic_vector(0 downto 0);
        hardoccalen     : in     vl_logic_vector(0 downto 0);
        lpbkn           : in     vl_logic_vector(0 downto 0);
        lpbkp           : in     vl_logic_vector(0 downto 0);
        nonuserfrompmaux: in     vl_logic_vector(0 downto 0);
        occlk           : in     vl_logic_vector(0 downto 0);
        rdlpbkn         : out    vl_logic_vector(0 downto 0);
        rdlpbkp         : out    vl_logic_vector(0 downto 0);
        rstn            : in     vl_logic_vector(0 downto 0);
        rxqpipulldn     : in     vl_logic_vector(0 downto 0);
        rxrefclk        : out    vl_logic_vector(0 downto 0);
        sd              : out    vl_logic_vector(0 downto 0);
        slpbk           : in     vl_logic_vector(0 downto 0);
        vonlp           : in     vl_logic_vector(0 downto 0);
        voplp           : in     vl_logic_vector(0 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of sd_threshold : constant is 1;
    attribute mti_svvh_generic_type of vcm_sel : constant is 1;
    attribute mti_svvh_generic_type of vcm_current_add : constant is 1;
    attribute mti_svvh_generic_type of qpi_enable : constant is 1;
    attribute mti_svvh_generic_type of rx_sel_bias_source : constant is 1;
    attribute mti_svvh_generic_type of bypass_eqz_stages_234 : constant is 1;
    attribute mti_svvh_generic_type of cdr_clock_enable : constant is 1;
    attribute mti_svvh_generic_type of term_sel : constant is 1;
    attribute mti_svvh_generic_type of sd_on : constant is 1;
    attribute mti_svvh_generic_type of avmm_group_channel_index : constant is 1;
    attribute mti_svvh_generic_type of rx_dc_gain : constant is 1;
    attribute mti_svvh_generic_type of diagnostic_loopback : constant is 1;
    attribute mti_svvh_generic_type of user_base_address : constant is 1;
    attribute mti_svvh_generic_type of offset_cal_pd : constant is 1;
    attribute mti_svvh_generic_type of channel_number : constant is 1;
    attribute mti_svvh_generic_type of vccela_supply_voltage : constant is 1;
    attribute mti_svvh_generic_type of pdb_sd : constant is 1;
    attribute mti_svvh_generic_type of use_default_base_address : constant is 1;
    attribute mti_svvh_generic_type of pmos_gain_peak : constant is 1;
    attribute mti_svvh_generic_type of sd_off : constant is 1;
    attribute mti_svvh_generic_type of input_vcm_sel : constant is 1;
    attribute mti_svvh_generic_type of ct_equalizer_setting : constant is 1;
    attribute mti_svvh_generic_type of enable_rx_gainctrl_pciemode : constant is 1;
    attribute mti_svvh_generic_type of eq_bw_sel : constant is 1;
    attribute mti_svvh_generic_type of cdrclk_to_cgb : constant is 1;
    attribute mti_svvh_generic_type of serial_loopback : constant is 1;
    attribute mti_svvh_generic_type of dfe_pi_bw : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of adce_rgen_bw : constant is 1;
    attribute mti_svvh_generic_type of adce_hsf_hfbw : constant is 1;
    attribute mti_svvh_generic_type of monitor_bw_sel : constant is 1;
    attribute mti_svvh_generic_type of adce_rambit_en : constant is 1;
    attribute mti_svvh_generic_type of mode_adce : constant is 1;
    attribute mti_svvh_generic_type of pcie : constant is 1;
    attribute mti_svvh_generic_type of adce_rst : constant is 1;
    attribute mti_svvh_generic_type of dfe_ibias : constant is 1;
    attribute mti_svvh_generic_type of dfe_adapt : constant is 1;
    attribute mti_svvh_generic_type of adapt_sequence : constant is 1;
    attribute mti_svvh_generic_type of lfclk : constant is 1;
    attribute mti_svvh_generic_type of hfclk : constant is 1;
    attribute mti_svvh_generic_type of hsf_hx : constant is 1;
    attribute mti_svvh_generic_type of dc_bw : constant is 1;
    attribute mti_svvh_generic_type of lpf_bw : constant is 1;
    attribute mti_svvh_generic_type of lpf_gain : constant is 1;
    attribute mti_svvh_generic_type of hpf_bw : constant is 1;
    attribute mti_svvh_generic_type of rect_adj : constant is 1;
    attribute mti_svvh_generic_type of rgen_mode : constant is 1;
    attribute mti_svvh_generic_type of rgen_vod_max : constant is 1;
    attribute mti_svvh_generic_type of rgen_vod_int : constant is 1;
    attribute mti_svvh_generic_type of rgen_vod_min : constant is 1;
    attribute mti_svvh_generic_type of max_eqa : constant is 1;
    attribute mti_svvh_generic_type of max_eqb : constant is 1;
    attribute mti_svvh_generic_type of max_eqc : constant is 1;
    attribute mti_svvh_generic_type of max_eqd : constant is 1;
    attribute mti_svvh_generic_type of max_eqv : constant is 1;
    attribute mti_svvh_generic_type of min_eqctrl : constant is 1;
    attribute mti_svvh_generic_type of lock_lf_ovd : constant is 1;
    attribute mti_svvh_generic_type of lf_offset_step : constant is 1;
    attribute mti_svvh_generic_type of hf_offset_step : constant is 1;
    attribute mti_svvh_generic_type of lf_offset : constant is 1;
    attribute mti_svvh_generic_type of hf_offset : constant is 1;
    attribute mti_svvh_generic_type of macro_hfclk_divide : constant is 1;
    attribute mti_svvh_generic_type of macro_lfclk_divide : constant is 1;
    attribute mti_svvh_generic_type of hfclk_duration_value : constant is 1;
    attribute mti_svvh_generic_type of hfclk_duration : constant is 1;
    attribute mti_svvh_generic_type of hfclk_edge_lock_value : constant is 1;
    attribute mti_svvh_generic_type of hfclk_edge_lock : constant is 1;
    attribute mti_svvh_generic_type of hfclk_lock_for_adapt_done_value : constant is 1;
    attribute mti_svvh_generic_type of hfclk_lock_for_adapt_done : constant is 1;
    attribute mti_svvh_generic_type of lfclk_duration_value : constant is 1;
    attribute mti_svvh_generic_type of lfclk_duration : constant is 1;
    attribute mti_svvh_generic_type of lfclk_edge_lock_value : constant is 1;
    attribute mti_svvh_generic_type of lfclk_edge_lock : constant is 1;
    attribute mti_svvh_generic_type of lfclk_lock_for_adapt_done_value : constant is 1;
    attribute mti_svvh_generic_type of lfclk_lock_for_adapt_done : constant is 1;
    attribute mti_svvh_generic_type of adce_atb : constant is 1;
    attribute mti_svvh_generic_type of adce_reserved : constant is 1;
    attribute mti_svvh_generic_type of bias_rgen_enable : constant is 1;
    attribute mti_svvh_generic_type of level_1t : constant is 1;
    attribute mti_svvh_generic_type of level_2t : constant is 1;
    attribute mti_svvh_generic_type of level_3t : constant is 1;
    attribute mti_svvh_generic_type of level_4t : constant is 1;
    attribute mti_svvh_generic_type of level_5t : constant is 1;
    attribute mti_svvh_generic_type of phase_steps_sel_dfe : constant is 1;
    attribute mti_svvh_generic_type of vco_phase_sel : constant is 1;
    attribute mti_svvh_generic_type of clk_source_sel : constant is 1;
    attribute mti_svvh_generic_type of polarity_2t : constant is 1;
    attribute mti_svvh_generic_type of polarity_3t : constant is 1;
    attribute mti_svvh_generic_type of polarity_4t : constant is 1;
    attribute mti_svvh_generic_type of polarity_5t : constant is 1;
    attribute mti_svvh_generic_type of offset_ev_level : constant is 1;
    attribute mti_svvh_generic_type of offset_od_level : constant is 1;
    attribute mti_svvh_generic_type of offset_evh_level : constant is 1;
    attribute mti_svvh_generic_type of offset_evl_level : constant is 1;
    attribute mti_svvh_generic_type of offset_odh_level : constant is 1;
    attribute mti_svvh_generic_type of offset_odl_level : constant is 1;
    attribute mti_svvh_generic_type of offset_testmux : constant is 1;
    attribute mti_svvh_generic_type of adapt_en : constant is 1;
    attribute mti_svvh_generic_type of adapt_bypass : constant is 1;
    attribute mti_svvh_generic_type of speed_mode : constant is 1;
    attribute mti_svvh_generic_type of vref : constant is 1;
    attribute mti_svvh_generic_type of atb : constant is 1;
    attribute mti_svvh_generic_type of pcnt1_bsel : constant is 1;
    attribute mti_svvh_generic_type of pcnt2_bsel : constant is 1;
    attribute mti_svvh_generic_type of pcnt3_bsel : constant is 1;
    attribute mti_svvh_generic_type of pcnt4_bsel : constant is 1;
    attribute mti_svvh_generic_type of pcnt5_bsel : constant is 1;
    attribute mti_svvh_generic_type of adapt_mode : constant is 1;
    attribute mti_svvh_generic_type of adapt_vcm_op_en : constant is 1;
    attribute mti_svvh_generic_type of adapt_hold_en : constant is 1;
    attribute mti_svvh_generic_type of adapt_limit_en : constant is 1;
    attribute mti_svvh_generic_type of pdb_odi : constant is 1;
    attribute mti_svvh_generic_type of vert_threshold : constant is 1;
    attribute mti_svvh_generic_type of v_vert_threshold_scaling : constant is 1;
    attribute mti_svvh_generic_type of phase_steps_sel_odi : constant is 1;
    attribute mti_svvh_generic_type of bit_error_check_enable : constant is 1;
    attribute mti_svvh_generic_type of out_to_nxt_ch : constant is 1;
    attribute mti_svvh_generic_type of select_1d_eye : constant is 1;
    attribute mti_svvh_generic_type of rx_manual_mode : constant is 1;
    attribute mti_svvh_generic_type of select_testbus : constant is 1;
    attribute mti_svvh_generic_type of clk_sel : constant is 1;
    attribute mti_svvh_generic_type of reverse_loopback : constant is 1;
    attribute mti_svvh_generic_type of to_jitter_enable : constant is 1;
    attribute mti_svvh_generic_type of to_scale_jitter : constant is 1;
    attribute mti_svvh_generic_type of cal_eye_pdb : constant is 1;
    attribute mti_svvh_generic_type of cal_dfe_pdb : constant is 1;
    attribute mti_svvh_generic_type of cal_offset_mode : constant is 1;
    attribute mti_svvh_generic_type of cal_set_timer : constant is 1;
    attribute mti_svvh_generic_type of cal_limit_sa_cap : constant is 1;
    attribute mti_svvh_generic_type of cal_oneshot : constant is 1;
    attribute mti_svvh_generic_type of rx_dprio_sel : constant is 1;
    attribute mti_svvh_generic_type of bbpd_dprio_sel : constant is 1;
    attribute mti_svvh_generic_type of eye_dprio_sel : constant is 1;
    attribute mti_svvh_generic_type of dfe_dprio_sel : constant is 1;
    attribute mti_svvh_generic_type of offset_cal_pd_top : constant is 1;
    attribute mti_svvh_generic_type of offset_att_en : constant is 1;
    attribute mti_svvh_generic_type of cal_status_sel : constant is 1;
    attribute mti_svvh_generic_type of cal_limit_bbpd_sa_cal : constant is 1;
    attribute mti_svvh_generic_type of rx_det_pdb : constant is 1;
    attribute mti_svvh_generic_type of counter_0 : constant is 1;
    attribute mti_svvh_generic_type of counter_1 : constant is 1;
    attribute mti_svvh_generic_type of counter_2 : constant is 1;
    attribute mti_svvh_generic_type of counter_3 : constant is 1;
    attribute mti_svvh_generic_type of pcie_qpi_sel : constant is 1;
    attribute mti_svvh_generic_type of rx_manual_mode_test : constant is 1;
end stratixv_hssi_pma_rx_buf;
