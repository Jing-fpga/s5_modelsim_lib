`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mM0aXFoMEo//mgs5NCX5l5ewcrJGVZ7MGbBI94Ma9KtZGXro9Qyil08DY5dSCiwD
csc/1Do6Z6UmTwJcUsE91bDal4Zpt/jGj23oB9fwOuFpPVKJc0h4EZHSL++XE8cX
M8Vu+t8DIho7MT1XdkNclAOYbRCW8tfhbxqK9nZnULFmqFRjOqmgmhX8kNTgfl7C
KfcTskKkeBbRwQvWZlDWh1lfmVNDrmwZ379uNZj5mHhQeUqEtgsjiRnppSw05RSJ
ZWra7SuOcHwx3KQYSLdeTCHfWLcIchJEfKuiuJJ/Mfp70cQQ3J3TW0MaDZAuxEYR
vM6vGW0xYRz2uRVNYi70KP07diVcSNAT+mAnMFtWlUvLHkfOqtujowlR83QZfxA9
Bq5bvegxytCymN1ymz5pTQPw7lt1wzYVLG7DfbRjI1ilNeHGidqYZJJaCGotjRMm
fmjM5fm7WP1m0Fiz+8csGiuDe0JAgCOj4LRFxSEcRRE0zm0Nf6zhktYMH8DO05tn
yDeobrzv+dZjML7B8TmvjEw+dIhFMLqHDnBhUUouvUNhmFc86dIMCeRSc+xspMv+
zu5TVitlkSVAnaPzexbbkkXrEaxH0i1RckkM9Me5eW6rhxyoUVe3GHNvvhwDv+8c
9I1uHSRhC4F+4a6v5b3RzYmtpmVR2HJxoIoElhFbN6Md/0igOKy3dWIaWUvCXXoB
lyRc0YSIgAAkkTCDKZIIY0g0RldULL3A1X7FmI3Lgh+IRX2MSMii9HV1MQzWvuAL
eGeCzVr87ABeI+AuM1LH+VdIwaKY06xgSNfC1B1s/hK2gJZsU9XyXQjzw57IhyL2
mkVPm8Jg3G33wgU3buEO7qKhJW1df33+0v5jFLszOn/hTlBxu2CESah6B4wR0t4R
YUNvDTBJTqh/Kb3lPR38t1HBcDUyvaKTQY59TFr+0U0=
`protect END_PROTECTED
