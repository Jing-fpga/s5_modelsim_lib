`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sdpFbpGuOoRQReyTaD7jzoklofwQIz4woO82O2gGZ8LIRNvBW/TrDE1Z9qTSYOLQ
1R5ubG9IEaxPlwlhlFkRqdb3fN4uJkZUSBa9PjvT8jVqfbi1wuudJl4WvhIKxxTR
RFQXRVcMUrDmptEswPiNxPQVVueadh6qno7aFwo3XRx3ENAKXk/JnpV7L61gUpaU
4JQTRsNiy1lnmu2lC7h2FUqHh+qzAjlzRethGf3n4bGHKNxSGSu34QvXQuRgC2+7
cEYg3xpxq9HyXkHA4iweoRoYPy2Dyww1lXOMPAhUURahOHVGDHhLDXpU+5bPMl3O
IGlkL1KFbyoaqGuL1CITBupGP2QZQ3mKQJc6F952YFgH0aWrVCEBa+jMVUHICreE
yiJC2x4uWOpqaX2UfzK3VGXL92KGk4Lzy1Me883i09/7ENVZDI89j55b60QOMRUM
N15RR6vqUjWFDyOb/yP2sHwK0roFRVdS7dLo/eJUYUSX3d63yMXUCfhiJoCpu2j6
obXL15X4mztVestg5T1kjyW3X0oz1z5+/OdQji72aOMvOXxHlhJEYeLtyJg8k5ur
awrVWfHW0a7H6sQ1t2zErA==
`protect END_PROTECTED
