`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T5l+0l7c4I8U9TNgCJ9XvIFLqcJrZTcFgMgSWhFnYbeRFoD5Tvl+9Z4/EXF3Rhhx
w3EXn2fjpN/1cm8q11EnMX2xhf5KBqtQFkyVxwDKTjc65pNHk7elOD6B15pfh6aj
fEZ5tCqF/vrDxnCcRgThVMuc06ghN6qLWyqN4AGYR4Lm6aa/MkGfuzlXitKclEAr
ZmZXcrCB2xDtOjiecJvxqE92NzPTf9bRUH0Xiz+T3Vv9PlQ4PD/uMIINmW8nKsNk
brDZ73as5pbsy7xg3aeXRmO0Tjgi/EjfG3eCe9xNJv8HE/ZFsfU644KrgnY2z9G4
qHVwCZQpqBJSMhaOQDUzr9b2d7HjZQEajax39kycY7txEMkEX7uvtmnSopPKohNi
O+WBdJtYHAMgQgVQ3mWifKqq5rvg3+sGMk/YjIfP2aFN7YIPnUG8SOqdAps9GFaD
LdQT4XrgTAcZs1idt+TaksIQanv+iDk3qfstQ16zK/wM3VHnt7qdPzMBOV2JlkoL
FVAXbu6KrQ6HdalKIQ7k5VJN11Ase3Wg1uYXp44Yi1CjLaujsX4BmbU5uiA+wDTZ
OWbEjHWBGfrsOOtFX/LnhdmhwzRObMQnenho6tVx12Z4Q+GcC2dNNEka5Qu1etzv
jJSQXcSPo7s4hEH1nqistHpHtUajIkz5y/2nABOjv4XFP3X8AH92MHazM5fpoP+x
spRjIWyjjOXwK3leEHGP/wNWsyZWVlIHZWc/za2/na7mZRSYHuUugS5zuL4scq+t
WLHLUdxbWdaGdlIBzibqKPrPKnMVrSptmWYero1P3lPLUoEbvkK84ZqK37qpl3O+
VpYBfNt59hPxZm3GA2yVjOzxZuv206O7QyinBrqogh9wmt26U3eVgNouVIlShoiR
wZO7Y22LP0Qi7P8MuHm+ZTNJaxHPA+F0ygxKf7cyCmljULqzrHODuP2jsKazFC2c
lica7azyVX29ATkz5+8xMJQieliL5Ib0VeDejkBzf1qmoOejuly6VwbHPn7YSxnd
5KabMi99zLH24Li3LwMOUHV1/ImDLuH99IDpWVGPsLj/FlgdmbVXyM9BBMbsyxP4
exwBjGuCN8t0dSW1w59jASBFGsPtBO8FPo/36iwixAt1s7/u0Bn9d1rvSmmFGu4j
MoJGb1H28wh0VP4vzsSiUkABAxUkTEo28hI0170QQd5r5uPVs2k7VvC5hqXZgyNC
G73alGNxfDb/AbIudW2ZIm5NPMkjVlF7xu7AGXwp3A/HVGX1yGshYaeIba5WHJfm
e9+bDr0QZRYIAYj7zFySVJMoTwCVDjVjmdVaOetAHbC0A+ZvkKwSswA3+e3OeFLD
/8ZbfJz9fP4lc5s4bptOMOGs7GDmUHZy3EsbuEj4ROuFXgsKj5M2FFXY5SaIfyAX
SIbgJfdbYvGW753nafxkB8T4go9fMHpAsFPXaSII4ClxWxfMdfXXAxgXRv0R/ASW
yjcH6h0fYIoKJ/arjOwynxPjot2LYm0GcuTlpRIpy+cQ+iMTF/d8k2dQzTsi/7xD
49SnuSvdhedPmr3B2i/gnaBEnFASzVIu8DbaILMch8cdAUdDNyJ9aL2FsQAAbT8C
c/ySuKoP055jmPqAtceG3E/vyEn0f3EwOLB8U/oZxWeEIwYg0Bf77UF7VWaPS7ya
CIB3u/yKJiSgyBUksc0tLMJ4EhGefbpW3ZwFwCTiDyUB0hsk3UamYjC3Bl6VCEso
a/T+mdlqBOF/Se3cI0qMUlDQNevs60w+EDQnxjzwXOT94RWkBTPM8fr/zv8auyfp
vCd3o6TQVY+6Qn3lVt1WCzspdPwTcFZ5/rcJG5x9GiQkI679uPDQSqyHOQJxvlRr
N0AZ3EuJ1ktAfLuRkkfEGv3WVcBBgJaEr7/2GXtYDWNk3fkPmvKM0/phMkLOFrZH
b87cF63UzcjSdp5O1AIzZSVbiTfYK9ktdRK7gJP/JZvXHrW6wDh5ajxdfUYYUW1t
+dysW/jiUsamZZzt8sogC4HpfaGswQo7DqC60QFhNkgwUbUbYQixTLHVVnpXTHfq
ZmORI1VEKUUwCq5shEesUC+giudS7CYc5wr+SEMmEtzD/HavjsulVIfsHJwRhNtv
Q5kJQlS0VgHbJLfKwBGykU4b7e6j0hs1LsVSqjqDMZVL/Kul12BxEgSbBVgnhAnc
pYb+t4kSO6xrLVU/P4mM8abEnQ5vWXMk5gAm1hGKqIFpJrXoiE96oGHDNY3aOZz2
YKqJ4xuBFuJtpYha5Ww5Z5Wj0Zdt5jbdfgcN4U6poQAg615GyCCgR4WwpA17qOJ8
tK3HeLquWJSzNJ/KqYzrsmQB2Ndsve6Vfhty2kot+PvblwSPhzhxcZRrIbA4gyzL
+dn9fOpu7MXFhnV6e9Kx93622H5F6HlUmyFMwCsZJMSIvZQcZo9qUiyjB7egX38j
wX+wbN/4mXV1wHIJvrDEJkephS+SUkr7PAYYc6SKFP/hcjdJqd19jRzWyeJuYBdA
ev76U/3+fjuqHpSuXGtuqt6Bj04WnRV5KiZ6aJMggYdZmddk2648I/dYL3m6L2aY
9mWi2ZxfC2heRqaOe5pR/IsY/8kt+Ll0f9P3POxRBJ8Ee1ZiRlrlQIiUNcd9VVyf
lNtJJup0XXy6SJ1iWueFZ0L3ukv1/qDMhzGLaW4t5TS3p/Yu59QpgC+fanWvWtzo
dwyKiVStYQnm48tJRthP1O/NpwZKqU4LTUDdzuXUD+iFtKppzJxbVuqEWuWKPl2M
sVdJubpXLW/ivJ/fid9MmPcgJIcF3FVMhzv8Lu6w1BFftnvjLbQeou9LqghwqB71
xFFKHuLoGhOTGiEA559N0Uekaa0Uxu1IBah9BYPt6NHGMtQjG3vriH/RuXkJQvE1
n2gziVfJl9hURhHTQIM905as2xM09T54l/EHawsp94AgxsRJeFz5jkDePHShh308
C5+cqbvGgTDPhtYoYaxIGvQjUuLaV37TWoXbKVRJilgb395z/LHKyvz+Mf3gKGEJ
ebVMYboGOpZU/gjZfNH8OCv8MXFSlRSEPBuQeH73W0WmHhRdBlv/uXW9Sd3OTKzn
eDcvCGrf4uglEOUtow9KLCldeqxoE2ZgVQK4LJxDppw3my00XudoRBA5CV36W+ss
U6j53nCrJcqgTSnP/3sssTcqG0tVK3mTMPvs0Cxhh1R6fzOf6vUql49pmzj6VCx5
nGdTtPSDNe9rh3oHiZ8r9bIFToROC73nGpUqrmNZQoxxWti1aAW7fazcjMOsGTU7
zEeNhpxNSRwDRCtDeKP0467LigVSpoaD/VufM3x1ckzj4jqAnYTWl/+V4r0TMdHe
B7h2tCiDwupyH0BrdvlN7URN6217m9qIuJiMnmvr1Q26G6+TA2AgSoSxzE7uGKid
PojhhnhIrxwWN/BX6rVSjlYXhZN1YhUAEO7p4VlO5c6l5dRZrPk66xzqoE03TGKm
5QQb67ECa8xyJpjULioHRdrC3mkk80cVQ2jPpvNYiGt73mGMKxM6DK0BRQ1/H3qo
bq1WW4QpiYmYwoypjlxkmB9Dlj80+5leG4CGt3oWGnB2aTGEdZhKnMhetj9N4+/B
C40Z4xIaFBswAyiwqCV/Bz2XVVYpIcGmesHLKcahrfFZ753aY8RfG2VZOwbd9Agt
dBUo9u2J4bCaENuSWgRB05biNsJqVxH5HpoY6z+tEbMJlXF2UTLhEGI32lcMf8h9
088KC6Qt/3zLYS3EwBDJlNiNmixQd6hb7Y0C2HiGlKNCQfw8BdsoGWX1iV6HWsnF
11L7n4/ozuCu+ogPqe0a6IT6bVnQy3TDYTPC0M+hoiCt2+HovEBJ1U+ZepYugn33
V8EyGPO1rSlJCUiZiJI2vhm1sLQHm03FGo8IAAfVUPguXulgFzMJ1XmdFMLX0zcm
`protect END_PROTECTED
