`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hhfawsb34n1+ZrwPP8cxKquI5bgmkJi1sS60qdS2PtgggS+bfV7Jb6Wv9tC3pwNr
xnGGF++UEhn4w68Go+srhsCJ+0v6EAW/u6JXbLcMTN8uTJnq98EjYu6kZ+eKukj2
HkkRYFdglTL+hjCWOMDwaRrdjSiyog/aOBYO5m4fI9SPrdLLcZeWiC69hSxIKil2
dJzCirRsCMIBW1uUTtEownSlZbF+rsDkDq5umhtZACdrrD9Si25PyvSYhjF9rrQM
wJlcGuvCH0KuCyzcrgsAVycd4sUjBcxebApLqvNvQ9ClZTrG4+EHPryPmrL7xQFK
JizwZs7wyLSmnBgOz6d8oLu+cLiDxSnLqU8o3UzLb7OS2q64Q1JiI8c+QudxtOaY
HpNzD9xL/ju1Ed8G1uOc/4SvYWxhUHBcZ0VjS6sfcrTLm7BWAKt6TIyP+2r8ssdq
9xmMg/mhEbTEOMTjOvOzY7hLpFKiK4zWd6LXk8VNicAYDoBbt92n+NhPSWxfAi4H
bPQb3ZsPbxomQmpHDyeS2U786YybprTANNvaJXMNYGTJHdHQiOLUb/8gSy7guplC
RlQ4zfcVazbiKe3CD1dEq6WAPZIDEc9Sej+euDWCY5TwVjEyAxZiOFnPktyGZI0H
L6xjXnE09gVoll9rFt5d63rBuKc4ruYaQYMxnX0SY7PEu6gqljQ30MOUIe7AqFrJ
TyVjH9X+RU/ejl0iM/+d4Ie1vRo23k/lnnlaOsKBSE47KoogF98GGGMn8NYb577p
y4+nDbJR4CTqUXkASZHsH3/glVw8tvfRSxKESu585sHSNKsaRFAEgKtexnnCDAz7
tQdvkc9s4uea3DmJlJ8Wr4ScCJSPwFZ6CzEphyD5/GXkgKQAEekI59B4IwfA/NHX
bAtePwWHB/O8fMbuaD3VaeWxv7wu5z2kynTfExWF1qk2VrOoSsbjhRt/J0DSHKKW
uF9fnyCkP0gNCpVyTPY5MdWMTAe4PbpB05xjUSBO3vgUemzMKzP76j5u7PrIVZDU
6s47BUE9K+44tEZvgYFl6RiA9uO/GhZftylYjcRMoT8hxGnIjMqlFGRG36CyvD6e
oZUHTobRmXv+8/yyiuVuXnWjk6bESPlcvrsdtX2zBTe4g1doujGPFXrFbSUeOctL
tyDe0O4YmvvBBXvWlAio8zLblvjQgrXgTUuoVukZLBCmKMNqk4N6UvEcIqofeVWL
yrNGMl2JoxFyB94BXIDfPen+fvn2SAQDii2GwOlM2OtkPtCo1axiiCueOydu3F1d
Et7dMmI64NJaPCNGrXfb5A==
`protect END_PROTECTED
