`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BlX4qZx3buQXn9zYHRJV5DcdJfoAOM8md9L2x7AZmwzr05tqLwfNO1H5+gn72hR6
IU++ISX+UCgV+2nkzJigJB8QPU7zutZ8IdKINs68OgkXSF4wSEFD1dnaAKRclIoV
IDIY8YfxUcv1ry7Q4cdgxNWuNUWabwutEgo+0HfEJL6MNRU1GbfQ6mL57nwSsFzU
sUJYQ8CYQFe1782ySqT5lhh5bmBcIZdTgUvD13uYqZ8weK0HdngR6q05eSQrwX8U
hjirutJ+lbbO7GDjrTtnnQezZ2fU+FINwavhzHsqA13n231e/GVT51PDe918keuH
tuSwoeT8ap1WL9h5IeQjhNJq6SmCEgfXp4wVXTa3MPvUnfNH/Iy9AcWNFMti3Id4
ED17jmbJUnEaJxK6h8dHxk27y5htMyoQQw8E3xoHlj65kyNB/Y22qpx5vu2jLF9g
/6nJrnFyYMwBjYWstOzn+brcQ+WaaSVRh+GT3hkZ6br5vObEskcNMkV+8FBh89Pb
b5uDwXzdg0s9fexAAbZQl+DLaJL5ltpmqXb6EDl3Q6zoEi+669oFgc9cBOeL2ey3
FVNq68alR5u3nm6+XVnmNb46NXRQu5VAm737cEfMzhYIEyEmYlO2WfQdJbscFbwy
`protect END_PROTECTED
