`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qY1BslCR2b4WziQxC7zF4GvS8BqR5nr+Dp5D+NYrR/aA39eG8KKJRiPQdR5IL4B9
JWnb5yZcE8vM3CwlPPYzp0vNbbr/4yOX+cKNU+Ou3TgEJ1RxMuNzTbHCTPbR+TA/
oJHK6Pot+ga57yKyE2LSoVifqYDyYb0sAexG5PHidpJLWBk38yRSSZ4lMUP98w6P
UBSvsj4hsuTcwBpWO4in810Dog7I3EVej/7EPQRp4tjTsI0NLH6phS4IB8qYC/OT
bF7cOiTSXY/sRBu4kdNDE47EpFxyuvcfdGsU5wGfJGucQppotSq8/EVlnShtUKeX
m92ujdF4tT8en5HUA6O4iYUK7Ra/RSVs6nOkf6yifiAV77BSi7k8iSXv27nx1aJz
o5fQl8Jnn3qbYO1WsM9F26cZfBfaLjm/Et+CfXaIikDY0MST8zHL6v8euTgQ8tmo
vpmRMSMEaYJdYA7bjtmFFr0/nLqSJaEc2zSQl4hFhQwp47Y5UfctcR9sw/COOX2a
4vZqW9CCJxwvmE4Jtd/PrNXDAPNnlZPgk2q2jbHtn4Sm7jull7HgstwP4BDyN8tP
0Y0gQUt3iZ/IIrhLQZNHdJo1TrfWdILQu7XlpHD/WkRP9YhI/rA6r3v0fVTjyoNr
48/vZHceFEKhYlHOjFHSjja01HxmxYe/0UP2I+FX8DP6A/wWkMZA80ol33agsywO
bP/A50S5pIWKj763iay4FaVXJ10lJYdspiLk1gIi1VXKNDVhfhVCAJTgtjzpiLdI
3OOQ3gOk9JYbFyAC7zCN1nz/sxqyWvtOXMY1BaC4IstgXA0UF8vNPjOK9Onna7Nq
dqxIZEDOIh5wSp9q1GV4/cOsY1WeQMjUDbiUOY3wyE0l+WgeGrodW6qzo0ZZUttV
2hbvBOVp+fhwTH2gFPPCg6UhTJmvgG5WTY0cm9PHC6AVykYOQLVBe/iRW4Cj1SWa
gIRJLrYanD3bhIkGcPeSviUZzDZZCkCqtpVDdgrXzNpOGE60AhwYngjj00NEfmOu
9MJ3L+oaRI3yIkwoHYJyetq9OeTgJ01fdFQwg8PDaZbypPWE6y7ZF8tnO59UzmcS
b2fGSNVhiXOOaXvNwLtc/vw/6f6h6X2bFbt8FXeWuVVflFT92y8gQ4WzaQFenCQO
GDBR/PB7JBjKbAN3r3lHifCk7YxuBTAwULqwaIRRdjJNZnOhzAd3SdAjUz7g5tst
iOTZESZubXZSObN/CZxhvkz58FsGQL63oVFSQpk4zMD0cAVqk4f33XEFFQh1b/fL
gp/bJNcaZAhGL310T+Za7UJZGUA1Zf4obqaqy9En9a/DF7A1SHzubKzbOLRA5Hcj
xuvH4UYkGksNlHlLevQ1hJO5kFWp7bLvNYn8s4/3LaDYVYfq18vkv+78IGHODERn
hiUcXWwvf8e60MDgw8OzEIx4MC+L2zYPn0wQ+XKqArIWWXWtsq0nnGHn+SWLkS1W
j45zt7p2OZgM5DklF1RJX0xlkT49YwjLpz6aJWzj8703G3lcWOox88/B3uUoxf/V
RQj3nPfJ1h4soBye1/H1eCQAro9FltPlSPfpFOmk+XdIykfIU01hh++Z5dGQCAOL
eA+EmZzTh/zCXalA9GccMq4Pp2m151txfPO5nAxOzYOU1I8HWlouyc15jJB9i+NG
K2L9J/QrWocKvDtAl6pOkDKIrbvc/dKgsP3gI2UWVxDSR7Mw++w9QVeYoIkC9gNH
VdR2iYzKLMwyHCEiNMVevfHv8fCy9mWMYZOUzAmHtD9TDK19Xb1N8vNIblFHQL7b
rPqTJ+YEQVHTLYUhtIsoaSU5bRWue2vo+bD2epznla6aT7RSoMcceT85X97LYk/O
ovMlBj1P0+R7n6uwAwcGFltqvSpqKu5RrjBObGvXBRRnSvNyc882bmEw1tuVjbWq
clNxL5j0BbNqmTxscbxQsiv7kODNtkFnr92V8HicsQu4l/BuyEIExV442t24tG5f
lzExzDPBHLkJ+2N2ytcQ1MJWXzcwup6k3LiTpRealcELtsXVtXEQMn76UN5rFE83
7hdcdE4xBNjvdRHvDA83VYYVqC2TLb7pxqYzbisdpIe8a0g6n3yz32ZbHbKSyppH
ILOheQ2qNDsWiIxbh7/usZxmdKNs4zMXFGC+W+SevbtUxQGC7uDuflhUGjL5EOxb
`protect END_PROTECTED
