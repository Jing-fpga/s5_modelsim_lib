`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VoqJCQnn7x5prPyFpkCcbWAIRF9UQ6yXItTMOYKbqiMD9CFyzMuZNFZMryAbHmOt
gPg/iJCWDUPCVX/33XW8ResVh5B8WKk/ecw1VjTiWN+ktEU30nmYYLkRNkvRgbZm
ELZyDq0fMvD3CxaXhn0x7WNi6HE4T3PXkX/KR5rxvixOwcVdqvGxal08NjIy09Tn
+zEKvTcOnc2YleK8v/Yb9qpJvq1YapKiS0SLWAfWmUS84m/rSGiIjqjNdkfk7quM
iBMQwWBr0lTZGC62HeXiXgylvBDPPO1KUN+uRY4MqIMuFzWnOrUmMpHZwWCFkTdV
uqSJ9dd/BrLs6dLckGFVamJCpoeG7lIYgjXvA/VAguYEfSqz/C/PJjjJn2CiB13H
T9kqTeh+wXSGshDrhwNsDsZTbwwVHxfuCoEkTnTJvHl1S5v2L4e5asaY5mAn2J2U
dgd4n6d8o529SAkYJQuRkd7GlI6ZG3D9sGzEL2KTPhIkhxazAcD4sIRjsMPzFpuz
hhpgP40XTqTO9IOoA4k0DfPShY5bMswR+4nuybAsdRO43YCE8qQNZFZYTAk6ADlr
WW7WC9G6ynoEn1ey+3HB7STQguQHLv8gX+bRbD+qKvrWr2Rv0qQFnlScnzmexR55
qSXfCWe8VC/saWzq7ypq0SIrvTF11+pUg1cvLgR2pZnd9Hh8xrHiWEmylbXvtWQH
+6G4oABYc28JUYdaj8x6aHLnUE5/KUUCn6TWrHqaW68TOREEPDzYPTzpLy9oP5bh
tbVvrL3mJJIER3WX1AHuNUhuHrhe+Xa6ChdiIjd6ptis9d5b191bUeE3FKSALNTX
BxZ/s7oNPYYsJn3TqEl1bXPEKoZAN41+IeTPN7vvMWwperG2a4wDde+EdGbZ5K7C
03MddBqFX0UPu2cEZJbhvlb6zqpjEzxtdO4a2Oed+rfZ6vRJR+NYD9hI7WQl3nGa
esbIAEYhVgJMz93PTkOQAKpW0QkmBezPLDjqLnrG7ranEi8u6C19afKv/ZNsnwm0
tJLsr9kUdoVgysP1t0fepbPTYlkRH0AxW2jobcZ1+B3qzABOhRnKK5wXg1/R+itp
tkORCfFHElgeUgPMvkSlGXGHunWCub+/Vzty6hUs2TWnYQXWPsNnDDOskmJpOxyw
b94sSUveXoK/lVA7E3DbwNvprann+0opFac6weRW5EfXhOhNhy0X+zyPWsFntsu2
ZNQ/kc5Re0/DCsQh1CgZGX5UQXRQqKYsDKwUej2bVfsNvtT/HswrvfoT/nYWKFtX
pBUjjhNHyPNT/qYkTXgAL4CZbUrH/wXhjL8bs7Sudacs/bkmKF37mC8S4nRYvQgE
BqzHv7uyoE88xMJz08UP3pWu5nU9a+DgLYG59K93Ls4DSpIw3vgGusEwgcVihZKm
xmuXWWQdLBKhIxhKSYPTs7OyR3Zfu5y24RLo6Huoa5eEyhZQGlWoy0cCCMcBC/4w
7LSz6BlMN2espP0rGYKyel7TkjXGxHY11UNvm5Mr3/3tu/Pw/B1SX8IbvVdHFz8i
MrFt6uJu59lz82oO85M+Zzj00EY1pEP0xLZB7erZ79i6YoWX6iB8eGiruo4fWnty
EtEKQMKxrQBcIEU97mQ4FP9ZfxH8pUHE7xVCN57F8Oj9aWm29sVo0Ccb0WNln3Ev
hOdCXLKh6VLyKBf+YEWO91aX0ZTlsasLK2GHO5441KTgCUQSipEcAPShIDnHAuM9
P3Fo/MsZbFYhLtWNmH/xNqBs0s7EybhuK7dUPjiQsj1eVyAtm7MtpvzDcZntAkSw
5TeRu9pIFPYU64rkEDQ+cGARO3u+in6jeBhCxaSc/elUw1JJDah0+URN3wdkY7kI
PCej9NEkvFqBOlWqos3dSl4/2o6z1nSUZXeLR1Fh1yLGPFSJJOY+KxD60Qb12L0M
dy4DQaCSKezb2WzxxsmlcBOfAfPham/GU+ThfzlDObCbBovB/xmktDJ8Am5uR7FZ
B5NhKiFYLYiLhUyioQaHmFlTHHwGMxf48Gz3k5UCnz5y0frhrs5kL0AhcYZE5aEP
GQZsIRto9jzGso4Qzf44I5aPi43qXmLz6G1kldK489VkeaJQm49+EXiD9yKkRXfT
/4zgYbwsDL62h+xt6EIFANR7ev0544peUZEklea+md1CZRC7bgmki8VYJ5iTvD+d
HxjaaKOO8/q3YERy4N1zivSxXxeFqPWGlMT/eD6jlD8DivONBIyhm1Kgoj12IIFZ
Y2BKzJGHD1hByhA+rCW6hiEo4VCeiBwoZrF0hA9cl92fjFAQ+HJm1sIUNzuyZ5XP
JTbEWBO2rGNRSJidfS2ByqskBMUfn15ib78MvcWMcXE6LA+z9dcGAmkCXCyXvuYz
t242bfOUQOf3GGRR5QhitbwkeziW+sQmUysl5+GqX2O8kwgdfN2jJV2zV9g2zMNg
bCHiXNQlB4/UKgpzxSL+ifyS8MVUDElK9gw3HSZqKkbWzRwEWvDxJegUtI1z3KQW
O0JdVOLqFMI8W+db3H2uSMsZXUDK2mgXvj1GNe1LMGwJXo8azRoa3aqaIBJGqiU4
CWKrEQfnNtGOkLppAFc6swQtab3VNAGJ8MuplHHB0zF6AiFlJyNoK5B9483sIzhO
o8tu0/9tieVhDCOLolotR7CzdwDt8//2kx2O0sB/XPOVZbRcgbJgLlq54ZPUqjTZ
8ZkgH7JZNuRXJmiuZW4E1wkXzwk4yO59eXK9B6SxoxpShbDqD+WGDVq03TdRfJdV
Si3A6FTEOWIKmMNjv/C3IQzKIJ2YBy8zMbcqsPiuzS3nQ0nzLxTqVH2GYwT1v6cZ
svaISHriNAOfjnAOODoRdtX8UojJNBXWldXgimqbXBb+4wExQajeiMcelNwOfREi
PM1+7Rt05PA1/0dXiSraKEuRjrB1ha8u9hYpOcNLIdSZ18eLJiC0ChWf8SnRumzm
5LKfmFu0VwHTy7WUDN2Lf6NxpIbGNj/sbD7XX5tuT1ge8BCzMBReWZKZPdSttGSi
MM3O0Nvl8Zpxpscuyd8Vyab/lDrc8k4bwWBhFGwUTIEH8nFk+lLEw4c54vwfbEUR
66AGZe4us3OhLdWCPDWTYTbESGfVLR7L+3PvhUP9mkb9f/h9qJdU0q+D7ZaM+g2A
NAZU634ZfXcUedKm6pM4+i8pVSErKZvrqkJaY51fyJcTMrOog4xHjNTuT1eGcnMO
/bL7rQnpeCiryi5SAPFauRcKT1EHwritKgMnS4evJOZbrgretVnE2/PPZU7U/e9J
mh/Cx9ZYzBY+5y0+hIAW8VZVUHKKgYD8YaTFgx3vCYx8p0hBPMwn7/9rmkNmZn/z
9/zGMl40zad5eexcpYPbqrEXbnq2+OLz6EvtQExhBHzGL3obAo+FSS8Ks4BgGEto
CI2VZomoy91lgEF3+fsOKalEFLr1uoqnRH3wHHxmLeRpIrSscIVlv95shIJO07XX
stBg140bGHMeXV/aW2PPWM1IVwRPPy5WO0zwY+LUk56x0hKoVTdQlkwCf3mASp83
1CV0O5QWhbzc/+TfHdVI0Iymyu3dcznm9/0oH4xvZCDgzQRPRj/YRB70/+vp7XEH
NqjgmncSAquA6yC3JiA/pFBn9x63cupVZQLMtb3XhimgS01m2G2RT6Fb5wiDn/GE
XqEXmQue1zpGgBOWkej9WLoWo+sJ58R47eJiR00uEPRv036YqJ4fD2PwYqn2ZrVS
XiIhgEFU6qI+co/Z9Qr9FubaMw4ltIPwLRcCmOVXPgjruWmfSBqi/4Pgxk6ZBZIO
Z8SegNv+E+xbgWkAQPme9ODB2HAFZOaPJ/jLEQdfalx9KKdXaethaMtf44lZTOwi
KK0dXfsOshHvKMuHCV1677hgKtvW/VKnZNeiFxkY+7UFbndiA63b3luipCtVweMb
5gXDJWbguJbeSl1kt+/FEoa9f8/8Rqanck3Q6/n2OSW0UAY6xPzNlY2IIkBdtrfe
Ha0cSsHMsBTrKocFYXCNIk5zH2r5Qj3y45jhMFRpMaLHaAJH0ZIzyNTLdyHbhaQq
1+v1uHUibH3mAaaHej5SSGynC0r3LRzporMKvcRPpJGMpL4i/TtmHqCci73CPBvg
dgm3d5pmMOb5lcp1tkxYdjHVjjqyk6uS16ajxwsEus1xmuBXRrm4Ybe5SIINgdL6
FkToSY8gQ0huf98pe65c79twBm7zTL/XiZeUWxrotr21q9akMZPGAQKmaMqS21Li
GnKLuKcN9A4gY9rxd80N7AoRZQgt+0NLPb0vDVjQf9BhusQw9zOB8Vy4+tE5+UPW
xQgUjNcYfW5+2CNOmeJGjQPhR+ki6RkWMv50xf28Sc7CY9F4zYBXyM5E6rqsZR3a
eqgw75ri3l2O3q0rv3VWFaKNydN7Z/nhtk7npRe7zkf3t8mANlZF8uxZXSqrmqGj
PIU6TPzopozJL1zGJWBXAt6inkjX7SOCe6exarXuqumb1cmaysXoF4eT++JpN5rn
JwCIoiMymDzgPuUAuIavTMNpCqaxzEmRNbtEomHiX25WeNNpCDngG88RuLkKZaG5
z2hmobjzc3sdGxn/c+02LblSxFFKi41Kru9AAz1ftXHmoqDa0Qd9I0AVNhzaFNJS
+nxvEqX53ZMvF5/SVqpWBnTOT8SDfjdm/gjM0AgQzMP4apPsidGnNxQgzc9fFdhd
EGIoPAyehw0h4U06OQXJpZq2w3Hl9ylwPUGco84QbONzk9r+7IlnnV17fbhvc8C9
AJLwbFgEGpHT4hu1jaZy1GyrfCburauvU13NARH1WpBDPltJf7X4aWhFOicU/8im
w3rxzuG/qf2qxWCNn9rwNzASfZFfT24kh4ZE1rZZFOabSMUDumIa/GFpkD3n7aVz
bwLt14TRnfV6y5WI5zdCER8OsUbyakqPxbOlDWFncOHo1a2Z3vlqn9Kpey1n5YOd
ElJZ8WqAc0XbY45lKP48cabHpV8SSONbaQ3FE4XFZGTdek1H6wUzt3hTK2saT7x/
A2itCyfZMJ/vVTV7V2J2dATv/X0SI6DFulEmVm6NyIMyMr3K9/tEMFSopvUTwDq1
Lssek1ll70VtI36GiPSzBFVtTXmoErLib4FIzJ5JIbyNjUN5r2OLxubb9xOqmSpI
eOFz02ieq/B+r74JIbXx8Z1eJAiYHjerJOmNUZWJQG1P1Z4/+fWZHeoCEOHez6h5
OgWX8L8RXCmQzCnHtG2y5OLNh+g+J1KBV1BBNKz1S9D7J4MDHz5hwKssuCLrVpWN
sbvVW+DYJpk7oXZ6MyXpAY3kXwazKnAkA8B5l+EwR0e7kSCJ5acqFnlC9CCobHML
4fahoSs0dniwZlATkSx+Oz6ZkAP8B7XDhHhyW1TNv38oVOd8NZfF2hRIfH4ZQP0i
/MJbsX5dSBuBve+JwPevjsGRdVIOp7WIYvIqF7Q03doMT2VTQE4OOmNJO/H/ZMg3
WIBweB9ypeWxguYtIGlbqwkyox72g/fFdQZYZbtWp90bwXXkyqHrSD0VECZxSPsH
J8EwAgYh0wViJUyXdt09kHgD9NBJQ/vVbLG4f3nLOkjiuPjJWtrVuSCuAD6M+00k
QVKaAMDVbouLKswfJFcR6SwnwRasadr0BcLpJDjY/mYqjbKOZduu1hRDPEoEzMwt
NHRAS+D7e8OMXVxQQU5mRyimjH86M6tx+j3eXfhl2fbVTcDFhXhXpE19zvVVTt8A
qjzQPH7i9+uliUQDEOykApklzfgEK24O5uSwxBPJjMJNWpNEfKzTVrEJreyfbENE
3eJgHvrrdKjfVFfwVE4C4xDTeyQviQfaHLXjv7jDq16HT8YWEHOzizg3prx/LgAv
HawQLJbA89mFWgN8GmqdGsZqQB3uuYsU9dfWorMeZxiJ1PGUWUuTbLwa45Xa/q4G
sZdyU8N6edKASH6jHIUqe/GqtzTC2vajCatr/nZwNJDlEn5jf4vJ+y3iMNjhSxNW
eZ55cqCc11XDChkhYyjA11CePK0AHZCI7akTyjCpe86xC135WLRHTzk1mukNNml8
Vc/YGDJKy86CH9jayabpQH6NOworqfLbVbAzUiq5CKH2qDup6/jQlGriCIe5ouiS
nNp/0CG8i52LuBL3sbAU/482XjzxF7nctavgLL4S+xpype6RcG5Ndwl2F3RkQR8o
UsOR1iqwtgrLQma0UkD6PT8gnGTNgZLTUgHK2qr+zFgWDHKN5U318ay15MCCbaUw
87GH0XLestlXFb0IN2QK/jkGCaLlhCGW3nS1V3cLD+smW89nVOtL4ULUA5V9w2X+
EfvbYdEbhx0JpUhb6jSaH+3fiD3kNXdxFrfNq1djzKy+FRwRdtZtaCAm2KpAJAS0
lXK+6KZY05tkR4zzBi9aYn34lnuLo9CawDtzkPGGEqzq9b+LLWl1nK8U7LjwVRV7
ksFQULag4J7sv0PMTKUnIPVDScnRYM78at+txWJZPdAz9eNQW9OfClJlcJzRV4lb
sCwDy8iYJOVSoHO8YzBIe2JgvqGE3abb5IYXMqG420Ip1cC3NiZOxIYFbta7UArl
15MLyIXElLA2vMDMxbDAzes7xuPsKljsQOfmLNmkeQ7Jat8o0CN/dGpY0tfh0W7D
arr26CXWI/nNrmoiALe8aSxnrX+rp8QI0OVOA7bxEq2E4T+yz9280jc91VVPdOFY
A5T/H7prbjYO3ZC2fGca7n9gVV5T+i+FBRt9wUx/VYXQTi8KnHi3Z2trgHXizFer
5QBtRstV0l2nc0W3baxOPwkgbQECORHHSvGQbnCw6dPw9vl8arXw5HpmDsDFUMw4
gzZi+011ho9VKQqhkitN/Ec8z9YIQ3XvODfDcBGEHIEEnQsZd1DaGBKOUw/R7Fff
VaTN5rNGfkJPwahRHeeIuhcnh5hrHSp0UCFVhZWZbvbDL+JynJQlPmIi8fXMxEBR
ckbzHfvZTF11p+4gg8cPtPFEBXXQjyGgH4iKycEQanvJsiGMMuk6c5pz2p19+M7g
4CrQj0CIqOWn3Dsze9Bgz4xqrgiTUk+O5UqAsWMOGffiti/ch/YLj4qwX77MSHh4
y1p2yHIzRTxqIisN5IcqxBSOMH6duRrTjx8t85tFSYjAFyrdJ+M0sraBZ1UCDEaO
2vxsSjg88yNlsiq6IZm0WilkY/6GlXs6EZV5amdLdxQdmbEgt6y4FvXil0yAsci0
xMFNXy1sr0hA2e4F0+o0cVsQsPWPxc+DYvgULZA17hnzxrw+n7Eb24rnFp0WmwAV
/naPWrEy3fzf7FiL7ehu8k0eo5YdT0Ewdyv6vVjfhRv0PUcQrsa36aMIITYdxuQL
GKLUeC9AGuEpdJrPuXCfhrvUnnELaospPHuIWBc75QgM9vb2AJNL7s941syMqM+Z
8W/BiY6cU1PgsEYHyNGzOer+kxn2/n0pzy3BcWN8nYgRyUO8slvU/WcceBqtXJr3
HLvUm7cRmqUSnpkNBLPQzh2SNCTHqLO32Spwqakd2olUgrO96nqae5d/SXw4IY7c
YtNAeXzGt1k6KdOc3AWFj3I49iAbmPRpiefQ3uo4IG04ulhkArQx0MMWgPrCLmvZ
9zEFbVs62u3TP3aMQtaDNFC0hTTq0BTry2XuTccFz+fvLumX6SvgdiDNaaGBjPk3
UBxat9UkaP9yauI7RUmee/CHxv5zmwE5pLtOw20+9874dzBll1uGm8LIfkqhdCj2
d+LUtt8ffnGpPHk/7F3+wiRDRLNWbvovykuNPawhuF3JIyqAikSCQiAz2qtZk5Gk
OQx6s9l0NJn1sbdj1yNkB7oQYhBX/x9bip7Frl8/t7Xbh4xWcoTEEC9m8zVwXZiP
6NZFuglw5KRtau7w4uJSjV4+2tgfD4gcoDbt0N/uinF01XuBG2FTsAm0UPJwgc+h
PMgQ4LN1+UUcgO2UVO7GsycPhBslT9EbZytknvH+sPr/fngN0tSTcSUPAIjakzdw
9qqV212pKKj9/tb738mj0snKWBIRI5XhRViVH/CehquW+Nru3yWcoSs2MzBphbgH
RjdRiro3gXdRSoss4JS1qt/3/dgAL+zSrs95zsu7X0UTNsDzJr9+gnhwbrKCf5x2
nMxAIWKsaQmTC5+l8si1ezgX3glihD/nTW83LMaA3St6y1IWo/MkK92gwvLmjkrY
TNkFiNaZwDvt8uhbGo1AunJyQQvOvZfPqrKgNkDoJoTkSFLCkbfZe57bOdiyxbD+
sQRmoRJRi8myqeT24sEUzapALL8ZnHhbStwbxqiMnIGCmNWvGacyfvf9NnyvIdpw
inkzomjAOUy/scorPI482D/LwMZ6Hr/aYjUxxJ2s/LSn+Oo0CLpPVCIAzjoiz/sq
ac5HxIvuzhd82jZVvmoFV0JXmrIszsaYsuGNy1aaGIV767M41zuWBG67dE9CPEoh
POHqxJze5uNweE5yp24Vf9NdBmG9LIwk4bhB6pchyd11QfW6y2t5WF0GkddBbp6C
2CAsI2nU0bowmeP/6nn3BK3FgQn+/VeY077J9eefJpmJFZW6AQfOh9xQF0bGH16E
g5rVj7BobiFUGiTQlpPqH3w0oNcAfs0tdwqqRGyz7qC/bRcD0uQl+Tx185nSF3Kj
tWNwe8Z04l9frCLfxdCas1ueIdMeUT2rCci2IdhD2U9nVVVKZnarbge0jGWrl4d/
IoDOTl/qQopyCp1wKkJfvwgHSW8opD8OMo41lcIIh0OPnLKmxplOQP/BKFMYgD4R
QP3vjVKXOQhUwQMX7vF+V1COmWQIM24TwFO6AWs09KONoMBJ77fz6Sb6C1OjSfgr
NKkeRyyvijgueBRMUnel9utHpkC0wy84/dm88Z81aO43Pg64TxZsxFQBFRW31Kqd
qUqK2aMCgl9C+V7p8s1aaLHmzq0wjwuFs/TGd87c07ha4W/5V8ScrikbfhrtMLid
+1Wb96YC/7kmEzHkF2kOAzYFSeRobJle8US8SSaudYjmbsaGSzBCrpiFB1wt0NBO
6KcTc8w92yLqrpN9IGRfhb1o1DtSjTMvJTKYOcAqvCu/xhL8lXBCPXk2eh3ZgkAU
q5lgJRdHSM6Xhyw/vRtt0H4MytdEVsVrKxdQfvnXbJzUllxZVgZzvKnHaN7jNX1Y
3Dfs4VJ29aig4BCm+69RhEfnhuXb5o5Pq5d6zbFlekfQpSeujWfj7DbkvCnh8Ry/
IM3sAwN/hMpiTa1yV8/nM7joah8eZIcFOL6WHDebroeXIMF27timXibePWpiVHyD
2wcGt2+B9g4TZ3zrqoAyF4S0YI7ORLO9dG3Ag2PrzgIXZJIX91vLJ83kk2W1QNpU
6lkrXOczEt/TjSjPxsKfuOdHNNk5eeoYg/uQTlBYWBFZ8v3uMyRI+5JAte8kQPef
Ki9+T0yZnwviu47l30XiXvTGaU5wUpZscKeqB743D756LugVg1kZzVa3TV5eYfeZ
SFjWzPUnsd9zKQBVo3fv3CKySc2O4BhqnCmLiasHHEceSgBa7tpxrsGWQTRBQxqu
OoC5s6Fq8lVzyVOAo1omr1/cKFKmz9152F8IQ9E5ppygWOr3uOqz4cQsZ1jau2bv
ty/v5QDoX6cXCyiN+7zLBRgi1R9QHP5/1lkPIUnSpNiVLvb2RT0RKZzY3LkEEPvj
F38F0sFW7N1X8f2fNA+sNpCHOinWlDhufSlCsr2V/qPO9GARHW6rQzVwm/6E+zjt
jPE0GWL0Jx5ZZmKqL5BtbaBK6EeOfThyhJkgw2NneD98VLkFcIOxnX6qx/BMon2p
buKT5Ur8Dwyxt7rfnX3MCofJmjfTrzu3wyUY+VznIXxpbvEWvmOFQ4rxHN06fzuB
jbqqg/TEJcaTWOLiTwCpSQ==
`protect END_PROTECTED
