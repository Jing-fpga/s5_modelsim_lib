`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZTjij3Jkwigppl0I3OpHVpa7nYGS4OTfs1Kcrysm5OVWpwaiPmc+7HWGMDpJ7Qn8
zTAvmr9kC4njxFGpkPTMVZDUBvRg5FkB4fE5m0C/pj6nU+VTIk+KgMTwpea9pJWP
JLqgUcUhVmLkX3cEgVOWeroXTngDZARkPvAeGObLOvzle4qwDi3C1ZJ/q0EWL0RN
0CszfLt0TVQEzyp3x94S48Kc1KTNrQszVsWx1TApKeDI5hxE2mXPR8y6qC2iRPXH
z1H8DQBKxNbSwyJDpBEQYE6sAJxn4I9Q64L4mdtEqcz1R1DSYKLVSsd5CoAVMtHn
9wB05kHo+uL4BEGlG8YZ15WiAFEKSiI5WYEvkDRUoeMuk3AkqfMk4Xa3HbKRKUZI
687aLv1LmFORaTbggj2R7fgnCpLi4eyC4/PtXeY9fJCPZwzHitamDHUmThAw1xub
M+VJ4m7WsdKYQevXlMP0Rt8HIyIkS/P9pMYTYyBbhL8dQP442ucsHWVMkvSx51AI
j40cEd36c5tgsamg1NWhAcQ8dqqaKd7uNPKebyiK6pSLqhWVNFG6QHIW/RMwPDBr
lt1m1BZ2SrWJRN+dhZ/iu1wf+gwF2TDIJH0S4HwDTkTi+jbFamHNuNjeBoTLBvtQ
GJSlscpgHQWeQHbJcA7wVA7bGHZ4dhNK+ol/GHqoGTZNpMItIT63JlCnPDlWrvtH
RLcWRTQ5FPf8cxP86dT3XKWRyQS9vCByMNLC7/IcOdQF7/o20seKBkpr7MawjSIn
VAttLQRpr96LtGSGeP1JwPBtOjbZa0sW+28IjgEg8GubCe2IIA7zVAdmJxADzreA
A3D4CSh96CU7ucpQElJqnYClAUvE3VCAuN8QA3/ef2ru/09GDXMqGfKec5ERT3S+
r9Z5WLI97gaBSG/0+QqA7O8plFkLbx2FCIPH0Fh77Y71k6UQ1sO7E8Hcm8gH9lQ6
DFRYAVykXgwXzGqCdMYAAPeLeC5Cw6NkhXN58VBBWiHYNc80SXm+iAK23C+cfy4A
mQKOd/TH90szewD8NXFtoNFZLsZyVIuTezwfcDd3EPlfWWiTR3HtZUfPBMCo/CMa
icVX0izYzp5ALr5AUPJRYIEuF8dKZXtx4L8JTU6SAb/y2umF5ASe7ao+qdh5RAnD
6f/TQSiI+7FL2iSST0jG7S7ZkAv1UqgFeut4kV91LMlVmLVkC1hJSTKTJUdArwU7
zOHSQY1EKpyD1vnJE6PKwzzKkA58fq6V9kpRb0SBKhu/ALnoRyIQ/z3dlkLXNB2+
kbp41whM7KJPLIDHH7UDzdoXFqFBBS0gN4+ouhK5CrmTm2oTCqKgkLupS2wJlV3X
d5Ow4USVWDJAxuKnIuK/ihQpwN5MHIkpD8umYfbdEdJGByB3S6h4yil0owYJVhI7
80phzoh+CiVybY3QvgpL/rOa2qpB/6X2rPns4NTh+jhtJjiY9frfIJswxJeMWELK
2Em/82NlSAbINwzDxBvhBOft+UhWJtfB/YB0mRTYGtZ2rNSGL6A96RfLvzOC0PFK
XIBwIvlc3abLrE/opzzzWOBxEW7bt0PYfax5HmYKsw50FyrwpYlmnrmbbwVdN/LE
QAdiDbnbfLAdGDP/5ya6io5RzcYGkosZDxgYdEBZk4/IxgRMCiwWhL6oGrzGRujM
UUv0Ebs0TSBVzcZyL7RiGIwEnsnlIuwL0Rg9rsXCdM/Yxl+wwJS9vzL5w4D1jojf
N72piMiZRCdh+Fl2D4C3wpP66o8+/JOnxVTJNMlKvQ9WDh8BPTETx5v9YI8F5Jrz
kdjRar/qs4fdQHVWS0cFTGDJjsCtkUixfPAPCf+PQuk=
`protect END_PROTECTED
