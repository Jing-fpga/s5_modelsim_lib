`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DY+J5a9Ug5uyv8Pxe7XaGRcOyBP2vsOS0D6LlYoRKtJLxuFUxHq02YRkTJogOJL6
9H1I8TPXOaFylPHHIjY3yeByFLxP5EMPty2rJWvdighmGuywC08lCjrukvS7QsEL
C3zTja0kjN60L0wJI6IVq9FQ4RVosl/XyH+tsrEHiRxCwNseolMM3fIxa6+T+Nun
FoznRuJ2u0TuvG+BA19sOAC9BZ8fgbZDQkn370GI3R2igHem88O2TmNbcN+5nVCm
7/emosH8pa8qPvP8tF0Ezj8XmLasCA2iwPEL8bRTaXo6A4gxE/yGXBS8z24quy0H
8wgwhm0RD2QOsn/cP6Wi9ZsOWraOoN0JIaBI2p91X4C6FWdSZpvfLjPZVlxZ/xJ2
N9qiqSyLprOp7VuPg+9PSPXLud2xLwbZpj6AtoadbukU0tiscz9gRu6YcH6vPwni
f52KqTiOokR9fKPf4z3Y2SluG2kwZPxFtY33a153qUP7ovW0F5mV51/jOnSUXv5V
GdgmOdDUuN6od4546vlY5I4GIyxXZHzkxzKPY4YzWk7lPP+rf7MXjIL1vy3WCEol
/Y8eE7M35FcErDuHnW/o1a0i2oeM8bb201bAhX5UxPJHyY3XTNp5IaFHXQqP0izR
AgQohj6v+/NHdMsufefI44FiSiidQcUZZNWEOWhAGldJN49OEC6rm9RdRwnaUFqp
t+hNULTQqwafiP9quhTpOwgCfGoaeFMMS4LFdXb9AVLNKPgQhnpPWIWiG2Rjp1Tw
O6DdKgj9W6kos6Dz/5r5G5nhY6tlZtIWyRIKqI1NqEM6GtkseGqDgoizcXj0T2ap
zecN8yeiiWsGzMuFgpKIqtXxymXGspklw7CYb/ORdzn1LivA3bKi66c38Fs39b2w
96P5B974tIHK/qz5J6BuHR2Mu/aFCUfWSRgMOGYHgEZ3M9auDqKKeIRpEVMxpFTe
pS15mtWMIKxbJbKvW4UGFN+3mnnY8nOSXCXR0y0KOTGQF6oOLNXiSM+Abza9RHP4
61LewWJOQM5szmEqcgtdnJ/g8TLsD43KlzyjxUoHwVHWR+7ZdgpYJFHBKEQ45lhF
Ng2V/pUFtJrbqBJCc6FKJ5zdobm0LfC02Wi1/Y8tZTpanoUSZCqtUZNRZxaDsXiW
3JKpHsiqbNN5n0SoFYrwMMUvTbrfjE3ybVy8+l+5skl8osm7rDjh2s/31g7zMTy8
8DdqLwLLF7+mP8hbomIE4BT4o0wwqDelhZdaWnWrdOcmBh+n0AfT1uaT0XfIT9Wc
4qy3Y4ueNZZFoE4QjSQXqMVITqb5v33jygVvEGW9s89XcBmqMbMOmQeWCX8XpXOJ
CmPwHf8T8eQ5dt5MY1BykTZqBEEquhqXP6UthvSr8RGO5y8iVDlWTnY3WUs2tRjp
SqsPAcv5wWJ9VBASgo4/0lNtJ7qycCwl65UvhrkEh0ING/U9MHaFZzO5r8PD8O+k
HM8DAhJEWvDViQjWQ9Eyd5HdPruQnoJvcWYaesuQYQP9qh4acO2cLzEtigocvOi6
MzosX/zJiQrUp4CeXKX1ili+nePrhguwAOMeGlOb2IkXeN/LAE+AJIRjAEWbLTkP
R7MpUP8S9L4CFMbTEmzEcK96E6cWcuRQKrICxqGbfpXe14cH2LSgpbI8YPOkLn4b
w5js2PzQZavHLSyyjLL4qGo+gsYhal2fm6IB1U++5Ml3f9odcToqpmjH0G4lWuCk
63RAVAkDfcyQG8vzMj94xJbrsWVk/bkHPeIUvVS6RfZv5vY6o3qJZiMdZUdUcjxd
rY1ENjRGG5EerifH63NshUAY0ABOAMWazRzXGBH7uiEqmJhB+yMhnppX6ReQngS6
eUYLWDlsOquR/zGst/c2msPlWgiQjga+kFEdbrNt/9NPhFvzQXEllu+ddjH7degZ
W5j9IhUcSmTU3qTF/sKeiYFVx4KANqxazwqlJg5frXuxRTzFdBzuUk/fDPsHENH9
/rIeZzMt9l3mv1JwmxflbMQANkIhKCbvoIVekF34nNWq2QQKCS0v2SpPdfhVD1W5
Df9jNhXbh/SWjXdZqOekXGZK7Vsvml1Vy2QP5khEUBtHbFJXaHs/Xzuk0pB9PT3C
uowG02/62fDO2QFbCC3syYUCze3f7QYokvniPZq/Y8+NEj+TPDNBjkn4EsOyQqU3
xrtUDEJ4xKafvNWXjMO51VulHiUBAqQ81islG80GlxgilH853PZRO5ZP9/nNeyhV
DjyEREH+0R+6Y5d+DCVqWhPw5GRC7knznDTQLymHfuB1Etc3ThehcRqL5sgq7r/G
CIkiJmI+BiRUhohBDfgsJdgZB47Zg13wEo2Cdyksx3gXxydcqtTaBN7H6/kOg95u
m/xs6O8aRjAGMp7lzoWNVeh5cEga4JRRNZJp7KLWnmT/cVrarKlf5ihcQdVfa/Zf
S462YqVRYU/wqoH6Gs6MvLWEtqpQgkEYh8CGI3v61HcenKIn4QstmwNO1RSuCqpE
zXtrci+sqiACi/zxpYhLndOx4pOeDxt5JbRXqQDU8hRmVW2UmIiS9jfU0mqeH4l1
D4XIKKv7KMzuyTc+Lv8bLkuWn+TLTWkwLNCDbqyfqfgydC2RacUMKXBs0/XIUJ09
wePfJ3AUJjMqS5xyKYFQ8PE406aYJwlpHI9YxxoCxPyfHkace5QWo8E5swnDDE+2
/7ZY5DBnSu8+71DWyyMS6p44pRZnWh4pyUw75MqlxfUEdh24tKUvBCQrYKxV/kTk
uKf2UhTEWJTEaugb0d6RMuBuqxhNAICSOoEMU+DUZzChRCS2/teaUaovwGoppMFl
sZnvHoPz6huvRNf9ETJ7YjWq/mZUTaGT5Od4xX6vaPFsU2Xce1XN+fYVorIjBKan
SaPVIj/jsK5tc2x54stBjHuEvdO/B16/ZefSKRE2Gade0MH+5murQ8fxgCTofd44
ah8PWd/TI2qbbJlN+U6SMA3lFXsukMPaqup9NvkOYCSdg6zbCPYzG0g7J3sgW7yQ
vEnNIDZ4IW7ngY8o5F3s/MgVLJPn5DOx1k/fb+JkM9dgMk2zgTb/QRBCDGwB9Vuq
3tKuHSyUh69zcMuvAXLahTqrzG7AlHdtG3O/bbvMjvmcEqguj5KLGml0jLHOb1ja
oDQs2mrgpVG5xZWr5M7LFgUa7+uVbLMWSWu689/7e+AsQeahpXFa/jRgqV5S3rmL
WpSrQBp9NAZDOL2MOViK377QnUJ7k6wUgA2oqVpjxysfwiNv9kkDCCJMGB/hs704
HfjYCPFpNCG9+lqyXQrKFE16cNE/KDfET+Wl/v5qKVtLKU1Xb2OpG5NJ8ENGG19B
drWdeN9ERq9A/lCHK/EqIQYTk+C4JiFfY23xHVc6HeKQuNoPzH+Ws+weudBRYDjU
BjLJf4C3tvuOkKFpo51xrTZmJ6L6Uh7o+yz8Ia1xhNKo6VPxizlRJX+Rn6Lo8pEC
RRw3hHycDl28X08QN+FG+5DnwGIxPF/VX2qeywwEdCbd/NFpN9FUTe50AqXMdSCi
1oXOP9r79Gf2He+bIoo5pIbYelmACwqt4lKFxo8to+iroduTWPQ8m7eri89xhnU4
2wPYF1S73oPHf0BA0lLutYV+t6aqDwe/7ZMHjqf0pTi2T2HDHY8kdaZRHhaXC8Rk
NvWC3OJiAgz6BEbEoCbGSjtm9GUDFV6J5zMLhMbbtweKpsVB53Z5pOUMgPLQSCtI
xkv1gQCP2nT0RYwJZOFHsQnBQZ0cokY99ODbUVIEtAW9nquXbVKMP8vTsPOlGavH
Cznb5Ya0k/rCcUqlAQPCsab+Ox7bja5hgHGjgW/BHVNZYLPnz0sWmSycnaUESpMm
zLCIZi4vpRMfnqhjKmI0xyQYao62TUjP+NZes4DiSNPCpe+I+uSkkA2kf1Jo1nOi
gKK/DW8vqep3e3Xs+qKl7mI5VUMjElaFMmk+MbQPP1Gj8/+NO9R+ZREpjpMK6Ucz
ddGxZT7EerZGdXjhWFjIJ/5gVY4ZvdbIUK3xHN7laQ5Og3GITe2gf6IsgGF6KOZv
8MR/7ndOBFEKsQHpBCY2vdQQWVDVayDT01/wbOAuRMrfnm/aJRaFA//BbH7c3WYM
+sB7wH/UB9rXbjVJZOm6en+y762fP/mVb9s8QESeubHU4y/jUS1eUH8IlX1wNmO5
`protect END_PROTECTED
