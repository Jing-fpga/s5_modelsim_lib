`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d8hOcYxCucX+mMdTtrruzFfvGVOIB2R4nw4wOt+EXase/HIza9VTtNLDhoGy32EJ
y4Y4HCYWEXIO+5mZZ1FRJ5mDj7LPHLRzAnC5tVNA59/mGQbBmdmihCMnmVbqhtly
ghtwzfJ7puTuEyYjwC8FAjDX8/OiQ9AzxlS2AZZ7tSIQ0JJfvmqEPblqaQzuD2eC
LcJe3JH6tSClkkirOJd6Q/gqKEH3JmM2LUp+TgxU2Q4NGMhBnK5N5D5zveHLrArG
h+mG46ksGzC2mYMU7Nty0fu5HOkYmQGJ4NpiPS0g+tZv9RMz7Q4K4NRaYZe+OYKn
iUmDvdOozYP9AdUDgFSdWzVo0o7TQ9H1tc8JmRyrvopbQaGLp2dSCDHfWKpEoPjt
WlYAv20gfh7H06HROrsiFpkaBhOZjEj2CN5EsXgQ41wWDDgWfMRmKJdG178YUKFI
KTy0xbX/u4SB8SiLeiOFNsBBAukRFP/YGN2CdoQcS+feGLkSL8hko2xP0NOZRp0v
pi6uLRoa622xt5Uxo2H/SCsQK6ALsFgXu6DO3axt/vTuzBv+DsYhhD9h4OnBT2MF
dCpZ4lz1T5ypO/XL6NA+iIQoFQCH2G9CK3d4lsEjM9qkUGIkWFrunamAxMlfEX6T
Ctnlv4y87W4ukrw6T1Nok21WwesC+Md2DbmY1T9YKei0BoJGl3A3CZaNgBd9RGpj
LbatxPbF7ikLb5sGKauH/FJyOmYPDVUbBGZPtUwAyPSrdvqeuZuR8uB2CIpyRWsR
sn/MHOd9Q6WozGMFfFCMs8FllAG8CV/Snh/ndlt+Xaq2+NO0D7i3KSnkKGfRfdrb
Q3RUt/z0pPIS0IknM1kAU/4/OrJm3ENEPjUQ/iZA6UmueZlHDbZYAT9zW1iFm837
vaeosG8IlNAlj5tAgwGK3PxIAQu7jZLUESjhqRsxC3IJPOusP2ceQu2UCDjxjBxX
bZYSOQvnTQFKuPwqHao0AcWFKRuAX038EvUabcjmpSgohHcuNCYrMlineqnoj0Bt
b6C+kndqyr2wkVoIvui89jrjw4+v3qHbiF2tHTsZe0cUU/mWJW2hEzOZY54LAuTO
XRJRlo18EXDp9KLPgW92YNcT2mII5J1H/QmEyYEUgwl+Lf04Tr4Km/XQdCIsiavR
nsxVmotKsq31BnZfGkeBgSejMIkbSePKtdF/I2TYVWw4fF+Ruk2K/dN7vpPIwgCh
GRBnc5UOUZjaN9adZRv9+lcx0aj+fDmvxnfjrUkj6VGNECy9o1q18arFkOlXC6jo
6h6J7wCtAOYOCD94LXp4CQxbfWI3Be0ldcZj14bifCmycOCAlLgLr5XO+t7hk4NQ
vHuaCND/YomsyOLQIwZ3JZNOY1cjC62KzoY4xA0qssFvzpkPZPlsCEZea/GtW/Zd
d71pcLGOUN10cOcmbEjEQ45OGft/mNe+qdOx0hExXY1eTY993wzMjmdDs6utsBsK
GgVRE+iq0ONqjtG2XmnJfYawM5XakmWvEumStGAwfqEIIq5JlgN/WHO4H8z6tRXn
63hm9zfTa88OiCdK9bkRjCvhIoPBd3LKgPBvLcKdsK15DCLIg80jZbQp7+7L/EKx
Vkc5zqJQQcatvB1YOTC3bAS2leOH9TMtsiJybzN7oBYSzJmdrykxHOnUJt1GOEik
yYD4twyehjWfs5Fggm7mX9RhccwhHxtQNK5OLmiUqb6CV1mnW+2YolMW+whYWgSN
D4dkFqnQrB70mwsYXRQ/qnXnt043XklB5rsQ9eHCVdZaNP3ZP6LKv7mIs/p1Y+ov
vOLRBqHiMH9EkwlbW+A/dA==
`protect END_PROTECTED
