`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
maHcdRl5xn+J3sjPQb2GrR3L24GElF9HQFZPugRbXQPaLepTKAiqF5ALhVoFjWU1
ZD9WNE9r8Is0uHZ2+ys4bLx+CANMwYpRYYAeu1JGQ83MSMH7PLLyz2RRboZZDF16
3M8kIPscICKfiV2emqwwo0bPf0TATuKA1o6Z5bQN7iLqwptF4X98RZ+iffFvJqFr
BTRDVyijghl99so4ZaWs559xOAIg44ydtZPQh42VWlKuPjQe9nz/ZtDj+hnSQ501
kIx893b4T5d7m+WLb5TPpAEsBACZ166D09UMeP3YjOTYkxYwWdSoYbzj35iMgvVt
JRYbApcmknXS4ei0rbnvTWYN2hQ8HBd7ddWi922bhexC3xSDGVpRs3f5zqB/udR3
jgM50GwHyui9al2IiKxrvTHvSJ5m2EU8iJXCoZ+yEmE/jjLP3VmaoMh9A6uAajFU
0depmqF7vDmm2FQVWI0KbUc2x7dMT22S4P6LjeHazUTXVtJ4AoCBr/B5jElkUw6O
nVEXCchUMp8kKgvIfxTEi30flNlrHYPBgHldoXZm405in2V+fo3KRrbk3DwHRJxH
hoJxlXRQ90lF/twESxPRqff5yuxJmsePYP7ucCktUCrBo+/swSW24AVTJmV5+XWZ
6uE2k6FL07AK5uq3+pGv0wffNmQJzRab2izC3K+swYBWIZ31jJpcFvus3uAYkR9y
UKtDpTmAPmeOREAcLMwszJO4uBSUnW53RYWLwc+NvnNb+8rWefU8Lqw/qrPlvtnt
SzsYePUdRlaxX0qoa7hEiW/le5Cq16tUM/23Db+mv8bespS+9TDAnULd4Du3vPtG
R69B3GTm2VBhpHdNBq3YQeEOmNPJmaSNR6q0ynfSbQkKgI5J79t8xpLF3cp08Rst
FFBJDnmU90mE15wlC9Pt/Wfo6N0xK4ELWOe/vV94GWmFhFhdJsPn30BWDl0APdd5
e8hCyiiSDnKSO5rTRiqie7XUsr7iyeEw+T3RaYaRQy5PelkknneSBYbfW9S/+ViG
b7qvvGembqsO6T8/fhM2aZITfQMeiJNJcuImX1AucewtPrGR6LqaUAyCM51rTSTP
cPRFqi9iz10vRCGpq2srVwLEt8bNRU9BcvAZKG9pyK3O9sb/ZZa2Q4+3M/vGe24e
tdaWOnKClXhmNJqUpc9X/AxlB6WWox7xwcaNWZe4YG9EG0JvBwU1r497TqdZEYA/
DYPsS81n3C2gzWPUM/f3p4GiSHDpWRGEQ2UJ7uIXBt5CNIKfsyfejPSsuVvnASZB
oeG5i93+B2VxZ/zAat7gBzqQKksiZQLxoQIDCCwlw5QWMHxbGh6UOFySD4WbBXUN
ghal6z0DR7zw8iO+7qGIGjNl2/N5FAgXY6BQhqTa2FePCOAmWbvFoZHus0CRIDwA
PLVmeL9rU6aqph4HqgLgptdehyjBBRUuFcRtTdphW6wz1MVKyPDYON64Vc4adptl
WtPloVrr3jhVX5KYNJpv3hxmeOPfSHPHL1jZHeyGC1KHFGE3HRklzZ00WDoUJeP7
InXDsjsvOY4JwKV+uaYzARNrn2bYrhDhKkUzJt/YwdveqkOAGzEkh5bZK3hVYMyo
5Qm2cwC2JVSy/3UTZsJKthFfI66xev02Bs7NHpJ1QONRAOb5/lnYrktgQd2F56EM
0Kj5NdzUecyfj4ZFLBSuiDIi98vpoXbaaCMQtASJ8Gbo2SCaISI0NI0+L3c7lkVV
AWTr4cFUzWp35kr1QL4CY+lQiGkf1gwGwPafwBX2S0HvfCqBDmLP+DpxW8cL2N2I
CimCS31YlJVyqNgBu2pOVYId0HzTf8EfgKQ6lKTo9l9tUrX6e/mhLeoQfuaT6COz
87WgJeuLjsD/6Ip8mlqDzdTwGsflcBks7fINDMRb534pYVmg7cPgVt/tHY4+LpHq
TyWnX8l4/yUGxkHVv/3BpzntBIezFBcWdr741gakK1KFB0strbKdxqB/dC95LHob
AJ5HUtA7y/9vodIhchEoPm7isiesnmCV2sOaFTD6DjDWbtxGnYyg6QLvn60mUtyH
DMTmAcqJhw29yua4/Gg8r66DQ2KQLUxvuKR2iBVorCTt9/vcYkAXEP/TVjerBTpM
RvGNqlzdJ4EUm0P91fkwip2NW0ApOmU+qAljJBCcFmAKQMeEAZLi+57EYUHz3gK5
VBpAUfN9Q9kbyqQfVYN74Nd0cKuavdMT4BsU7Gkc3oAhhvBQt6aujqinYbHwUPfP
uPMYCrGF0TiexK9jpgayKMA/nQEVpS4LcLlGe31Tn0VhFMFC/RDH03QGHAF+8OTY
IWprz6f/IMYYUKMTtraanHW7mdpZfqPsLwDOlVjR/5Sd8YvVZYx6ioIt/INz3MCT
x4yoddIqpQXvhudr3ikmG+WSvXwExTFVJA2HnC3f4uz4eQe2aLZywjR7fV9TF/rG
z/xKoEZcJFdiz1/+k68sVj6Q532u+Qi6ys252UCsZ9nMnsyXJFzK9oxnXmiQC2uV
+mojHS7ftU93KyvmiF3yWy2ewu0TemHQgwNG6B1YtnTTjIc5LDtynNKDHQwjzukd
4LzOg+wv20+Qkii48WmPWiaBHCB6QF275pE7up9Y7gych9hXAALXK9fGNytRpdcY
Lx+w92h1LprTSb9blg6FvZ6tAIMkBaCbwDFAFs7ap+8Ten1xEQJ8qpwnOo+qVHIa
yWChawmOxRYzhWxIxqtHW3kOm8APVBaqgKXZ1NEmB87aqo25gTWhoGHHqU6FVzfQ
4ZZZkj8UmYqXFqbQMARR7yXefAHzkhJXXxR76hN4rN5v41wNKiTtFgaaVG5SAJKI
j08ITpRrtNm3Gesz/gP6ROgcOfyDdXe1WQLem2xQs5ZdZ2BxbX8f/Tyrb2IZPI5V
FpBw02yUtnPrf9yE4SMvNf+6MTSCZSSHu+KuR7+tO0ZUcIEX/kevwyihSPsZ6key
aGu8Im7W/T6KdmDMjiTZkPujo9ldCFitrAaKzP7qORor0PoPedXTBEb1vA9WKcFB
0Muh9pjI9J7HHDi8H61bscnv9lJmW8/l46RjGW4T0LiiSEHmvSYs9deCY9PkF0p5
22K6GxU2yyxz5VAdRaA5Zn5/cnoNPFt7VxRMh2x29lOJVgPxVumAFp8mqAU1rf5/
vuKGxjS1wwZ9XY64eybd9WwBFiGbk4QrJJ04AfkTbXjRyq5PE9TvjR7zsTiapZz2
bqzy8tjion8pjKpHj01t7cSYUq/vtDP7qE6cPgbS19C+4GriimsITmB/rDpAv4O3
igNWu+PFj0jCBQYE0VvXCsc7cGjlqjSaa0A6Xqaf1VX1usDXBxDzqGnHZNLfT+P2
zzxP0nxUaORcsDqcAc4orAsjjjlNCp1X7gzBsX92PyF5Qg82T7iwIGkJ/krTIiT3
Gfv+qdlx/Dml8BAYtebrYu8F/gH6HPLQgEk3yA6pUBYoZTEAqSwSMPBtbWOtculP
3jV4ahp1DFsoLIz92fYhl9o5K7/8Id/cey3GZqdA6U46OrAswPlDAEX6VMp8t3yZ
p4IGeVsq31nAMeRwLxjhoVz5L5MFZcZifAj7VHYaW5rXMQgl6yR8MUsgQmmPMs8Q
rybQgS6Xurpowl4VXoYhyIX5eP3X+HIbqvxQOwSDPLYMbMdmnYYdVGG7tP1wcQbE
z18Hwf7hqnSmRc1O/whfnFSRCGhUDg7EMChQ/KjS0EUlG/BHLnzAZL2I4+2BW3Tt
yiZWavpe5KbsR+NvrazxgcjLgTOfeNI18WIXsmiQXlwowH6pEa+ckXttvrMZy4dc
f0gRQQdceT0aQVEXEifZl502076J6fcVhYKx8TkuIcEzf6Kw/lSJaoifXsqi6e19
SwqrcaqBVA1n+WFNpXJ4gH7+datIkWdvAPNGbLHHJXq7pDiY8VSKpCYgZofZNlXb
30jDOJsgspuyMtJvFydVGJ7JtiWQB9/bYs8A11GHeyEccKK0nJ3ivkot793FGodn
CLuaZJegAus3DnHIqcKZu2ut7cMrxVTHP2vsayyO5Xz+6ZQHOFpnbUE1GyDFtOix
kqTzKp52Nd/gdA+AeokWntMicvHxbSAavcFxIJPbABZQ2WFmBtUILKnjguk4FW/m
kCZW+r/p0FDRJBcBWUUYdEc9jR6QLWlJIES80fDvB/bjvSJ7C9M4PJbg/ljWG34U
rDsHSiIGfYLm3oLP0p8OWrwKZclGbV9GCpDEzWsa1nqWhdj6e100qD2jvGBKuHOw
PcbSkvD6zY2jufHyeVW+rofx2MQykG30L1YM0aRgBIQp/Z49bHdyOayHvhQWvDzM
zKhdu7zCJ37q2jl2vDBqtizZECQ+FOuTFGE0v4NRfenpdGdg3ZDYHqO7PHgI2/KB
tJTtcRE/MZI4c31vnXx+z5eHZ7bfzJz13Df/l6mqpF3Fomd9hxGfcMkUVwIwIldu
QL37HRV2QX3oxZe0OofU3lS4b+uVAuHlg8Cq9u9uXPqaJwLy5P3f/I+8Zk2pz32Q
oqYmL2wPYHgQ0YUzLmHYT7ankSd7zajUkbDnX5s1e7kltwwvE3iBdLBlVKIOpaIt
IgS+HF5z4mBvR/XUHeIbK5vsFkGRPj4r+FfQEGWGp9akt5W9FmUDsbRbfntVBUU9
/M4Sqw4Br+rgwTv86XDAyC7MDKPSzQH+XYq/QA2SheEikMCwecuvQHHs+HBwyEXf
1xwpjdC4rjlxd0UFeMaHC4prDYd9KJgiTNx5vkmHeNfsLH1Y9IZSmdjce3CNBa0V
9NMV95ZuizvlASS9l4e4Ctvgh2EvZLBiIXPER0Hz1q7ha4YFj4OJ/DIbDzPJsTwK
Mm2XUSRtcG6iywlLdR+vRUMG1burOgl6WzrZWn4JOv/vaaBdikRTW4JAIgVM9R4u
s+UaKRgUeNjJS67heum3HNfOwlpb9Ppgik6/MlphfdONu99ghiGI7hdlUNdVLxLc
MKeUw7ylu84krZoIo4WFQS38+Diq/7ntFSSKAkYU7/PlTKr+J4OMKmx2Xhkpllmf
dnvTaGMn8w7Epvpb1/2YLfoU4XYWbLoT0zDoIWydcD8v38KuqrPz2YNXNndaM2or
URSRpVBLwJdLaklYD6Y4qIu4qNPPzo1sAxu4QDf9nmBwh+d0GbfdUI/LuUqn9ct9
6KvwbO0mmZrBlfFnaZa52wUlTYyyOhwPfUq5z37R74zUc14LWu4CzUNvVLgnZeFC
MYTJXOsLGL2fXVKei3O+cz81fDvaLsJMjB3D6tXYW5Qrelh20kOHC3be3wMcM8Z/
iAllakxIyHZFS0PouuUZYJX1arJI6yEttxkPkplioz3NaTzL9V8Qgxx4ZDONE+NA
yIzKUedgAeszW4Kk3AOQg9rh6C5PVm+oLy4iqXB67uwChVVTCKiqqeY6LrGdqMw1
sEruNsYh6oqBCzkihZNVUR5GJqxbsj09tos8HX9GEi/uxmRIwUhSn2FTsj35HHCL
C2zGEkHWH9uGBhIrHdD0FYzJ6AYyTBQbcRDaYJK+OgLGepWzhjCWVK9S5bhPWc9V
ilYWZ1hD2BYcavO1mLY3DPkw3wezzaxuCuAwcGhGLNDP3ENEQIKCgzM2LeIxt+Hs
g75L5x42lU3gJT8MU2bHRN5DfqiUjsPu/BNa5v2fDOKe2FsqtOm2UQ1anDmXULZV
mfKH0QWU8+1IxNms2NHsuSlKYMf7cr2m8bJNl6hEKa4PawNqGyGJ8YnyU+oooaxn
XjiS+w/IZoAsNrSWlkLN0N1Gsgi1Oh2vqM5Zj/bPxDYsrAp1r5WK/AvOw9iJlFzv
7Rrrx0pPCh26I2rksNyMIL7PFaBbPRjOUbzHkeadRLI0J9G/bljF8gVFJ+9KBkk2
Nwd1urGBW7Qik/G7WLY+Mu2QR0WD5GUDNDNwwcGvVwhrF3IJIt2V6RtA6e4PskQz
VhhNNiXln8DDLPJgOxM6pL9C3HnuNEe/s0K7GygjVtadv3q+xUewXKizl5QtQPte
K8rR6GvpvknkegaMTuwDOT/KPnqFz4BbjjQ5666c5zrlB6V0LscsaLTCr9PlyC3G
gMuMvd1mxrQxnGitZXfW9CXzatOjBIulxFe4Mpon6uBH8J1lgK61MgNr6KB391Dt
jmOfWDFh7v2/sbS6K0KzRVoFKw7/tbGH3fpKL6/2JVSCMYGTnTNQN4IYRdeIS0Gr
pyJLv77bIOVHaY7q1J4K49uCCaFKjTqSikdZDCD2s3BYnuOgAq+htvC2mHja3Kqv
nuFM7gtSWxka2KWGgSD9BXlJ48XaMnY/t4UX1RKGRuk9VMhas1WTIo0MsmCTcdE7
KV9K+7MwKWyp1cugMeOxhKj1Lm73RDTV7Auw2ql/qqYTZGM3fcp5O58qKt4aWhps
jEYO8HgVqlrzsT2UUkO2/srQ6UcN8qZZFC09zsW8Lh6EVV2KHEq9WR9XjEa+eSCT
vwXPo8FLq4YBcF8kk7N0dSRZ/UtDQoTs+aj8scHZfx5LeySlh6d1koH9afRhjzdX
CFfgKdsPgfiMxTwWFMAYCvmpl42Jwpo1xZujOU+CT8CkN3PShB0aUjgp4+TFy/o3
MdHCiq15H+m4KFC7Q49YW02iW7W1CWefdiJKcM8EO5uauPiez6J2+NCSAt7j4CzS
u2ztZW7isTUN66NyuR0c+ZMCcXslBLyXl3abANYzoGyeDUoSR7TOt6vUiG329BVr
oWXrJJATic/aIsMJmb/q5Db0BDVgyTtrbaaBKcocNprIGm32VD17ejkKIlK0AY47
/P46OpWcwU2TBaKRNa63068bKiRg7CHT9C4IRWhAuwcR1TVWizw5WGL18EkMDw54
Y9UzIbsnVy69bI8q+PKbTBpeznNSPULxRwvDzFy28ASnN3Cy/8ABSX7LifEnySUU
ggGYUUm0UO1LTiiAjmLilab9KszEoFURfx+kkZhoq1LU04Dh93YcUp7ZZSoXwxhh
JyBQmCf2Wba+ttgqeGAUWvQCI61fwBirtGIFN80FeJExZ1mNd7KxiZXgyCx4QPF0
UAY4arolWVkPFWU0oecWtP+2H6sPHiQAVkgqXYR+7gss7cdWMJXZRwc8z6vAqdYm
+P92nzx+SucBayuY+FxZbfkvCwpQ2WPHi0+a9+Wp1Gj7hEmE9tpaOe3f2KijmJeQ
DwAUBRf0R2Usz7yfw5YtKS9hXD3X46bKqaS1si6ZrjrgWdE/mY2CxxPKO2vFKJHa
2kNf9YlNMXDb78KhV1ufPGgIYyc7zuTaz0R4UHQUloG8Y5AOVtZbMQenZDUNrcuh
V1c6zwf8y869Czw04G0NHw/YqjYmahZqKXPyKbuvtAPfLtAcefcgOH0ZOwL/qSFL
9aM1/tRavWRDrItn3js/ri9mJ9ROVRFlmjKKa/apF0eyv60+s7rojtj7fAX/eZBI
6TO8KiWl1g3UDqkvGEtRLwtVRllTwk9ZFT3m88JDw6rzNzChlKKdPInQm8Ph+DEW
i7kD4k3VfN6fpKhKCfkOwdx5AJdVK8kquZUfpCU4jcUEZ5Md3eeMtsanOvLeOy8f
+KfhbRUHNvb0jTYsKfr23ots79pePIG/WwRnQqJtJX8RuKX1U+E0+1N7IfxAwH+C
S7iEQuQy4N3M7tWQQAeBq09KYf/gDI5avFynVYLRiz1/viiRN+runO06ywtdoh4n
GP4TOsinV0aUdmusAfDpHuIyt+oW8nb7yHeu+XE6DatRjVP0xk+OLRafYzK7xAWj
dqz9NxgpBwvWYZYYrhTWOkOhu0n2thq9WBzbtpQ5VxypoVFJ/QXpS7aIqRM2SlwU
vtDnAcG2Cc4twPQBI7iZN8nmsshFO3EZYcPOHSASsMihiiAurzFMLrFbsxlSYO11
mCIZYJWc/u/ntnVGkXIvAkXv2cJmxf5WYZgSZYX+DIr7fQ6vadBySitEzHTYGpew
cxACJG+QxuhDCNfoLjMVt3tVqaQIjGEppFy2H4TQ/VT7Z3azMz2lOfbaNTIw1mXf
yuMKVgErZDq2sCcYhaqv3FIxyiIskYOGudDShQM/f5FNRv/WC8geQ5fpK+u9gp6p
iMsxC0DY4s1gsWT6vMzf4EtS0tAz9k/gir3tgfxvnSimI8C9zq+lFxqndPlBNLNR
a/eUF8cJztQ5B8fuP+fL+Qdn/N6AiFVVfYBDa/EAqZlLzcoCLcV+xaargusPomk9
pDoTRTqN0ka6J5qVLkbjeOi0tPMyEYE4CB71BOlQzKB7Lu8LZtTQ/97bNziIfGnp
DFahDDLz97ja/5SNWx6FWei+iEp3li1fX7fMNqeCBAxKtZYKjcNf1KNNLgdqa1YO
u2dmRGYSaGtCf1mL0ojACdnX7mJNHGqR6Y33aYwR4OsyuS+Jz+sAgPfF0Ap0ctav
TZuW2EUzi66x9W3pZ01PzuQZITNQWiS/A3q7jlBfhMQpg4ij1Lju6SZjYzwCY0q6
yd4c1s1Tb23wR9fzskGQBxuL4K3V7xomb4U/G+FKd7G6Yd80wnTR48zxcLsrCfpe
R9M6wgJ/cckr0GjU4ARuP47ucgkhc3glC0m2E1FZh/eIswY6Aj8xds3Lg0bq3zhh
NSLXdWjlta0vSQDCZWf0QdK9+kMy7wPIzDFnMo8xCjmVIYZvmNoFK4C8mHhqv6Gs
lT0IiyqpQnd6wN/L2ZhHkAovMOwvFWzv9q+AK1/sNM4MCXGms6iF14VOkGa4kx+m
vMnfZ6CtG+h01ZWt9WNU2xPlwhT6jPeS/Wijy64G7m94s5r57oZcAs/HpDTpBS3h
ncFx7WexVlCVrp2mcV0QsyCyYJJgNtd4/jO1KUM1cxF2G4/F0rWRgaVvNgoXJws/
rIe187CQGco65+gAWSPaR0/TTOkaqzYzzch9dQixwZFw4G8vCToibFsVXlA8gneM
RTcy3YVEYbnETrV5wLUlhl2v5mY2dIjrBaWdtgd23Tgli0NyiULXCQXy54RiIkPZ
B4ni3jvdb+f8ImCqc5TTieMmq9V89KHpQ+VD6Jp7VmFsCLhhXJa3AspNw4LA7Mce
EWyX/XlxhuDZ0jE9PoedWhTisN+I326LixE01QPlD7Ry/5ZgtuPrqcXvyJY+ui1S
qhT8ObRINI3+rTwOppT7GEGdBLC8+ycu/AqSHK7Cn+x0NgD+NOSL1j6F8eDs8LFF
vL8p18n+VEBJMIpONHNRQAg+6p8t3YjqV5IMp/Yhlo7rHPeXA2yvV4CcuVCDmR9o
B/WwaJjgXJ+Mj3UHVjS2oe53W5sn0yDPySYIAxd6Pi1YEgdp6vrqpiFt+rHuh6ss
LB5+yRvEuVa3wRxKcKqejrKOhIImBk81tIJrz2V/SbBb0X+cek+JBeVDyHHHiZGv
BMF/Ok6P6+z+4eU5pp4Y/81bcZRDYQ+3C/kYNK0vWsfGqHLvTcy3/AREUtYzrw0O
2LIPxOwNZbuzgJ1c1oh26mbY6rADeMXqbnHEVbYMF0Kfbg3O8JlsjheYJgTGTR4E
rMinc+XuBL2iti1MPtQdDLIQaCAldFkAN3sHH0PYzY9nOkxTUOQR6yUBcY5QJ9H1
UVSJ2ZZVeluDj1YqGM/vsYevKcX3fpNtFi6kYlzC+vWVIzdcM0bWpEv9qHvUgUXO
6nIJBCqdzI/lE957s7vVYGX5IFu3YbW6a5m+Oa+AE61iGadFGh/K+5fbHvWVVU+E
8tTnmMtbX6NpdxEEthd4rTwkXrqSXAngN3Tqzy7hNBI7vuTxR8S4u6ut9AN5gLKo
uIjE0Tumg473hz0xvEL3R9lz1HEH0GBndy3fXB7bmkeD/MxGReCPJI429sdkgWMx
`protect END_PROTECTED
