`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H0O8EOcGPEEsnNaupnsag4mZNZX1G+WTqm6t+kj5Qcpz1FqAg+/VMqZ6UBQej22z
7dllhKp2xEojy9lkp951YN/EAJrnj4wh3CXUPN+vXh2I59QIcN8g6D/fDpqzLhTg
EaXqZBf/vKkb4ezIxiNAY6VqBDpehuE4IHBY60QEIdh3hEELJwI4oIsbNzqd/aE3
T7KJax2tnLsJoheXJJ2T02IQGrUz8SycIkn7gZFUNmbJ0L9fiMsnAvUGHygzl4Eo
tOyCmPG0dH0jzJPDy/EFXSU+9khGoTSn1F1ofGjGSlk6QOoiie4O+e4UXjFh4JwT
Yziwv6ZX/CYyHzj0o+9nqZYClaByLRpSyqXU064OyaLeskPnlN9/Va+Un1zCLByh
s6X45AgljSTXvjuWx1uLmv5M8q6URJFA6RbQb+dt0U1N+YLna+pKJ/DkRhFMGeQQ
ZZO+qapeMtvCKhnkwy+gRtglyn+pNBEbKcSSs//j8sjH5Ztjv0+eQ/i/rzTuuaU0
qZ5zZf2e4TRwGXEX9QzFv1b5cpKKTD6TZCOkv7SJ3GSW5aL0xMOMv81WLWByuczY
D0xyC4X0s4+sXUnvPP6yfmr/XByqAOAMs8xm1BwcO+Ck/iPqqcL/GmIv96P6LmCJ
vqAmLVSsKpbVPkztDDvuZwhLONKp/xM0QTzCvu7OkmZvLiQAzkLbg99X/V/DHdWr
iFJ5WCK9nXDycfOW3bIKn1g64rwDsRNJnJBgKQpLGGutrO50vuQ69EN5lL6mst7Y
BB3EzB5d7RsbrvcEfMvDyOl6ZIil9AWvL9f/2q3J7zgZszMApnCf1sS/7ebU+kK4
rvjDULsEUzRTTlVR7rhNfo33ds2eTJSxQ7gVQ8NK5EJYzU2ljVIBDH3j/LkVRkao
ourN4Sq/s+PiiP/3mN5V6SXNnTxCpeT9GFPUIT+BVEERnIlZFg8WUmQDVkBiqj78
5JIRvsjs4y/+qmAXFTNZpv5GL7l4hQd/Z8p/CjfI6tyD6bPqviWwgJd1F4l/ETBO
aza9yxo1g6nvbX+83xxkjq5yDOaJGi6dKP7FsQCkwv/kuobJ5zGEhDJ4W5wS/KPI
XvKJgNJdtl3SxQYA1nfrAIo2FIg6G7eAX8pql6Yy5+WFId8sVBB6lCpeuKPQtErw
TLt9WjHev4KhfsCizBCMTCGN5+PEa53I/X+Qf/VQ0KksxjBm/NFSRmiQ3OZjErF4
4bELDiUwwqDR5ooKlDf9QJBtbN2gBIUVOX92T7s35wtyQMasVN4N2zZZfBw4I5bJ
HgaBOFw1MQjqVjkKir2nqLgbhoHBbItSp8mvCOJkE0Ehq+bptDPps+SF4JWztn9p
v/2u57TbK8Pg7fzgmCxzsBVZYUnksna3eXlC4VDeRYASv/qG8XAlmAQ5Gn0StlzM
3BoheALbkE4S+RoVneU7/WQKhsbLHczzEWIVZSzJFxG5qbBHqG34DtKRjg4urCxx
ZuPyBdFGs7cY/oBOuULuZrdukvaTJKP6cVyGZLrJTMyqxz+WvInRy4p2zrqT8bGA
XyojHZY4lqTiV6q7BS4PWuNr6mQluJ/6hOvjjB7OH8oPv9e/JLpfuYO84birslUQ
4wpdIYkKYS/Trs10UlBVOzeIzrVUJTVnizYHajqlKYM5a+3e8t6OLOFPKZNj6VHy
LMlwnXkOT5TEq5rXCSHY2rcThq5tm4qz2oEpakANRdySxb4tN3TeOfSE/OJKifH+
7KjifC8w63xMqd0fRoIT7eLAh89q8efrQ3EY4Gk6zuuns25trUZm13n9+OSdgRBH
oHXslmUP8wkP1/fpclD9uipadCrZ0Q7etmlqjkWoQVGmGgvapNBVu6fKZAmakV+1
a8qzGzm+KvIhST3qAHntC9QjmoB7R9gzmu+JF0Zu73s3uepGUPBjanBnAyxx17rb
ccRPcT0DW+CYNAlJKsjEcQ==
`protect END_PROTECTED
