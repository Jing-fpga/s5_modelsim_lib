`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F4I/PNt0DNYsnm6a0BZVbwwSMYHcAhwz7hhper+eKsOfkbxCTcjm+1B6IAOiOiFx
bg2m7S3cTHMN49/GMhnVtlLv9m7+3ySto5iE+HhcJXaafDIRkXoT7bS8GgSWcabq
W5YVeT87jZFo3t5XV2Rx+Kv3JhqC2c5DZUX4D+wrzleCtOA8C3fUkqOKkcwy8ZMd
sSxEL8I+pbgduXwpKC0Fpi7GAXofe4BL/Ig6bYROH/rMiq6w9nihyegrktL8OwmA
ChZzXk2c10NOL/RBPUEMPOX03K0Y3hxRoHl/AxXnrGqlJMCYrhnai0RWAqJbc1Sj
CT+fM0M0FpmyWaiMAbPN4vPlso+XLXncrcJUDvzN2hIqakf/puifEeO5k0wrjpDy
qdNx7rogKzgNpf+Cag+qbkVr857BLKW73q9ZGZBkDYSFfP7OFoxQ6XlFxc11gnp5
aU9RTTEvMB32AxwkUU+gwOSxTeF4XO4HOlS3lkcZdSyoZYkze2UC+NpT0iNVtiJ0
h6DLin25MT+8ge5qA+j6JBf0DtcBjjdyFDPfylO5d26l46d+oLjNkvezW6Ham+l4
IifFyXZOg/zNbPUk4v+TL479Enkwaewq9rkl2tGVYN05BFo6oZj0/3X8uZq6MzoT
U/ySTgfafTM8uAzj2bKxK3Vywf+MZ5TAdsvBJLiUSADxkZhsNyTn90oNhxpECDAU
PccUJDAOn79EzLQvMJgvGrnExSuFxQk2tLfsvgPU0Lw+1fvPK5UveGLR35XsJCiw
zLBgt/TJU2jsznKz0TxSe4X4kf2kMP3gEZBttFV2i3uPBQtnPb9Utdxwkm8H9Kq+
BNAum5yFg30m+3HYTS93dwRir59yORyWaMkM2M7TCj3BN8JcXfh49ac1AklUtFRG
sLL72QYEgVMsMHuKsBTJpRSWrCVXiGWOc7tEs36UQLMk9ls89fHz3ZbMXD0yjpdD
DcYcJX/hc/slbcmFb0BOdjsijC/qSb0O2SznujUzItM3SaUQptrTV9M3LopiSVrV
jCDwxRe/FHtgnB/u5/LQgxCDX8qK4McSBL0rSAuK+fOjoZ9N3cXJf+OEdCb1mmwO
oq+o6NhgHtoeAK/CUMkQyfoFs/NZhIDx8hh+2iLTIJ/Z5mEfaePqDJlCNbYaIFkz
IS5L9cqt+NNrdvaSHGvyaTz00RtEL91JKmz6AgJy7M60us2YAkCNRxAFel8dqyEp
GfYgFTkGcrGW2lJYikAqZE6uArAZSD1kc+oO6/C9l1wjg/4CMBtosOOSBLxhzCma
8tULuYMJyxIL8J/1LRXdAeuCQjVxECk2KouprgN0/xnUKvAnXfKPB1atTc9SNP3e
aUoa+hZ5avDoA1QzG6o5/yECjSk6j4JdyAy/8TrUss11PShxwxyEWGuHR3nZ/yKP
9rgriDYmPk/hjm6ez9ilSGnk7XpLrlmAh257LxE/gH+nYYqhB3IccYHqrHv9qsuN
H8D8lWERxT/uWMd6Lr3TzeEcRB7KQRI+REf5tZ8phavP3oyMK4cHq+gpILsw2xxe
ovfOKhxxTPZpFCfFhZRjXydbkG4dM4Cg9YvLrKC6P+eRpgIu8JHM5bBoTMWUUEG6
8qCqNqabhmzEY6/fDrzZyc6nusTZrKDxwcEmcARN6RXqy5TDDZECQ+gURGffktRR
4fv8YEhwizDksKv5K51BeN9438ou32+bDM8JJCVxv6+JyxkzKvDNur/vUqoU5Zd7
mEoq2aRlxw1qjonFWOH4u7wUuQTi5YIsxsLjctNSq9r1LaETPY5jinUq7vGcjPen
0DudZUS5eiRcmu/NYZtONIF9mEeS99n4F+8uH/7i4rxCNQ9e7Pl+LKXnrXaebzUh
ruBDhCqhkoJDPysH4WB2OIRebxvh2DV04IzepGTe9+8heqwo0SM4YtgdDTP7o6a6
ksaG5gO8BQSNa701XKqaV83PwReaIa/tK7BijEBImbFLBEnuN8ddSd+j89w7NZJW
dS/Od86GM9OKEWu2bih68MkXFIUCEuHonmLVbwKh8MB8HXl7EhZ0ow+A+oz2c64l
hKVv26q6JGJ+/dEC1fYEf0inbFT0hSj6N1QijGThHEJ1AsoZ41etRdA+LZMCPx48
4DBWICrCOFJH5S9kb71K3Riw11NPNAxMYeyBme9ZUZzMRw4jrElsle5ZXfS36XMt
KDUSFV2rtMGgeZzxSR3+pGoSezlYtT3/xmuHiLlv6WWutBGASEGlESMV+8DiVjkC
+NnNZv7ZjwkW6LPH1vxHM3s23ZRgm65PbLR+bEvL9SK7mM6KJQrYfA47tobzmAnL
4boTTGfSjfxKjzyuiYiqBqfVdCi4klAn2OKBXVkSIpZrm0sP3mcPcd/O6su/9Zee
E6E4wtGsTZMZcEjZYCP5RUYKZWRpHT0N9cx7LiOJyltYPxDduEEy49xKPoZ1Oaw1
bJJWffd8HD2X2YZ/Yl0nPg9rFoknYX8e3vJLChL9BnhZydy+ry1t9ECS8FBqtuhj
L3wO0FPNmMjROLSo2FiswujfRnvrmhmH8wr1hyOqIpjRe1R1waD9TXdYiS9HZ4VR
XD/4ETbOm6MWQ+duVnp29A+GCrGf05XXWIhuYIHs5gXopfpjvUh4N9OyGjKoP5oV
TnkfC+znIH024CYCUt4vd0Bx/NhfLFSr2IxHTgpy2o/XtGCKrxadyf54RGplxB6N
lNHaDP4mcd0bbUu+7EHed4oW2UMqum2/I6SOeyqHJMxV6OhfOQOcjh9YTKM3TL5L
HfLqjFI2NcPc6OQ68C1f+aY/ODqLA+D+xG0fCQNedJmFnGEiwnKapPkJrwBPK/4v
Q/4PkHAFulEA/nP+sfsgUVNyQrpEfXFNIs2ZCgKmyH5PlxczAQ0SsD/YW2mGUdNC
OdXn19+wP1HuKikGpADf2iAb9Kgxg5X+qMFifH9HAZ9m7u9ExZxW33mksVEgnvop
XqY6eRAhA4rjzg4dy/xnCaZEHWX0saGnBHjArjaki++Vir4R9Mwje4QmV46oJzMh
LYdVvb+S1gA3uYUSqdEKg6e1frPGfGdXlOCSQEcZWFv6C7+nTAURJfjyogjR3kkg
B66QzyaYDsRGzKj2Pv5FM6qQfF8/LB+0O2v/KcRyHe2M06ljwhFpwC96kCjd2y8M
YLwsxHcgDMH9xgq1MHZZE8ivLybzqTRPC85MKgdUYWx8kVGKGi2wNKHfuGuMmUKE
xSb7oHep8AAuturUFXEQI7BiSeGGXTA/MQXasFIJ77ZDVlZISjaZVcuXalub68VC
RmbGr9jfXOH8Vi1O2tq+nI8yqQN7UVObpDaJl8SvgaC2tt7UtbxppXJR00XUe1oD
litSUkHkfdG2BroSdsOfr5x12pNXyigRJ00AXOQSG04cvBnAqn8ar7YA8PrCEh1N
hCgXX5eimVGdjjEbFb06+fyQUeIsFyPbd+3expWSkngUl3NRnrKuaCjfGQRG94p9
`protect END_PROTECTED
