`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ptAa+/bp2pOIfW42Pdih+r8z44ulIICler/O/R3qzosOG8HB4QNED8ZFRPijbAAb
iq7rJ0J2zPC4rcC9OR+zT1+MeZ1zlURn1B8cnTMSxxw0F9U4FW5BMY5GSZJGmjCO
iAQZTqamwlwaZAUghDX3av0B0WqC4mNcRukasy5DSONMi5rY06RX7OBWRG6kEywV
uVsxF3gcR/vN/Vu4gjFLKzkKCZnXG/e+oLJe6Bt5cJeTsrEbr75cfK42aMnfOUiH
OntnI2tDf6Dk9QnPgMeLAptvy77qN9t8qRVFyYSXiXLaN2SG2iPs8Vvzvw11PJkT
Ri+NIvVo9H2lj6dS5HfEN1yNzJM1poieKml6tRdgFJ12WWmlrOiYcAbrdkYTNpoX
Tv7SKvcCIMNK/A76i3LC3Vi57oMkIllTTx2ZqKxF8f5Ayqa9LBndPb0HCxQ3MfrR
feEjsAtfGGa7bd3Z/5hci+9UwG/xOOuQq2V1V8gACFRDXNahu6vLDSW+jChJ34VE
dU6PRV+FRyFNC2r3Y+LONlr0VfoT4qovjuoBjaMyPSxnMLrxAHdHw4QR7T4G3tAv
waR+AEXaRyXfVMVdFbZqMxal1gWIGxtfHw7CTag3FpBa8YYvJzF7k3P3FQrmgknw
zrWn4cDAyajMIKskbe+laSL9riK06seAPfGuJEZD7GaYN6BZqq1ZgKYVxH9l5iS9
sDCHrmZyDAU9MzQFIdBIx+FSRmQY57xT8f5Iz7m9rUB7WZ0ghEYWoOz8QjkCBm3k
RMvVcBjS01IY3cO4AGuo6UuUU+HXXre8YS6uJiYvAzOuZHcNmfwyoxVR+lqvnKbe
N3iJ/cRgv1uBAwvjR0fgTK59wg7f5PHeS+otTkWe38j4bAPI2axCB2VPt7Cj1LJw
qjSEPAD4m52rjD5qPllGkyNyepoKCpRJJ84f/+TYf8U7ZCZR0LTyDp6INZO/gOmJ
xJmf/7eMzuyjLfYAKQfDW7yzKXRQyV34AkZ7UpCMEGnKAg8wsQomY8Zdg7oMOKtT
gXGqoCDqBGVpCdcPbiUePRitMqExW7A+MY42fxtUuKEmabPSnpUa/fAAy5iytHkX
c5smjubjv2w2FX7Inhdi0/Qf5SVsE+FwuXeSxhq/QXkdvFZ5GmeTGLcCAdqHE3gW
OvbSM9dJiDl1KmKZZHmDfzW17tQ06rCYu9jSs3iBPcBMxxM9hbjgeoZa/9DNkbtN
zfcOwWGeLeNmDm2vkzxX/noCWCz5lskTt0vBUkOPWDMcMpCkn7DtqXgyjur4ZTUa
djHeVgMtBYXRNjlgFN+DMgn3O8jY+U8+Bu8bocCNr0CdL831uvs8wp395WjPdNTW
7+AY7CuWZhpKrN6jEpLgV9BMsuONUj+WeUFzvjeCxnL3AGW99VDDE7+0irCd03b2
NQ90MbKRDtOuW9pJgRB5vULJvy5LKysIE2e9DU77sHg7nd6YE68o58ihlfTZp3FV
6VQhxzAHDwxhns4og2AzJVGRocw5rjKldMWzag7eGZdw1BJ0bwHlxx/QpMRdGPYL
fPhVC8b0Q4+N7fX9RKCqX3yrhhyMEjK0wWJ7h8Y+ZZ+6mQSlz1ag/L9aLQXI6CoL
XACWUUhH60YscZ5hgECwfaiMB0U7PIIRux89Mc4Vzq/mhAUC8M/Pvlx50HeGmEpy
dsoI0JXb/c8gHr/tP9H1BAKWtLV8AM4YWOH4IDmTefWEyHUt9GEYrzakUjS2CIpp
naSJd0wajJQVlNGOE3Qer2/nPuF4s4Y1rPrDPV6gdNosE64jkqjCCMQkZr4Gp1t2
nCKRihAsD7egSyMhhplcrWb1AjdO9jx8//N04GkAftFGFJQrHf/t2Et9Vi9+PHWx
KM34iCAP+SeFH67zeG18B6q5YElYWly0TkJMhC7IrievnIBKzbXzW3PtB6jq/Gjl
OzcSoke6kFHIv6bG0joL4kFC6G1XhBI9jfPLoNjB7ELTrtboFo3xPOdDDPz+MrA1
vVIYhZuxJlg8KW9bxon5gPTjyENkTgP8NFa9Gz9hCA7JG3G5oBAMH5ygGZ4dpG4R
qAFz8hGUc3JrVgjvfxhKY5Suoopm4WPyBEaxYiwjybA2XLLj7gfyjp3JG282Faqr
oww1MXufgdBOVUT2mDGUVn0CkKYS0c8gMZtTinJwM2cUexyGBZNV+QlqlI+HCnP2
0ARWcIIA5MiuWzRtqg3LoTMR9dYU/LIuNulqmdQxiG4i1U6jUKzfA0uPbHaxtx4S
NsRM4o5hCPOq3gVXb9fW6bnhjfzwxDtXZQvxdcfZv8PxX093AL26/jStH9pcOluo
3tCuyzKReLJjp1EeZFDCMXCyasyPQeWh8Mkyihx7pVz8VfQk9OIiupuTEHcOj5te
c5aztrbBNwrr9L9aYHFemTgin4I9YnDZ3iqbdDAbWSVnNn3Z1HYHbw4Nd8QFcd3r
4kvKZSfPuGwhakYOnWgHNQfQ9hF/F+SMePCm4TR0VdOeBpKdeTCdFKFbUoYO4FOc
tGQZNmhXu1y3DWXR+QTvQq0sLPRs3F5JtVyY7ziWvcq3e5LPstkEqYMuuouSjvR8
mg5oUqPU4aG+TwSBEDHC5f3hTKdM9aaoXzb/ikU3W8vu3Qffm2JTNx3k0OoV3zvj
V8zcfuVOksiyQBj5YF7l0URYmzmARoq8IVJn1aYVXSxuyXyw+XFI+MgW8k6nGOMJ
`protect END_PROTECTED
