`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6UBmIYZVnLG410+XQk7IaeCHBlDF3BGlHKSWc8R9PgZRbPdstxagBI1UsW4es2s7
gX91ut8avKNAlb57qKQaizVmo6lRAvHLf02W/HyV0fycuBlIMZrsSZnB+fJ1Vr/a
VGe/aBMJW3D1RtiDBxOtN3O8mOVH2fQXwljhg79lxCoynQ4vPHGn6kja9t+18fL1
cJHfZpO6iuaATiMC6ThPUcB6LXJUala7d3jgPoPrVlxyoGqVJWINq+YY2oZCojLp
dtYBv3x5uX4d8LJ2IKLKVzPU++Ygvv/6DDRnfemUTyU3BCnl4J6WGtrLeAbwkfZa
8Kyra0y3cUyrNzQ+7mYIBY39koXTkOmDL9g/Z/Eh0g398HJJASSNeNGeu+TYiCAu
G3B1X/mpT/3autQkzSjCeaseu1lIzj8lSQAdUmtClihzJVQ47Cy880TL8ywVkgLW
oWP5XWdDNEXNZse2xw1Lys0YodSI2NSXgD+q4m0VwsoN2yKGJwMkAcVkNHk8W6Ud
QeXcQBH9ScXIhthl0xgdW2FNsW4waUuBtiBu9PJAzYHfI6phRt5ml9FkvMq8nnhG
502PhKwfvlM1yN7cNPc5SyDURF+kXb7AJalAt0eN4JaqKWVOkq7352zjemcqBFRo
hvyO9ibM9nJswiB97lyxZVlxiU60WA++27uvhTAya4UYyL73z87rdWrm8/ezo+ko
C8dihCn9VYejBxPddpNCFs8LHPhWUVotobEfVPWeajFgzQEx3tvNKmk0Hkd2EKFB
SRUOHCEzNFASMMRemS3h8BJdPsmfp7wYI6yHhLGl/eHsXIMqQU0Oc+JsHdzACyfO
YibhaQG5LRJkLzwYAqK8gpvLk8888Ip0i2MvV2ZsPL4rXeurlWEKpZWyKw3Ky5Yu
nq/4KM2mdInD2DmKSXuzl11YZ4yyQpl6719SfXZX5zIK+SYH1QNJdeeH6sg/UH0W
/qIrSsbGi5wZBUBp4GHhK41gM1tDFY0S03gj3AuSNcUGsAKj+XEdboxat73kCsSP
9PGRDM07eas304Pdvr6wfbmJCBoCuTO7oOYPRSo/k1FxnOH4oHqyfDht396ZXVqE
KNatgdknI5My0xIkBdSnWRrtfMdOdFH/dS8tHm7OuvGq4fHhXUN9W+bZ7l25FvWS
Zu4bt3V9KT8X+4MJ6wYZDwtSP9R37whurn5mF0buyLvNqngtQlUFfL8Ybcacql7s
Im8HE8Jn1ZCit/QMrKoELPFGLZg2gw0WKL99SEVgZiXbfXmASSf/V15/T+pnu6LC
+XXovtNR4xMK0Q2MQE9m3mRFaFZrAZKGpe4U/oM/nF3r1Kcoa5syPJ8/jml0pQMy
uWgcpUzANDCoL1vSLjhLNdkGpBeBWBKO75hsfOkTAT6lEyAcUZy8K2ff2I8JTixF
dTeKJPKrEAyreL0N8eG4laU2zU56BniUi43pe7X1/VwZFJhWJaSGQfZV/wTzgZD3
tc4gV4v0eh8TOHUIqDuStzmhQrHpAI0jxCtXs/cPf+ajoP/wpxaY9GZukPWXwJzx
bL7wSN+O9m7/ISUP3tlYRknQVN1rzSBst50+elxyEGtn5J+KUC2rcEOpaupHFpTs
e0vkbp4imSkoRfZNwD3AE3yeTVDI8gFToCMM8oWZUObPuNmD2oCLosWEpNJkAtBl
OwYvq4fpdMQQObyTxcMLOvE/RLA5gY8kCO9BHGuQwDcCcQWKJxBAZaLXzDbitX7N
Du7JnKLewc5Hgq4vDxpglwKFVUgE7fzAyzb5VpGHW0Z7fQaaXr8KVVhjaCJpbljy
dg6QvzhWKqkHnjmIrcTW5AbWnbqfkWDL53PGPBKTKN4HAJzBV6f4NYPvUhVO0WzU
S1zdUOXG3RsDlb3rSgvBelyWC/RMIidkFGct3SFMvgo9AfpvtA2qVxNagAYLjqoH
TgyMPmzfCb0c5Gq2nJpKtE0e5/URTnZWxn4nS+Z/e7WPLz4VQiwUZnR8oF+zUrmN
60Q6Un+onwrEvR3SJcibMSKgiVTGVhAXwT7F5Zg7lvriW3pXn0ybg61770rZM9Q5
/InW9WNVSBy/PERGZBOCyt8sCBj6zrGyq05hLjKItluHLaQtYPaGHJ8E1YKagH/v
AZJSEs5fX7mnNKMEvP1S8SdJVUwaacQHkQfqhUejPSjFFnFOARZ1yOdaP4e69RNC
n9uNO22mBVIuCF4EtW32eIOlyvw90biCSSEU9UnR32Nh+Q9Ik/RzbrwCks/DXKTR
9zdpWheQYCjCp7MzfjAjlvtpjGronCRuxBm8vGdSHpkmmxRU3x6WMn7Duq/s4SfD
KnvlDQTwHA+ArXff7X2t+J1K12UpCqsQltXlfU9XsxDbwXpHfHkuDH2EJitVh5Pn
zwayxPjCh6PmZcpIZCFdcnf+xDMiBo0bsd2BTQE14ZsZ22eY8xzQHnvM0hWs+jxr
0ZCLe08LCSaFxfN/b7HlxncHW6LlZCzRe+rAbQsHbas=
`protect END_PROTECTED
