`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
79Y45Ay1uVLPgLYy/T15VUNoCSraiqA4x3/pr3CCoRRVW4aUswAcKSnNPCBIVsoe
bSGatDC1v8cDb5fXPQOpOXKxs1ggb/r3C9DArV8YsNmxao74UGJPSXaEUOkjBt7U
+rGbAt0AfbV7sVTjCryaloF62Kqe9lwDhI82vt+T34Ms0k2R89tZN5kJZbhc+Dg1
lg1nOIGHUjRrjs7lExqm1KR3pEivN4EDda6fnXuDXi8OwZ+lCfPMXoGT4JG/kHv6
oCcLIz/omGiAeP7hg2KwpQ/ZZpDRFFJPcoSA8tWPsD+aH8JgHVZqZ1jHabmhXoIN
0/hEFtkW35znA9SM9EF/xRYXFzp9kLkxwKyjcyHstE1pAGtrn6OMG2WBjUvlSwKK
Yq3CYIFHZ/WWlDCSfvWNx9aaxbddtlZH0A0n4ov0DrC27z5pwudWvXqE1xA0V+Me
3tnl8WL+45PBJc9MBUQxP/s0tDy1Eln1ISPYZLj1PaCGedaCb+Mx6IjnNmKFlvKy
j8dD7FruBKbN78hoHSgeWxUs2Vi2XJp5pvIaKBZOZZwNAPKzzeJ/4hkWdKoF86Ft
9qyK12lqcWpn688mDMDFDBk1ehthBpoMU971EhteCaVq678wR9b252CGo2eUBC2F
GRzStpz1ap2/saKnvL076gJxu9g2BGCp1sdt67lD7Fx/HPr6A82lCy/0LPuCz0hP
W2GgOYSAcWRIMLtL1pwrXV0pJuz/a5RZDnGhQ6PTwPLURowX8qwvUUmIsu/26VXI
R6TmmCVNwMS5WtHgaxQRUy+Jgj5D18xgZf6wo9oiVkdCSppijA2yCU6Qfcd2gwv3
VxK5NIm5F2SZ//uNFTTTISuJI0fvoOmKSa7whqtZrKfrIwnDcS5QMwULAT/uJHA1
bqESDl/KO2diKYwfh+9GWyPhhfTXdwJ4iTODyOWgxCkLOD9Xrbr2bljLT7tq0rwV
uKiejD8X4DmKufNis2Udl54i+jpC41X8JmsAL7ZOqLZq3T6lzP1Lzj+hka8tu79h
hqo5AKASsWRGk7zIKJz253bXBXvE3FTjYmmbnLMnPJdpiiVVhFwtmItaEVEG0XWx
6G6if6ieIwsrwHhGOV4RLngJCKsBh/CIlnstLx0lDNZdH6ljf5av+EElfw46ywgM
sU7gzUdObpTBuVPmNf68l6TBc+iLOHAQyGJb8tF33c90Me15+PfPMCafJsbeKh2K
GCpUYL7IEcZR/j3bm69c45xPxU2WOG5265lrFsee4wYxD3AJq4+Q63a4+4aTYY2m
kpZB807MdEvukDNd5oqzjAS/M9OPdiZYOHvShfSedOj/se1z768DJ2njlgUPEr+K
ngJ2pMv2/7GkUMeDOBIkjKdWhiHC5YXr5M0farhCP2ijZ7uq8mLFZPGOY2bSriwE
YfDeMTrgKLVvBkJBtZh64kmD1gfBT1WnNA67aHbWUnKbB509gPguJp4JARJrgQXh
QXyaHNWe9C1nbCdELAuhnXKyq8RUMok1b41XvNvjnTZfmv2payFTwebIHw6w1/fi
XXo26QI+HCp6FiCpA/++dqLhMmxi3KSHASr13pJfEYkYGN/z84umKAMxGB5lhuDL
3MJPLeWD7AIdtGrO9i726nBYb3skg2u4iYStPnzC0m2h/mnSQB4ml+bF4lmYCXvR
cca/ap1QvMHOz/gbnPX+Z3wjtGIiKyjV7kWz7lMIC41Y4AkMiaudjaRM7NQXK22z
`protect END_PROTECTED
