`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KVFVVfOmF6hU5zzLh3xoExwIOinq+Z6ZdzkWCWbGq+gC6OjJQKGlEthlJXLEyvCg
YMtPtGFdiPaPjtHKl9uG77Y1SIKR/2c1cUpye5XGvnxxsyKmlXBkTrTm7u+p2lhz
99o7KgZ3N/nzHwCM7FDfFpius3jRR0jZH+0KKfBHrU+wcEHFY0vFP3aSy8O7p3sE
xTzBWHkDxMDziwA8mFSk9xwfkpBFd9eA9uc6Y05YGcIT6+P2qRm2TpopsIzEeMKL
9dcLerkRDW5PeP/UmgtIXFeUHspArYrRyrjQ257MtsrUENsjL3JdiBvK9C9CVJcV
aC+N6xErmjrrubhvmrPIdaBSa987A868IWCS3yFtttiOYQo+Yzd12nFg9Hq6Cz0Y
7szXFQ7cbY5k4u/Z9Tpt0M4ZQMeYLfDUQy07wN60U5AyxNC9uHsCQ1vWnaEwk8su
sugdJNLUaIYW7JBY+JMur+dzsOXUjbodBFGbr29iVS0A9Qk6oceaaqv4B8yamWuM
D3W3C0Fmxts/i3rJK6V2ShlCxEsATd2W8zXM1hRMTO82Kgcn2/nn+QwpObhbUDZ8
5iABJvoNvxmyI+LWRxcXBWChJSoteQxMe3hcCs47epkAuEtDaZnz9Eorh1LIz8tO
xp0ViPVUXuzguVuOh6NdHqxHmgScXiAEwN8wv+nrhFX2wUxq+BbferexsQjy3Obt
iyWU+ZUaYsJ6TVwOflqwA2BsDxaM28P51OjbiIt3D1WZXNMqHD/sFHYUdayJ+CGU
vjrQ2lXAafLaUb1SankGfnaELHrN6iqh5Jj76QPfWJ2VF0VwdXh49OgMMaMX7NFs
dyF/2EmsIk8DbhtQ8LR6JB/kA+1rwWiqaUIWlJa0g7QpJ+OOr+fIPT8PnlbW5K6N
Rso1I/MTBgK0WX1ekXQ/lTLN3dUBPTCIF4wYhp7HvQRAYv8ZGsMFGFYB+YS+2gEN
B6GjejqlKX6+DJ/husoQ4HZUIqO5+sJRtWBcW3uaQQeKhhtzI3WGSrPcCgomEDsK
n+9dQ3hyFv+VzqfwPGRnrC3p85h+E6zPPinvWMINLwjOatinyU0svfxys8NadiSS
RPrjUuummXCtZreNWhuqV+uoC2qxfSsSErKeEmnPyTM=
`protect END_PROTECTED
