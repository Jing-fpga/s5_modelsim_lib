`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xRkOhgRZ2VFT5wsx896zBrIwL02Pww+I5pwJX7/shv8zpiLQauOV+TIDEdMXpjiE
dRsML1roj/Vz3R53lFF9EjONegI4Hc/eI0avo2zSg5hS3xMrArd/1KTymgYuwyEG
cPwT3fYwlN8JXh0dWZoh6m714WObB1Xl05iWqtJgY197BMpizb/Pw59nN4hp9uH6
uwJy7jkcvhYw8jJHPKoaFexY/DaIg30b1yRQFCQ4NBCfOmA64mZOHBe3FldM9fn4
S2yOLQCh/vv1+wc9QfLHK3r3hjk1dqdtRR6zlS88hw8D99L+10TFhTXUi005pEyX
uGoFx6FBuhA8zQS/t+os3/nGRrDYk5s9Ls2esslYK62yakSb3LoBM6eMGP2ngBOd
cLu+TEuD+SAGCAHmqMIeyRTA8euxSPUFksEeLwyyTFt4kj76o8xRZW3/MTaKSIxu
7eNE9XtZJVjwOhV01rjam53HfVgJU75VbqbimMpiAgzkoKPsmW7u95k9zyWqHRTJ
7BNVaE6yXG6c9rJJTU9Pdgc6coVNs1qg1coqDVRweio+wAXf+gYF9ddP1ud28hwA
rmCBfB0zs9lJ7P8RMpxVJNDxwg9NhUqDH1+NZZFd+tB3sZUbrLWgmCVGtCTZG+s3
nxdyrYYQeGvTYXUH4kD7kL7exns/PAV+SfYxNRAkJ/UbzXGHXomoJjD4niIgColf
tHVcKqd+BQUfBEaqBLucWB7e0zCziD/qnnkJLqbYCc1oJi5geDs//hUmv6T/qoSz
7YXDLgPxGpBcVqj7OLv57TKy5rgvZQYMVFZlGGxUnJ724RtMzBrVlEvETENAajJv
YUXKCLcAHHlEU9klcFxh9/elIYN75MVoPqngEX9YrWEeiJIgKdz6hRYmriqum51a
l3z8dKDTjX+laQZn4A7p0CLWms08uZNvJqJ2yQ6T889pw1fyylkb8rZTYYvkINN9
/fHiW9htsdtTLjo/CZuHJSC3ffLLSkQ/A4WshOOYnoTkz8KnYBlJ+Y1zgHyQMD71
rLdNS6obinKa958qTLUxIiUzjWKsiFpuynj/BqS4lqrWUSruwZmOlyDo4Qarn3f9
lDEC5nvWcjEqv3N76RqKp+AxgwIDRlS76+Kx2ZyIJbIlNcwCAh++M19x72VDtJQ8
1kik9vnk4q9qgpteXpOvMEUjqQYa82ALqqtT4jEMYB/zzon2J2v+7AngHwhtNcEf
mgZo8LbhqwazIGwuMOzWHCUGTllBEyC+zwx1bAV0X7c4X0nRfxHwyz5VpmVugrIT
FiEKPleIY6MGXjUzC0Yy2a2GgTTzLxplaBtU21BToK8qJABs/A6XuqC/tK/E3JPE
1eJgZLx9JrUJRFxTzGyftOGvpznPsqDSP6tM+TZYkI1ZhVxig47Fonw9wMqgKYcV
bju2O6WKRVBzSI9lk2w8fBKybDOXv7q4Ef1Y00ejc34vBQ3JYrpYXkYC2XV/oq3R
RsNFOTDX5iYiOuFUOQl/BAB08oML1UOMtU2nquHDtwt7sWMrqTmr5KBlJcoW4TyR
CqE3y1P3gFSVlaxeZaoiPpL7dhBpk1xnsbU09SiWqKA9gQ3rG0PrX1kahD3sIohS
jT5O39zXlDIDt4Opsb3ObVCq4a037V7X6eyPR6GA2rfN4AhejXhbE1zLzTgQoqgo
XGEeJtwysS02c45C2h+d359T9muKGGFw7jzvoyIktI9rJXbCqtoLWlHeHpr9l2iY
1ah7N8D6PGrGtB7i/5+kDYU5WMD3AqOBM4jxLxLDb9TGCsTvVSquZPezm2Ob1X5o
t1FDrbmMoGAqW0dxnYJDeLC94gDrePiLSQalmpUwo/FmClv5flg5fTOT1P+FB0gB
3uFGLhsG7Q/GAHdQ4GZjyPtePZrFdg46OFeUpQ51EEO2pXYs0pGjLaRkI+/HOOYD
B8lgO7SisvZ33s0MUSEQKSZ0FOvRijuu4m8qMgKwdXSowaK/b31c3u7LOwHTYqVz
+8xdeePJLvORKKNyGtK9Xpk837ZnD0KcPouve81Ct+JQl6Sk5ztTxSVQm0j0ezam
QBTQm3TD5u5rnpug37L52W4dfszVf0/YSmF568xaFPmi3rOx6PRzkysuWAdOZg2K
hpereDn4MUB5JiAra/jEL97lpZSSLyxcujAeKV25dkko2GeuuNlbduUm4W0D89JV
0Yscabc1CtqlVFaAza2rPrsmvOEeTPfNd7NCDTZ0g6MC423yhACkQae8gwHT+tHw
qsTOBemxQ1fbyZhv4rrrzecSn8vS4idZfzA195ngYYW7RBpnkOskcFkqhS+YvBbt
a0HXW7DBwi15FQcQo4KAcm95AG4e1ZkfFLJGcLtZc38htKWqq8z5ZTvqVjGmItiv
TbPP6o/XN/rEpqaCYGBnNQQzwiRHa6oI3eewa7pEkZfo3wQofn5uqtn+86oVrtYd
iAvwpYcVLG4MLOH9Hn4GO7Hv1A7vQ/5uSDgLL1GvK4Vif2lA82zulm4TL/O75LJ5
yn+9PlAwsXOPWLjZtqZQOfBqF9UEpFG82YLPjC1A4r9c1+YG04w4czw8Lwv0GwwP
jcv3EVyI21Q4OKelAX7O8uBjWkFX9RNZu6u/vIpdCS2dJEG/RHvh/V7PRv8iXTO8
N3Psj74KOuYUUEkvSz0rV/1pT8sr3nGDA/mdV2ffPYMpJOZH5f9CBd2vA5ak4P8g
61VdqfB6iF509Q+nciriyLlKHuEj42geRyJcF8077TOMkthUKptM2ylQX2gcQT+z
NPOO1nhC0+DAV6fXKz3vX45xLIzhtmmjCHcEPhvW7hIW5Xu/iRi2NLYLW/NlO5c+
FCH5bYd7atsUZvPZ76znJ+uW+AXkV4T2dNLO0rCkIB9/nNhj4XqaeNMc+v467QDM
KkOIaJhdoneQ2NntTATQ3HifHT+XPRMUTzzjVN9oOX+qOL4lDBTMts6plNvoVVfp
HRPTuJq5y73adMbfEkS0yGNbtbscGMVg0eN1Wc5+rTu0Xvq8TE9TmLzTr3pymhOx
t+xp8XAeAk7zj4LApYJj63z8b1M3+L4sWeDKHbBrl5lii6wINsbZdr3xhi293aLj
lWtJFOrajRniXmnGFUNzhip//DQvaefPvzfBKdX8Nbm6LXKpKPQ0VjzHQn9L1lQY
+7bkX0lP877otfYveUhtPS6CI6szLgEpnXEB7fEtUsCpi47ZLkvkO9I4LTYEpSy3
/UI6VX4+5y30Mi4dYnBlbIBnccavc94yjjjCSu7/LQfxaZkbid9Q86E9unOs3qzT
fgFbD4P+9Bqho/ZOEAOQGfUb/3iZEYE+Ol2VU+VN0pO6AAo4/exNJ8BTOLTnL9oG
uB92YA5ks9tuQEolDjNN3AWKl+9T/LPBHSdWtCuUIhOdFPpjRVJ7Dun0y2Q/va8n
t6xJcJgkGsOY9AG+DGWDcKh567JpJ2WvT0kMHqDL2mcVsXIhRB7n0eVAPsAnXxTD
ZaENqMcXdwjMVyIKwe3qG67mOwXQCbfcIXIsn5co+3TYWfYxoJaLYWZEmiVgLrl5
107wF4tk6/f34/pen4YgEobaXHiCrkp8DGV5NSMSGYF6JxZY7CjW86Zot3ae5uxj
h+sVOHAQ9ak7BHUCV+o7M3e6AMP4TVury6fr3N8yQKQFvc0yaD8sZNw4sLt6klLi
0zdsh/lNCFseZN2yYfieZblwCAeTCpXjprMfg6vexyII5WQeKDcEZ7MBqDWZZoEk
rlF2KDZvhg586VYh2WCXIHhgIOH3ecKPqM5qoY8c+bKbIURezbOaCkm6xif0lcxJ
XFrVz+qBItgWfGsYZeTtyymrWdLTTLnybcynwvBukgWZcTJDsCIDL4XcmLWKnaNf
DVCeKE3i2cDc+AU69GWAyTAyLuD/GuAYyvPtVtfwhMqyM/Uu9HRvd+N+KanQTy5o
U3OwxpqirK5YVdv9nq8Gv0R6E4OwdbKC3a8InVWj6sg2AN4aYZwVIBdvJEq3U33f
h8bn5XabU3yOsp6ZQVyxaq+4TJyCQkS9DVs5FNTDO6ZsPQwLxrwJt1L4ncSmilvf
m0UH9krJXkygZx+QyLTVJ8EjG+HGPRw+MgVHmm6kacmLAUxwX+t2XQYuR13ebuTk
X20FR/UK6b2N9RVDF6JJC6fwbUML1JvTRSL1AOGuow21WpquXRfvAAIAjMZAerXF
YJKj/GsFpRrISeQ3lJlVvwCXtLxxrt2GuePWC5y3JXrCWYglxSPOOKwBH3ZSKIsC
BUCocC0e7NYO26W2H7RoTeK6pNasmYNXNicgrNtihynLWbLppXXhIeNj6e4yD9dk
xJWPFqVIUuJJLBQAzA4Tlf0A7hd8eLNL4QVAkmiaTpaIyc7jRQTCFVOpoAoNc6/T
cm1SB4n6vNq19I+3ijzFV29C8Llb9RCPgGE9hJJdnpsGzlwFFpqwzxZU5QDfJEoX
HX31XN867oERKnn04fMWX5/Sxq7dUAVzwEzdCvpcEysL8gEIll+/Iy2jFv/8drJk
IYlQQfPnTDoUMVey/z0uAyFLwgxD0D1BEkxUntXCUw0A9C26A8qeP3O/jmRz92PN
nDJ8icmeNmx5SoPwbvPj5Lk21OMQf6hxhWW0wpfhxuGevhuG80ZzYzDgri24noqK
4sAkbPFla2zLU+GdC7473JVKuqI6siHlTR0I/wx4oP8oWZDGk++2nWueJXuNHSzF
johEUMQ3omxKLeVSumh7Ij+5AyEGWuft54WXs3venMEYWVnOqWxszF22Sazw06G5
dTyCdKG0tWIoNPqU+rnKdMDvGSN4Qe7Tyu+3h+0JjYQKaT/Ob4+7x02Z53wLPiQM
aMW3Ce/lzEJnAG0u+mWRYEMz46Ni6dRip5nYfUBrR/1FiSS3aKTp0pFsrCa0+JyY
D+rw9AVH47wJaInXdk+orRGq4BXYObwagC5ba+N9mt2uWk8Iy5NjzOQyUZMVXDJk
OkluJaGcj9Gju7E21dnBPVNmCl1AfcPhrWLw5YXZQ2IeJmRwJicg1kCxqdtqEfrB
0jCAQOSUq4e5mTzHM5JIRTq31LyklEF1hUuJjATMBIQ+ZKD5LK/xzA9RGSzR8tFH
t+M6rBg22PAHxu9+DJM6MKm/D81nzhxfJk2ce+yLlwmfpA+8l9GUz6SkSvVMetto
XguB1w89BpCot/Z49Zq8Md6J4p17MsNdNIMspEYcDbqqcGd98OQmzVxnfkBMuGCL
Xm7tkrhIyNs/+SAaotWeTeA+kmmzD9d9ImyiVfxUfs7eQ4C8YBk/YUIXu+TG2INk
7+deTz31nk2pPJc9hk0WwSUDmQfwZ7NYItQLcjGAiQxpXx6yyE76vVWJmVBxFqjS
JjD8bfTyGopqzKxPURizTDv0pDEsX+CqXcBM4KEbB0uFy1roZrIQ3lOEfsxgb3HI
+9cB/dTCMULMz9ODK5lDJUOJdgBuKJb84FcF6Y3C9Hql8M0+wUN+VAOlbuRu5rQ6
mkfnnNwxH9rcCbapR5qj7YW6pup3LdUn1vj3dFCMKNNHMKtfEsurwJv7XCC+Cd/s
mfvp59BH+5fxLMfSUl/E86MPU8glvamF0ggmBpIkpPPCHEeyWcTfM3XGtrz+TYIx
00YYUgrMhNe6WUaFfgySCC+XVr2SPZD+Kq6dzCA7h9OH/Lpq4hAW78toLd7A1Obp
BxQRUxFPwJAXTFImN480p5cfU2Y1sBCHSdbLvn5baAkCQSSoiB7TJcSdONqdIMtT
aqKsvQpN6J8o75STY+YTe/W37y74p061nzZlWtRHzUBVPaDpGSgC7z8QJjV7qhBA
tj/uFmWxpd/PMAXMJlbiQUjn1JGk3zDJTU0A8nQYJO1CKfNGlw7rzaJ7Fxgn49XW
J/LTB5zYy3Vr1MYKxxvDEZPlJN3mxLTqKmOKWXYbABCIYL3Zd2NC0NJTG9eLUb46
AvMFchpqAeeXrbTfn1slsZJ/o8nUyIsxr5ArDkybRAB0zg23InurfsPPXTDeHZAW
SOVMd8fNhEmT+sTDXy4y4H8gfbJBfJQX5k0CTVRYeX6+sL7kkx0z2Xowd+pWc8/x
ruxYkIFMGSkTJdyQNYmdqZJslg+qw8SpPb8UiEC446HYsBY/qClg9gwGE5HE8eFH
7Xt1/xGx82lqbPJiwP5Mrw4Br9SfmsZ7i5Vpdh9A2wjUmTh0t3IwGxHI0pIJWcfX
M74l9zGqoi48puqb8Mh93TUuvoETmD11i5mDX966lZ0Mu1jGvVdU7hNNHDLpSgXb
TEVKjfhOa4oWQx+65xenXUpXkpPhQeYMPohxrpCSCjTiIxXLz5i28Sok3XlHoU3r
fPmXICGNicP4xY5/inGa+bZ9Tns7E8FRuIZpk8OgKjwjCNC1AN6ht8V9ULblEyzd
NdL2jXPTuPu6dChTMHtkbXws8ZFzHdAoOTEhifW+VAOvFxeD9ltSFXS24IF9Fcjg
9JjxcGR/azZ6csTRjm9ovlWO5KDLjz7jwLueus+EbxisaCgvPMHUXsNzeFx8hMdX
9EZ8Tf+ZdzKesJZRB4FIgC2AZbxUkEw55+r5m1o70qipJJImV9+vjeOp3sRtv0mU
RnwzI958mwtsVpR81L9A1J+6I+hHhMWN2yKlgd9x+o8TH0CfoIVO+z3CjwfbO46n
HDT192T/4dC/6B/m/NZIAsUnIKx900zRH5EFuFH1eoKPx+mROpI2A6ju/PazS0za
itRMq3tU0P8Fq4M+sQsmbOqFv4nN5Kt/bNtVtqJ27FIgGWKmR9EIqwE8oJlJ0nit
cW00i+vZO83lfXVxEuXCSFVvMVDlDrp8ySDpmDAB78y2J+i3c9P7T7cMa4z3vXsq
z/uIDqVR1ZhY2gleqSoO2v5vs9Gfyeae+eU1aVovGyxRrqGbQLgiLn1OguegRW00
nvamwC06njwNRPBy0XjRAZGVnfKEhTQTd1fPJjPmA0oyR/UVBe5N9fGRNyWVdP28
spCwFkkbGvf9jChk1iMv1vmsD6ijMh1fZMrEdnkAh0nTwh62LLgCbS2Br4cXMTX0
N+MlOZ+0XdZWvl2AVSpGR3bb0pvrWKuI+ZdwPwVaQNQFnShYVSJFDUp0Kuqjt1WP
IfaeavBa81w00MvynkJMiMzDZCcynALLyuxg66neXmm6FKJvObESUeMcb+fiWcrP
QhkmghZShO50IVD6wCMz50d3g3w8NxOMFkMs+p2y4Z0StCyCnDIC+Tnx04YZPSXv
s1uF/TIrkG6VYLsI8qLpmBqaGZhUhdjVGPHipHiQ10s+gGkSUafgDS/Rvpl8A6Y7
/s02hh/WvfBvFLR+ufEMxFQcPTgpOhG8+uCywIAz6o/8q4++255kR/sclVDYB3FW
ySa2MC772r4L6Gu8IvB/sl7GuP1OdQivR1h1libvvC2xkYVgmE4p7NOmk6Rb9WgB
sFfAjs/zm+4eGn83xbQ9l0ikedq8RyZ+L2/RZXmyOiHwtYiurs+kStO0mXO8Fh4A
I97qJgGVi7weEMA/a0M/MDoBmB4PHG71qrWI/9WxNAP0zXPuaptni35RD3mex5WZ
84TdmeHVhm0TBKuthV/Gt9+6+wEpB+v/YM9kEyJa3zhwJ8QlJceKgP8++ONAoRVq
ZiqvMeLhR1hLx/1BHolipUci1v0Lpg15R33oN+vJltDe06wjJG4L/2+EwWwoPaz0
C9MJGqUZ7DRcCoV3/Gdfy1QcMxoWkcncjrwxUktziDD4R+9i0iKX4cqKDpuGWv7a
dywcfknvkuvWC8Gcsg/ct9lPOC4+SMzjw97gB6AjSDbGWnAFIerbRmrp51UD5Wzm
ajbtewVEcC6veu5OEkZk8nWPO9GT+8gROxLhK8fTaKMUq8Z9TMt8/tw+NACy00Gr
dvjjMk3pa236zdxZNARSzj2gkDjX7M9C4oRagI0wSPnSzwHA6ojChcFwYu+ZLWxc
J1SP6dcwrVgH1JI7wKYU6fxvfnkFdhbJHv3SBJ+knXFAh5OAFe7L0JPif+qgKicC
2ouPK2TFbMo/HTlr9A/UKntSGTpsrGg/TYi6dn7gQnDgkWA1G1RZFpevI+23y1Aa
DO9A7RCS6T+X0KpTvsEPvZLD4Bg0ESJ24oSI/6aMxHSkRVbzigOksajWp6WU/tMJ
11xJqKkwMJcIxs8OoyvoVCR12cXCdVduiig9MfALSuAwgGHalnfTZhSFt7T2KexR
Mr7B5rjOaKN6u/4atiwB/JGmBbhqJY/zd8I8jrQIa9RFJQB6c06lyyyI+PEmmYry
AVE14rJq6V3nZLLSjYvN8F57Twc9cD0ppv/BOkmgwlxCLr6v0tTjzU1mveXVvfzy
1VFgwWtFvtBhABskUSpPXD4klqzOoT3H0b5+iRUqdZmhuaoWPFJs7jMA2+WVTeic
B+siaL4s/Jxh3QA8ll0PcROgQL6VVZPkAlX4dTFsKmDWbHajdogrihCJLBC8bkzQ
Z2oX02l8sv8Czjm2ikjV4S7RIOXsdNS9Yi/Y7XAz+AFDazgzPpL8GSL7LnOL/P2B
bb+dhsdHhcCWfU3qVxn6QHg4nh0eE3hKxcGgQ4lWKfkQYQnKHcU47qrJkBGaOU8l
c9Mqd9uGM81knrmmJRCc3BJXSUDFIaHMhaXM47FvORjkDhdYGTiONCp9gr8C04Aj
y964EWNdHU/l6CzE4DK8KGWWjISnaaisKsdnsBx7okYY7kNCE0eraP+bkq8l8XJS
41usQT7zTr//x4gd5sxvOyM8+iCrLFZhkB3ph622SteqX8h8y2MzFHucvSpfU8Jm
ipWWuiQTPEHCMDxdhYCysN/edlHIhIWsFLHQYGWzPr/9/XxF8iR2/g2Ig3dCm3OH
GY4RqZtLkP2QnkU53fZFhoniMSi5xuuvaezPj2428N5l3j3UCkusoL6HGlPbMmoK
+xZWHp1reTg2uwm6YucWDvRXbf5JIPmCPEjQGUllcWPDgl67MS/YAmoA9R+xAQzR
In3fBl/lv1oFREsFaFFpFD1S9FEZETxdAuRFI6irLFIZ0o1hysHpOjuX7nb4JFhE
dXbUeUNTveRTdqMsvPNdE5wQKrIwJt3IgCQeFZyk6LCsI/ZNsPtJz9G/py0vWdVW
u47xR5Ul0LK/Bt+9NebV42JRajbbC5ZCijkOlrwXMIVW7tlbFpGdqfU02ehldzrB
OQ/O3h1PvnT8JY94/eBayovvcpSXQVH5ajGSlhfdO+YWotg5CUZKbbPexxzTJauR
NamGFH2ZXShHlNCua1lmO9a9bnvAteioAJkYAoawcQr8IRDHdSKBvLX8NlRKk81V
gQ8uvaXptF5a9ov7JIL2fBoMqkYY8Ok4kphCCH4DlBL6vLyyB7pCQlvDmv5x+Dfo
N7hy8YeyJP6/aD6ALNN6u/BHabD81J3mdVGSG3JgL5BHkaaEsEll5iD8JzYFYc11
RiaQRNBiYysFMPiBjTtoMZqgUUHk+xNM9rnl+7l0f2fglv5uklkDN+Uk4ENfZtRI
6GHoRqGaooPHCyu16xxwfllmfb5T7LgYSCdgR9KBNLfzsfzZC9H0Xu9MhV3ZVQPT
fjU8j/TBYWkLUxKqRf+uKl5lJRscDiCUxERrXRQWAqBPfXcERt3y/RETQxTpTmWP
wgEDMU8xCFhX2ERwa5Qg8EDeW+GK6KIHP9a5CIN4vA2d2PLBruIpi8o8qyBet7jF
jR6wkkWjNoVyId9W5BL5vZ5f+fgbVg8IDCy7/WuPVUybalgpfzd31TDUtS3lnPxa
Q3ssU10PRmpF4PquBn5cQ5aKBiHW7kQVP71wORAiAr26gyk35hwKIxZt3h5HFmzQ
s1DKBPkF/DufdsZS5lNamhg9fHfI4BF5r0dif7qf7JJIhYqeWzVOyap7oixJJf7L
s6CGfU8XAQnQzCHstRtTSSuJtTPblnm4yIf9IPvAjbppGUWcgumbfrXBVK0Vt3k3
v+Xqhcfbm5SLVte6SUK0FwcZl3XvmcadMaHCyQus0uNr/ys+60ffL0p5ulsczSlq
`protect END_PROTECTED
