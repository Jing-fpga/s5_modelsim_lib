`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j2RPZAKtF1k5SBA5SuIodvn95+DkMVHfXSsjmxbV/W7vx95tnUufOSJK/5f6AXnm
hFfkpBkP3Oxgw8fhpwPHIz0FVG0gmYALLcPEVJ7tDtVP5NwiwKuxcwei8GnxZ9KC
4EY/eQFgwhGCLCXzduEPjyXZMgTKNh5/2AsrMTncVUqc/J+OCwM2IQTiALbEApi/
kJ1HVQ6REf9BlefumXTpNu1z2g/CePVT3lrMe2XaY13/ZHOPib0jVZOyOTGPsw7U
KOJC4cL1nNg6upD8jXOIRiDo7ddtKqevgibd2nBW/Jm/kq6d3mXaeEYl2RR0ES2b
yYBPa0DMdYpnw6HEQRSzY50HUijdQKO/EoY/2utOxEyyz6DTgWSXtDqNAeuFVfFd
GlbllbfEPcKE6yT95659xdYkrxCpXPm74NOs44rYJrpUVrAsZ78j/7WF5/KEa2W2
CUN5osNwEkGnGUD2Yjc9xnosEzBWhERsGG/rS3/U8hhcVOsKPnixTO6wTKQ+mPzS
eAWN9m+7y4aJasrs/P0ZVff9kQXFtpwkguwXMf9/xMwM9KtxCrRFDVr0ZwUjKvxV
a0GO8ealgOM4H+jK17gcDobin/ettHWs4v6j9M4AtdLtwqeXZLHQXjqMVCFiie6t
kaFLDZxzrAMZzyZpRZBQN1SapEAtI86xc9dsWHhGsY/cR9JLSe+0GEWUpl+boxR8
CoecYZoHxj1LKczbkCZH//lxOlJ7lVf5T9vATTHC5YR9rukqhBjUh+rslDnaX6LK
BjEZO54QrW7XZD814nci6k8wCbmBDAf3ghhBhdBN4XTNVAw8yuUp6R9LvhanvtT/
gkUmo5JmsQ1YLrXd1xFtGxJloHvZkgewZdUnzKBLSpPfzqAgUuuu7FCU7seF/ppz
kxF5bl57t8blm7M3QBd898xUFJFWE4Z8OYkktr8LqKnn/SQKYnaOOIIiUwiNR8E9
ycq3wAoKhH3MhvR09OqpsZ4ArWPhITIpdfjTyvlSdHnrtShNdii5QlWs434X5NAb
VUoLJUflE5TG+DdTp0NL03hxKymo5flyOcme0+s7eHd2Ub78++Mxs41hknJMXfme
vVqPrlLWIUKzHzGYKWHso/UZszvD+LEnArZ+g2yMtM01ZwJsopj+l4JGnpyFd63X
GMfvRyhJblzw7UCOx88MUY5k4yNcSwUg1G2zLzL1ZGmstSCIGBT/2OffeSXmQCwd
HKBUgxFrgigztTA7hqg8BqonCbARTRx/eqLuFOyJFV+hBMGqASXP5zoRmkc6mRt/
k3opwLi4uoyhmzPgHYlhFjEHi6vzn+iLp4sV8z4PvwZKmpLQfFNV4euIfhwVJdH/
5Wr3+bhqKLEp81kXtr24Xw==
`protect END_PROTECTED
