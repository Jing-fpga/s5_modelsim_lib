`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wnEp/d1xjqzDG42tz/AQrTtp69n3GN9lgI6i2jSj4B17y8l5jgql3+f4XCWGZxzM
58M73X/mcC80FQQa2bxVSSl8DwaqB3lYnKuVahHDP7IbYShrnLYnFo1iUMM40gW9
IshouLoqXpd5aOSsCtL3IUNcr29HPcqLcKwypFz84q/qysrB4MnJPpm7JE8kypIi
m0nOmE77/zJCjsXzVy5z7ljuJGArYzSF044kb+OC3o5ri8O+SeT3TY53br5GTQW5
iEGBtVKQMjU4ls3wqj0ZFBp8yM+kFAi5mulBmERaDro1aZtLULa4ZOKXyT1Wh0FW
Aa+0ojwHM2qXBESPPIcWwqvWODrj/dO0UmT1proLduKVjN8S+UQd+sC/wClnXmA3
OJg6h0Tz2PJIu5HWS/PXY4XjexfT9IFHXtCvqAEztqTmjF/PY8gUGcjdQc2Xg6Fy
O8185EeOz3mkQtTFVghTSJCotl3I5LWJB2gvbycvYmuEAq7XiZTqsTx9P6l2lvBv
qasvm0+6tR0T4kZtyY6H+ntDWT9CrSFXaxbcAv1oOF45aLZwBHJmJR559hjugqRc
G/zFGR8QcosE3DqO+Ut6h67ukMQucB2tnz06mVvc1xD7gxt1Sbm2e3uuS0x3VaWM
NbEa2oE3WpcQxBdryAl3ps+Hji5rn7eD7UOK1kJ8DAMmy0MNIkzY4felD7chhUgF
mwz27s2lbM8h5ylzSbQEhaqs+yZo8CR1ysFudRz2gezNfYn+efnpwxRJLi9SmBq2
DBJBMYPmy4w/EU1PvZbTSAFO5/OgXx/4JoHUMHArc9QY4hp9K9Vk2aMs9nYc37x4
4I3zKjz+5lQSDQXeNLE4olM1zENlufHKbWvje7EWQ3AXKEl67gBjiC3pB9OOKR/9
YpEVywIz5aGn6xa7NL4RY7jtRefAhGrrtGPw28PLw5ifhBG1jitIiZF57xDGGvtK
dcs7IJfQKab4tSdjUfKewzTVwJHrYnQQWugs2/rtWxAtGYraIel0mD7WPpMcOxK8
0wO0U3WVr42J7MdbDi29Wyhy0PG/wYxdY2TcP6Ix2YVYVO3aJ0QoIgzTFJalO6r+
xi+pX2baVnw56ovuSV9Axr+BhceINDCGspUzcYRH8jlzgrDpMED178zqAyLOXo2t
OZhr974Rei2lGSPZ1mKfP7uxZqAOFtwB06dxfjbAiFTqLVVXb/Zf5yoSdkDP9JJG
9H2DAldro+Mz5x78yO5+L3bbqIMhuCpDC2WmI/ouLx6Rp+vjZP4m8f88gA0bMcAL
AEvx0EOQ2Xk8w2HHl9oADENJ8BJoKIz/CCUbfuQ6MxWiq/89bbHxwVQcEcZ2x2wD
nW2D9KN75NYXph+hF+nGSBVY1VBolKT8NG8SJDe5Ogvg+EYphDYJ2TShekM/3Kot
fIT+WZe6e1v9naMQFhvVSUJVlN4ZQwabyvM22rPRa73rapeeDDVXViO5RIRDBNDy
meRz+v7jXc3QSw6YHrTncVByW1ZLHh7TA3xZbwC43+0GdbcDpx9oE4/0dZV6denR
bFSGnZKx3kZa9lbZUgbJM5o0I5lE3PIg6NvDtl2NePLgwCzdIunRUrFGH9CpEK1V
aKbJkeI5rjQbLljdDhysz/TRVcnw+afJZ9Ee104JeYhzp37rf5UuNAJQpOgTZxjb
VRzUZKUOgE4DhSKiXNrH+rhhmXT/3R6g2O9KDH5359Xin5KerFfzAOmljVUqdE/Y
n1kDRkWpErw5NN+vgdXH4La2QvWY96/HErWR5aOFIZm38hbmjbLIk8l0Ee1WmpdL
6Uu3vUl45ubmsZc7DSXkpmrhz7Cb/syRAtmAtRNhdRPaCxV9JZA9NEqIaMJ/1fJt
HKZt6mmEun6lMcjit3+7UeXAt/SEChTt1LddQLlcfDlkRcYco7ooJrZjXrH8tr3M
Xsd8OUqMu/PlrWfsdmWzMXmXwRfn5TICj4oerylqUxAmQ/Gvb4Tpl+r9FZn0zzpJ
dSTtSLkncMLyhXPMlR7O98WCYFIAdM1EMlxFZ/dz7rGOP5QxAiWopK4/4HSprdGP
zFBqmVOe9GO+LvxyFmDujCfYxsUUWDFKNEtCj48SMKlQUfFBVLWf0wTg368b/v/Z
C7PwFsSROjUhM1KJqwkCjmUG2UABdumabsq7xQHxdXPaLWkWATeaPli/NmEdqKaa
TCN9KC6DPrilLON5atp62pL06KjulE4WP5SMncMxU6wh4oiuUTWN4La5nVJcPVdG
CK2FS+gFwQN0kF0mpFHGIrU22fOvPS4nJyl1ws4YF4GMmPBoqLB7vtPcK/PCeeEr
yb61pGTagbn3DLql6v5mT+5fdLnTrp6uC+ls6uvMhZflvVVYOU5LsV6OTbMpc/dW
58f+GfthK3AB0eLq2UMc1R113tN17Bkbkkc8DJJl3d5bc5pPcmmGULXSPqF+30yc
bQcoA6wsx8U8SHf3NowgCK4+0t/+ns4V8aZPJG1r2AwB2QQcVNglfKs9Utg52DTN
vopZdPMz7U47TTi/fTtssErAgKuWLa+msXU4MyRlRpVOFSEX4mnBzjrIjqiFUsEJ
SBShtrCB38esX36/JPtAA/g2Y702xHrdEOH2N3wmieA5ZFyJokA8iI3JUOW8Id6w
QKXtwEvj9xkc7jYt2037ZCnc2ZZ39VJTylG9V7errmmRGa0jH5y5DUGey5K5zSNv
upCjUsGHjK8eSOhojdh/JQgluUpy48WVsu2UZCcBg51nf/gZIlEUDXyrscXG+ipu
eKyg4Lstwym0GuBvPcmZYknXM71dkOndNTUJNyGsa6Kx2VuhbARVoe7qQUVuHcbr
H1LZLdr/Bv52gf/UKKYkegG9NHqtSHKdxWYhgl6eyrINU1I+H6Ss2dUPCFiQiX1V
sj2uK7IYhKVyYnGcD8XegqNg6PTshORGyP27nTecupRx79hnAxqtUKLeitwxANE8
STX7duToz1D5qw9NH/0TTF28JcX0Lw18Xt42otWUTOQYdSdd3v5+ga0N/SW0jCC2
+DDsXDdORk3wzpp2I1yn3yaWnOWfdjjSuPcU5xBpzUh6ZROvdtj0dSMJnCc+qLA+
y31UzD8mCfOUKtGqwoall8W1wHjNfqqNkdvZ+UK5eIuTSDtklAd48t77evNmSNIk
vT1ojHV7Frb2CNgL3yUtMRvKyprRoQ/YGRhp0KDxoP/cDIXo4klmNx5tDce0Xqx0
SBp9R1MbMoOa+PJYJt73PczquqhmWXebWC1eHrUwEsESA7HPAOeoXukM9TqP+yaN
9qQF5ineE3Fk0xZSjshv2Iz5BXvT8AzXQgSOg4JGWTOw/NaskHSi8/QSceOXrHai
koXbraS0j9Hi8F+nEiMtvHxQXYeThKjks+MsfMlnnly1yv5Igqw79FMdxahN4sAZ
kCi/nhzbrRWsdTwXz0OE7OS37e9PB+ME92EDRd8wyQEIO3ZFOo0BhPgmZvgiCBxa
zeeg3tttgU6UxPB5+qZf34M2ZWS4nNQ1QgRvL1aVNx9XwEEZXotGFL+cTJ0DkQSR
AUmNpVwEyb0QkDWs/UzReamsw0BI1bNbE5wmhby5ZkD6BSMpYa5Pjfq4M19dzswT
Ubt4LIuRRbXVTQKfB4zdVqTVlpuHhBwY8z1ar6QxC7Tfy6Ty6I2f3eWg+qexUZj4
UvVmailDzW2UgE92lrsIIN450cIBypv9ms4R1vpAF11QmRSynhRmBJ7PX7Y88P6F
UcDp0Ii+KlFCZINyPzvTFj9hyXIqwzwksI0ET0eUwgcZJUgRkNuj7WzceLNV9jla
GZ5UOxiabUKkYnjn/HDQUS7JHE4CiHIh8tLEZEu0BlG6f/2JxWfasdR55nmnhWEB
c3h8Vr1/QXZMwQFWGY9tCgHT4QqFHQsbdYpdMiVXEWfGbWeIt+YRB+CZ3WTYV6Jh
AIZ92ZBvYGKFVU/FC2E09fo8TvWick3rnxfoDD51qNnCB8IECD2zkzDGWYfd8SjC
IUXB6YbHOoHlLW21itdRcTJVVxxsh0hA3kSfZui9CEnQXjNDwWm/MvVm3NskH0pM
lgm9DfgeCIELrUWDmbwPEbGG7rci5A9ApWydzip7XS+1g/SAUMHvsuUYtuxbst73
BB9X8/bJj7aeO8H7c3q1ISEitNsMFqlo3eb5nVEgreCE7k8JRZGqr8sMxdLluLJt
TWKyxXFlQbOjCggacRH3Zy9o5jN7LpekdWIWmBfdT+KyoAeIhLVHCfQ8kugccUlS
8RzmP1P0JQH96eq7GSPpCOqsk27zer89ScfmOStMp0xstEvECC3JNvp2PjozCKrf
kYEDUNrSTxAf6FGfImuvz4h2GRodFx3IoaZhcMMsREpMHR3uB06m2/acuVK5GXoI
fBjVnA7AoKSchqFLjUGMw1qscSJwegwXfRmxzpXT2vRqp35x10lGJWCSD1o7qM6e
CUvl2fxTxDBvTrZBmqVS4sEZDiGnb0ECORrikjX3WAx4+x5hU9U+4LkxHsqAlaOf
j+zmjic5Bjrgid6nPJVNzfoUEBFXzq/yAFCtG1sBJ1C2bvypsBxYhMC8R2kXDLTK
oXxJyaYl4Oo10JgYeVry4ze/+cyfnOH2VwHOFmKvZOJD5EGI29Ue1YybvOWIOOUd
ALv28AaRozHCOa4JcRDnQMOg6+i60M6rfenOr3GF4npXb/7CD8SY6YoADYYAn0Qx
M+NZrnCcwvpfq6+gAjKmxCuiBARfrKwM0y7k1RYexqKND2SqzsxkCYPo3+NV1WnM
zVNvPJq104dpHH7L2Bz+WY0HjCrJ6MVieWrCri6O56ofFfdTPo5UExl/nvq7qeWf
k/GGLhI+W8QOFwQUqIcm6zEBnpv5+9rHzJbFyN5eXxKrP5gQag+qlT0loBDEFy4q
7KvL4kVvvIXrT0JpAJEJUcmtk7uPrG3f2M6lNoLN4gG8HojWnItpp/G5zMBDv/iy
glDC5OWlAkD0HbxlAA2sgCwb32NSJiMw0aeJPOuPB2ZZdPdQNqrkAxkFeykRksF+
ob+quc9BJ6j6bEwRMpCQ9OeTTvT/aY+98g6jqqPOzRev7ABBkUf+ZHA2y8yLwWs0
HJEcmiBSfSQP2rq8J6ZZ+0DTt/ZiQ1n3vymunYic1A4sxuu48Rc8loIP6/h/0WSQ
DtxopIUnmFrGE9SfSingmdjggPzryAtxY7wufkQWKzGxqtTAxJzH048DNC4gP0o+
2BtlqtfXzWctPeHkcqUdNN5LP4wCSEEmUEOxeNxQvsjrZKLNffQRz6JJ5Nt+O5Et
zzqjCvmRsdoCUnKtCcTjf0/sqyQLb3jpm3oM2onqwcJGT7PlbLg6+Gpx2J8CoCHb
zoXNBT4x3hQ2oPaFTCUggMQrf6scPNAm6cqck+x4KSe3N8SgBtRJ8kvnAivOI4zU
LuhU80M1baHZHLwMmdtNPg8CZZzVEOUTDefwJvThjV05JEWBluz6VErcKdOZSO50
0vMJKjEjZiRVttoSofRpTAABWA6xJxWx8f5pE1elU9l9+PhwwjZikvxqcfRqMiih
w6Dm9OGq5V7y4wqgWsDQoviLZo8pEY3DTZ7AbqaLHhEmyhJu+i33llijUHPf2Ird
o+C0cwkvx41ZLyzzfxn1GnE2cMlbCDVayWI/LoHRidNnhAf0IbN08wnVrNIM57Zt
nXgi3G4KkmFSOjDtGL9veAkpj0vNM5LoE19kMR69zrBMKRHGt7bolZ99Tt7RNn2O
pqudJiueVm27ARaXFeUFAIDwKPy51Cl5egROZ8D2UTop7CyeJxoYSwLlH+ZvW+42
aO2u77I+8txa9Iw7aYtg+ROMpjFSDUibSHXKUK9rcoAYcKv2XMpoMX0ciEu6H1vf
G39hB8EALOB1lGUJ89fXZ2Ml9XB8dSIIT6IBDvCDWPXq+FNH3Wm8fldaXgwDlJ77
HXrCBh/fvXmsmaL1uLYSXN13MQb1HQai4IBjP5exupY=
`protect END_PROTECTED
