`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OFA2ittoHxYC5tQjpe8gQNVL8WKegDKCpjO5NsDSQz+1KdLB8eR9hP55QPkyiop/
h7u7V7JogK+ulckJjeLXRs9gNiN+fc83W8+Zo4Qt3vejg2LbF1SW76tiAPPjLVEW
4yMmLPWhOEnIUxE1c3/yZ63+KwqkEQbONfWHN5a+z/NgbX84ZoYx4k0R3/6K/mII
HzAKtcOOq8Jr+KpitqaNN6TnrbJnXyN/NIdYDIAXVG0UNQFzHnGhjIJxCwpQTLg8
w/ymW4AHBeHoQ3qFGBM7j21wkaRGHoWXjKPKIzCB9yO/l0qILTCsK6dJNaKiwVfM
RMWQjORM7Q25dfL6mMCK6Xu0nwH+9xS09LYP4WpW52fbibbIcotN8qsN9Pa5FSTl
Q8pdkDili1vKA3igRDdn/JYMx7u/NuBfQPv2gtABMiE/fe5t7vdpLTG4OHXCLq3C
Ug7HkppoaucD6fqZeMisMo/BOUCdxKL3+G6qiRqzeYcqTga9t+oABg5LynaiV769
YkNzqruPmR0MCo3upoPf2fqlne1IMgVV/MOrCuhJXl7TK3WHcoOzn3FjKu7cGEP1
B7HeSprTBQcpUqX0Dw2fkm26j4GSnW2yxdq54u7D7hCOoqsYQtM/IvOuNWcWRdIe
xzH3TEnsJfTvYMj84Tl7dCK67QfmRY3pAIA6w7+FeLI=
`protect END_PROTECTED
