`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OL3y9OtIQkSYEDRli3f0FShi0zvav+kuiJm+IJjvX9yUgjJcupaMtJw7GGF4o3+U
WfvbBjxhQqnWEThDApFAVBCL4m4RwRznwdJLncMJJy676cJEnSlFhkGNF0NJYiox
MVi3mDzkHVdOf62oPfiZZ5Uh95F8PiVUdUEXGUz0Y5PSpMkHpGtZyix70DrRofeL
YX6ZGx/6kcX61Z42XaW6zWm0lVBdvLaw4kpXm4moKwJVArmFhohiWvstwhXSdA9+
nd3jXeD2Y2H9a+mjioyPULGt6eUJxTvZn+c0xU8Mxyo8vyqLmtdCxCqefyTTzkeu
uepf7o4IwdSccqu70pn0tC1WQ0ZAlbFJsWoEVX43uCF2/qOYIrVaat5j3cjMs49I
B1C5OEihxzzv8Q8TV5SNW98lLBEkgV2kCuDI163x3cX3tKOqe60GJrBEn+wTVocw
4ksHOYx3+3YeQgI1JDtMewm1sg3AqSiyMg7Pp6gFQIyYbci+6E/IUJD6WM9fOQuZ
cwsDlSjRWPOne7DyaR8SFBnCIppBVXo/kApMss3mIqIimO/NvLCcVcYj42XSCOzA
0Cfzdo56JMhLzDVMc8h83U9xlFTSLbeGCyYW7uT4LK2bSeErfiVGZBFIXEdZZOJ5
Kj9YMN6aeMoEvB530qgTdo2J/YZ6Wf2u9sBa3f7hJ44sruuYPvCvSx2Edi+rh7b8
uBpDVIyrrvgqqIxOGMFE4D/nVs3uYes860rcyUa4yTnwF8PglAkpO4OOxhBlrlEr
H8w7/c13mbZN73TckyOW7JolQY8HCvCUlAv5hj8u2gRQu45fTUApndl7I33uqqLA
c2CLqtJWa2uQ92wsfhf8IP6oDwabEtoI9pILaNwKmfJS0nKginUlqdhfqtJVuBbb
DuL5osOp5iTuIs73T6A8RD+MyWoU2pyue01Whe+R/RIseIsXgejpeq++3B2t+rUJ
YfDiOV9uysUoKfRweovBdqSor4XwZ7Y2mh6ptrXaej9To4gPwy+IdI6wiM6l0u0s
HNvq8OTPOt297R8jOTWBL9cC8YoRnuRWFwJ22ybe4wj+kZaWR5nD4srfP3mNQBXP
wN9hA4QTIJ2vfjfpaC3dcc4QCX4WHVZ/E+3PKHFqE/o93HwCjRxTtW5jcIJl/HWS
cjgE3B7HX5aa6xrsOUDaxXZbL9ksBwdIzDf6kz/9oROXQfL/yAsAnTu/CNt0RF+3
CgcH/jWdoroMndTo+eY1uY44c56V/jYoigvYHW8oF0cCVzUFy1BKN8ZSdn7WtzvX
rCQ7iWVmc7bSSfmefGAUuGLR3p8v9qFwh5q+mpX7dxEG1pc67Nmcajj2jlAsDpYy
ZTDhIJ9DBwqZf7H3DzWVfh3KPsT/JJ8GJzRjlGq2uy2dyF+yDf9A0rfVapKwNo2Y
k8huofEdpEwWJQ0OtYpE1gzWN5s6WgJekciI8g73fP9nMD1L5RNyVopplji3LqaJ
jyAjKEHRHQuMpJhRNU+tu5IvCO1rd2mBMRJHIwWdSSYur2YA0bf8HaqYFIp4F9E0
CiIZ5Is10obHdkbxadkoDGl+WwDwxoOM3P4xKbauKe35dK7/j8TPVDV0IZLBfqHy
AlN2l0H0EPTQf1Hw/Dh0RvHNDsSOq0Ga7xGnet/BVkkD7PoFhtSZrTQk8a5m8D0+
2fFkv5XJMLJtuNLtAFEfw+HNZwxtICbOOvDIpsuVO+u1So3IeXWnnU/iUQTc+Tp4
Ppti/c6d+90m85a9A/fCipp/ULdR58VPdPA79BclpucU21vWxtY5eb9sxFgf3RSc
E42RhjNn32MWZv9g4wtSAm9K/2sGxr6qqD47aOUdd6635BSgeBv3pPjHrF609nHl
1bRvECe5Cb31itQgbal5I57Z4mw1xcZY8E2Ad0B4+QXjS0eXWlZOBq3E6w4j+CeN
fpUds62U/zYKrAcauVcORqAmsak8IogudV20LPgfP92KokpR94f04VchF17mZDDq
xsv0LGqRWHa+NHZYhOP6A2dhASTQgLvdZPXq2bIuh48Mm5Gk5J+NRq3bnAtCXzyR
4rSLXje3XWEP7NP8N3rp8rA8lEfyUmHZ5O+SCbxrGzUeQBEXd40sHYK4WYEBY3nu
qAYBslSnuCSMuDwvBbVbsPafSmYpFxYcvJ/LdtCpKXhQX6r0sa4TBEc6zrwI4a2Y
aAy2QDZekPSPwXzsFTdF6u4UxSwTa5QG8Xf38a7gcQIhS6HKH5z5zW1AcCwAF9xC
ccXF9Ibh/wtI/KI7owexFmZ7w4iFboqw8ZqIDviWJOuYtBPiCwVZnPcGjU29jBot
cpHkIUc+Ml1eUdf0tXFGEp2JjFEm3e8wkYXCmkgpVgjY4HGRbPl5dZ6eGS139yrb
fknerIRZcrREy1TzjW+Fq+xnEL7wty9TyaZymM8cr/9O5AeNpSnp1EFfgdYuw5WE
Ffcz6QhlmaMW6aPuwx9KvEtAktcMEw+ifNigm66OUvjZIKypAubazZGmTerkehLs
avs/TFsXlR9mDU9muhQ4MIkUadD6sr1BKWIityk5hl4a0qMS9o5BUYRePqKarb4Q
JaPqtXtjaKpYVPnCo+fDrFbcd1gclPBxZ9uJAiULY7UaGFv3qFnOoumHxzO4CY7s
TtB+d55QTrxxWBVkFjOn4uNzrR745R/Jb1wJs4n2g3mG9vswt1OOkZxcJUakNAOC
JtC9eZz0CjZHdUEdD3DISr4kdKC6IjwD38jvq25QmmKADCpZJzpL28y/8ppAaoKU
0kBVZ9XcwKikdF5RZlzsicVxgym0mwO/ZLYR0hYzINskI6b0uIGmfAZREL3QsxFw
GMjvVy9liNHwrtI1wOMEOm0OfYNIsvmhegz/bwiBejTiujOZTQl3QpmVbpWSNnJe
etlt2+3cmZcFc74bP2sEgDH5Kc8iS/Sbd/pXdo05uXhnXtdv7V46s/Nwsh4uKq1/
4VY8S8UDcL0Y5H5yDCQAEyPfPYS8K34D8/ixcwC8T6VoLs8RToH7dT38aOM6K1Tk
tH1X9c7PkO2Hvd807lBE9pIxlizUFssSczlM1kIIwXdVubIIKst/J1lOrhJKwndD
vsUn3RpRa1DJuxN1ENStE0sr95Ntbv/+4+/CjKSv6f44+4eAaeGT1YvSOrE1ChcG
kGIAz9Klc4xZoBjJAMMDiXZ3JJwEayb4dffGSAl2EUPOuSne3QB12eta4kHyZ9Fa
L9RD8/CpgHoVfftbgWlMUejIWkNpbu6eeBxbIZ6YGE7oBQUA7TbCtHuaNAVulnZ9
M3olAoXtxTlTg8NtrrnXtGKMqiMna0r3gRSYAYH6ja6kGNcsU7WtCh0fYpgkHiWx
ZJP4dFrAW/acERTiKYtO31at9yISTYDkHd6Z5JUvuHc/9fzbmITo4r4uiLU9TrcZ
sC4PgRkQ0Vooku2pwkdcpzOtle7a0MgPcYf3NxQ5KeEbsE2MsfxcC6EouMZEjusn
u5JTxL3mJX/UnrNOFYVOViLDHh+aM+luImfgahfpVeVwhLEwRNn6dvygNHP85Qtf
LhedmgoSooXT0brJ+4uJz5XgK/FtrxJCVy9z87SFwCOeQ+Ph1Q/wVJBOOgzFrW/G
KvSF/V/AZnrZw2EJ7Y2TPEYlElCZRkInLyZYgVPbINCtY8rsLCXBjHVXuyHDW+gi
gtUkOdWiYoJbMGHq85xuTQ==
`protect END_PROTECTED
