`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l+k50sT8jWWOTZFgI0tIKrnQkHqwOyVGfzRTMIJlE/c3XlKAvLaNgskX5W6ZjJPn
r03SmtPF8bdtjs8BDQLwYaTvH/8+gZhSxMo4YvQ1OPmyQ0I+WllPPekRd+HBR2eX
SrhLCeHKkjF7RyboM0K2nXzKCBLgLsnqVzFMIn2ApRU1y7JGdyAmxyUbLKSj/0mp
GOegff5XCzTlHmFLc+Kn+1y4yBnmFimjDOjF+xjOlSL1L7UmTo0Pv4FyA2MJ/6nO
2qMM4ntHHX0IsUrtXy7sXHxS/uYCCWnPTDtZYCda6ecL1qSKZIvNunr0tXPgRIkV
WVzhuLgZi95qI9IEmOfiGD3NJcZ1+q2vOTCMgX9pXarGBNyGv+UDcR8LRnXrQ7xE
y0t8216+oM31k10iELUfmqaP5qiFbkNk9HUR5kLETAC2iYHCJFv79dpgJsIvJYlL
yShs1Fry2t97pP04bRtTJcDsbURDgAYWI/hpTShe++3+9xtot4iEDMw4LVvs6D4+
8dL6RAyBGXFFH5k31UPjEZ0HeHrv8IAUCPSBUjRGvX+ZZJ1mQTVlogHJQhZGrCcC
UflhvjZdgB4yP+Cjh0dqF3QqKsGOoEuZCRbWDIBtXQ+C3nwoLY2wuBcDaWtcgbW7
GowLodNXJMgtZ4tO+09AhnzVIJhp18jLNlTHtkTAAjMbTXrh3mwzaRgQBFYZ2h2s
9wnUnprY795XQrvaV2Wscwj/UR9F0OS9U8YuFmU4tRxaftvyh3JJiT8gaEV9+zNv
TbP7bZ55KnxsJwu+TShQdIM0gKbDVYJ+EDU/lgmwQiemXy6TJSa4Yml2Wmv+aF2c
zTEuUc98g31mJbr/jFO8zw2NACyUpE7CzrIEI6nERCPT5EhJroFbd2HBfsSFJdR2
1/OxuIB6NaerStQqoBdv47mM1ivy1KbwvGmlTAuvx10/EaHGBKRBNQyWxDhlcBSe
20GLh1003UQhNkTk1NkuR7Dtv0BfxRIJTf8u89q2kBfPMl0XQU/Ey6UOSS793BYr
PpP4Bdzw59pe2IygtUomSPABG8bCDQ7NhiQJVYlPsKUaCr5wCe7/cCOB0KsQQi1r
OYJVQvFU9CcakW2o3P2mwSkuYRg+dD2k21cO1nag928M36E9KfufczK8eo9fvT6z
iyzKOHe4E3AqW9TTx+ZRDaWS0xssVG/qX7QPE8V2695mVpYkVMW7lw7EPAcyQqYT
tBt4hM1w3TyqAz50m9b0KA==
`protect END_PROTECTED
