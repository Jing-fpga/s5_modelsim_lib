`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NKLQzsjRlmgNKfdwR5n4Y9kPD18oz8gWQWNWAkTV+rrEZtdpjKp3oDZju0lzXCfO
7a/g2ChabqE8sqRa+YNQ8lj8kcsvNMmHXMDTgcV0+Hfpalw5l787igIFVfjR3nYk
jo9R38oK4QeC8y1WussbrDn26QMOfujs5MO1Q39zzYaIkoZQbqDYQEd/TYyshUcx
iXEsKE/Yl0/1FjWVU8MUDzgyK6dLX4LquEF075NlbujYotUu/BTsDFSs1kgOQvrG
2disOzbLtaO4tIJyzquBA8KuBrtiq9cx/APOT7tbsPFAuFL4b+rxOE/njhwtrwKS
ebZpIOjL2LgXQzP3kIkjTgeuA0hZOKL+yxWB6XAuqLuZqEqB72iH7pKujXAjmDpw
rUM8M3bsCJSTO4GfVYshXykx6PeKslcvZvFnhA1W6bRMIBZSCwnNjKS1WDX+v3/4
yNP+1ixlaZ8uM6sGJEXMPuIzalEH+9cTvSM4Og3btdpw+iaNdCoqp/cBLfhi/ftw
XzYEq33UKVbqMi+esvZtMcKDaqtdLKzKS4757IOF9MN581aQsJBnlQLhXe6zj/Pf
XIEmqalUFsRbX28nDWb2PivrHdC3IleXXp4h7Ov4CHaIDcfrilXBRYbVwIig7k4P
yctHmMRjcH30WfToOIEpGDJlJaR2ogHaB1+u+rAI8PvTI14co3s7TKr4qRp9NrdB
ZldiIHjCgkHKjVELLH5GQiTY90LgAwRnLverFnwCU3sW5JIWrSUys9/HXMF5zG7D
+H1eju2eMdbhJi1WZeS6ULd7WQQVaGrpXGAzTtU8ehV8b3v3skeJsEycbl829G9G
cVunDNIhB10XrmW/m5R5KDXzx3rWbX3Wz5DyOR9cyhdb8TarXtn8TxdNLPDTwkb4
yOwJSDu7oNN22xDKUSUjV7buy/dhs73wrn3KmHpOwbaEpp43LVXz02lNHRsosAyl
GvtQ+u4LPfHXHH5K02t43auiB1VwnDyANXouuTkM0QYUG692zSzivhFcapoa3AmA
l9TVgOQQ6LV1xsxAAX5M5PALjN+t5Sq/2cpiIElkwLmd4COW0j5SL3+67Hi4Jezd
cLuDNZ7mACZfDpY5egHgr5hlUR+hSQY9UEKdb1hTB36j5pB0lfzwsS3VUZLkFUag
uLNBf24g8EzvtesShHwU07jhqat2Vyxq3o+ANrea6fDOtg1/0lZW1YNhVkQBAMl+
usZFzj7qPYPKtVjjVC5wqMxOJX6UZnW/0SGnKlu3a3msDfyRALFT8bqok24BUgd3
BGsgUvIQEpaP9ObzpblAWzwwQE/liJuO2xPKRxKqja3nkXSJZZfWd0N3Ey3NOJzv
mEw5fEDYKmPFJGPdyfZ7AccCtob/GdLWvdYPLt12lVb+q4TV4YrjzRVoBSDF65Aq
3d6QqqBWCsKTBB0i/2fj+K2mMMDVn8WOFnOlq0zSb/08ubHSmhC09txIis5bap5t
UsUP3o7G0kxo9FXF7NTZdQFV5djMqs1q9Y6WBN8boWxhmtIS4cEm88jE0jNFl+nS
WlGUQpp8qcFTPne+6HoRTRSN/TYdA7SkO5UqdGwgAFePpFSxWdvjN3VVTpmCBXPk
I6l34TxxwR2vFEkDlOJFLDNgkSsB51A/eS5dzZ4FcyDaukmZBPSnjsrp1vejZALf
r/Cr3niU05Lvh8dao6iY/Ayjj6JftztaqfjCw1e3TGO3q5WYWhSKs31ce3OwfmE5
qXh4h9dtLXVn6HiUTse+4lP7Nje6MWqOzeioybl9YhpgiNgHmasoW3LO3S+u1Jhj
UUABXFUEz6v5aUGFm58A47W3gGiZZ6zZkWTiumGDcRwUamtCExkWApDAotTLIDv5
N/w4zEGxt/bNjwWBw99Spr4omW8f/zjAfWyUXpNUmi5AY+dtdeSfPLAlF67vM9x4
Ws22oKm/uaKdjHEXKtiRxDhAgsADlDrBfbcg0Xk8p0/XyfcQLtwMkjGNa0APjSrw
8RTnK9/xymiCqZhyK38Ed/xhUYoGAOixbR1ZTm4KY+8enMgicxKjeJa7jsTaX2Ey
EfUDvpvNGlFjrfsA6dLvb/NN2IYK2ylSD1UQJzqT/fACvt3n1+mTNc7PIsAU94kn
Hw6LxdcPM51TWhcQLHCDuoow3Zu+VLlxg+k8j5sag5nGGMQamxUgTXTictu/JkMS
aiCUWXVwhglFlFmAbufzKKBCIm5WAGyFXlCYiYk9Y+Hi9Y+Rijf6vvE5JLoNbPgY
kc+WkiZWo6HmxmVHaSXpEBiZZ6UVB7Uo369AZX5CZoD67AERE+1x2jkQBCJL88nI
GXB/OBH+rbp2BTrrGfncIcDvxNAO898k0HiUZTZSmIgfHmXs//M4lf2wZcmyscnh
2tsgjaDBFdSS8F9QFljAOdMvWWVb5AmpS68A0yh/nGYZxo6ZQcY94Bm+eXj9JLgw
sUC2iM+d3FhfZ6ddGIZUrd+9nxie7E/orSm/KKacBcH7FkDmko4ojKIRC3sbpLjD
0HxKMYrxkynP/HJdxbvcEWAx/9NW1h+nlgndHPKW0Cl02y173YXZnyu4kK0pQbrG
hpLkY1cYWYofVBGZr0k9ceoiufIA5ZzpuO+1QkC+fZM=
`protect END_PROTECTED
