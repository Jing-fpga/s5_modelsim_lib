`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1mgpds/pIkf7Up7AylKdKuk8kjFUCuUswmHYHBF91V0zXe8kOaEIyH2UvIbTI2sN
+GsjBnd3WiZKwGHkTv98WBJ0wPniBHyECNpwi4cf2l4EIfipDOy3ZbTeYZOxfR+P
OK7JUmR1weNelIyKb9JfrlxJ3JkkM/aSgon41JsxdoKq/4YDXyRzpD5WEKdW/IaX
Pg08WDbBW9xampXWkVGwDMH36AMzrkH76hkYS9z/XLhC55TS++H+tC+Xucx2sNyY
0SXeowfGvVAilDXtkKVk7m5ePl5WHyTgfdIjlvMVxjs8Ha5xVOtbqg822JFiPzB2
KCm5wYeqRiKhhd6h3CnVaYZCIeoK8AZcf2yD7Ee2Uw2rx3ht1JpaKxSuf/08d2gL
vqsNqvLOF7qjv6gQSj9CaN03+p0uSPUxpN3vJm8AZvlaWgzHhzc5csR0vAvVSo9o
zdnxafFHJya79c3DtZWWP/YzEVqmvMeNu0TShAyLweauxO+4FfXJpphfBIUbn9W5
r5UVVu7KfrFDgL7pN39S+66dS73Jvgq6E6cHMbirTyQzrmK7mPIYXBrPI2InOC63
cJU+nHleEsU6CiNwgZ7ysCC6LcNGzgJCHPkVgFTkLeIlpjjx42desfh1z84Md6KH
afl9eVrYH6nUR4a/Ml294b2EkF/vgg+fBCzpP3EBJzl4euju0UTipwrUWaOje52B
5jyShADKTzABju7iaY+iUFPRaiQKZaC4ysS/sNRLiPnVIZAQB++7uxEBNsClgCqn
nzonj9W0VDp8W8hVmSqGZuaUuWwwn9242Tlzoq2QL+7Xbt1aq+sMSOFA+Ll836pI
cxixkEhzcpHidhIs5OqdroBPKjVfLaNmGz6rO2qI075LzlYtI7i6c5ta1HI2I7LV
hUkzUUrPT88kyrQEitbo4v5zBO8nteXSJsS98Jxil+Hvs7yylZloDZl3287HIb63
cT0AFkda6H6dpiP6j5gUHiqXfr8brr2wPLeCZjumEAQAzmal0RrAmo2V6Wujnfbq
`protect END_PROTECTED
