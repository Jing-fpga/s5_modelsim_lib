`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Elfoxfu8h3S1U7n0zUtD6TICpvZtBm3/Cpl8wZ3XDZG9uOMbP9sVkstpKguTp14G
qNQGU/jli6PVIV/SEJtnslRsRDkEvvl4045FlRX9G3NF8WTZaev0IcYATBKCSC0W
LcQsgPcPFtdd5PnSAo6+WHleOCIZyoJLQ5+zwHh3TurtNyNj5hjcrzcJK0nYYhdz
0suiynADBtP3NqiTmzQMtBKeTUUVM3JStuR7dSob6t/ioL7073qWcvwnHE6dRKNW
fUqZCUd6F41bEC7Gl18Fef0gthiLU2Dyp2HCtSRpHsc0+I02FMDjB0aerOoYnjhL
y87skPM2qnKZtDR2OnquBvo7xR7G8uqHbxE6HN1QH4E/Uvi///fCu4h5kpE49wLO
mO47R2FZPkBgGG32c4yMu2X05EH8SCGrgGSyRBVQabn5um92igNGwut5mlIazqvM
+gSnp/i7COF3m1hZHgSqXnj16GRJrpOGURW2+WwIjnmaUK8LFpqoFJ5YCO6PIlDR
qgl7yH4GadQAxcjQuEiae/qJ8q9CAI3zOOfijI4/8OPcdiOO8HB+V2CenrV2ik6r
6an1tSO+0sgkXcaQYxoSMDp6eabYvOj6o5t8I/MyqneHIWtMkZvC4FfFWRRaZf33
mLkRemR2ZtCE3UAE/Vxg8KYFgWUeAduY1KAEjoEbr9qk54Mo75d8PYoCR6Fo+weI
bCy+17nju3gkJJ1zwx92ZBN/VPN3xxcPjSDWGnZ8BZMFo/Sc3BughHU5uYd7SAHd
fViYLgvpjRfN3pro6Vi+yyVIG1PJ0cs5O1YRGP4ulvp/LyBJXVD6+8x7GiRktzo8
tMLCC+nYKDkufOvwyIwITL9hdVhNkg31Q2m59CcmACCYf5aAbbbwdtnAcmyeQbEH
QnOMQPfHSAcpclyfR8S62RA4Ms0UVFBv2o0pbjqKzSs3Mcw2wD4ZJPU048EnMlDW
/tSlnEw3CqtD0w30WNJ/8A0Ujt2WxYmYMbYJuCvrHquXK/QTxRfCNpg5pXePLgd/
3W99PoG2Z6sWqSDxHlczNyz6i4fsmaE/JlG0dClqq/F+VPNmmYW4VV6XTlye4oTt
4W6ZCSuJ0i3GYEES8qPewCPzYQ+Wu7SoRyO6xaS9BsDaXkjKlq8UL+BgTwcMP9UZ
VTWFsQaXSeIWidMFfsKebkxh1wW/PNvfPGVW/l9I8uHs73IrcIp+mt8RklftWWqH
9WLIr89bK/k2JUkDpGx2PdSF1G+TeDhHEtuJ7mEZ/uvGYlVYRxGPMoeyNZIpC1No
j89vfaPREJen4W7yyK6BR/gimz2fjhLKyT4EIcuRLy1/wKRe+uztjFttrGRJh2gO
oOYLNR3UP5l+N8xU0/ZKDFJG7WziPZL+96FClcsJPOdCkbow8u3qHWX9AVXxqbzt
xny6XU/TedwphlZqnhM/+T5LpvH4f+EinHBJsjMes7VuJHjvZBAwfU6FNQcMMWnf
n88VG7YcxMgVU7aGAWbY933xHfjsL7B3nLBnIFdt5ybNwErboqdF7fTLbPPNDmHT
I+H51yNnbOjz7ACMgsIgft8a69Jv9BulJXcTq0JP/xRZp5GDQ06cESdp5SmtYc5E
y+lOM2UG9hFoFama7JfNrUl4p44Cgi3j5LDqAX32iAi7GT39sQje5b4dnJdPXM5K
rUxxTa2NjqsyJiDgijWut8ow20up7aAe89SE1zq/XQDTeMGZkNRiRsqdRICcrHJD
aEA2YtpMiR/D7Af61RvwyGigOk8fCsfHrqYrzkg2l1Of1eeM+RoYi/MxYgU9xb0C
J5x8jPdGs9JFzX4J94ZP29jLzuowXev6x1n0LYTk/n84V9rypcXlrnXnFdRe9emr
vyD2kixVC2MYRoRnhVAFgyBk4QBUkriHv02MI6j6vOEmH2UzAAV59NywPgoNFcz1
+ahcIZ3Y1PT1Cg5EDr/AJhXst/uhvubk6vnkeXwU5Fi/fho2+VAidg7i0guAkJt/
k28f1Los9oLeei+8TyF2GysHo8Cgmd9nfPT5jE7pdqwQ5U7izmn0qBapJ/FholS3
JFJyF2Qea40xrtMuwvOeOmMgyLsIdceOF/yomo0HOq/7P4VgJTovRHt5ZcuTcmgt
p8dfcJmbqHmLJmEnOIWYrHikyCZkSS/cdcuR2kX0ozizI2/pjQW+XodxEOGDRFhw
lVcZMzg4g/P9+WnmzTU90YRmZv4zD4IXTKy9fWLxDyQD/3wyxtJCXm/GA6E9CC30
+ZhnD7Hn9ZLxtACjnvz7Z5XdomoK3qJDEArqALI4j355x5j1RebLw2b8B1hAn5nG
sxVYwpAaO86uBFfMgnvkyKosEWpmQqA42YDP7GnykurjD7jWiOV/ubFfDyhp2liU
iSZhfzrj7Octr1gs9blUCpv/jDCod/ns3oncs1hAAXAA0mbMs8I8G2WovU+SJHbK
gcU8NYAosyFacHmHVbOvTPT4v2zsvoZesx5pcNSFLtgSIocMCjjYLf+7ZdDEu+hE
RgEMS+z6eZdPmIRgJP4BlDVSmnCbZY5hWdekv/3iRtnZXN75JGBRk0vMUFgupzdL
qav0S6Gb4fLs+yE9v3+5Sum9BrGwZjkzA+Xzb9WLFkEAZ/gg0RrheDTxySye2oW3
mucrwVFw0iSborq6foBWS9CFa88ppeyvHgr8cW9Gw/eAFI2QOuaCmDem6yiAzxmp
xy+EXK3y/Sl3d/xzw2+L/FLCVhO+LPTDgzzi6YIavI714rIb8HcvJl2iNSxwpNvt
WzYlscwFZ+Ib4acKMU+uva1oGulsrZQpd6ktbw7I8aY0WfySwaHVXp5uOzJHTxw4
cyeSHKpCnfejkZem0aCuK1pZOlpE5Zub+lozdz6XBE4Har2ef/ZMCXHautOQ21eQ
VOsa6eqSs9FpD297sQTmJcaGl5kqtweUIlrb6UsQB0K107mAifCYSLcOGWWf698l
NmH7jfzJUWwIiYtL37oQ00H/JJlbxOAgq3cCIIbJgBNS/F+c43ZwC31tHamyJJZ/
OL1m+guww4Ai7CBJbUJ5GQBGFC8Id2SiL4XTrpPyYf8lZIFYYFe4XykPn3dDZGPQ
h3F558Ueuqlk2hRPrE5t7dR6VMaC5apjpWqYqhnsj28ogKR2qVQ3gLIoLIgyHbDE
QKq2ToTDh7aHlDckqhQm4617eLXh3wbLXaKXx8kTitkqJFyDVHq0daTT48Pk08uE
YaFgSxkqBwwLSbA9Qaw1oySZ1yR04jZ6wDSlIfoLENQIHFflXicqEgzKv2sJF6hb
7mjb/4ovarxmzqmRgb0PfxQwDODiTd0+bknl3KTcj7hBfig4yrciTPd8oRWDQMBG
a71TOJvcEDRk7zyiPq1wF11a31tgv8vdpnbZLNh7wb6bQ3jEk2bwFhZoHTmr4CNA
jDs55yMLBfChV4JShMZHaupLqGUKS04WZgWj/obvCscThfsG8pHwZZHp7wVC0Adv
ma0DKC4NHoM6wftFqUzf8eJJSdfmhF+NS5jmMVGiBf/csdnBa5Wpmq2Ku36VlaEN
WsdFJ2eG3VxymdJJl/KJqbmVC6fXJxBEJTqQASAdTqFQWsjWbakRISdn1wFMrpTj
WbfgWZP2FXNvty7yheDtzuiz0ioP5GOIJJxcUYDTYqGXFLPkeKS0z9Szmp14nwM0
WFW6HKiTecLQh06stsAvTpAka5y0Saig/behy+sAR6k1oPA4BRKHwwYffqAFlov1
ehp6hBHEbZ9lKcMwATfK2WwL7VDAatMJ6sQ6PSSpR8mkKdAbr32gvhRt18wQfdNw
cAKum5hRIpmHVS7Xi16CzDcRzXqT0R3mybr4pJ527S1mJoCnfe1BTK9YIxeuxI18
t1vyZ+Yzgzqeh7Jpjsq1Wr85mfJKtQ/xvljRpkpCJnsKZGDM7c4QAUC+uF2Azoc6
DG/VTmq4N7RliXnZUcof+J1Ss7Y0plcSxSWlHhRkUpqV3/0mUzA9CkbzgaZzJZTK
o6RV61/j61UkWwVQ/EvybKZHmtVxYuwkhiPXpgaeP1sgiRtkZ85L9KwFuyKffcG6
TxRgqVa2DUwLynC8n3rxrTzwaoLY9qMyT7Ox1nhzNwzoDXMAYktWPb8jF2zAQwfX
9aahguF4XH7bHZc5xL9N77bRQWzcfthB4TxVdyixRPdmY7AH3dTrVXtXUmqY5wL9
ncbIylqWqcZgZyOd2zlcUCgGyC7FczFXG8V2e+wQP6LL34VjJMXJGPGNmZ4q1lGt
LDAZQBLyV2OzJti0gDS0VYHxQiENr5L52fwv2HOa84xicwMjY4wSCwZuPpjpqsNa
OHNdgTcvLkFiNLPBBP5v/xg2mZjM5xaSSSMJ6yhJ3U3fCVBMxhjuI8qh/qEmHWhi
H8cRzg1EwqQA+eH7FyfMmcMDHJGkK8VwMaRfKe6pbCayXW+2dA+6g1G+lnHkmu30
i5rREzJwp3CfQoo7yEjqDJG2kNrv/zBV+PzUFtuLzCOH0Fz1bDgOcM2WQMt59I7S
`protect END_PROTECTED
