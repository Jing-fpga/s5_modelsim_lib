`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KNjOVW0JBNINX+Zv1rRETpW8f5v1MtXKduqAAUKcxkqXrP0wmXhqucX0pz0Q92xC
rX8fTcl8rl2VZ+bJ2Rm6ytiXjmiQvd7i6QUpbglJW/1nx008ovMUTBvXUDUGewHW
Di9RWhPwul7GTW25HO3i+XxbtN0zPXy/Re5eJjC49m3DEFbARGiWL1VZPyRqAE3G
aJZWuBpgAMfF4ArG4TZUOZFkG2hMAk0FQISWuh4r/SAS5/MoAiyt3As5A6g32SXx
Mq1OMCShFDpaD34rWretmknY0Yd6sK0J4cGfjrKG45TpKEsgaN1Jk5CYKb6bZ5hV
fCyt8FfOxIqaF9Oq3Cd5Gw1/5gE6uOecA6q8vThocnLllhUSWXled1t4BD4KBFxS
4J6ChqLG73aQshLE0ZVfjOI+MslKpjjUEA+ZPNt009eZ6sm3UIIAgKX3nuaVE6Pu
YdqHUVwszVnCMiY1RFUfDDGjuCvWI0wDDPHW3I5w6CMKBUl0ktJAcb5XmlhP4LFB
dT+cB74PTpNEcdiFqODcRExMuCyxLVWEltw0L6v+aRNBm8lqU/gAeW7fZrdBJhTT
A84Mp8/IsdqbeEfgxUp+GBHmJ2hT27vWyNfto5BQ6Zy4kvfMbxtXwxyYd0Ppuu2M
1HgnVdV4fk3BxQjLSe434u8ab+iaVddiHrEPiGVlCAjIxFUz3LY7y28W/D9Dy1GK
8jQjrI/Mi0aZdrTC6rOacqNeHI05kNvRrvddVorR2NPk8FGZdk7VDeLujghRkcjw
EgLct8ajmr1wUb61uz6v0zLIsANc8HIq7NGvzm3gu3DjZ29LVOXTiIEClUNea7K8
oxM9Sho0N5R1i5Dw6ab8QM8XN2mkdGzhvK2uYjhneEX3mEV87BGAWuFM5px+T4st
S9lBbuI9yfRGqy77x4g0Ql3M+PyCOG67+LwYpabrlkwClP+N55hjPY0Lk4j6L5LF
E+CHiisgdf9jfNTu5Bbt3LcU/YHWcbjNKiCAD1htvLN3T1FfoXTYwnRUaAt4v9gv
CZXamrXYh7A7g5QMWN77gbQNycUU+DcpzOnuHf8x3kgHXI4/kFFh7ek63myivnpj
V50RK3+YhKFiEsoFXy9tOJJ/V89XvNyHWmBTIBHnJw55DjCoAJlZHlak2bobNv7z
ZXTfLTaOIzsN7nysW6K/L2GYn1zvLOsbQi5cu08VtSaSLSN/M83xf1xT9x2wTZ1c
2VORo7HNX7UHJh+57mvS7+iRNtoCHNNpLVFHYhDOjXUazLPxT7gbfBBYq8V96EX8
Fx8xSULALADf+kgzx1FYZzkUk4LXaqbkrMO++5fl85cMRHriW4UH9Z91MYHthqz8
lVygsnzy9QYUmI/xnDqBf3LlGR4QqUZgqJCN3sswcwOnP394XzK1gbgaG4SqfKWb
2qgY6icG7xJUpeb3nrZhrW73gSNPxyEhYFxe9RkkbRXMNjvL+RsY5RiTLgFuSQ7x
gfL8e4nk1x1D2AU9RNq8v6LEgGXb+eLMTEJZ9Xmt8gFJQrUYZbAkeccsH8R+WrCz
X0mDYEpapHGuta4dtT9PjtPG+vR4c837YeMJrG4zqx0sYdncEA42aoYbaNRJQ7tz
Iyn+JJBPDvqehy9v7pnHCUIsIqU3Lj4EDnlVhCvW/OFBjJVzwdkGPY6FrOfWYVnm
TU1HNwc+6T9CjvWBzDmMTcrHIpEunrPKN99EJ9WsXWzL/fU4Vz4Yc0wlIpLb0K0n
z0A9bB/YnJ9osuJ+BJAWVTGyyDLqkREexVXbzvkfay0OVrWWuVCmfc06YIcGy27f
t1UiMKzLa0z36TBwzGamc/53eUz0oh1U9CMdPSSmAbYQ1scGGMdmONZYfwk2uNfS
07oQA7uWOO+q4bJxTv5h5zh4WVM8tFvauCsExHykTNe1S+BCGyWTG087MkMaeFRu
bqOm+B4iziaMmH+sRa/SddWqZbh+L14zXxZiGs5YnPAsLdfAQ9UkZ6bBL9uo37Wg
25fVjOG+xZJgz0JSx/ZjQNgAIPZz55GFtSunQTf0deRxvx2P0CJ5t4XW9H1yUKAI
2l8LbiGYUFmKDzeGixsqk78XDwXcl1NhCaFaKJq83PYvUiJKtjBeXwvKDac0rldo
v9ZtkoaFxHKe6wR9kwwqy24bjeI63OxNePpYAUXqJGyE0N1vm0e+jUhHF8AabnU+
p6IZUfnUoQH9idikPXIdNV2WrfaWxGTTuQ9mO3JL9KSAMmeqq00Oh3/U4TnpzaKT
7H5odNU15pAeSbrosdNeZUGFJBRK/MNxaVAkczyu0Ryxrv+8KO73nxw2OzaSpvGn
sqlLEKre2l26Khs7hHGIijWHE7kDW2V7NQEiEh3alW5w73waSYcShOVTIDdUu2gG
sZ218sOUyHAjauugX/ux7g5YmjlPtggA9yfoNITWQ0TMCy4r95deZ4zpAneFw3i2
AdGZnD2VcX2yu5zw9IgJ88NeKkcaRkhtO2e8rWlJ4zbFSvmgE70cAzdq8nUSF98z
n1LNYYwGH06wV3RPH+epPi/M43V/VOpOiJhC3G7UikZO/nrFWA3IDKZ0lFG/NENw
aHFuTEWOFtseDeBd/W+j7xqmtMy+x3Xysn1pqH/8hGkiwNKQWxHIgL2Wsegl1k6i
blIu9ycP9sp9BUOCmp3787zIcDZ+2X1SC+Jm5+EAkMKhUHC9uxJX1lvAlLBVez1U
Cz+oIO+2M22R2iSeVn1pG7lcGU8M301nR256VRtcOOVTonlaD/OhkN/u+Ft9NBjI
fkLaElqjt/lkLNGyDKjfgpimnn4COc6oT0lCXkEMfDGZpjhUjhSYVLcG3E5pOXod
E1l8llMKXkQwNuzMN5rOlEfJL2I9Bu3+VptxOOfvMoYbXJ8tVlpxRq6hW++aRgxf
inng+i8b06g9J6CJKBPa4+CtGhHZfEwmsEA7RqiqcqUZ+ExAdMbWurKs/ezg8FEy
R0SkTbCHc7fm45hOpgji+6QxmuGWK8EIY76o2mAtR8ab2BCFPklNSBD+/GMwZGDd
obiuQzH2WmhW9pNf8JMmFMh2eInALRqMmJ0dYG0MfrEGJmUdAGySzqA5T9lSmcGq
ViVMZV9px6vHF2LmhFIi/bUhMe1Z/sCQ8Rb0iPcw88j3Vd78aCWKEbyGnLrLLgGx
Uop+oC2a1XCOsgwPAoieJrscETnU9Ii4vbGr3wmVrWPhWQEHchPLaCcTOKpKxnA5
`protect END_PROTECTED
