`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0k8jk+6Q7ybaNqgZzAPPR5I5lC1pNW++f52D8P4HlYlTN5GQA5TvoTZ4LwK7qPUf
YzZNIDXwCHtWi/B9pWvusTi2uVi84RE0dGTaJfk+/3i9JquAuamf2WmeBTg1vcm2
mcxxn1IgK3cban4TPKy5F3cS6VC9y9ugOTJXZ+xt72bhtQttiDPUQdHAm5D9InUh
GH0zOYGPlyt3K5D0+PhPDt9SrxTZOlC/t3VurNgD6I72OtqD5htXY6C1pwPQAqwp
qmW16Il0DChB5J8dQUa8jMUuDkYRuNXE7YOZ6tCCLu+JJTjq8kWUgJv+/2YmZuQE
OQZ8pjCLVwgZL1lr2ID7qrb32sMP2i9niAxBUcEWCQovFOaxMsTn0/hEmIpoTIo5
9KJoWLWXUnPLre/Y8MDX+CzDMjtZtLf4xVNMh2x55Si74m2hwQSOc5hwjNe+dKqV
cBzVI+pEgucJG7ZWzdr5XZF2s77SnrQQhgLvZ96EuGkVU7UNtNVYuphunDuqB58U
tgvbm79k4ytubHfjxuEoEKs8u4rwlxwC6SB+LOgp54lBn0Us9yaBbA9rs1hPr/s0
/yLHUDGDtnrbbMPsKwYpKO9P9bYR8/bm3h2+1xsgVVWfY9ux+ukV5ttTF8+cp/3y
dValNuMh9puEVOXb3fXmPbrA6foHzDrUqxc+fDYHIs2SJFfsFvij5efBdYMTrJzT
2hg846udrKxKIpp9Q+JNHArrr5OzK66n0Sdpb3XVq7ehT0cgFwudfOWHyqIxky1H
HCDUgnc3NRfseeQq8zwufi/M3ooo8FnrWxouAFgPIOFa6SXcCk8kK/79f9Slc2CU
a67jeuaz7NBjRHDS+8GQn2rL4XOr4O4SdufApDkxdna/rVyf3mpV5eDZ7Sv1kztS
gdVMB9j8FIGmpKA2biVJcCApjjMYYqQkqQSRbM7T2ymdM+wU7S9APqoOaYSBt6me
rgTCF3/4hpqdvbFyUCNPFxpoRQOJ1X7pbRF2aXbotzbTNuPTdmum0Phb5BvBb0WR
DwdosumRlsYYRAhF9qDCpvuiaoWtXNrVb0QElv3/Fe1PRchIG9eeexvM+5Tvhruy
d33Q4RjaKopwm1NHb7T3oSc2EDlddcGxZu20JSIRB6XYuRfzFsBTwgEGMpRCFOG3
rNq1s+YJzx0Kh4kNK2AZYmNCz2SrW5mpi5NaOISQe4KxUnXy9Cz5WNaRU+B5/jsE
V+vWqvkPyKtG/WtnT1MDFpSsL+ozb33c/5vcLS8qMKlt8VROoIj09wUO1PSuSbHm
6mcam+G6JqhJagAe5Loods1uNCN3bfvWybZCxe2HKkSMfpm2CPxIqJGGQvwJC9bh
PbqAyiAiFBAmQinEZSOkcVjAPMGewScHyqMkqMs3CnbnyAsUjROYZctscyIi2Zgy
IsOhW8Le4Pp5jw8o5qQfqkx9T0p7GD9GGECh64s1MEPjW1BTJInkf5nYmfTNZDwZ
b+EOIfc+oJCKfVlUOCXJrMyn7PAvPXrULLiFzIHUZbGoj8Qf/aXNuPya5rAeJfKa
A1WJxXWWkzCtp1YraWKyKhfSYrms76NBO/x8iVCc8MYD722JskvJX+0IR9GdMSbQ
dGbWUiZ61UrFHHxiwgm1ezWissB+vYP9KoeocHxiK6D3NDOouuXOziUTqwTStA1n
zxtnxJ1ye2QjvM3bDN9oSOBC52eOSCdl5ac5790h2lTlG3AoCvQIn10WB3xRqq2d
ghomCyvNexfCFVeJuCZxLe+LIDYpCWnrVTe4TEge/oTwRqoin5RTU6NZalK0fLtR
Rjw7WpKmNp8y1/Xy+AHoi4JoXRJwEviIoHqh1Z8bTgiawr2iA3rsAVx8Dw/jD79N
jMbl3p8EeSYA2+wW+mQ6iYdMarDLyPmLw/PnloGPcsHYIakSckD03StWPx+8W7d7
MI68I7Hq6hD25zuUUGb9/aiVoWptdKE7yv0W/XD+tUZDZ2p/i3QGfHRDR/X0o7Id
WoGsf6LDlicIchRFJ7pWzXyI2XnK2nefHuJ8Dpqm/QteMjG38/ZDeIfkoESyXB/V
hvDIxiEKGCnkC7tXhEHoLl97GiWqlljEf+5QmmIsHNVUH3OJeAbIapq4A+H9EmT9
GwlteMXeDR3ikRGIA61yco+Gekd1uj20kx67nd6U9mMsAD3AZgRF49rsYI1jCpNe
QjY94L7RD5buKuq2kF9SlYGN/Ho3Jd1UftppBUFNp/vUeDJKyKHtk3e72odI4Z3j
8A/L5iQ4ferO2JBYcMDw8FTvk4vx04qTPUQwR5UZD7eUgOzUGOLSTwQSDDamDaPD
lV+N8WFfoTYB6VRlY/i6uoRVeIYF/SdFnyKaUiZP1I6evt9VQk1qx+bbyeTECMx+
XoP1UehBmgNCYo4qmOIFiSgsJfI7r9qb4ksVWxhH8GA4aIjYi6By0jXDzoO8/wn5
LyhKqiIGwh54okmPFemcvMWyWUbGOlsO7PZVBQkfhfIo7IrWtORhqOL8lhJk67Wo
22IPlYHpg2H4+TO4RxkGkXyH2Pfijki7hAwBLT5SH+w+RSRF2Gow/pWISOLYoqdW
hlz+btTGMvAYD87D7nWxcZpWODuu6KgDHoYxAMsgD9/zGhhOTJhWdszPgFk59QLr
KMlvK7mVOogHe0PGj6NNN41H/96jK8FVYQJ2OhUvI8X0jyU/W12x88wciN8zFrRu
d9V/Q95ArQCnt+LxXFGSrLr6Lpfa9wrLGlsO9qFVZQfPsoFpSxOTpXq/LFhNPvgk
hUZ70U3e17OfSU3PrAaSWyaS80F8/AfeCJwJujbIt3lTs/EB2Q2cK18yonO7QMpc
HzHdqMqoS9fwCMuYGJkvmLPSzdDX8Btss1g2ddNx/+buPOQGakBNYO13AyqGsWai
Uf9qDNGtJHm6c/hGDDNbjJXtN3xWej4neXr0j0PbM/Qpb3PNuQAu6dWScbr8Pz8R
zyDC3dRAIbcomZRjib/98FCN+2jJ8iQ9luidIGVyqQXy9IGgdyKW5tVJMT2jCL0p
1XvbrYMtqly+Qe9CGwIXBjQ/v9iH66eu8VPw8o6X0S95NM+03UAydTKbXFJlPAny
CYtKza+IC0z8IktGc4NP2bsKLxJxUCy3OZeHaW5FgSnCwz0zwxsnUkIdgbW8a7nd
6g33ZBugaFkzmHBe411fddlXmd2XAA/FgRi+j1IjOyY7vORT/IRAwN0A1q6uuaCl
xUwE3CyoPQIVJasKuCNL2mbsKGHBfPIaEk1Q8FBDt3P6avoKmNptXXe1EFZuzm6H
fMFpIK7ythacBHgRSO8sGKPCEl+aT/knltjcu7EBVVkuRd41kxvrznuvDY4Q/SNV
pRS/eAxGxgQbTQ3P7B8kOfA7E2s18c5x6JTx8b1sZ5LJJ24MnQVlo8nng7HszX7F
StXOh26DX7/NEF2y0ucnwQ0qBLNzDmrZTCOzaIJozXl43RO8YNOapwRZRNpOoEI9
AYpE5dAxEVCzX3gjx361pVDHbpxpStV0TuYhUyzqOLAopa6sf4/D/oAEPfwBlIAE
w5RpFM6zKrgEwoNhDtTOjJV9oCJ7XYqBffU/QBpTpss+DDJMskxzHwg2wHhPAOMW
QJbIp4HYpJ29kizLExGV8KTlSASTdN4UlbAtqmFAKzDYV0KwWKGeIYM9O7jpWKjS
8S7/KfrQSDXGiaZQ4Thj3orQsb6YafhO/pl/ACqOS45/YWEQltJuhEIHb3Gt9JJ9
DnTnuYzQ7lYsBh3GS0jTvTkq20px/Yg6RFGyI8H1yVZH8RKCPnythtGaUu6VdLjW
C+wjNQDiHCK/V2pIDzouVc8lPJM2ch3MDgsHrqrKuedV8/zARCnOD+YAA4k+uOoQ
oWpV5DGyR4X4DlbM4LlTyjsOLPeTrGt5bsGGoUN+MIxC4iWzAh4gqzLmq2LpPYGg
OXvX+s18dUWO+vipraXAmGXKDCUO+/X6sp77AccwYT3tQ+b1Fd9lQ+Z8bIIJMYmm
0Kl5m2ehN+V4VT+u9YKDL8KXUoZ44ZjxDh8wVBgYwH2wUll8UYwQ94WFW7z0hsjZ
HVRZ4sTrta3R5oswTG1x812FNRntr0mAkWaqgco16YE=
`protect END_PROTECTED
