`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DZSQ5gNZr/y47bypG5ghiKvgH/YMuGAtHzPgPRkDRuiKKxBv5A97dKE0R1kYAvUV
i7Ia0ROwcCkdd/QWAFC8e0DpUUdGst9sqPQ8oZkq/PaIHtiJcjZUyeVdS81A2+Ns
SuE2kjKwMtckr4EzPLXrdp5FjhUk/yV4bjSFL8/kMfq8TxrDSfGV1oUi6GbzvCjy
dERtlyHO/RbxRWBJuSFYRW8mckFGVzvuI7XBiBj1pXk2AO1RCgpzrkSaWbNY6ddh
jvGjq9mQqLzAQfbittNvUqJ0vqFzBtHpYLT9klO9iNiLmRFT4Rp5NLW1igY/p63L
TmkoPWlod1cP0E9n6N9tReyAeDGLt294xTCtkIOFdL+KZeIQ6u1jR4L4Mk2kQJty
qsoNo9rFkavXB05r+iQjdagN3u2kGmtJrg3P4LwrY7AR2Qarb3bt5ec9lmAuIkLM
xx1aHlA+AEwlz1Gt5ZlSeqyB0otQxPfID0RG6BU3Y/chyGGPr7KvRTcqU0m6OYL1
xrrgmLb1Hl6qJ5jTAtleXr/JhgeX/kEoq/6dBgWwpENEiL53DL9InI4bG4IwEc5W
PqGVIK9pmGw+EQsTQk0bEwyKNJJfXcs1Mwbo6v7luwccwZAqPeRQnLritNnYGmCD
qITSSy3wgNvXZdd167E6mQMoEgLrZbZkkNC61P5So4TbYT5YZ289UNUxOxVS90gX
6A3sAFIeo5Bf1mk9e3B09tp95fqUTO6P9QDuseBotR94RtNbcI+g7hfM6Cq8Bdvo
ihlQwuuk4pB0Czl1fKnSId5KKivu2aPu3OM7Cyf/WcOPI9srtAm+Nu0rlg7h+ZRn
BG37atLrjIXTkTCjjxRfc9MfW4vUwx5J3Jo2+v+79aiuecyQliAh04I2Tc16h/UH
CWCZznZR91CgO4cA8rHTHKImFNnq3lB7PisBr85UYC+NybFGGYEBjBZa8CT3KY6D
htEw8UqnsiCBhe7iSDl6nO+AvWflpU6YA3KvFbUZTy/W1dkjqUlpGfGMyGBHc6ny
r8GRuLwlHpce3O94XgvWltYmeIChg/Es65ZoYJN4Ve0J8krs/KxGiYCKnZ/+Q1fs
//F3rn6T5TXfIMueaWM9b7PwBWWF6ZAx/EdOq7Pglbf1XH5NoYr3NV0aIm3dgH5A
iTD3GERa+j5IwnEoMRWy02Tg7c7rZDVtG3gc2yhhBy+KqlG1lLfF4AE3MoZZUsIW
9zLK8TAsOM8NRhfydPSPRHyYGMogMmF9Ktfz95BShjhgr73cZ/h9uObtFq7uK+ef
CrEOXOx0YGgneRBnEd8WHkg1GWwR91Z1dgf/PcJOZ/t0aEEX0vosGFr9uxcb4Cw8
u0mmwt1o2QRlD2C7n5y2YumtUBAZcQhx1f4Bxyam3tQwC2gfU7I0Qs+AtK6jcpUe
p4E8k6i/wcv4oh14YMBfHH6svbpC6xrZK69780WZnzc5WW5Mxt1Vj8Y/hY33cSK5
u8B/tcJYmuDNqEwyoHPFCG80kxaCNJZ4br1IHMDd0dFof0jzFgL06cbWCFsC2N/L
rnEIGPSCYmEe3KE6STuKjTDCdsHq7FJnQNuVPmOEL6JaWStW7dEtfEvMR+tJqtez
NfZkhbLbn540Tr8zrxj5gFcT/q7b1uQAtRS09RS1bUhNJkUpy4sdsUnyoM3EZmiJ
9/3gPmQfDZDql+kWMwXFdxGUIp+8Vcr7Odqalj7s7m7u+cYvkyfdC00bgDPO2Uv3
AEpMiMG3NJLWAaPX60GBYyZh1X0k//6KI5obkYh3oaQ3bRKnWW2hLrU6+qzBNc1Q
0Dz6x1BQ1rvZFioj0WcGF+tFutA8BcPFHPFt6gptpRT2z//zT1Bbm6YGgXGkYTTk
NbJ42asm6gZsqJ2pcZtiTS4e4tWzQR2qHOy+b1yPwswfmKgEa9z29C4qj4G7xZJQ
alvTZecFUw4CmSrZ/Evmh9YVi/UZGo0feqn/nU3BaFtcD839xDEWxQE8De549mF6
G93udglrKbSQzzlp5QTPJSTHbPfKoM/Etwx7CgEaiXhfBF+FLihGG2Ke440geZQk
Vji8k6+//9vAgurflsSe1TkL4oVAR7o2qljQqbf1oyNOYh4rsRqBe+qoX2g4EbYb
4W7I9ooNWo5/MsABivut4e1EFGWGnrz53FmdhkIXmAPdrzQRnhLlGiVDK0zIIWjj
GdOgqIilNMI1I1oiMI+UnqdE32tjjMEjF57XK/R2kLyQraOoHONLyI9N/d0wm/94
wPxkGaOnK79dW6J3aIpAWZM+OIy9YgVqBknQD7ub8REIUTLbu3zdMPZp6yxsAVH2
1vRSSGZNTaY+T6WwIs9kpt1Rts4DLFgPZ84+RD5DP/VNv48I6kgSNdOQJAHW2Wlo
pRTOwKrFQ87qdakXnurSwbfgI1cDwvu6RXsZH9gVDWhsZDN+FvJokdyiSpj3vdWC
JtCbrkmDnvfd2hROITubVv7VXIC/nd8h74m2at/zgadHfE6IG/0Ye0ThNLjvE+ot
6s8vYlI02fhLPEqnGAhWHlI7ArLUBD8igsScx+yG8OtYsGBWL4ykW18s0gIkVyZM
lXPNbikgusZJHiJLXJ4ZNjMoq8cq3ea5YZm+gNAsam2cXHWRVscHzW8wsrAxE+NJ
qEH7X3BhtepsqOCkHnO+S4ONgt1vcateobdlN4TbMcPGXGWCiowc88z2FL7Wk+0c
kFKmMV2rMduX+rrMiC17H6TgJBbdJFpaJgcppHWhw6igPIVAnIfCqzCRgqMz9cxk
380P3PEHZsWCW9I13jDvcM2MGV37CUNgjsR7ySSsagqEQg+hhgPKF3jtm1i4h0Js
Nbbo29l/31udf5jmpiBqe7sp0qntHNTHyNzuLbeOtn9XYTx1FrP4lRSvo4rA1IgG
ul379pqvEqU7747tm+H5PHPcgp+VywGahdXMv13KUASZBknBk4jHsIMG1EA6iw+7
YgSpfQaHpj2utN+oMbR9eEPmkimAoxRBLoXaK0jxCZMTWQ82nsiHFZliemsw6Nj9
hR1P2Yd9KxdNRw4ZLVtdalWhaiJ4PUGXVZvos2GNO5XuGm4J78eVWpam5zNMdUKJ
R+xDaTAQg/rijuP9f6HOMxXiNmSK4S446e855WjC/af/K6iA50NwLVl1Z5m/98qb
7Bkus5QL5Z8Yg3fcXGzot99tkbi4x1Gc8Khfb44OWcGeXZpd+7702Cs3yQ/yFeNU
AxIBLm13wJOxgelZ/A8Nhqx9STbAD8urvr5B0c1CrUO+EisZ8okjMV93Js6hydKe
6FfCX56bE75GUSFfWhquLrlpVFJJoTTyIbbofisHX2hOJcm3L6oOAKbdWTo435u1
aukmWuqgiA5KKC6lEIjNR8I6LRj2mFsC158dM3pdKOr9H/U979IyREttXP2bZrMw
MjguqJpHODba3fgQsMjJfLucwwi1NKMvclcdgTfGlhCv21BoLcDQoqrnj89/SS19
Y6wWlz5jEBbsEn/2fA+PhfzG2q5gxNNCexV/PDOA4FpdEeMsZJhctxYNnZDtixi2
SYlaEA1vqZxdUxUYqJMMlxqW+gDRDO6D85jOHPNnMum6FocoAOf3Ju5dZ3zB+Rai
CK6mC7kC8HWiGfatbYRxvBtVdIALk13W+TkuWPFOK0Xo7hlVYYevYS9PpjGFiHtd
5pcpLfu4wmeVh6rHn+yqFrvgjvAi2STuJ8ALVlSXnsTdlDcriA6XS/IeQ84Xc9b7
cmibSWsRDJeLmSZwX77Jr6hs8MmOxlH4/VbK7IMECyPtEZt9eCTu4w6ewdVkH9Ag
tmk8YGjNaWN6MvGqjKa4YJNxxlK9RXxchwEmn+DtIoJxAInAUKXKzmk5x/X7nol0
/u2ZryyTN1uwRi6rjwApUsVKyZut9dZa54awKjQ2wRUrpDS1BUKrnqqUpAVD79T5
8JYBddKfku6RElJiLNNYMvJOJl54ie7pYtGw1Kal+6cNlsibOES2KzAQn60yrji+
LodZHv4aetzebqIjoh2CxLBN/O9wP0sn0hs3Gpj7NS3RLVSyFTX0RBYHWRHb99QG
VsJkhqYWvEn0GrDsVc/+hQZ/JSSzRoE3EvEjluo6LkzxdNssIhtelCTOL67ssANx
jIQbautIQPgpvY5Er3hWQ5KZTsw9hDPWNZ4zPOPjdMiYi6AeKkkqkQJuoJj2rOKa
dodKwRLKIyGwXJ3fTaPOlyd7s7u0pnN1JHXCHkSLoXi8N4Cwjczao5pHgRaukpDt
CZ4aHuIqiyRUcpZxlpVlZu8S0/6tFpOfoATiwUWTTmHM31yBh+YuzqkgEnue+PHd
FoU7pXfR6iOksa89gIPJ9C+BwbiMU5+BG3PMBRvkH3SxYELc+1lU6ETvp1pXZb8U
F9qdTF4wPZZ4cA2LhY7WLm+AjKOakBr+k9ni5/4eDPZWMEEfF34zuFmIDnTnT2CO
AnsaKcVWBX4szcQTtNrEv/Be4GbmCGAtinndVYJsnJIwz4fOIAVmquXdRkP4XbzD
Qt1CR8vX3+RUg8qXraiZiFkaP1yrHhoMXJYUh7GwTxrbR/Le2FG5SCPKKXMatFSb
EcHuYKgPyZ0RMFfYUfTvJN+LASSqUI5oPIGB2O4VqcR3KpbfVB6kvsJfSwxlA1E2
+iZWM2gUQFw2T19XVG5IqGpgn4Xhy8iSSOGjnGB5nlVeFA2Nlbf6GFTegvl7y7c7
qFvLCe1fl0pTDZ+ulB3sk2Z6xrLGxqByHsJyhm9PjM9YwrzSybYS+9W0ojoPpLF0
gTn8pjJASnTyhk9y+Auqe0gvlclrdU52W0ERTbonYK4SXTSTkfw3tORtJ8RxEBwB
6xNyr4ygEVJa4jH4FzSXypW7z1u+uA8pqHQd1xuJOW5YQNau9bOMJiQo0DmVhW1x
iMb0RtYauU2rKyI+QhFoB/jLvFCRP2skdN4G7NlBGR2s6u/9y5ap2wGGi9CUO/5D
x9Q015vjEgMvqE8IqYtN+qn/yQb3c2UmDJpAEHb9VxIR9RwbO2oQ+8W57CQUzDH8
Ye+oRoImoOKztAKiK0btfK0qW1TUS+lygu1LMlE0zc7cJY/sW3rkEzRt3jOsZV2m
WUsVp/vLj27zkTuhdKCUqj6h4nh03yNuI51RSqwpIHkgYmFoXYfve2oz70uCMus4
AdAlM21hecPirG703j0QJOKo6ZkmVQllznkdehOK8glzHhZwMXbGuzURotZSPDRM
8oIOqXDowQEe6jWaDomxinnORxDx0fLC0mp62OBS9v4+SeSIr527IdYmN2i90VKN
X9uXrxCoULiMa/ZxyVzjAMMPX2A49X4CeeASGB45AItYCXVexZmUkxqAl6xT6QJl
lAiIvXPD/OCaYFNPU7lpUXAkMoTm+XsKjVAwWgoVkIcb4Xh2LdoaX/5ud9Ej7cqm
i8ipz/cXVBj8jiyIqWUuvb0t5v0sFm4MOznwoFcv5ZOdy0ApD4yu+ync4dyBGhV/
HO71dX1+9h1N/aPZiWCzEFdDWaW7Egiqg5/O6OYcWlDynpPuzEqkkiJYUogg7eAQ
IoPumBmA9l2DUH2iVUuOFqm8h2YeTfq7Rtx4+y74pKNRnwOYWnLA2+Jq9gxwS7Il
Q9pJJnDvKbUcKGzEfOMilQ29CkM+NthYm979ZqFWV5APuR/YZTNp/a1OE/B1SYIx
Clv7f/UymZEAMHHNnaKCEoov4qCZv+9u9QkoBcSx/nuN0i2lchab6rAFg+vUWfsK
gjVjuxx+9Tl/iKMJHeFKibZcjCsADV4/heyaltvlFRbjxWsXSdqJxL/o1DeU+jy4
ZJXL0YS1RW8bZSzT1ny795fJEz8nkPRZOZzT2K1yWnMSpP+aldKgtHzRyGcwJTZ7
gJZAXm5JAkCvqf/eR/Uvka7F1tgkKbFg3endeZykhHO6hAmmQ8jzKqPPzATw2Hhy
j+RHB7VqWdt38hf8/1Jg93v7lTHFrp3ZGB6RqfqplS3At1kUkJGUrct7pXtBy/dH
PmJ7MtuCFVXoUV4xjNMi4LHPTc1auz6KxDhs+LQt4/v7JgsnW1uvR29yc9Tl6yuX
fUIcCn+/JouwSlHf9tuFQg9fHnjQt4wPe6R8sR9TigY9eZ5oRZHM4fIhke7HabDx
ZKBxI72jEr/eFR5YqZWbVE+TPe7VRhnU+Wv84JgkZE8jGBe42EWn20GHE4aUM2xA
uraWwMFVOtg9EQwlOCXksSgJPXvgAImahYxQjJyVdGOvIIYe95uhpxODWQowhzcQ
K6L+401sScrtlghcmO8PV5PYqih157GLRJnviAwW9HEu7WikuMDkqg+lCi5yecrY
DgjEhe26LAQXTWiunp0Ez8Xih0PdqdNBOuQS6rL1yhu2O7OOKsbaiof2Z/Tdoj+r
WMmWUY9Cp1FxNng2GL0tR77JsNUeB6jqcfrX3duVgm3/glF00hAjsmVAOSA/SuzL
/VTeDvKJ0yJKFt/H+JVVATxtLEu4wOvwDpRsz9OBNJyl1Q27BtjFLDriTlgWI3PR
fGOqJx/vW2KJ/1MQJgLuguRKc0KabqqVpi9Aw1ZgOjldxGlnxk0LQ+Qj7f2397iX
I+50NYVfBmVUhVSrHhVnaElyPGiobC7ch2hNnx5lSRBEuun6PzXNs5ui92ha7kGt
vdpJUWilnzorvMKNiw+3nCHebGJ2Gjok6XeOuE6K8eC86mnkjCd2GxVEoKzEKoO3
Dm+vqPNo/Cf6zdcNBhM1dLcN3VQjrQSkqGGtYEg/6s9wrC0cWXzT2LArXVTWgodv
YZjfElxWHzSoDi92prqkZvESfSU3B2FflJhRftOBESzPw1l7Es1a/EsnD35yqMyj
CLteE8EWuE7e4mSzxhaYdDM/VubrtUoFXatdBXusI99s0tydXV/7k6TsUDg3fhgs
glfcS5gV0YWVDZukuchAlUSZVD9xZdR4zl2SBEWh5xIljTZ7Qk2LfOq+ytg8kaEB
X3eM1iNNa6F2kKLFwU2caZLdw8InuBaoj5qYapz9083KQh51FhwIFTI17trnrDyX
4a443Yw45nA1AWpHp/v+Xex5JP+Fn6nZTTxtTObO6sVq4Vd2j3I2pRp9217sNMNQ
PGUYVW6r4TBHLVDvWzISV90VWkxYllGH8HOXTs7mHoUYSLOPmb3hfTpIh6Z7f9kx
XRd9WwtEGa5HzpMtT6nnM6O9SCPn0iRgnvU0dG6nmRGCyvk03egQrj6STG5hK6YZ
BGzRw4p0Fk38i10JJMeITEgKsxQMZ2OvAUJH/v+HRJdaS20eSb/du8j586cH2oAf
JYF0jfLWdCvGjR1MniCrO6Ldn2hiVT6noQrZTuUEWDnSwuC9O/vmeHOChhmCbAJC
mw/RKAfWJEo2rqI7AnZc4kI6zeT70EkxVoZF7+3QBx/jwNfzTyxG1pLbx+jG4gcZ
5PdkKNMqZftDYYgawoXLM2dQwvn3/00+8B71sFO8PqZ/lKHioSUPuzDLUXrePo2E
TWRGdMsp0W33I/BLxKgNVJj2tQZWRsz9ZYChQks9pOQqgBFH1h3n23FYvh1A25GB
7Z07ZIHpM5YAO4WqMFniYZI50ryS+7Ify8mnjugMuweeubpcfK5jXo+syQnLsfX4
oI0qizDeZ4DM+yBL4o8W3LL9KVJmBr5wlQrl7/0wRav8apGXumICuTr1YHjNckAF
dinR+mIF9h4C8ypZO4DkjYfkfMXgfNqLQxhXikoNFEyf3tEwFfMI+joeScrqD0ZC
yMTl3WJ9kxnZe2g6GAE3A+Z0kFRhn69gGd3CmeBvXeEyL7aTKhBRPQfLo46/Cimf
cOpfVEYJkZFT3YXn7dFa/ARv0Zpq8IJ+GDZzsPJ+dKGJdP4Ivi124bMcXEbUh7Bd
kEnxaZZq+oV31QlWO5KTil3LcmDsOn3Cl2rqQ8y+I1zgDIOnxdJ5+jqdxvgrNj7D
X8QMphOIg8zMVU4SzvHUg/ACWjBNXn8qy4gIrdQQqykW0159/YNzJlnqghm3CPnc
T+UivuADCojoKH5hRJsyTfhsMraO61h4m9AOR7mDuFfhB8BQSyrSktCoyVp1WXZt
KZYDVn1VLP+wxNhFfRiyRTKM+kvAsmTEVwHkm4uC6d0r4MzvGJsWm6gzlw4XOsI8
mnCMUrKD7szIAePc7aZ3i7fz/4nKJH+nvQamsVBxTZZBM97UV0fRAkFJuRnJsD14
dzfNxtzBfTyRHCbRU7rJ5Rxf2v+Ia8rr9SfbKzLrbRFphxI9Q16BPgMbDOHLcUBY
9jJiSOzSC8AW59jWFgdW3f7Lcttg5rDI7axrJprYUDa/FA95JQRGu1UTdAJpeTo2
cY/0PBqUhEki1qQ228fQZKZuYyzPAh87WJd4hD5pZaEiyyeW0bZ9ukBDqVrPyHuR
EOGtKiRqNFqy6tfwQCaCW6UmcFu2eK5Dz3OmIIlhsu91zgzuCzSrSlD+zg1YH7wV
FtlIOY03Ug6OqnqGuf9p6KQee4TOAx5cR8Rgp5qjcZBAqlxtN1buk2mMkTv/7ZAU
RFqIkbyGsN+BCtCrFOrCHL1Op1XwhyOPa3qjVyRBkXh4gRFuERXRyvglfjzcZAY/
QkmQk4P9bhV9tSfJA05Qk6NjFZPT52OyMTv7ixRdVz7nijcxUUyfOadGlTSfb8tu
M9xU+2gdh4Y5jcNozNsFHkz5IdPq4QfZUfFIbvBQNlP/VviZjIAFe61JnqzBvZF5
Kv7u2Neh57Lx8873JGJ4zfcXTSniwybZvUMwPHwOIuozwMDTuPDIxdc0nZP/5Bom
HerFzSnY7LtJ6jxjaWY185kVSzbYzb36S352HS4w3srT/8aH4bDD0PZUusEMirzz
NBuLM+wJvKNN/6ZZ/q4L/lGgBA4nTHOt44LKTUo7WW9iE7eIz1ZVoHDZOen5ErU0
EHiA7GFxSlICPyJibho8gA==
`protect END_PROTECTED
