`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mKc+rpLcbV2ps6vQfeNU2g8h2FabINiVRdQnr6J/7n5PHIpd/X/OmcX8cJ+LrtYP
+1VzR4jz8125kwF27bMK8xlUbGsIoffG0nxq6mFC1MFS1w7Vufkjf+z7vXJ5nsuD
2y2QzqTxrOzXqEZZanc9qjAL4ykJ6tuNs9vPeSRLEuUHtLEFOkMhXlZQPs+knkSu
7wG4N4ARz1iGvzwzyJrNdQHfL3zZ3NPKMgqxtP6X6IBNA0eqeV6JSCEVs/MfCdQL
kWjtZRvftMDkPmUKKtvZEMLWcUnYSCuDFsqyC87kKTkqc2DF7YA4OOgMoi4eSWOi
zbDBe8Fxr6stf2XtaBH+cDs/+KNcQ8nRgk/oa5UF/38wfxqfM2eHz8nEezgWSxJH
D1XGZXi5PwurcgJ98C+Prq+QNPfLlX5kyUpauD8FMqypJ46dIL8nJGfUR5F9gcMq
VhH7KUO7M99fsBJ6rWr7CAZjGpS2Vo041YbZnp3xk5EMdpQAH63KgMqTxYQVrlvh
OTbB7NxwQWCMZLY2CLvs+Fx0eBxydNMm8xVuc6doC8XiLS7EDfjH/ax9MsaluaRM
SM4HOHutDz2sG3VUgDChiQy0RX2F1QcxtxA6HaMrmuA/iIhLbhkrygHIbjqNzChh
l6hede2EdS5SDCuFgPHrkmf1ogJ8fh874JU/0xR/5kZh7ar4TMneF9ssAam7L+wg
8y8qrPy9othM4v1csDmMJwpXDVIo+C87R6aq4v1KJEtB8xAoyZC7gH0dUcAjSA7d
Ir55UValYRm55xf0zYnS+NL7MnLtCNW5hG5hqEJGtKRvki0UWdHz7LFJkkd3XvL1
X8uMG7WyWcZsKTrs7gAVBfItaibzRXD0wooHHRlKxcQzrRop+obCR8xPtxKbtF4v
RLEWUlcrRFVrHLGYNEXKqoRuyBC7Xg4dkTSPCpT3mr3GliwgHOz5tCF+RKcyfP+u
gClgzbI9dfhbR1llN0KiwfMy+nqzNk0Xr3kAyrnOefGwkbNS8joA4eHJZp3FbIz1
3OT2x9JRgCVu605S0l5Vkdtp19ODNpWn4LMhdclscwK02GoaiTxSES3DpQn52gXk
8rCKhov34c0TWNYdSeT/DWmhPhf8j0IabdkWm1w1ngxngMYGSNwWudLDcWzvnNlZ
EJQ46R126RAoh0Py5rWw+AB6Ja8LxIvWdCMw6Vp5jKqlUAUBduMTmz0u0mmaHCQ3
RlWW2IA2CVxeMUzEyKKeIw==
`protect END_PROTECTED
