`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ddCAW7Ih8UCm6UkTIyzaGUp35rlF5PV1ffgVJVbtyCjIcLB03VhkynvTVxTmwQxg
Z/1xothwCHdwsucXrlj2wBpa716Paxdj5knD0YTC54aDzJn2dcRbUG2/3JresOtr
g9FOVHpIZPRuN5Ib8xwA5Ewh5Fg7CdicA6CmbSSpp1UqGZIhl8zum8XWX5WZDHSE
s89M8B30B8OdMOJSAdWytpPypPx0J9A8aHQwE2B0R2gjA2lXWmtkgPuBNWyFbrlX
slE/EvT7BiXKBcaZzu3pkpzzaGweGW7hIv08tix9Z6odU0Pz/Z3UDoHNEwDPGNVZ
BNYlERgTmDEJJQks9a5HADVEUdSividYoADSluiLJYV4KT5ps4R8xm83KmV0cVdD
+38vXBQG1UCKjd8T4yD+zPzw9KZgPHIwnv2G45gNB1nYiNslugSkER3dj3FVZTVr
8+pgJzWEApBO8Av5oF3zy37SDXz5EXK3F7H/rLFSD9ot55Z//HCcIVa9i+akiWkW
s6w3CYvC3pgkSprxHSw/zsJodhglcKTGnt9i5vglEfX16zS8rZRXJxhZ0PW5uH8u
jc7HPWG2+KeKaoedwI5rlMeJhnwJrnTKT2YeWBYjZ2rK7n2hUTFsdtReC9F/jSSU
1x0HY090y1Kp9KtpBWX8sRb66Amxtc0Uc/OiM3G3yXRSDyN5fXOH0NrXizBW+TMI
CQV7i+dO9aRyabxTVPB1hg==
`protect END_PROTECTED
