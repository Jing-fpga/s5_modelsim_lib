`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FvaPWo3Q9D46kR9iGRr9ku5Irfv0eZ9Ezejz6uhguVEFc2/TMidoUazCflyk4EgB
OFDKQiz+E0PmeD3VPM32d5nZsr1lyXP4WuwXXWDaEAT8jpfJAFYRKNoLMG8KHXPr
hHq7N2BzoMyKMYuBHfqFZLB3G4lAhv7SaKCBFrxTSNXY2GLihnjnN3B0ajUgHRnz
/q5KF344ETju0CyT8H+qGMigPlSB2sOrIUF6XINRMIjp8nfY12Aeb+CuTIgRkc5o
vuYTVTEAcOrM25+Uf0J8IGf18EKPJX4fpgfxPni2lOGdxfeXJedfHLGuXFwfCDqv
mHnq7GUTIqAK7TdM3RKDfoqdJBBXd6IX88GEAUZBRv2ulrqf5arS4ysLbwnh3Z72
lHedlzdE8LbA6xsh3GZt+bLPCQDqEXPAq10o0hDOvV5XmEhwW9R3dGpOgEqUYopr
DuSFXwjC5QBAMHKvu+paEAla1HiGJAFjaB08sSxGfiuRO+e4KpgSjKAiBL8VuRdJ
q0lDCqQX0q++Li6P97F92Qv7y+olIMyi7eKOmptpp8xvHlTmkf4CQjGdSwD4IpDa
jXolMnHAbhbxjqeGGVJeIP4TPMppdPAnIWILz5o0uamFREmuBUWUayxPElZUjwlp
5tcHiLks5KGt86rK8Z7PoagViNlZdnS5XgdLETMI0PE=
`protect END_PROTECTED
