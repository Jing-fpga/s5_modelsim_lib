`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zSmIdqbvhqnZ8LoxfjsfVA2oOl4YN34xhp4W6xL7Ey0EyuAr1C3a6LZQK8bpDn/D
F1t9OEwREWAWc57fO7FBkkQzgtZCYHleECkfkXealyJAf7gf+bPq4vM/Ks58LOVW
qKlkMvR/CXocNGt35MAXUn2CYXBn3wtsCsAJ6K00zNyUwSaTu5qvm1qzLEXXEAKR
B5SpUDfY4/+xl502UbPXuKWOT9gQkk5G2txzcLUkenkQHoIphYpFLtI6tT9KBIJH
OtVXNHsRhMDeyNB+Jc9TrN9It8NQft+7KnELS7BArbOb2BNC0OC4JcFbGc5DzOxd
93qPitOdPM1luVDJrcwXkkL9/I+3hUP4cOmo1zY91vDJOPW0h5JiScESstV4vlrJ
UgZAea3ioGTDYspyaDPYh+XoCN2xnc3htNYzpN+p3HNwcIdhyr51lzRWVUMQdko5
3HhRJ5zkAYGmZNkdmzPgngjqICTFB6ZHxlr8Be5PznMMsjDihBlt17NRLzdgBJ4E
YJdEdqdhKWnXRTMqS4NefU8G+MNgfPvPj6ZX5MFUO7Q=
`protect END_PROTECTED
