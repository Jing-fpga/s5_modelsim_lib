`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x5MvYzO3xANkocC4xbg/ZzLCGuPtEFbe8ZM7uQaGl46IY4p6AvsNbjosTzbbNDQN
8X/HgE98Cq+iDLKZzzLHUs7UZT0Br+Gncia7PRyfRwhhkMUSLznmQ+jdZC+h8uGK
OlgN8v6gOlObrEa2wldR3KUpWJdGKeaND1xX2lA+P7BMQm8w/khwxMrdiFZFM8Ut
QUjNA5UJ1rg+Y31jwP7kYC4jcwSPUR7rfLyR/T+5/Gavv+iY6yr3XGMMwaEK8B1z
B07mmE2iKktYHBenvcs1+BW1DkhhEQx9drqiWgg5xd/XjXpz+i5fygf3gvunm/py
DHTL1lXTWP4MaTcJ5ECwUQvlF8l9r464lmCgAb9FvWOXu5UKj/nj6OWGFthElu++
1ykyb+Qy/6lQJ2vDw3DYgXNjxLe27UFxXDLgL9pnwTD4Rh5UWbEsDb0tPFWKGawZ
PXMGaGQu9XWHUZgUVQYnZrVndk8EEFPBKvvneiwJzVumZ3+Ef1F5DA31Yd9X9CJR
ryCuDiFtTTWcMeVWA5X5wP4OjnYupIsBYmhHZ0EIeY6l6XMNpIzz9f5N1v/8JgxL
JC0nGY5loqpL8vZCgHx9j6aV1JsCwOWfKpOJOApFzh9kOykV24paJeoXQaxtVUTz
Y1Y/wjJGYr/dETEOu8suW9T6M9gtpsvVlV/pxHSpje+zv1BAsOu1O8b8sfCl5mJ7
KJblhs96YvEIs5GNoVx3+emA86hdnuwhPx+imrkOfsubqUn0Ob1WKmYDT9ORwJV7
iMj74Jghb0puIocbFAPXK2L7hTNK4RTHgSpmTW/0Wjo1rxhAib1et8L4QITzH82n
rqRqIMPwxi4vmJcbCOnVtJljSmmRpRymFTrQHpupI7KWvjpcyMq+AZOouAXo5VQS
fq75LYXL3W6xpmC6ozGY1JKKMCOnXYnNYizNeGKhk5Spitb+9fwDJYVN+9n1ISdt
gzNHezUFcNhWHINHpDAa2wUsTKwrKXgwl7aVAtzke2WWPyP9r23N0U9tgW4kCgXT
WzfrNE/gp4MYb3YBsAwANfh4D0GFijmdzgqxq7DcnM4Y6TaTaqOKcWLLPkC1fWSK
l0pIxxrWzUWCmpgfaC/Uut5m5OxJEYNtQS55Eu3BjG3t/qFjqFkPaW2KPtwQelaD
xOIj929sUXdApO/IntJ8i1QiO/3KG1NH4BZgu0FityFausaAdbU2RSxE/w72Y2eW
nT4c19eIQjOy5MVIk+3Qqmr3jnRb1GrM3J9pxCI9f9+fK6PYgLOz9h5Yz/vVNKB5
ITlsByX/j9ilwVfB+PVAM0yo/k01lO25ft3IPWxIWjdf7145GS7QScXw1i4m02fd
Huqd/TtrqbuHX0Z1qqMdXDOOxiiQIztDtAXDNA4lw1Ocj9iFUrXBa2Xqp5Byj0wH
Mh0P0g7KtDMYl8zkW+1uaaNv4aepS2XL7foLy9X6D8DkFRxQSyvXZyuEA3xNSLbX
3gITcs5UgsOYFnx4dFHcV0ahd7R+dKPA0oU0DXl1E31pu868OFRKBBKoRdR9Bwm8
EwR9PdqTyZLwSjNZSkapKstalpdTSGyK+u3ekvC4Kwcj2DvkvFtug/Y5IqlhQZSQ
9Y97+o3OrOmEP0bQ8LzCSbnGwyo+Rotw7mZIsSET4DaOuW9yZoUM4mELA6EeI5Fq
zmnNF9lH5VRlEhKQ5PDQxPgkVREhS+N891mqAj2HgEy6ULxTM1ozmViO4dj6JHSi
8XzRec/I7SDzH/7bq1dk3VJ0MWMv9n4/YtFk4/vvUUfzm/lQWnpEe3g/llL/lGf8
x+JKVaKzszU6qtPWoRo2XFi0UcijhMTXOKDQr/3pf34sp7ZDOnhQ13hnvh1FL6Hf
UAsMK4qZCJiSABUa65HPcVhaGyVp6ak8gMwXfEFSjtl/+Fx5K5EyWml0VjoNhTxp
3Gcxdry2jgkTqOXJuf2j+IQaZXmo6AwZmL9C0xfnEvhuwJ6Vluy6uwjJzkirwqLi
XbQl8TwsUZPHtELBBXvtMyosZqkHx5OboGgf08BF1a+/tWAnO6Kdm3LfhFqwAEiu
++0UZsN1wfXOMzSM349y2yzsuHQTvvs2yfMqXEcv77Y1+t1uh2qVuILRyEeeBRAj
sCeDJmGyCh1CngkI6krBfn+1SXT1xV7foJq6pYMOr+EUjREO4I5i3zRZGAEX6hwq
dOAAjQcWbXCOmKPpV6wrGqZMik1RXMdaI9zFGe5XuCHqrX3DImvdzmVsIZ/yY9sa
QQ46QYZzZw4CFFcSX8ndDgtdh8REjH5xm00ZS4zNYYym76tFLZvSyK+L3OL1u4Pq
oogAbSCkiPppRAI37ZXJZ9v9YrpIgAv3KvqK+c/jkRf68ZfHDiQ1AnGP1/yMF7oR
/SA8O/yQEXeGuLDkGjWo0iEIFjxouaRyXGaRy8GsbOp1PlchDAUcNfP643IO6rvs
8VKjXw61kF5qfJ3fMKNTLqoiHqdRL8+HIgXnWN+f6TVNnF5xMZH2vFpyQEzdyZ4b
Q8yOSww0i8O/J0Z5psMXXe6lI1Vihhmt9rlRw0dAUTPyNspXhpJcLjTx6MQ8u0Z0
InNVg7iOBemTJio+f+e43K4SGbOtka+h1qYuJ8VftcHEY01xI4alBN4fD+jvSQuG
kl+3u+IzWCEv1Di651+30J3WuSwKz1uGtZ/ftvrJSqYh0mKJu/m2YJV8ftjdjzCC
hMVlO3KHrB3Zc3yAvBxuql+kWalqrdFq58ggAPiG7sF62wHhRIankVWMrmlSAyGn
C2zlLItDKycx3YdHga4aZrbS410ZDNbstj+Tss+SVA2Evljho9t6O+cNAQdvXVTf
brXRMrsAS6/vTN85CFZB/Hw7xqzKV+zIY8FO+inaRxozxbxEn4QjhWHnUufm+5nC
CpA8SR8HyjBz7+yTOMYOs6MRJml6yHgWOwOx+a/+gMe6pjnFfKnGTMTtn1W4p+dY
9IsDnH8d9FdvwfIP0gx2e5IpFcP0fTD/JywaWJqPPhsiGfc2TcEW5eaR92x6EKek
4/CRQ1V2I2lG6DmoT92MK7OHILKrfy70NvRy+lAHeG0WEVW33jnMRasWTcfLPanX
EwNiPLcOiuYNtpxizCm27/273SZDm8Dkhc206OjkdvJwBMCtMAxwLwUsl6ok48cI
OfnP/Kc0VnxBSEwkqFPUeP9WSu9vsGpwvGkhBsps7FkXMEFUoRVp/JylYn8ZHzJG
hDYBnTvisvbRRz2HX4UOSt/P606lkpsP2qgWG5zfXZjVnAVwgo4vAjTvFBs4pLAa
t3smO7tZC1Bqlh2SR+OAhTYegHM+e00FDs8Krg/MXh0rUFQfwzfxRzlE69GlyTC8
lY1QGvjc9r8gnfidBErvQ3e2nhdlt32sZiQapetenbPv+i6RuZdtf1GbRaMJ8pF/
5WmyAA1DsWmFhb4NFGb+jx9kWs4u35AlNwtaRdg4RY1/EsyzpuD6aZRO8RNW7bVh
ngbbC/dk2bpkqJXKl/GYitEZhLtR37ZIs/Xr9sqyi7QgZTMKdsPQ3T/K3sokPUXS
xsMqDtvd9dbGFfDrZrsgpwa75t6YPMHgSsPOahKrHNnxkveWKp7W/kwzgq1x5slU
FLD4OUx8gwhw2xZ+yrBWnVSHsz/bKiA2n+xZiHm+paiBLBT2bqyATM7vKspO+mlb
wjE89kMKinpTEdC2+H9i9Lt2iMLBdlNAD7fbwjBw2uLtfSST86vXxdT/ThwmPbnV
B3NvVKEznwxhj2KEQX8DCREzh2rAZIaa3IQ5pBNPnnwnpu0TFHCAU0++g7ZSza7A
ElXpdu2/+xSp0qq0PQAc9L9a+HQj/yZo/OAFnGRSyunbDsJPTcQEOe5ole/w7ubc
RnWNiOAuCoHmYerDGyNwOsiMrg4sG/New5wxHTr7UnRIVHvzLoxYNzSpITpEnMTF
5Kd7HAvX61rSgs0XPyzHvM+C1LlZ841vbEcqCFQJcwJikch7KEdvH7ooiXJvO8UI
9OrN+HVJ2O2wXk3HDhKvitTqHFx4rfCHt9vdETYOmv1qoowFAu3V3P5qWKI/5HLV
boPsuH9oqlRDuigd8n8QmWcirZn+O2VYfIff9Nng7HVNpoJoJ7Q7GmXLEMKTES+Z
SRewo6zEXUeUax/vMz1fAFLOguB7S8xorhJm90EKhP9F+u12m+9oS7VFTIFZGSpH
aw4AN4jup+Odek7bspIk1lTavFulxBkfn9w3yHxMNXrzzz7LGLP3tjcUcszfuKc6
hUY1sz2l0kcv0UjXUQF/4LTQj/zbjrxGoSeoocpMtYZXSF0sLn/zkXfx7kXHZiEV
qt/+X2odmoMaefeS73KMFIuls0BJaDVIYZoIFfh7Y79P4SlOsgefaan/0eCvjUkm
rX2M45GujTyFxVzrXKmVVFR2y5yZ87Jci5ngHwnKKWp8uouIy6Dj2NAuK9XUK5j3
VSsX1h522ht+yIo3nskOGZWIaHJLWdaqJ8nz+dXgoNJoTA+87kKRS6PyaKY8xe44
oPvGhNDrU22VSzkCkbqOoMXj9t8mCLOOKP2WtpgnbqRJVNZDQrnToeoHf/GXjMcb
jSYnKmVw+fbnVqSBDkOUbZvtBLLbOcTl90jPRxv0/FYFIpowYL68NHtVgHvYPF0t
cWRHV9aOv2aS8UHNFetxRHTnixXUinRp7Af9XG4kia7lvTbu58FR74vC5VfTKUPR
+0M5xPUpOZ52t0s2G3S34ii4Xc8/6oKWNUo+3EecYz2w0RmDqDSypZwo4osUEylB
jnzWyF6URTtIiWItdOYZ1L98Nv+WoqSr3Wxa+b3WdHRWu3w2etSS6ghjL6K7FalD
zSs6T/YpxjERC+OCBIflpLUGY+qtnLl4eU60giC14SeQyPfjIxupFpUXOqbV/ZLN
0viFZzx6e/tWs5BKyEhB4XFHT635d4ZrS7nxcNEInY1ruNx2JT1wj3S/R3IAiLLD
NNTq76CYxU+j2bm8jj01Zff4OVg5ptdQR417B9n0nGrWIYT8rEPiIt3GkjRB7Id5
Eu7w06FehGHzc9sK42+uD9Jl85CR8dsK4+TwHcwl4OM2c5V4mOUi1snQXLiNmaBn
YiVE/ncj3xC/dyHlH+UTnDo//nW9JioW8dHQKniCh8QFXhk6ivFuxD/5QZ2TzjLQ
qGDrds0XFJ3CT1PbVOVXAX0YoQ9tizbwBW34ScE9gEdJhKMjn+CIOm8d8XVQk1Gf
Rc9vf6YEhQN+UimSDE0aTuslupDtsFOzlSetscAfaduOB+D2vWx0bjVLW/NJK8VM
B2nmbTZtYsXIXITX2/+JVikTGFAmx4osVH1BrePH6V6x4PbYbknIIMoMivD9f+uL
hiiGQAu0gNbGs+zwX9KNVpRbFgskk/R+3TWDqgx6V+NlfB3zbwQwZ/m3kyW4cvJo
hHnBme82T5gv8J+FtPipWQbDdkwAlgX5Hv1sy2uH7dPaDQqYUkARe6mLZ7V9Qe2M
p+egYQm929WlNxCKqvFllKcwBoqNllVhbFtXQ/T7LRQxgaPcmw53pRAir19+bl3O
UpSonBk5sfWuX+FPIiK+C2+sdm0DnG3De+ss06qAeeFLjtAoYnzsu+ZdcSEP5dEB
Z1Hy2EWdpjWLzxTOUnIRLlY7oZDPApXUIfx+JmUu0YAUyhjEyLsaWAHjMpJvz6m6
ZAousrl9gbexk8CUkDJ0vl/XRd60bU2VXIV+RKPG5AptxIReR48fbrJcT9jVGnp7
QVVa+Vxq7uvCckA9hSMpPbFwW9V6RZwqPLZCjtXokJ2No/ESaydIP74DV8UxJVNB
/DKVsW7eylgwXYqisAqKPEOh7KDs9sXAWqqLyxQX+X6pdxCxe3hBUflfIhW8AAkX
6Gcctxg8BW2dqwxnWaXvaU1/vUDXZkVzsNJwHWN9YHsqAfCDfHpUG4t5aIzH9Dyc
aYum1QjDXK/qkm3wmkb+2+IML+XyDQjnOY4J0Q2tV3w42rh9WJFBORUkESA9mczi
o9OUj+VPkyzqy9+XvtH8ceCtxQftUjX+4SnXZdLbfEbTAaGl7tMFbTHYhp89GhPm
y3tmc7yorTKizMm1F8CgNTqf6s7wqZlFo/G/3R4A29hlNbNo9GSB7C8OZ6hnVj69
YlE0END7if62Dk6iqZ87GNmY9np1kmsWvIWL78GXMoWkCpcV/ogw3RAl+EFwchES
fb1HUzbwDIe2NyP6HUCc/E0wP7N3VLBfq/78KA3lxyHnvhKXjAL3h5znFEp60xhz
JOpbo5UHlahXxFWph1Oe3ZHec5DTZ/eRuBnRlmh44s1YyZWnkdSlEZ71kR7sU2Vs
VYkGAU2Sp/0RQPRm1/VT6c5QTG0R+CrWnl868PLoKrHr18cYPihc9AZZE5EV3pDi
SMRhGyDJleT3hGLDlbmSTA==
`protect END_PROTECTED
