`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sPdze9ys+JqC/4xf+7w9idzmymJ02ij7ZMyaKQpZcsbbMnVqmDV8ZZwRM+j4/0E8
MT18add8lrM1EZv4mdBW4FMm0N4BItfqBLckGUwl0t+dCSXVgwJdQjqeURGon3FJ
18D/u4Hi6yDaMvOgpJ0siGxwHuCBha93iqgfofPGAtXbD1EY3N06pB3+QnNqMssJ
EHu3tM7XI09x/W44y0NiYaDNbYgo7MfLXoU1+sC8oqI4UQsbjKsT9EXKBEwXLclA
4a7oziZtkJOKfg5+bnNItM3LUiLKLcApEccRR413G7IcqaSlkpXncN22PP/fMxnY
dYcDX8hxEeMrWkZlTdHftMvBygXFKHDVmO3fTV/nPMTCKhf6AEdwh7Y9ZPz7CWYh
kyZhcfvLMqSCsf0z5T/6qlevRIIkNTVaheiOcj35NDx/wkA5H/s+kcZOdgVbNGq+
lZZt2g0iBB/0NRnX3pKmtPdS0bOTXN1rg5yR5WApGJW81gnW2l689H5zv+DHYTPi
BYLyvBPMuyiZBwZDNXBzuG1AqSznwDtZgROZVx/KA4ljqY2XWBkeDnB288VOL5Bb
csAfcCwgbcV/eZ0GgzKQgL3ezUiLeJ0JWc+rHDm0xl6NVdT/zyUysTtJr2hnUDR1
`protect END_PROTECTED
