`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ok9Dmk8UlbsngMiMd9KqrTeKvpED7VuHsnfSsm45OMQtW+vjXgIxBiMGM/aE8JHJ
j9A1JhNuoz+Fmcq9KGHT+m6Fp2iGwKdayEdkYFm54uT305Ni5AZsfizKYRZO9LQ3
KTbAvRLZVwSvW3HTnnwkVnKJj184jiyQHklIH45eMOTKKesRSdJBbmfbjDCPTRdS
69yPv59Y+qaiG9SQiK/JMuDZLDt6fd9ip+GCyh6g8K3ogKlLsDixz8TQo77borAy
K3P1D9ERGqyl8y/y4oQWw1bbh7+ci0IUSRLk8ETfl2d9bj3q+roa0ZeHXvwb/MwV
Rf16MwO+gPgaDxrlmozwC2uhvJRxkughUe0pXcHF6fA770yCLi8OPVU4nJ0cnffI
ZhvEanuRoFMgl0rw3wv7OupkZB1Wc86otKSJjWt/u8jSxO5aryG7iTG9bbMAPUnv
4BxkbzhJEAyIHAnKAbKZy2QhYwcv4TN5qT7w5FtZVwZxsyBhv6+sM07S/UT/tDzh
D9AfV1DgXP9/2w66EfOwQ0ToMXUdqebYHwfTzM9r5VhyoeAVCVcbC68R7fseE9gA
WnOUZbGmHY728gLrc1QOjyk0zW14jeTxneR2BTc4EB7N75PD92v8Xje9rtNNw1ny
ZgZFoxHQvtIJ1s/qa72psw==
`protect END_PROTECTED
