`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
66M0pTre0Rm4cobdvV7SEvddGWakDM0dZXtVJ9Fne1bm+XF30JpemqVkDXl1rwt7
aLzTpG2gSTEQPGMEnyB3RMfFa5SO8om7rmb26x8+9E39ymBNhZKdCK8lxuyVWEnx
+A86Y8qbJDAbjsHh/d8vzgUIYBgd7KHrs8ruJ2OU8LqODc43DeKAM24htScxPvB2
TkwBHLVP7sJX/QeqzTjtnTxvGrBCIXEWZBKSt0jbL482QWF0cG58OOwSGvdZ9/hf
jXA85dOJt/3/f3yR5zbZFDuqLelaFNfeXHbDjmZcnJIlzNXbOQQXSJw43QsApip9
I1bumII0EhQ17TERWW1wEJ++RsJ92pObuyIA1Dmk3GD5JPvGvIec5Fuw/4aOTReA
Oq9UyffYLEug+kiUyghS9797umMEjiuBkpkloaP8qwoqXfSA3kcEKS5vQStnoZsU
UPH+hn+mVK9zCW5JCrhpgoIy/A7kAFrcL9s1erb9sD0+i+VOxZwNHDPoC+oM9WPT
RH4Sir6beWGsX4lUjl8VUEkPbjeyrJ+WFksSCopcrEnP52xEl0eYgL0EZP0o/NuX
qhBZGd0rkS+w/JGqJpRGOiupe/TVWzJPYZ1Eu5U5exc5+tCfjOyyW9unxdQ49WnH
PNGs6To7lhK8ufeNFPu4TBwvwoEUh+K0mLJ75EYdjl1UOED9mFwQkmS/IJZu+A7N
TOaYSOF9H96XOF8BQBBuwIl2cY5EDVlXY80o/wSBWgI=
`protect END_PROTECTED
