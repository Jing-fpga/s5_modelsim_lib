`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2WhdJ6V77my+YKmrfOpLkEpO7MOF++brRg1XEbzA94RFel8+FKCOP0BuWCxaz6SE
c14gsxMGccaPptDqy8IUzrYKViXz8W27/i9Ugyq00PQUM6GYAfZTVMvJWNbjNU8C
Wou07p22yNVJdwFmNF99yXtxbhuzZOjJ8lkmADludXqJFwysIE+lffkdX0EivovL
M92o93Xfg/1vD/WOzNorNKGjgJbW6BxbyGT0P3mhqg0kPwqYjycolvJMPbtgEQHj
8pGojuyv/URgr22CRhzTJtLTBHX5k6WipXRaqcZGxUP2/s88eoyi92NPDWq/Xp1r
dz/Yjm2SKA2bzdguvjpiWOQr4f28JZoha83F6tM96EiXskHbOED0jlABj7E1Pa60
DbwTdN861AZbl9ZiGmGV5d8eDXew7oYiIIcIteKKTSwhFwxHQQQ+xt+yR7jkgHPZ
EeEFn3qtISqYFwEKSlNWmK6txe5W8o4t6b/DIFqQFnX/LYyL+M9d70G4EZ2+Gt1P
PF9zEFYBJEFWWkJ+MZuGrioquruLk4yu8ndTElUq6rNCJAYEXKfnnPyWRAuFOg7l
hHkJtNE3IIkeFGo27N1Wmd2rLFRoa/dEpcvJek+8lhKAIFzZl+NBEv2Eh01WUgiz
ZGv0HB3t4OefOUXNxupthWF3NJaXjdweWibf5Qscoj6rOgnq0wxLiMphUEbF6zhe
84oU+sGtJi8J76oRA6rYuMxuajvkKvhOA5lKikbQZ6yrpJWoJmpOhLJUV5qa//jX
yAJ3FOKiLxcjwlpLF3A5D9X2Vsj6+Owb0AiplFr882cKVSS2aly986yulxxe0vvw
KRbjwnp7BCmfbq1t3FD1YxL7H56T/7kK+XzCaA3I/PG5pEBepKxQue/FxpJGb6JC
9zBOzf7dEjZFSSrYjiDNKcvYz94CQ+GFT5rDmK8l41oKyWiLEah9pe1pRjLJRZnl
P6gYP5rrH7csvYqT33B4i/oFMoJK3K0LGUlYGliXI9SV6rj0+yLRpqTxbhIgrfr2
ptA0XebzPDtypHRsdH/2XElhkccvwZXyc/l/z2uNTvWhOgN6qHo3gUMFbJFfE4th
K8+HS0+H5PdqDQAYO8U2xjFgB7VSHHJ+kEdaA2Uu3bHZPX+t5AsdUlqOiW1Z4X5b
MQ7VqUyI52whZ+Ex4CJ8ekI20f92J125Z/R11rpta7p3kCXex3sQ9V0khpLyzzZ3
PsZwINQMuR/crHo1hDNGzsyQOeoa4Eh3aSEJ2u9FrHnZ/3yg0/9RmWDiONUYN+dr
op5W6YXqLV4o70/3PhxXtTYsMOGcMKj9mKGZPICgJ2/M6BRYlLMNCkUiHLB4oSAM
vAjr3ABua/3m+Tp6kkkFJbJ4zu6js7wPQSJbjoywbDXjUl5B3XQvSrw4NIh4nk8I
LompShmlIl/vipDgJb510uLZkYKiCNCmgfaNjxrP1KbyQ+4VL3uvBsmYUC8UGuKO
+2B2G6+m/8PtlJOOB0o6b0il4dnnjN9uydYluEzVLe431S37LsMYJADTzdvO4oA3
isMgCy60y00YjuTLvzEK+H62F8JVJGAVszpM62KUULmeZfxg8o6HCdsqNCyvg+PK
9Z4VDEXil26+muwdfOC7SDWswexnCw/nwvBzxoW8u9TR728c+D+xYad80+kBeeXg
X84R/d3D9Q/RnwenvGscPWpaN4sXTIwdTAMexXQL+HTjlEcvn6kcCEcCE32mMnDg
L8P476QUjVLotFubS8dGWSmoqGcq0KzdK/CP+Nhz/by1Xe4XEkZNu8cju0KT7hYG
1OQOZWczDTLjQ3me7OjIonoR22gsk4ttAF2EcQmbaQpQ6sgg6JquzomrZ19FstEm
aRRu2uQwHBs0fNVlJC+D7W5L+pYvWClFxBonQIBVL6P3LCz87D3TKzpk5aLKRtWA
78+9LJXXrBYjJjFfeo49h0ktGQiF1KTz2Eb8t0rhazb5A/znelguZB9gozaiObmv
ybvgIwaanCn74xo9bvI36T3E5Hdn3lfSLn6LsIvZ9tPNBSNcC/hOLBaojtl+Q38w
SXVbeAQbUkiRDM6ckz2D2trUbzk+0UQKS0xQflEk/VCuiIhdH3c0tM1c866jER96
UMcYoqKvlzRpztMLPA/gjxX1FPupbszgsHJU/cOotNWz0Zu+Cb+TxMtMsG8qAeu8
IgKKKbYYznpto8ceakgTKFWSAq2EDIn2YLS8uLD6ekO6bHKkMBQodfgV1T/fxBU7
hB2+lNUIJhtIPHxSj0NGRkEXsovYDI2P7QkgEQSdaTIWAPoLE4R/8yfUtSgYu1dW
LBkoOkh9WZ73p1BzlOfe+XRcXFTgdE+hvgqZ0W70rWioPxzouNDjbO7WwF+td9bk
WQmG8rgcCMjZ8taOFVXgi2b5IDfzohNUdhLyW3yY0D1YqJXS8WCchdd9K0mIirjE
A3s7MP4CTK1v+bq4DWPiSih3TOCPe7S5uEakrKG5+qfiHRLOf+PfI5u6E+1v5HAb
mJAX+u5MExiOjAddGnaKaDWluLLlHxPlmhrUhvYABF/7oGlcp8Ec0k+eG23L9ltK
gSOAVHFtqEruyf+K8neViSp2cRs2WZuqZmBC34xyDXsmufjzz9SNY/pbGpx8tCmT
0qi9IS1cO7+XtD0uiSauYMiseaLVDkL9wAUg2QYzt6sHnKKonzHuwghnDPMzUFnx
Or58B0pvntG43HU9A7bYbJ73aUxf8cAYXgW3iWTdpUaHK3JPYZUaqHM6k8swB/kb
SpFeTimjlVXzo5SgR0ClccuB/PsZAFhZCZr651hCftWiJo74T2P39e9McI+aVX6D
sWf1uiFupWuj4KOXcLs0zYiOTfWHJIEkHe6NcIkrNAEcmEjzIqZkkQig+s2LiUeo
o/FdAh3MJRXvoE+FnfFOPupouSuIl7g767reYp8KHL/lIEQH711feEsSdCBpA8Ee
Or/nUxP/8G0cllChvG+qGtjQi6Q1RuUjL9KHDYr+I+2QEmWuAMb2sQkeuXbAh1ne
GQMIKAx92EH2DLiSUqBHk/ogB1vah+thXyrNMDvfdWWGaNSRGLvo4xlY9mwjNx9W
a5BniCCgoO5zNB0h16BjvyXpJ0PxvudLBWZC7X674f1M+OhiIvhZhTVc2qaIEZnS
zirbtudN7BIMXF/eP2MOAM+hOQImg03gAft/8AJ6b6FJg76Dih6W3MdouGw0zuxX
I8tx1lydG6erPX+OPH+OR8sXQSHGHihfnm4F701Yum5vuvIvPqPtqBdRcFZyjFDR
mJ/Wd5WdakSOzzfJxuDg5q8jhp3xKZqnNswSIT1CSxJvD3UUcYP8bYSj7YaJfFg9
HtVj7H7I/Y7u4NKPHVxu++Nh2AiBpO+HFEBM1FQEjX4AOdXr/9Bcq5PopoPXdXvB
vx6FZeLtwBeJSwUql5U2ap7+WOqJgXVyftUYzrjG6GwJwpVE532haI5dhN7ePfOi
u6lO1sXgXDuiwQCwvvXqXWv32sJJJKKsFcYdJPQaMgFR7Z4uvOTLBt+ReutCtI+G
KKJaRcuE1LkkUProflMWoYTW7ZbAXAMPgMQ6wFQhJdlTnsTkC6ChM/ndE8r3MVIZ
oDfp7nqZ5VeCOrP0IX3xgE7MomTy8wKLknJs9DePWK2H4K0tYGFpyF2ED8aWcCi7
eLWiiP/+N6l8Usiw4EHdTCIVX4Uu3w01PPP2DPQ5mnjRsf8la1oS9VoiWO5caT66
Io35EA8CF6Anfw3ZPreN6DPJI5n8XLSPYv2Jm9wrbLdf+Ok5IS+lAeKvsu58Lc9p
2gQtxY5++iKfbTntgVCQ/t4Ss58/0EpdwDaA0jUVX7wNvwVcfjIAZntgjBZJXk5a
J192IG+SZoLT3/wWb0OP9vrxEAMCeCe1V9ZYr9pQED32/MmZ00Tjsra210uyxKP2
NKNaUfVH3uSBC3EvCdLOd+vJMhW3P9jtBAKOxo0vlu69JuEBXTPDtW7aNjok72yZ
VyBIMYqkXEF45H6MZQNM1utMYu2F2yJOzdGToO06HyDkVlcho3FYY05KXumBKfi6
wSHjEO5n+AXCK7VSyAUYrpZvQVcO6NzLfFNbsyFEiPnW0ajlugCVQTyE3FmkNRI8
h8mK2dtfUwoGm7YoueVcHZbF7F9bnVzWagFrajcQcM0ulz3z/IR2+bN6aVa8PM+W
//sHQj6NIF7JOju/68Pk+Htn5aVfYVqQ9IdDgP8/vULPqC8PlV1wAK3VVpaxVfag
jSQIizKfrW1xeQc4fw942LjXTPCyDyyJlEgUZ3/x66OoKLknUs5bO26KnROze1+e
fNyHOXcQo0qBvoUnVgzhlKWzMhaZcV6BxT8o/vfXOAd7Ejkl88vh4LqmoYWjOgwj
KwsdtmTj+W5HfFl26s+pQSTsWJC++9bITZG8L6m1qFX5o8MYH4Okw0laMcbKjTMu
gtShPiMg10qWvYOTq0pmo2Rxgv2ltLt5Oud92vWQxCHmYdQcoXtplnVXjHK6mP6n
vBjR3ToKlULS5U978Io7nUih5GcH9UkXA9TI5R21HGm+CevwnclVA509dpO5sLzk
+slUIy3w4YiUboGkypsLvkiuhQO9TgE7gViEXZDU09sG1FPjcHiqnFDahiMidzOU
D/QCuGCYiWeYjFsoWVUe7SRXqeUaybNU6ZL+zCTr/aBh7iy97pZHcxYSB+SuYEiF
WQ7ACo9Mprs7S0OFe+Pm49hhsw4ImH6FypA2tW2JfxE5EJZD5IhFBvqijXqnqLqH
3ODAzzCd1WUDdjsnyyW0RiuqpEMn9NdajGhAj3HYKPHJ7fjfYmWhfMFgk/Gt2fu1
OkMlRcbLpkQuHKdh0CYEg441+fR1Kj17mD8PikNAG9lxMbll3eFccfYeiXZSp4jL
eBmcLRXTGNekmt2p6XalWfY72IiwA7zLWRuXzAASukBSwdKCecUvm9kbWGw4rt+I
aeaxgJOKnITrbxG1Hnk8EydT8qvazeCIbPLjZCPeedoZl6snQ6AGqf0G8I8h5GXb
nM3fJhag0EzJ6A7SjOEfEpI2uU/7EGZkjOFHOnfvmc/kZYXP96NTdy8t0GEZ0BLK
XgTIzPZ281aGd9EW6HTvp2rdX/cQjXCGsXCXe9D/Lih3a9UCeZ8Nbm6jaDP9kfr1
TxLnFi78ltvWpsIo5P5mzfi6AKgS2Kd3XhkVV3EgvlJ0ZpZZkVCW/SPtV3oFBsve
f4/LBvydTOIEmTz90Ij6iRx/xwNnn8TCEovuLmupPmr63baIF4pjDVyYH9PkRY3/
LjuUlMxRL67wopgBpanZemDwjBYtcPbSGYGHC2WFh3L/Xx7BvmTf+xEw5LYdb+l2
YTI6RZw++zp5sLQ/OiC0YCO1U2AC+TXd6+p0GPHnFOwRLvktMuLRBfcSqvQeXljO
kNWKaWS5GIZfcZTYrJGeH0u3WJmnc+1sdxNqCBkC4wbJSNaR5/yyopZgNUHRKKGS
BjXPNVrn1OyP9vLRPMpnAmxxUcL6lJ7AjoYiIsM+X8bk3gxVdq3McrdTSmTPbYqB
6EiafI1hjNITx5NRyAa2aYHXEt/jVs2m+DBLM1v85tR6st5VVwFBWdghHRNAqM0W
h0/BVCl+UxpCju1e9Qb8D9HGtm6JHlVaN0JUAiYEIkzVaw6/DYkULZWIrNivlMny
qkLnvtNj3XCftEB0kJK03jLbmDAXXxpZaHR8eQPxTEkHjlXvWqzf6WZsKjfpjJ8z
wv8gatVG7iSMbLued9CIqVij+oVIejuP79KkoNz2i3uF1OynguXw9zupwacQIpYW
wxp52diTa3jAqEV080waKyNFoAhBdBGkd6Ub5tDQIgBNW31GudPkZM/u9AgPNlWI
RB+I7OT2FsqdQF5JgOw594sMIPJS6qPTop13kcPE3TfbjpsX32z/fX8G6zau7H/J
YU+IqpXgJOa/Pc9ALqer0N1D06k5zsT/1ipZSjh6IKr7o8AjCduWiaeN0p77mVjO
jWTe/bE1CU4mbKY5kOJaX0TOTBUyrph71c/uV/IKy8A7NwZRaNLkxUodIKUFHH/V
GcbnjKKxElaJvkE83rZZpB2g53VedQQA0WRCo3B8kszF6jxoA8w3HB1gUsFErKca
uo7g/ZIzXdusRoyvtt0d29E51E8VwGT9/hqq+87DeoM20EBQJ79CiPLGiX96FrOE
pEAyLT5Dz356fNjdi1ktCwix2swE7TNxhK+B25oXhJ5lVa2GblbXgJIViGVs/W2v
zfU0UV940pHq+lfx83ReaBXLmGW48ryDYJAUckjUCcg5Wyrfj95tGNKxBgIJKWFI
AvyDFA/luQ5Lx0cs2qnv5/8d02WLw4STM8e16BjgLi08VhNJsSphzq5z/UgMG9iz
kg2zqux8wguaI+8bBxN2IQC1wEsFSbJWVq7T7GbjlcV1qIzOgVy2DokQO90FcxWt
mS85nQqc6/6EytuX+eGxYULq+nR0L5Izsi/jIyOnB3M69Kc2OuA8nflRPrkHiiFK
qpnqASzXxh3+e1OVQ3wAwO5KSdMBDmg+DDsQr+WJ7fDO8H0d48Afeh1rbGmi80gX
7dHNx/DmBTImCDJNbckS76QOCD3tgZAQ0m1jKPENC9ZwxniUzURb1e/RyWC5SIQ3
NcPjDMOGddCiS0eSU5zy/TnGBSlq+Vsiz/fzXqdnoucEUXWrxLUmbKHX8OTJsM8Z
UYXrxBHpqzZksIizljB1eRjF4bTcThxX3Khy8gsc4LLZ0L8FnwcEU+ouf/u6OIF0
JiamGxZLY1YmjLe1duOTHS2idMkupuKgsLh0dkkozbvdhavZuZgxdwh0BGXgSZkM
s+WJxSt4BLsS8l6Ga7tPrjLOnYIw9W03dQUoyzJfsB0SW1HQ2Uz4sbmAiAyZoETO
scfkrFar4P5eg78kQMnPOPx2YPyMXzUOzniekLxWDNI7OrN0jLppp0BtxvybrQBU
wl2+7Ngb+3++dWA+5qx0T9wkRt46yS4B3zUpGiWuKpSGxXSzdKi+1baL392kIHR+
R2J3X4JAj540Gzqy6dkkOOH4iDkiSZDxXtRoQHJsnQv1oaWCVHbzdXxyHJK1ADz9
REQqKpCQ7OjtCooH0GFGvw==
`protect END_PROTECTED
