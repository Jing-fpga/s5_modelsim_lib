`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7FCzoF3mI13eg1YTQd3HJ10GHEFIodOkaQpfo9OMnacSZ6by3EDrt4SDGnETVxoq
T13RufiDcUaOq+CM5us/FBWCjfW9MB5rK00j5bLUTCpB1rxsxtuPQc8C6vx8ahHW
XUnCbA9a8IswIk2Di2OIcrLxoURMlU1APtpAWRXHlOSCZWT19TqDEojAby+QuT6R
6OXmkV1gTvGa0ng/91P+LP1/mqHRjz3FcIFGwIHsFP5ntHLWyt2YvEVWhvIN92uN
38HsBwTxbrOclwaX9H8ubWGZHSLUlf6YaAuhiHzkvCGzx6AQ990zEVC0ofghnYcs
FzJKMik5rDiszCE0deShBUCdGh11e3lpjKCOlj2PvHC8MkQiGkNhtM+bIwOAj7qL
xTjaarS4Rur5NivYWUicVqBLbwbpUORJbVYQkbiBKW9a4LzvclQwcoCu+2WSr9/l
dTosC703BIK5DrlWW3isKqxuDZd4LydR3K8wbZ81kNQ5PThhUjGhoB4T0L5+0Upy
AiBEY3ncMrhewY4tmU0txBv86ADhVq6uzAOpUZmabyOMsQZTMtDQqcPtcsfxXUU3
Yz+fzw0w6cb8qde1sO0dLZrcoL3zLH1UtvOjE/3NqH/kHEgrGElRDjwy1daTRddt
YeQ2Um05P2T7hfd5hajCGH5WSYaQ8l7owEnti+abrN7gqOLavyGC95mZwuLFoNz5
WnosyogREIqkno/0a2LEnx9/ro2fZPEd/cghpCWT4VyCcruGBF4REduxwIA8KpBE
fXXos1DUuuD211QPKplv9T/liSfYPTZez/N9zTW72GB/dENUxE8pNEYZIMr1ZVwp
J+MJU4hzhSkZAVKMcTp7VqW2Ilb0bLjF+x7hGDFQ6cGO9EcRKjLorpkrUfJQqoo8
RWNfrHQCS/jOwxiUvE5rWe99YwbaCe/UhzP3pYdEL1b3SJdI4gQhN+Dg3UFKkFt/
oGLoHwCShPIc1sYzURsD8emwm4O8G5/S0vkD6pYPrsG/qX95cBXxO2z+dlyrJFwF
K36vigLiE9EKRnYbd0F1XWR2MupkfxCVorr1moMQRu0s1iZaOseWqNbFyThJYkLD
tyNjc8ZOdy3/wpxzw7aU/Uko6Pdr21uzu1y0Ph96IUlLWEgLlDHn7UnNSwtg8EDa
8xPdEXYbjOYu0NiRJNlGWf4ppHou4NUCbrn2R678fm1PAVQygMZgu1o20lfrxTh1
YwHDI8xpMvlLGEoW84zRm8IuYYkwMwl6ABSFipOkSX/bi3LjGQJVxVeNjvqjhll7
mDXnsv0TZnwQf/velIzxxJukyRioGrVkHgd0RnmvvfXuHQQiwV0MEXWV8TQhC8D3
6O4Kaav7mrdqLUgmI/dGwoCelPDcP9PnmB/ZJ0rX75+1h6r4Es7024XRL6lVLvmC
e6eT+CBQY1NZ9dYg8mfwJXYP950WXNjyg82wIlphcX4kXB3kGbrg3WKCCjb2Teep
frpaO900Se8YFrn1Bcjsr0HpcgKle4b1RF4K2XZat8PqVtscggpms5kl/U3s3YhX
ifvNB4n2CyI5jFbj/QxFupyg/uWgIRz0TvFhVtDMBFRUXH/ZYYRDw+L7kulwF/qo
nJVYyI/huZEum0vS8uuqFopC8sYYeGnl5NAgufsoLStmqJTCtxutTJGi0ilaUW8j
/3CK4LIXSkSutwxcXtwRjtvX3pYYJdA3xhNpSPzEEQTFWGcxIEFZmAB6N1/qgnxU
gXjsBiB2btLkiAsb8RcIvq5EElYVsw/1qhIN1sVlV+JcIhiOuu22aL8LzBlKF02O
y46HYi1fF6QKI4gFMvShmUHeOtT3dD0ozpu1d2pj+1Q3tmHQl3mtdg+2we29Q2xI
jcvO+iN7vymGsNWesoQdWa6M3UYaQExouXzvvNRwK535cC0rIsJdF/nUBeZQrcfI
oZU0vm4xnkOavSJEs840/zPQpWJTDTRc/D4MaXpXSKPB9NNHo5hpHpF/oSIus8WN
dX8C+KlMN4/ddwbQmpY/oEkMiyoYH2o1n1x7FCO4+hAFCy7J9CVOXcBqICRPo0wl
qdsB599r45C82hW7sdEycSZC3M6XFHBv8atLPeEZQmxCbCNa7tFCu81Nt7ys/gfw
05P7wB/6PZCCyUti2cxLMPWsNfbPfIkgnl7nlVVljxj9DG9Md9JytYe4it2qkMJl
fd32FNLQmxTomCNmWJ0HwrhxbuUc4n6pnRbBZ0j6LyKrtU0KNuKY3/eaDSkFkNuV
M0xFJcSeHuKXePrb3/nqU5m7ma6WwcPZByEaqofovz0jsn/yViFw8mQkhPRNLVr+
lzAScZ47+C2PDttTcUF4b0ktV3IweM9rMkXyEYV1NBVtPjSFV+fZOKE/AACLqj6O
bYKXO9wNDoP0Y/fD1oT4IdbgaUzs1HQNbVKK3MMtP0XbqwX1W/F76FNkLn2b6Yuv
+Mjtl1GmNo3iK6GO0gCk2aAWECZU2OvTEOj/upHVCJZ5q5LoDQuLii4dmT4PIfey
4s56Mj5WIn9+nHAsxaAMz7ty+XC+ez16GbjyUyj7eBGwkFV3p0Ww6ypuV/Ii9xUM
WKgCDoAORddQuJu7fjqp4hWZ1xpwZ6F4G2MlPkuzuocx8gIWkntADJzSxS2QUQ0i
cwlNIQdj4lGcjFdKlLz1slBNGc6oXUhHBWJAU9t5KVg4XEE/16BZav2dPVvP77/Y
tmwvaxK8bLe31iM1fizea7nUcVKhLsh4xxrAjN5scxB6frHKxBD8RbduZoTPFFKN
`protect END_PROTECTED
