`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J3qfO7Bm4CuO+0mFIVVHqyaPQLvek1kP9mmwmr1/8FWHj6NfIO98G22CD3CO2Mhq
LIBMxv6aHBIOGENL6nCzAm9dZnKYp7A2wlu4VVX0e5L0bB5w7LNlZAihuaBEOEk/
Id0imSmBTiPkrubqrzn9mcI4J3pR1IUX5eokQzp/IIu9OUCPRwuoBJsNg7arBj39
Um3yagoAD3O2A9TOUIOMgt5O27Zg3Uwlx3Bm98MZhpk/R9ZKc/rrVV4eEVoNV7El
9bzX/FiudepzoSU18xX2hwRJiBBeg+9z2X5weRF4701idOsp3IQnbOJYNLlpxGxY
w/Rkmc2Rf8szjLa7jo2JVknnPlv6VNS8f5hVM2EIn/2aN770iBisbn2siNpOBKqj
ZKQwlOy11t3FkUj9syV9IY+y2eVZsAJZdGZR8SdtxL+3Yz/F9FHi1W01j4350Kne
ppg6Iyh5BAfMif6oUe3y6BcHjQrr4QgssiIQUnLpph5Nghi9G81X++uAMvBJwyiJ
ZoW+Ce09htYpFG7M5/iOfg==
`protect END_PROTECTED
