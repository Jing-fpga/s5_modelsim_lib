`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
No5jKJ8uL+kPrcdy/ervhxHXqnFOP0gWwjEmHWxExYjGu6+OutEpUQGGTDB6zf+f
NfSmBfQf3v0Z1O3D/onSqZ9yGKiFtjSGcajLVxCOe92dylSu7+I3YgCh6lYuM2UE
hXMiZW8zLC9AACDOfJoFJbP/k+jQGxn9lX+ljNLfMzkSFqNGKuZ4VUeb996mFhFW
5fl26o5jRSP+ekRsFzUJgx8copYwn5uRHTjL4bnBGcVdrrHsZ5vL9VOa6tlN6Xmh
XMwRajuHdxjVpm1uX6sK4XbYB9JwIJZ+rL75a63bdnLI8y/iFvlWmAFwPnLO2vIM
Ss2/121rRrDj0P5BkrQyFA360pHsWrQ6oOsw3ow70VnmU4uoSSy1ifjvaMyJhnDh
sF6in9a8qhzTuoNZqZvQ8gvHw1AB2+uQOOKcN3+CxpRhs7FQ+CRuSvaSvt1FWz4D
dlcQkPHp3r2AKZOJrK2RyanDOkBfnVXceDUIBDfYwJxvB1C8Xy9WGAoUcStfXN+O
twj4+CevL74UxziQrudFZAXBRpbju3G3Qqo/DM93+ISw9t12sK8y4Bbwtx9Fj7DN
+rsqHn71uGXosTSK6nb8kw5YbsKV72Mvy2/Pdzdf6AmQuDt1+NYv5QDt9dnV2Jfl
z8o3dhzO0LOH6MHNvxZx4CsBtwmiUAUNL6DVFcmOF8z/PatBvaZ5ww89RmGm67oy
kAZuMOQxkD693OPNgCi527pBdCEVhWITUsHLoC/WIBh4Utj7Q0s22q27MLU1rnZ5
yHOxgbuoJj+35xekEWUp/hAQ1Jngx9QONQH8Xlq5sW4=
`protect END_PROTECTED
