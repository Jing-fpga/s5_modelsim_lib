`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nH6xOsTFBk49NToAIfC9t1tCzD/LXRKz1pLDEN156GBDgy72KRTlIl0ZBs37lfcg
9OQJCH+Aq5mYiwIFfEwjj0P6wZv7bn4rUrsVeFV3g3O6wPTBQne1tazE50wIC5o1
qRZKDpJzObIPl3KylC2ilnvi/d2eHiuqUsyad9FPKu4eVMFV1F3VXJs7Qv8inPUu
fweUcf6PhOkS5AsyX4FyTktiK62HjoAExslgGBj+IDJ/e8NCBhQGcSMcvInob4T8
qVK7tW/GsFwN5dAJQ5KyXz7neWlrtpFdTH6VPzKpK7y4EDE+tXLHKf9wzWZH1EGX
TalWMwNZLAHmnr9d/ddjMbT7+gwZ4VQXSuvqT9A4MarCwMGw1RfuN+vOl8Vgvqj3
BB8+PDjQdrIEc4pp8+lTGxQJscvlCENRFkY1FOn3+gFWe9Z7ndAE8ji0FOVxr4ag
Vk0+ABV3+1PmK11SdIFuJGV7RbZqTuAPyYcm2ue8Lj0sZe4Qke6wiabmaVPXC5GK
s3EjRLGtzN5L9QduFVlBpDdln2OeyZX1EpCzKLYtAj80d9xZrufItemK1wSD3OFr
MVKP7X9qinlMBnH1+UO1NkhMWhOQk1bZA+fpugciYHfmoteO5lS1PY+aTrJpFA6X
/DnFAe2NsaGq2BNooHGKZsM7EMqHQ8MnifMLwM5IywMRX/9RJJmf/g2cLoUIIoVj
s2PykRMPs639kNTFSqvmvnnC2qZtZDsBdvB4QoDXewhtc6lelA4jYVAtvoGre3gy
2RSv7P79CiuoRel7H3Pq807/YS6dRaLvlCCzl8DSWKMhVC2JAlmmFW/sLvBSrRQb
Vpqd7aVMZ1u+aI8g/VDtCjjynSM4t1g+zWx7iS/dD+dDYm+Gi+AbM2WHqsixvPBz
wmHwz53NGfrxDL89ZCG8aP+SsTKlbZ6nKZKvlTl9IEwpLp9/hwDDNfIAdTjf/Eas
gIA2GWbUPQ3QQoScOldsH3aiF/xqjgXjAbUFwSf39YhufRkh0B7mm6NbnQVQge8x
5nSGtwvr/AGIyRDfPRX2yVptbN7Qvqll0sj71NF66GchOCqzgDF4jKOEFUz4A9Tz
Uc6ojL+IgKBAuMO7Bpsp+3iNJUHzA/ZUA3OFQ3pO39M6B+pRPsU3cEiBCTInU0Tt
Kj+krcgldHSMxv/NpeQA1X38vhvH2Ha8XEoqyHnB6K7NOijEWFv+NgFX+97d8Ehm
zsAD6XH6jMhJ+BTaH45Pa0Gf+vKlOE1YkGyRAbbM0WZFrHuGRuPPzKnPK5HY5bLC
NHZ9EU4w/IvzNF8s8JQaVwFnOPJ61pQ5emhxbVPyc5jVYnshdkBV5WcMhaikW7yJ
VQjESm50M5jRYarTsA7bXg==
`protect END_PROTECTED
