`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A9XWJftRoD+sAWn4fNBka2GEAq83onVNOfxx3dhxFJEQZ59sa29gq9lH9c1NvesM
W7rXJH8tSnDR612nxb+4mRSmSw9OkHzkv3KusSEFUnTh7T9XwSK8jarX58I4hP2I
0xBVx1wL566H0iu29+WwUc7glBnwahW1GgdLOJkzIfzd5GQm/oXzEJMkuQ/K0VOm
bezWMhcPFpB3NmRXPP61VKokonvASI9C+9TCgxX63JOHJuT9/Cc2pqUttSjxJZqb
6eudw8p/mcNIbiWCIH29I0k6mUwVOcEth8MfD2b2lnRCdr0bE6oLj7fFk441VqXi
E9gPqORm8BXXZLnBZOh9SmQtJGRpipJOCdPgTDmb8PPwtZw4EYjUf36O+ztjENmn
8Eb2ZSCDkfinfou7qRG8U1chiJ5Pjy/5Az0vlcoI5J8014nZ9oMqe9SCbFtJJtTh
jsCEwLk3/QhMYmTgzOi7VEuBc2i9jpqijpMC9rNgwd8fG13Hpf1RHm0eZxbRCCW9
cA71nGsoej7towP4qaFSsCz50f4o+zTwkon4hlojZ1t/AL/GxafGmzWy4Dyec/UZ
OibpTgwFqDHi+7hvNDI23HxdnI5r9WsHbt8+Hxcuo1bLJcKsRLZtw75cZqONGb0M
ARx4Quivo8pHuiFLU751L12BxIjZwgIxs9dy6UYlJ/B3SAlsxOEKH8V1+qxDvCFy
1VfyTw/J6BeJxRFfmuv/jiUIT9iOuB8RNmjmHe1IAA/k31B4MKN4MJQ++WxcT4tE
aIU9ViVwQ5heULYstkg/FwFfYP5rldfKgwsnJ4BaClAnIneLNRGoDpwidOKTIabI
JsVcrRR4lohv6ZBqLChPq3yihQblwHlx7TbWBIILoJkdn+YncCtFRjgYECz3w4Ym
hWTujpOT2JY0o29K1xyt6nNyMbYL/PKjsdglI/oaJvr2QOHmYsPM3BEkP3CI1Ztv
BaxZGy3+vEuaJWoVE/UxJWk4Vs6oGeAkkzXWCYxZQmrHfnsg+xnwbq2Rihc+xla6
xie2mm1PjyxAml4ZwX2LqMaqaSL8PWBysr49z/nU/w/v7Ta/GLkwyw0yE0p5awOR
P2YxIj8dPaS+GSnAR2MGFlN2hq16TCzmCUmGS3VZP/1wdTH9bIsa2ADcX7zeJrSo
AVeYJqri/+UNyddOf12cwzm3IZSXPALa6JRF0lyFfo5YLZ+S+IgaDu/+6WmV32px
oWpYcnKNcdzs0J4mTqVXek6iSB5JOuzbkZww6USLyb1JKnQVzmuyj4GHx6uBVMpV
q3vMKiQsggQeWsp1uqyHdbDBCA6eILde7Bsp7kSi4XO5IUNZZDU01lZQyxYrSqjp
udzISHgiD3CXtcUfiIBbVcCtCiXnHULQt3ysByapFE8iEOlvnGrH2Rk67zb0+G5S
3IeV1U8LDOyrIoFOodRRUiRs0eC70akUfkFwfjoDSTfBquuSk9ZZMc2PoDR+CZCP
zUQEt3gQcqrHZm3RdROYW2MfUly7wPDzkNqrLWFWs1LMuDK0Nez4q95VZF1MU2tZ
gECxh+vq9Rgsji7vHMif6hPQ04GUWKNNbKu0hd47xH3/jSdQcFnmq9kub4G1dCCS
`protect END_PROTECTED
