`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q02EscqUu8+tUoKislYp1gv6W/u5jfBB+UhUOjc3AeA9uLORs2qN6a97hHL2NejA
a/iZyVQS1GEFHYBGN2NlbrSvnLy+JB70kUZh36C2mkYvwDqlUwPHcIxG93Ty8lAF
mxamVEUdYGb8U1v7aJBgj/l7zm/xO1xFFY1CJCbRMM4qouXH1OncLAzLXLvVhs6S
EeUbd3wzxDmIAZucq80GoKOoMN+v18vXfA5lb1+cMmw6/ox+aOFlRhegLlbPdDDB
G2U3UMPkod5oBMA/LhX3tP166jNQrnW07LIGFS4xEUEZiGs5K7/hISfy5AItjnYj
AKDypotXmP7ylwqOpscgqUoZhLArzLo+LfGL0TsAN2VCq1IApuvQcHJQYMbP/eAA
UR5+ZcNF2IhrnTbbODPwylUL/kD7+W9Kr5O4ghvAbJaVbkeZqiAZyq0xW4kPdCPy
XKo0OXgQChxUtDhYkJPQVDqsMHW7nVO4DJ0nDHGMoMe1YBirausO98UiyOKc3beA
BbtjA/qCpNBPuoPjfD+0JFkAu4DdY9cbhGq9g6KhpomPwvTyyETs3YxfpiwAZn+j
wDU9akhH3bbRmMzxcchQVb2s2WXKjs08RXpdJspzn4wCh/3HfClmvQk8+OiikABo
f/zNKFqhrWZJQuG49L6+3gEOeKmGfeuo0lkkHpW7e2mM4/huyn0I+os2dGa3wGSn
/YfNPivWByBAdfIzo78UjXWPGR7i6KSMI3CvylSY8GjD9LP9fjnb/8XyjHJUbxtA
QqWSgL0309bZO+dWC6KgClt8TrliSnHGdgSzNlkKQUoZMFrmiZ8jHQ8/gElyNrST
IZ4C1SSv6hG1IZdfokEnCzGSJzF3ET89acgrFANjfq4ZCmszERM/aJsEd9Cin23U
fr1TqVTjutP3jOBdgAxQTVlWffwrhmel9rSlHQ//mAl3050QiecTp+VyMRDIoM8V
DfGf2uW6gYNanYObyNLerhKhk1cv/AyIv20/DlfIq+qvB7h6QW+muTww3cgmyX9V
ADeVUQqisZ5uJxsdDh8UVxzRmwm4n0Fu4dhSCoaeXNoyU5uMr5qGCE/8Y5pyNEtj
RiF0JC4IpUt/qTY2jCcn0K2G886hnzQ+V/r1ysaHyR7IvRlO9aIvDinYYWO/B3x+
kpmrDYaxTQPMynpDw0AYg1z/ZMXhksL3g7fOeOqYKfw0vDhMrI9uOkFFGVbity9C
zotl3QbkP0rS/IK8T2C6pnKeBXeoUSuviSRegscIa9B9TNQa3qBLLo4/7xfQgrHg
lGTWLQSdRP3qGq9eeOpgLNvBDNypLcTDtqZaidDDxkh0B+dhaKAGOGbpZoMAY7Cu
MQxyv5nsdWqaeMx7yWOWuo5mvLhLOdt4YA4dnERMR5KoyTaBM1uFuhvJg7FwxdDD
R2szr4BSkr0oQC7TRWNBp7it7wJqRvvz6Ngx96oCVq23zOtPyR8pzkqCUQuEjibs
k5wRnkUdjAJdA0aZb5t7gS0vwYfxgJtWWFLEt0p7Nd4N+uw3M8vrJZIw9tTk008W
cSAOc5ByIWszniz+pKRTzfFFNYnDnWVAvyAnxArfPcveRuRYfnvkiD0eNPU2jBC9
hnUMHpFajerSGGjX9ij8Vp6sU2IYqnMwbGVsqzFxbyqxO409QGIXbUHLku8fYQwc
68OwBH4MoDUCs6GFW1Sw3PGPsMgWu7utnd2Pc/rpwVYyzSyTMYL+pIRC585FoXiu
hZ7Q8jIeKobc4j0NN8Zaf7c4128Q8AaQXqf0EjujHoudM352tKndQtqf/aq9HV/z
xsaQFpMqZVVT/RoA8uq44j69JTRHfhN1z3zANc4MR+i60rlMCnvDWQu971UQl7mE
6I80v1mL/nZ88Zhxi+FQnqXl1zJrKi9Pt8LK+j4shUuNgh/Il/XRnzeLDTeTqhRi
BV94utf6G7f6PC7Ret02hMCneVgT9HZuOGxN3ShxnFMCjl8vRBdT6hAJZoon17t2
z9e/jB6hd+ZZimJsdMTOUEmuVhhswnupS79VXvKOCRYotosm9E+74ICkxzLPg5tt
yPbXRwivxutZySGBx0yK0jlzPZpySkaSty8ufl7maUtC7e6eMhv3Xi+B5xPc6zbO
uH+OAR64B2D/+PqZuJRw7vvTnfONikDAtsZndIRGKvMekMLP1qBOCfA3KFpRuNwd
H+UefN62i1yuQHaZgPbeIwS18VVFnRW01pHGLEJWmpbrU6tACPwwMze8OcSG2Sbs
UKiVQM9lLkotc0ig2dDDu5LCBLjWePUmfTqvxgvKiaclv1Gdjpgy5g11CaK975Xd
sa1Oprs6s7+pIgvonIEUwRMC/s4sA7vWfx/kBFxa0WrfqjrNk8iObUP2VaOSDr+e
`protect END_PROTECTED
