`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZSYudmPbMgCCs0FBrVsoWwcpB2Iy2zmm1wpXGcA8SLzTyCXb2lD5+3dyXbbjzyBo
clH1HTebJxaZXyPf+qqU37XeA0qKHRtHXK2/DWgsMsmiI/fgM3+2TAKu2xv7ZM9b
2f7R7DYrWZZfmULBCd4dRNPdhoSMCitFaj3ittXNS61501hOA9wsW+kJBct4zLsj
neKOliauhP6qPnwP3L8lgxS5ng/Itcbij2ZPUQyHiTJj4tmn34Qy1YLhDfPMiU30
IZVtMhrkXWw5PCPlPUefDcEU9kriQ+f1Cy56hvtGBS6Wf73EybaDAI3khcVLg0zO
7tyMJseNQeyiKJo9OWX2TMn198m8qfY0xv6bs50fE5F2lYKAqdEjiBkVNg37pXfr
ChgqW1c/5bnolerk55cpjB4ZsgPRrCp6DwPNl2j32qPb3V1f4Nk5w3M3sRj9JzNG
p/wbs3nkw8HZ5oajRU67lfkA+FBVmfkfTZnpmhS8fdNGQMT3z2SDtHO1mUk/WBKz
wdOtDW0rA7UMGETuePvHdyfPKprdvHbDMqsh87GXKS4RK1G0wtI0nINonFHeOUhm
IDfSv4QMU8rSpGBXONi8ozo3a1vFxl/oRQXyoVdmo2VSA6IdPm8XlHpCdoYtiyJ9
kbCVoHbqfirnFPRIFjZxl+dWeIlmso8Xalzbf5B33I3xpqidXqbCshFfS8HuDrQu
xEfkQP96tVoCNyYXJ7gxUDzkITK3nRNo8eHEumeldOLpF5V3I1QvKwPP49HuikIV
vQvsPAJ90P3/JVYRoTCqVU20LB8O3mYyUWRJp8qnbSry7li+7CwYTysKEmBy59Z7
YwDXy3zciF2KIq0yf0c/jnqMZN6S26kWIR6ekkg7YCpN/FWwUwVHgLc9Cre2XyDq
nutEfWS8H1+HUInxtour5/gsonZzhhcnH4Syyy7vxdyFAjrhDKuDJ3/eWbeI0hru
OD7VxIYF69s+xPtTG3WSskd5ey6jPLLP8GO3yCIGKDSlygYkU1oDruB22MgEXMPV
B8adHIIHzFqYIv52arYDb3DI4LgHzwa/mI4DR5wWJMSs7x7r208j7+oxc218/1wn
Idykm/3TPBAhRH5mNsJ2msSfTznQMV3uP9ErVpFoGfVYq31VZB7miwv6twhzwNmj
G9gQhXS89LHWUr3vswYy0/33DQqlya1Bq2/QsAlntzxPuC1S9w/B1oqZi1ve2o2L
gLk+GGmYd/5McMfAxTRce82QLp9umLljenLpEF066Ai7Ie1wmi4FGYu1NpSiHJBT
Gun5klftltf/tOPK77+WFLgBloRDgmgc6BUKguCBytIL6olEaxGBTx7C/KpssTLO
8w9yX7Q45d+9vzCa+3zWgE3ZN1goQYmoY1dL7in2KAiiBsI3e8C3ESuBnJsZ4YUR
tO0ShPecnIsIeGiXjBrEP+PmWFzrxHVrFh0rQZvuCBmx5mxctOwRmi1NX6I2jJa7
NmgB0RgrBc49+2fb7OTyMCiZjaC3oXN9VNevEkxU4KIKwKH+eNu8MGofJqn2CXAU
k81/dppfwtCge58g49rYeGtR7b9O7Jq/tjXYCKzW9dfRblSF1Z9QGWoerpleRCe4
ImapWBuuq+SLDT0rLeOkA2hBQTs+Is5T7yyRSlkdM0T/h1V0275dDdUWW+IJyjIx
IkFdXbnZmfA1Hc7iixborHids2rHthJ6gJuchFpHwyq/LbCb3mmzaBLjnN2nlffL
cTWy9rKHSc0QWxxnc39jMmGFju1g5gKblAxhOzqSo0prQCSA/m5613ER8BqE/Q32
bUqAwVAL8jnsHmMNC2TPSSCo5qniH1LuYrYMMmItGkTTOFme1yMvcq68zjWJ46Ba
U4IEINlWNNyCkSfadreogTBK9QYxc72FWhoqB6fuBW4QBzJOlkHIJhyhK25FlIuC
tHfd7cvkfIWrYI1IlyHge+/3PbVmTwrmbUg95sD8KQndWe3UXKZ8dMRq8Ad6DOaW
QyD55l31RTlzzdov3NVnK2YjLJvwOJwKQ9ljxDqqCy4C4gqdVbxkEhmrk2VofI7k
2i1T+gOve3XkAvl/JSZOPLhJ4dGt4v+vmOi1ITHJCCpn3urdoBSbBggfMu3U+psZ
GKexeIWtnDGoLTEoL+IkrC+Shkt/66vMIWOBx64oMsnoOQTQz0F/IOnNkxy76UIs
/vrzFdLcHLVNH5KchEIsBeAzj4zLKOF7CI39cXxCuXFTvmDOTFeAmobF+f3b+L7/
fY8lylwXGHy3S7LsUOvRPkWUpcGQKGFZ7u5fCpIbiORNNzWYQ/QxGarfllHVq20q
LakVcoJ8Fy+nURqLD69mciyOyFzTDZC/jx1lqZSc8g8hNK2AScSHwklxgLYHcCJc
r23yYKTPzWor1F4AoZnc95wQ2aX13GTa/9vDunoGvm92ASFhPGCYDM5HxIyOXT/B
7iWfC20G4Ef1EnjvRrqHvzAIY3LRpYfzZWttl3gnrw8W+0R5AINMPqlnPtO6l4KQ
vNE4N4h+P1ReEYq2AMSQqLwhUxGj8d1z44pCeiZUr4IMGfn5xsWqLapqq6PLDjI8
rXWzp2bUQ+x+/hkS8uNw2UUcDeFAuWnPcFFIc4mfFc29ygiC4wD1PESnKDLEth47
Qm+mlGx0Zu4Do0cBU37sNNxZ4Nx9BAi1D14nijkMqa+Jw9Lz79+f3+44FsXyhLjh
tYFIysqEdfXTK6BHzSfW2GHDK765zBB0CJRHdAKwNhSIeUZZxrMV6Qvqxsm8UcPk
Zlz+pkuZy/c3NUhnIFF9NTOM7YPgBiFRo1iJhcK4uchslTQA+0dvFyaf0cHhMA9r
VH79uuj3rTmjtbB+uQmwbCLB+VWSIfH2gZn0Ft/BDmHGwqMNEVEBe3EL/CSUWt5q
oPRqblTCvftKTnph7w+RTg==
`protect END_PROTECTED
