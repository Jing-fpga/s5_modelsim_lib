`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/JoP/DEEIEPsvxVnPhbxVXR1Ws+A0NcdC3dMHVQnCIZq2PbQsw6weTEJSGXIZXcu
f+2zY5PJvAdPkK+mq0A+isSWreRkllQKWA23q2IoizydAs0WSGJA+gWpR9sGQpLp
V5CSNEvcJs0SpC0C5zj4taPO2ypfg6Z06a150SKKdgFvdxwd5PD8CgVzpiM7YEIZ
K8D5uIOU4rXF6Q6H1kFfvacvWdURv6yr9b4b1dpS+72zWNUuTxYIJtqzlaoPzzFj
QugSspZLym0x/WkV2RjG2xXLBUmCm3ix1npao14in1zPvgC9Vn4hLMlMamzBtwdg
K41EPtAJPQ6wOqW5S/hhBxt0v8t9fZ8Zzgm5oHAMU4MPrEf3FH6qBEZbOoy5fI4I
UvNA/aI86RUeRg/TsITVNPB80ZxP8/8Y9R/OPsTsB+ms7g2l4HuER2canwvCJlkF
ChPnBV10rGIBHlgN2LTgSpNGMqR2mVvUwqjSr09jQLLH4cVjX/Xa0wKU3KrZAQYL
qFrLJkt05QUQjmXNLOmpK+8n0mdeOP6YlAgO1+nkjcwXBjpiJDJeFoOvFq6+kpPf
+y7+wIlIexPLEgTkZ4+nGiB7nfj7RMs6K0SSiomjGp+H8RErlAYuT1zaYaP2OaZZ
zrt5VGgf9H3ayTc9+IxkSZecnyg2TAanGSsntFJv8Zxw7dcqMn2pZE4ClbqxwbIg
iyzaHLUmC4jSl9XAS7Rn3/9sVxrefEq9Iw+9TPoByzMArwyov4CmQ3LjneqoFiWF
GgWt/VB3U8lhJBx3R0P1G3SnDy7uZQ4NGvJIf2Mp4v0Bz6qnqtiwin754KVv8NfY
n1jhV85TAGY9wvIIlSCeV3Jopge8Yvu6dviBh22ol2UXMOGqySo41WhxrqjgC71n
DzgJpGvCU++LoVfjLhSPrcCcNpUWcunXD6kzfTLURWidIdE526M+dclqfixyzDO9
JsmI1347FzX6jzsahDvarsVvHYJAoi7WjopSVNoU/l6eMs00VwDl6pDiD/oA9tkl
bZrnYdbhVoPAHET2Mk0xLvEbL2ggoYTsopv2zwhYRXbQyKIXtwY5vgEKAlHTo8w5
EkumXDXtmWZEucbLfdRJbCT4h1d6g+d1yNXDZqrjcRNc2Ke1ImZ0YKtcoVCOOr2M
W5g4Ty0txLu3cSf6mxhtYmwJPbo/AL1YfapLP7h04FMDtGwS5dinCRpXkdVyw9Oi
ICFF8QAxf215gI1JHVJHJjmGkMexIGYdIKLcp2p7zpcoCohdtbOFtX4SqIqSeJ5L
pr/iOq7ablWpFqF/NSPEirKLJrrCREzqVc7smSKGZIZkVnRU9u4IJWMUgVcrYFW6
Ri/PdnseqddK7zi844vJ7aVqgFCQ2y25CjYlNSB6lD9y/acMYCBvY/nIQgIZnP+O
7ftNnXRuppO/Pau1bv5L69L7WFjLjuPST/Vt6TI3GBCu9r5edJ4PAu0WWydvLv6/
R3YPZKDAP8s287WYQNyUQZMKGYOp9utdUqZNuNikqu7nD6nZaA63K7ykicwLQM8O
p3o9tO84cjY6QRVskg9YEkk2OmQGanSctN1sRTq4kfa+Pv8LRc79wmNIb899Gqiz
8mFdr5YnamjyqXAXqjrEXSrZquKDT83nRk9k/p2DbTf07caRRqc0Z0KwhCdsZGri
3XDJ5P2+cnYQ9tjmbE6eFjHLz1DhzmLzwCD9EQoVKQY0X8hGQ5cb5aeQiO3yrewz
C7IXYec8E3lQpSYK4kHTHUUEmQ7c8G7KsvwjAqcAoFbeqAYi6b6ZQjPx4ds4I3Ac
PQK+/qfoSvFM1hiBBoR0ejmo2T3elSf98xUaxsRWrUkeggCp1d8/PJIBmf7NxIA0
jMC8CsReTGQYSStJiM8AjeviYM8yX9qwjZW+7OGxgSMRx+mtnakTMxXmfkF9Yngt
nh69SSD0KLCN5KLJwRk4sFFJRlf8rNQJ/wlSmqbwD8rgcw2holiRYVlLEUDspJHA
xtB7RTUHZNdi7z8m7QTTwiGqHwxUyeVrWEp0sKOL0xJ2Bh/2gYHjV1+BWbvceG8n
LTyaydb8wwvFw1/2ydlpTztKb2o6hnPcXQre/1usFdPL4r8SraJZ4kAaQdZNPXo+
lwSY2Qe8Ei+mnuVdMMUNzRvfNocq0Bx5DHf7bApnYexE/VHmTMfveB/uVuGAVEd7
4Oe9INCLs3QPNFtWdVCdZoiSaFutfJGe5SnRgor4TyT8r+6B95m2KW0HMrRMjoqP
OFCOxJr1A+spHKgn/pY/fP3DyqkRmwOFPWm11n7OIO6zcZ0M4oGtwwL6sI514DEi
3e6ilN5liFH0uNA/G6NTaEPmwTr6uZNiXsBEW8t7wPrVKTzOgJa6gTgwPPXYNHm2
uvRsKGnD4AY0EQgz4qFkU+GLM2yeLiz/yTOykgfH/fOnFomjxZ3ubt10X1jL+2hb
pN1vcpzRMBT5Igw7tkBKN/0ZcfD0pOCjrtwEoiR5YtMezncpEv7Khx5dlxYSiUtP
VkjuGJujnrp7dS9QJFsDh+claAMymdTIYEpx7RlLh+4MucD4sm7G4pVbhEPudhYi
GZgF7HEDnEJ4WCDN6pLlqGqsN2sv+YgbJV+dsSG0fSJmgC92Et1DvEfsV+LltKSM
3sRfMraS9KR16T8SHbj4I9FhFkHFrXCllzRLulsl5OsmIWnBnZm7uZr42Kp+xKIh
10fdAUkpzAMuNdoHRkBxIdIQTksjZeqGOr+hJ8AF7R/zHxTVjTYS6qQQiRLOfN5y
A2ms6TON6RbwE2Us4mGW7yrXyvnw3bEitANrqoN+2CEtUOe3bQSFOy67lvc1zzHB
04/K1zAsvyD2yCIZWwA5ZtDbAoZGfXPZatQ2aJcUYP3latTTh88+6C4hIPCEMKgo
2ZHNG0fAafcjmRTw0pjh9O21Kqsh/TsXEEd3k33yV6ILDcNhRnVrDC+AkNDpePpr
gGRlCPFVvuRjl9D5h3U15uDr/iFOmw5zinSwB6TlwXw3BgdQ8XxIUZ1IqoQjPGkk
bZ9OFuNM3KIFTKYfos4Sb+fRdCj2I0B4fE4mPAmEV85Ph95DllLO58PXW/a72qKb
KqJUp5S0s7oA2b4mV1kTE9ixJjVqWjRZ5CmJkhv0EoWpX0ZB4Z1Zv3fyhPP7zH6N
5B76nFLloavnH0NKPzyJ/hGIyvTI4QCwNxbYQ5SyKMVRAjCPgPRR7US2VV6NgD1I
t942ruiUL1U5sMAn7g/x5J9BBzYkloohenlb1eH5D6AEIcgl84G/MGVNXpfV53jJ
xF87oWTtKFuFnfuFLBx71dy5tb0WmSQD6g29jWNUdXarko7C2xYESaHrOAcjRsEy
1FYIcjrwztuH/Q+Ec7kRx3TLsYtshKkpU50RM4iwgCpnaNAdDBAl5YjcxJz+v7Pe
H6S4hYXf8cIoy0ktCtT4foPW9K2nrlEsSm8YwNUAVD3qm9p3lM6Nw3TI5u93BbG6
w4hZgSdO3PXWf5tgzwq+NTPA31Qh4aGRCo/GwsAT5eYRj0J2F+4AYBKRJbgOO44Y
IHICZUwR5kCp8vzXYbopQzB19w13d0O40fdU7iySW0MqDEXVxsrlwZxTWgA8qJbm
Aud8OQH3Lrv7RAjfajRIFDKwfs0QaztnRgnKMWETTzCi+EZgsh/uIzY62FE5XeFW
A8LyxsTRLjUq0wckXg2zvp7uf+c7TssSsZhQ9tRniKnlt9VlKFOpXlx4nsbt0DgJ
GRUGjk9EpK3OZhGJabKdJRaKZSFAvHi5HnZpmkBcn58NFsxDUkVgbQTrQQkfRC6G
HJF3QcEoUM9R2yljdupGs91WpJct+UeQmheUBqnatIvI9+sdcN1p74Gn+PRtzxnF
FHS//K7+bXI0g3v5uE4+1GSYNOIqngOeEt/9fpvPzfjrOOnORTY9GJq/eUF0IuwO
N0KMKQCaHkgQ7iVEtdbISEQOFKXMCdfDTa1bSTtjPLoIiXgQP1VpagNBrnKCw+XH
VlPxVHbHODPMyrViR3SkpKWtihhvqN9OSjm6GYpBFV54NECmoKiA9qFfeZM4hKjy
yOJzSV9Dj1gYUsHpelHbkgStcV79v66bxPyHEF5cTOpd9DUbWJ9ovUb6YM1b2WFJ
2kyGjiTGK5byAgIhYWRNrb5T5CQvpM4iGUdelh5zOVIicjwyD749GVbz6R1HvOmZ
74Xx5iyGgr8c7aMdUiCwIJV64FzceU9uBn//chHtnkDCw2JNbIjjzzoxJs5k/bG9
He5rBaSKugFXQMN3f8UJySGJkaMHqmZO5Qf7nmCiLTUat29kelYp1JsCK8iqyJFe
fb6aRpTeyi/bjPxuIgruwI1qxsb43OldgBPU14swUkj1P3r7ixmj1+puqUhFBycZ
T6ggjDSsH9WCvLtqM5wpEcs3sdiYdvdeyNzsKq98kp+j0SeM9LSimNWdKhTSj6BX
ZxAuWQ3uOUlmCSjwSdX4xqsM/VLub9PhInlB4TsaTiEueE2GCfRJB5YVpetKWhJU
PBzqNpskGbbhkTiw7HodK2bcMt1dD+YSMeQqv1RYps/sTW+vHtbPo9kOJnppWntT
tcZVWB+hXliH88S72GcJ/YH0Uh9+n886fRADiOk93Fkar6qINn+37Jm+/Mu+4G9N
pxvbKeqLU9QENkLCR4wUUjWlN4Zh7+nHATcEkOlQ+g+dFwB0wrPy9o7blqIPQ7Ei
DINmIP+lCxvnTk6T4X5ZEdTBmVE/f1Y/fSHyqQczekJ2ebuEkpOg88H/Xe7vxvbS
MnaxPJ1uPTKdAmmE2l1uuq2twwN5mOXuXGWyq/S7a829Aiyrq57f2Rr8wuzkqBnO
OG7qv1ptGwh92wvFvahGulWWzd9QRiRK+AUAHkXKWtNfXJ/UYlhT9DVZCNZPWZl5
+w2HM5HZtoq2REz7IciePIRMvwE2vYhlqSEaYpCgE7Dl9HnbzN5F8Jvz+Pj/dS4l
7lxvWinBkArhMZwU4bwMbFsAxgO1+676lM7Hb0Ra6NKR9MIVOZxLHIu00FmcAS/q
vauLb16SDgENLR2qXzjc9kCDKh1xD8qh9+mgRBAKV7v6Zzdumkt3sK+ZWpXhPHEN
p8+DG6ejK5JFyDNRCRQDEuuIpJ9WthSidlrjga/p+YpVGlNJp0QbAYhcM7O9YDGk
kb5eZOvacWD7CESfqTUhXFmIlkSflw2GdYHGs2hHNRb7wbAFnwVvR3T5Ox7PlKnx
fsWB6YMlPGGqtiSMboCaFNOcza8HzrpbYBwUJW0zKnsXh5eDoMqCJKufc4kDaZ8j
HUEzgQonoqaAPQVKF8hw3X50kIJ3MyNIXUXtLTklbWv2tubnxlF9+yIgt3Ar7OLD
fdLbFMLUM/zo11g7tdB9CBVA7CnkDVs1SWbabl9B2rXr91aHa8gqfebTe4b2QcYN
B4R02mHBDP10ay4KaeamNDBjOf2FvJ8Zbdd+i5HcgZkrBO+qzasB7Yy0f9pPArt0
CHzFQ1dt+orwSG5b06gB156uKtiaGeXXkebxTHcMQwHW7+XYdlbnnQ3uPiG5Z3Ef
Y2n7+jhU9C1aZxuSn+H65gg7qLB6nlp3wPFq3EpxJuAc0yPBOfp7GFPNuYnEC0ja
mkBCn/mj+uk7FPWJuDWBVkTlmwgrdbhfWZRZHxrvhyoVq5Nch4FTQFjcUSoCNmxT
owUE3Ek+4qIYelvwodNN8TJkUpLf/9r7cG4i7kDfTlUIHVRffk8OeurXl+mDL+Te
3/sgGIGFTY8olwbo6jbXO+MvgrFcfVkzRfCr0D+XF4Jo7T6ZkU/w4sxxNOWNJEFA
De4voMzFxcCGapJ1C0Jq4tY5pKAaT1ReuWXl11an/NZTb/ewr9jTh0tNSBQbNTjm
k0ENc0pE3u2aI+gJcvAm3mJPgtjes5/b/YAm9+A0B7sD2apdXyWZijyE2NPg69tc
ORKXxRPALv5qgI25rPssxRIFJlfJpHD3DfQDmvEKr8Ci56HOw2KHMILe6Te9qNwN
ScUYVqrlYCQB0AY8X6ZkCqXLPW4+kpPNh96jgqX2pkKh8d5H4XSrBFNmxWLzOkmV
iGUgik4kitWmF+Nt19ZUTaSMC/ITCQStdoqsC5GaiI19FGG0c5vIWPCpS+/vxeQq
qIiLhn+YeLyK3Byy5TOv8+OaAb+UqdUT22TrrS3HgS+xyVL4Eyv4cM3zaxw6cH7d
Mi3MX5tiftDMuHRU1RtZ5ohZpxnQQtxsHVF9pxQ2AlWqZqVYMfkZyXNXhnpwgf+V
8jUmRvAs99uG1S/HTqb/4qcXpThiJCMX/nB/Q8tqX427hg+bOBZmqHvP8K8f5IJE
So511Ai4HT3tjLj1vqzhMxIJDS87VnPuCrtGpBRNVCA+8kuHMk7hOdZEldKL3Q4o
irLwliVz0aI00/HwAb1l+KpFDwl99LQxv+NtQVnERlgeBX9woh/4m3jC0bO0avY3
87vuBMDJt2AaBDgT5q42h5MEe9Wk9AmdSzqjgwJ65xoL9ycWGjuVXHgSWkvxEFvm
+VHaTQml+A9dKRKi/slo2yobkuFkuSOUG94lONAAWCR4/BQaTbb8oTgrMBOsiT8Y
AezMoRpPtAGy8f/lNZlfvshtkfAwkGWYFQkxmguUiWDo1jFb4o+iaF26xvXdeYLZ
HXO6xPOakQiPbl60by78CpAma3vlXNKXB7PF+tRULJ+CADtujK+KSoOP0yQYdvQU
xxztZBmhjMirbOuZn/SVg6NvIfeumKIo+srqutzHcIaoOftv83PRTX9g2SmFAtoz
faUuPOqqcD0vUti3V/AzAm/vccuy0AK/Zc7oHa2ZCuOPkNMJSLHHJ0czJ3XKxkk2
9OwR5XSuX6HHMtGvYV1E/KdW26qZl3KLR8ZHEkAhffHByoIYe/gd0aM/S9uDRxl5
dOp+gn/cW61t7hsamYUF6dODtwNCe9jTI1CShK+GjfcaFYmxeLcj2wVX3ZrW6x8E
QttlyogUaBILxg90vaYo3FtNicMBC3KDEPvxuFuTOpsmpSkUKzdVCXlbhgQrifi5
9vN60QKFe+VsPdOLq+81nvt4ybtYW4dGgEA1hXv8cgyTAk1e/RDtQCdW/D9MpbzB
sq351QKya7pt/y95z+DPlABAAKYysY1234OoIH72nAWzWkNxsMM9a7gji+jRl2Ms
UOw8s3GrRYwZPkYkyMIZP1WFaxGlHa8m0439rePs1NI=
`protect END_PROTECTED
