`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SK05vTPEHA45SQkyKRTUfO0s6AwfqcM+Z6ktIwq/gg/v0b6XrrudyBrqOOmPd7Cc
CBukyx/ZIw90KutTD30yytLKveSdQREe2ZesxchDfBnNPEUrWt6MYW9AY/FT3Z2h
iafSiNBMzq3qrlWkUb+3GWWxPFLPhp5csFWBbJ0UKcHAxhDJTk11YQbLIju9o6qv
Crauj/eWsN0nFq5K8m90Ti96qzlRNmEsMXTbFm192dd64mbu9xpMQktypxlgoZlA
QoEg3eJQbz72LTFPyXPwuU/RyD3bEPPYwNzgLqTCmsljLS3XUHl9IAWS1W/fEAxW
ceKJsiUErv0J+a54Fle5/NR849/PstHQo8ja0OYq0QvmctDf0h5LhuNBKy8sdVs0
yE/Rd4hWy+V3WWv0bTXOMPDWWok/QrXILwL/AsHJr4RAEEs70j0N7a1BjZZ8iNcI
aW4rw/pyndoc9dZTWrP7/1EuNhVX8k19C58vaH/Ysbi73L6TtAUvd8A2/wxVEJur
JogyM8XQU3Ly29tG+0D1FvAIFSJp7sDNOkBzJV1LDiM6aS7i21UDmRw+9D+xO7jQ
xQnzOpSL3b+gUzTtJXt68F4G6lSvqrYbqV97i3qBmZaB5NBKigc/tDrHVh79ZM4b
iJIcqDHgbbt+hg1kNojxzN8u4iiT+41eRtU096SNc4euMWfC+SvLMgCoN0dhNIUn
AlLFeZYkRU1tPTHFx9biC8cKIxqYuNPkxc7jwUi1dARqRJNDmTwLFrla/wYMlkGR
kqW8YCvUaOClSPn1hqhRYVmgkTLfbTfrkHHkrrsQwuk=
`protect END_PROTECTED
