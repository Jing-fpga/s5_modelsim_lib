library verilog;
use verilog.vl_types.all;
entity stratixiv_pciehip_param is
    generic(
        advanced_errors : string  := "false";
        allow_rx_valid_empty: string  := "false";
        bar0_64bit_mem_space: string  := "true";
        bar0_io_space   : string  := "false";
        bar0_prefetchable: string  := "true";
        bar0_size_mask  : integer := 32;
        bar1_64bit_mem_space: string  := "false";
        bar1_io_space   : string  := "false";
        bar1_prefetchable: string  := "false";
        bar1_size_mask  : integer := 4;
        bar2_64bit_mem_space: string  := "false";
        bar2_io_space   : string  := "false";
        bar2_prefetchable: string  := "false";
        bar2_size_mask  : integer := 4;
        bar3_64bit_mem_space: string  := "false";
        bar3_io_space   : string  := "false";
        bar3_prefetchable: string  := "false";
        bar3_size_mask  : integer := 4;
        bar4_64bit_mem_space: string  := "false";
        bar4_io_space   : string  := "false";
        bar4_prefetchable: string  := "false";
        bar4_size_mask  : integer := 4;
        bar5_64bit_mem_space: string  := "false";
        bar5_io_space   : string  := "false";
        bar5_prefetchable: string  := "false";
        bar5_size_mask  : integer := 4;
        bar_io_window_size: string  := "NONE";
        bar_prefetchable: integer := 0;
        base_address    : integer := 0;
        bridge_port_ssid_support: string  := "false";
        bridge_port_vga_enable: string  := "false";
        bypass_cdc      : string  := "false";
        bypass_tl       : string  := "false";
        class_code      : integer := 16711680;
        completion_timeout: string  := "ABCD";
        core_clk_divider: integer := 1;
        core_clk_source : string  := "PLL_FIXED_CLK";
        credit_buffer_allocation_aux: string  := "BALANCED";
        deemphasis_enable: string  := "false";
        device_address  : integer := 0;
        device_id       : integer := 1;
        device_number   : integer := 0;
        diffclock_nfts_count: integer := 128;
        disable_cdc_clk_ppm: string  := "true";
        disable_async_l2_logic: string  := "false";
        disable_link_x2_support: string  := "false";
        disable_snoop_packet: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        dll_active_report_support: string  := "false";
        ei_delay_powerdown_count: integer := 10;
        eie_before_nfts_count: integer := 4;
        enable_adapter_half_rate_mode: string  := "false";
        enable_ch0_pclk_out: string  := "true";
        enable_completion_timeout_disable: string  := "true";
        enable_coreclk_out_half_rate: string  := "false";
        enable_ecrc_check: string  := "true";
        enable_ecrc_gen : string  := "true";
        enable_function_msi_support: string  := "true";
        enable_function_msix_support: string  := "false";
        enable_gen2_core: string  := "true";
        enable_hip_x1_loopback: string  := "false";
        enable_l1_aspm  : string  := "false";
        enable_msi_64bit_addressing: string  := "true";
        enable_msi_masking: string  := "false";
        enable_rcv0buf_a_we: string  := "true";
        enable_rcv0buf_b_re: string  := "true";
        enable_rcv0buf_output_regs: string  := "false";
        enable_rcv1buf_a_we: string  := "true";
        enable_rcv1buf_b_re: string  := "true";
        enable_rcv1buf_output_regs: string  := "false";
        enable_retrybuf_a_we: string  := "true";
        enable_retrybuf_b_re: string  := "true";
        enable_retrybuf_ecc: string  := "false";
        enable_retrybuf_output_regs: string  := "false";
        enable_retrybuf_x8_clk_stealing: integer := 0;
        enable_rx0buf_ecc: string  := "false";
        enable_rx0buf_x8_clk_stealing: integer := 0;
        enable_rx1buf_ecc: string  := "false";
        enable_rx1buf_x8_clk_stealing: integer := 0;
        enable_rx_buffer_checking: string  := "false";
        enable_rx_ei_l0s_exit_refined: string  := "false";
        enable_rx_reordering: string  := "true";
        enable_slot_register: string  := "false";
        endpoint_l0_latency: integer := 0;
        endpoint_l1_latency: integer := 0;
        expansion_base_address_register: integer := 0;
        extend_tag_field: string  := "false";
        fc_init_timer   : integer := 1024;
        flow_control_timeout_count: integer := 200;
        flow_control_update_count: integer := 30;
        gen2_diffclock_nfts_count: integer := 255;
        gen2_lane_rate_mode: string  := "false";
        gen2_sameclock_nfts_count: integer := 255;
        hot_plug_support: vl_logic_vector(0 to 6) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        iei_logic       : string  := "DISABLE";
        indicator       : integer := 7;
        l01_entry_latency: integer := 31;
        l0_exit_latency_diffclock: integer := 6;
        l0_exit_latency_sameclock: integer := 6;
        l1_exit_latency_diffclock: integer := 0;
        l1_exit_latency_sameclock: integer := 0;
        lane_mask       : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        low_priority_vc : integer := 0;
        max_link_width  : integer := 4;
        max_payload_size: integer := 2;
        maximum_current : integer := 0;
        migrated_from_prev_family: string  := "false";
        millisecond_cycle_count: integer := 0;
        mram_bist_settings: string  := "";
        msi_function_count: integer := 2;
        msix_pba_bir    : integer := 0;
        msix_pba_offset : integer := 0;
        msix_table_bir  : integer := 0;
        msix_table_offset: integer := 0;
        msix_table_size : integer := 0;
        no_command_completed: string  := "true";
        no_soft_reset   : string  := "false";
        pcie_mode       : string  := "SHARED_MODE";
        pme_state_enable: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        port_link_number: integer := 1;
        port_address    : integer := 0;
        register_pipe_signals: string  := "false";
        retry_buffer_last_active_address: integer := 4095;
        retry_buffer_memory_settings: integer := 0;
        revision_id     : integer := 1;
        rx0_adap_fifo_full_value: integer := 9;
        rx1_adap_fifo_full_value: integer := 9;
        rx_cdc_full_value: integer := 12;
        rx_idl_os_count : integer := 0;
        rx_ptr0_nonposted_dpram_max: integer := 0;
        rx_ptr0_nonposted_dpram_min: integer := 0;
        rx_ptr0_posted_dpram_max: integer := 0;
        rx_ptr0_posted_dpram_min: integer := 0;
        rx_ptr1_nonposted_dpram_max: integer := 0;
        rx_ptr1_nonposted_dpram_min: integer := 0;
        rx_ptr1_posted_dpram_max: integer := 0;
        rx_ptr1_posted_dpram_min: integer := 0;
        sameclock_nfts_count: integer := 128;
        single_rx_detect: integer := 0;
        skp_os_schedule_count: integer := 0;
        slot_number     : integer := 0;
        slot_power_limit: integer := 0;
        slot_power_scale: integer := 0;
        ssid            : integer := 0;
        ssvid           : integer := 0;
        subsystem_device_id: integer := 1;
        subsystem_vendor_id: integer := 4466;
        surprise_down_error_support: string  := "false";
        tx0_adap_fifo_full_value: integer := 11;
        tx1_adap_fifo_full_value: integer := 11;
        tx_cdc_full_value: integer := 12;
        tx_cdc_stop_dummy_full_value: integer := 11;
        use_crc_forwarding: string  := "false";
        vc0_clk_enable  : string  := "true";
        vc0_rx_buffer_memory_settings: integer := 0;
        vc0_rx_flow_ctrl_compl_data: integer := 448;
        vc0_rx_flow_ctrl_compl_header: integer := 112;
        vc0_rx_flow_ctrl_nonposted_data: integer := 0;
        vc0_rx_flow_ctrl_nonposted_header: integer := 54;
        vc0_rx_flow_ctrl_posted_data: integer := 360;
        vc0_rx_flow_ctrl_posted_header: integer := 50;
        vc1_clk_enable  : string  := "false";
        vc1_rx_buffer_memory_settings: integer := 0;
        vc1_rx_flow_ctrl_compl_data: integer := 448;
        vc1_rx_flow_ctrl_compl_header: integer := 112;
        vc1_rx_flow_ctrl_nonposted_data: integer := 0;
        vc1_rx_flow_ctrl_nonposted_header: integer := 54;
        vc1_rx_flow_ctrl_posted_data: integer := 360;
        vc1_rx_flow_ctrl_posted_header: integer := 50;
        vc_arbitration  : integer := 1;
        vc_enable       : vl_logic_vector(0 to 6) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        vendor_id       : integer := 4466
    );
    port(
        test_in         : in     vl_logic;
        csr_hip_in      : out    vl_logic_vector(1759 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of advanced_errors : constant is 1;
    attribute mti_svvh_generic_type of allow_rx_valid_empty : constant is 1;
    attribute mti_svvh_generic_type of bar0_64bit_mem_space : constant is 1;
    attribute mti_svvh_generic_type of bar0_io_space : constant is 1;
    attribute mti_svvh_generic_type of bar0_prefetchable : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar1_64bit_mem_space : constant is 1;
    attribute mti_svvh_generic_type of bar1_io_space : constant is 1;
    attribute mti_svvh_generic_type of bar1_prefetchable : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar2_64bit_mem_space : constant is 1;
    attribute mti_svvh_generic_type of bar2_io_space : constant is 1;
    attribute mti_svvh_generic_type of bar2_prefetchable : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar3_64bit_mem_space : constant is 1;
    attribute mti_svvh_generic_type of bar3_io_space : constant is 1;
    attribute mti_svvh_generic_type of bar3_prefetchable : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar4_64bit_mem_space : constant is 1;
    attribute mti_svvh_generic_type of bar4_io_space : constant is 1;
    attribute mti_svvh_generic_type of bar4_prefetchable : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar5_64bit_mem_space : constant is 1;
    attribute mti_svvh_generic_type of bar5_io_space : constant is 1;
    attribute mti_svvh_generic_type of bar5_prefetchable : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar_io_window_size : constant is 1;
    attribute mti_svvh_generic_type of bar_prefetchable : constant is 1;
    attribute mti_svvh_generic_type of base_address : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_ssid_support : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_vga_enable : constant is 1;
    attribute mti_svvh_generic_type of bypass_cdc : constant is 1;
    attribute mti_svvh_generic_type of bypass_tl : constant is 1;
    attribute mti_svvh_generic_type of class_code : constant is 1;
    attribute mti_svvh_generic_type of completion_timeout : constant is 1;
    attribute mti_svvh_generic_type of core_clk_divider : constant is 1;
    attribute mti_svvh_generic_type of core_clk_source : constant is 1;
    attribute mti_svvh_generic_type of credit_buffer_allocation_aux : constant is 1;
    attribute mti_svvh_generic_type of deemphasis_enable : constant is 1;
    attribute mti_svvh_generic_type of device_address : constant is 1;
    attribute mti_svvh_generic_type of device_id : constant is 1;
    attribute mti_svvh_generic_type of device_number : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of disable_cdc_clk_ppm : constant is 1;
    attribute mti_svvh_generic_type of disable_async_l2_logic : constant is 1;
    attribute mti_svvh_generic_type of disable_link_x2_support : constant is 1;
    attribute mti_svvh_generic_type of disable_snoop_packet : constant is 1;
    attribute mti_svvh_generic_type of dll_active_report_support : constant is 1;
    attribute mti_svvh_generic_type of ei_delay_powerdown_count : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of enable_adapter_half_rate_mode : constant is 1;
    attribute mti_svvh_generic_type of enable_ch0_pclk_out : constant is 1;
    attribute mti_svvh_generic_type of enable_completion_timeout_disable : constant is 1;
    attribute mti_svvh_generic_type of enable_coreclk_out_half_rate : constant is 1;
    attribute mti_svvh_generic_type of enable_ecrc_check : constant is 1;
    attribute mti_svvh_generic_type of enable_ecrc_gen : constant is 1;
    attribute mti_svvh_generic_type of enable_function_msi_support : constant is 1;
    attribute mti_svvh_generic_type of enable_function_msix_support : constant is 1;
    attribute mti_svvh_generic_type of enable_gen2_core : constant is 1;
    attribute mti_svvh_generic_type of enable_hip_x1_loopback : constant is 1;
    attribute mti_svvh_generic_type of enable_l1_aspm : constant is 1;
    attribute mti_svvh_generic_type of enable_msi_64bit_addressing : constant is 1;
    attribute mti_svvh_generic_type of enable_msi_masking : constant is 1;
    attribute mti_svvh_generic_type of enable_rcv0buf_a_we : constant is 1;
    attribute mti_svvh_generic_type of enable_rcv0buf_b_re : constant is 1;
    attribute mti_svvh_generic_type of enable_rcv0buf_output_regs : constant is 1;
    attribute mti_svvh_generic_type of enable_rcv1buf_a_we : constant is 1;
    attribute mti_svvh_generic_type of enable_rcv1buf_b_re : constant is 1;
    attribute mti_svvh_generic_type of enable_rcv1buf_output_regs : constant is 1;
    attribute mti_svvh_generic_type of enable_retrybuf_a_we : constant is 1;
    attribute mti_svvh_generic_type of enable_retrybuf_b_re : constant is 1;
    attribute mti_svvh_generic_type of enable_retrybuf_ecc : constant is 1;
    attribute mti_svvh_generic_type of enable_retrybuf_output_regs : constant is 1;
    attribute mti_svvh_generic_type of enable_retrybuf_x8_clk_stealing : constant is 1;
    attribute mti_svvh_generic_type of enable_rx0buf_ecc : constant is 1;
    attribute mti_svvh_generic_type of enable_rx0buf_x8_clk_stealing : constant is 1;
    attribute mti_svvh_generic_type of enable_rx1buf_ecc : constant is 1;
    attribute mti_svvh_generic_type of enable_rx1buf_x8_clk_stealing : constant is 1;
    attribute mti_svvh_generic_type of enable_rx_buffer_checking : constant is 1;
    attribute mti_svvh_generic_type of enable_rx_ei_l0s_exit_refined : constant is 1;
    attribute mti_svvh_generic_type of enable_rx_reordering : constant is 1;
    attribute mti_svvh_generic_type of enable_slot_register : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register : constant is 1;
    attribute mti_svvh_generic_type of extend_tag_field : constant is 1;
    attribute mti_svvh_generic_type of fc_init_timer : constant is 1;
    attribute mti_svvh_generic_type of flow_control_timeout_count : constant is 1;
    attribute mti_svvh_generic_type of flow_control_update_count : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of gen2_lane_rate_mode : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support : constant is 1;
    attribute mti_svvh_generic_type of iei_logic : constant is 1;
    attribute mti_svvh_generic_type of indicator : constant is 1;
    attribute mti_svvh_generic_type of l01_entry_latency : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock : constant is 1;
    attribute mti_svvh_generic_type of lane_mask : constant is 1;
    attribute mti_svvh_generic_type of low_priority_vc : constant is 1;
    attribute mti_svvh_generic_type of max_link_width : constant is 1;
    attribute mti_svvh_generic_type of max_payload_size : constant is 1;
    attribute mti_svvh_generic_type of maximum_current : constant is 1;
    attribute mti_svvh_generic_type of migrated_from_prev_family : constant is 1;
    attribute mti_svvh_generic_type of millisecond_cycle_count : constant is 1;
    attribute mti_svvh_generic_type of mram_bist_settings : constant is 1;
    attribute mti_svvh_generic_type of msi_function_count : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size : constant is 1;
    attribute mti_svvh_generic_type of no_command_completed : constant is 1;
    attribute mti_svvh_generic_type of no_soft_reset : constant is 1;
    attribute mti_svvh_generic_type of pcie_mode : constant is 1;
    attribute mti_svvh_generic_type of pme_state_enable : constant is 1;
    attribute mti_svvh_generic_type of port_link_number : constant is 1;
    attribute mti_svvh_generic_type of port_address : constant is 1;
    attribute mti_svvh_generic_type of register_pipe_signals : constant is 1;
    attribute mti_svvh_generic_type of retry_buffer_last_active_address : constant is 1;
    attribute mti_svvh_generic_type of retry_buffer_memory_settings : constant is 1;
    attribute mti_svvh_generic_type of revision_id : constant is 1;
    attribute mti_svvh_generic_type of rx0_adap_fifo_full_value : constant is 1;
    attribute mti_svvh_generic_type of rx1_adap_fifo_full_value : constant is 1;
    attribute mti_svvh_generic_type of rx_cdc_full_value : constant is 1;
    attribute mti_svvh_generic_type of rx_idl_os_count : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_nonposted_dpram_max : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_nonposted_dpram_min : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_posted_dpram_max : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_posted_dpram_min : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr1_nonposted_dpram_max : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr1_nonposted_dpram_min : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr1_posted_dpram_max : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr1_posted_dpram_min : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of single_rx_detect : constant is 1;
    attribute mti_svvh_generic_type of skp_os_schedule_count : constant is 1;
    attribute mti_svvh_generic_type of slot_number : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale : constant is 1;
    attribute mti_svvh_generic_type of ssid : constant is 1;
    attribute mti_svvh_generic_type of ssvid : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id : constant is 1;
    attribute mti_svvh_generic_type of surprise_down_error_support : constant is 1;
    attribute mti_svvh_generic_type of tx0_adap_fifo_full_value : constant is 1;
    attribute mti_svvh_generic_type of tx1_adap_fifo_full_value : constant is 1;
    attribute mti_svvh_generic_type of tx_cdc_full_value : constant is 1;
    attribute mti_svvh_generic_type of tx_cdc_stop_dummy_full_value : constant is 1;
    attribute mti_svvh_generic_type of use_crc_forwarding : constant is 1;
    attribute mti_svvh_generic_type of vc0_clk_enable : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_buffer_memory_settings : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_compl_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_compl_header : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_nonposted_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_nonposted_header : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_posted_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_posted_header : constant is 1;
    attribute mti_svvh_generic_type of vc1_clk_enable : constant is 1;
    attribute mti_svvh_generic_type of vc1_rx_buffer_memory_settings : constant is 1;
    attribute mti_svvh_generic_type of vc1_rx_flow_ctrl_compl_data : constant is 1;
    attribute mti_svvh_generic_type of vc1_rx_flow_ctrl_compl_header : constant is 1;
    attribute mti_svvh_generic_type of vc1_rx_flow_ctrl_nonposted_data : constant is 1;
    attribute mti_svvh_generic_type of vc1_rx_flow_ctrl_nonposted_header : constant is 1;
    attribute mti_svvh_generic_type of vc1_rx_flow_ctrl_posted_data : constant is 1;
    attribute mti_svvh_generic_type of vc1_rx_flow_ctrl_posted_header : constant is 1;
    attribute mti_svvh_generic_type of vc_arbitration : constant is 1;
    attribute mti_svvh_generic_type of vc_enable : constant is 1;
    attribute mti_svvh_generic_type of vendor_id : constant is 1;
end stratixiv_pciehip_param;
