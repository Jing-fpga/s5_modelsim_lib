`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZuCivGEi5iVSIaFYKYH2VIfW8iXQJ9y5u8weR/dxpUFbVgvY5SynHSjQ/d9cFpsw
O/ygoe8YLK/VRXli3YqvO3Q+xdQ8NeL9EWCjYBkZ/xmKJ1s1Csyb/RJR88U6q+DI
SBWRfd+lLxd8caZ126qwr/2sAv3gtqLg6BVwYYBUFWu3tITG+PnOyvYql9j3sITR
culrbhC8Bxd0ayUYes7cjonVhJs0beFzBMTEzaVgUUsjoF+r2fqa8V/IJnzNXIUO
ZgaFCcWaiPWZgl+mnYE/yZyQWd/0McT3GInoEE96mExx7DzzZFtCCTdv1d3CJxIV
XMRo/sKu0Iyrk5E4YA+8f4/n/Wc4Ls0KL2YI6nc2U9o2vNFIQ0tpsLUORuzoHjqq
4bSWGPE4O/fJa6LJzkfevtZc6vz8lCEdgr9MxIeY4x5iqnYRFPwCa0hDdIEpbx0U
Nyut+dtDzp+nULzjjUR/VKPp++hmX5A/cfRnYZXoQEoPfGNj9cAhSjuQOoYXninr
+Mb2GvjdTyPyUjZDpl4jTturGxHSooBu5gsu+vcGzCPgxi888uSeoDdhbQZQPT/+
EYSqwsF6UDwBkMBvsixyS2NhS+Qca8txGl6XKSWdG/ECRV7IWfu/Eet0S0n0b7hR
W2sVVwqVtvVShkJPA9qysRZD1yzxZ5UvCh8v6I1LaFurKG+NZAE2L1lJ3ibaN2ik
KLyNmqL7KoumRbjkpneILcVaHwcrifpkFe1W4h5ozH4zaHQ4p5W9T5UzDhCIHkxd
fTsZ1/oSZuRZxQ9SoCcl4RivNzumG5NgAdYoNCZoEpACtSFRFbvgacUK5k++LyBR
zclDjK3t7Dbk1/oqlpdKz+7oMyouQymUktkM5p6ndPT+JUmInhFkKK24ndGvf2fA
ZFZgGCN+j9I2AmoL7aPV7fFSOyM3DXVy+gjnE7AQqE2cCGz/WH7AalTC5ZVho+ZU
fdzHYtCE124fTmingIUKf9PtbH202C9TXTrBSwoZaQpo1pj+xvzv38XM+N3OS34q
MzF9anrlLD8yoGRivpfUjyYjJbwlP2KSipx2Gids/jdxjS6TD4rlY9Lxnw399MMg
bONffK5oXrq1JmzfK7gXvHii9K9zTCVtXfXkFamlfPmyyBDF++P5SR8F0pHutxiO
diVXLldXDiv7LAmVAU0qdxWE6XpuCmWAruFNX4IxwXNLf6wntpX5h9Jr1wYy8XPS
ND1pOqStMIeJtVQ0taljq1gs1wvXvsSc+y+FW/1Lw/wMBGSFIf9ASFoZRCVw6Hxq
sxod0TEQo3gjAeBihAVSH7k5A+bWQcMgpCU1lgighBk/tPRlolwq1B/hwIn67lfK
nAyAphaZbGkWEGPBrn+Og35o5zEYQUZEbZnoL8zjBxCJh4zAncmOfdsI6K39AGn1
`protect END_PROTECTED
