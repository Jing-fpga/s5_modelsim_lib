`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RXn+sOpWLFK97eThQWW6zyGn47j6KellWg2y/j+XZLuDdilFNpp8jNjE39Fs9WSa
46+h7i1BS5QQKbT+bI8eirocWZZiYXaKRZlWdNtVnvNV/JHGdTXJjSUydGAeERll
BY2QMcj5c+JJjZ4XHAiaRM3ueVWgHqw1HPIgbysAgR7goaUOkVMai3xVAEGn66L3
1I+oEcgYOL+fJCA7Kxd195X/g/NQpwP46+HPud5Qv+Fj+t/JDrdS8GvwAGcQg9DN
XkfAYCDTE5ewRj1F4J4TbH+A0xU6qFOCvt8b7sW3QiynE0eDzJLlEdDMdAAoepLl
+nOhiqTzXmDoYgUtAd2abmDUqc+TphCRToyvWWw7neZpPhOYvvejc/PpIMbeCy8N
TPZs2nByO7kzFmJ/ecik2AFVQt9KBhBcjAtapMacZpZzowD3WkKMsftcuO6Y9pNp
8N+A6HESV7q9VaJoevI2racERL0MUmbi6+Gxwh5t7Z/Y7Fsu3gAd//GBMfGRq2ws
aFIJ6940vzm7s4ttoBbOWdR+CplqRdprb1e8EM+d4ym9Y6MGPGlqgZlzIVKEh6i0
tK9X5oIXQl9XMUQYQJlXLeKmV6Tt5f0WLOaACDFBVRq3ZIzSnYZxhS3y2VwzhZlZ
O1s0uGH7bhuUu1kC32Q1YUCTs56BxuZm6ZqGvNUMTkBciY9SqIiWKJ8wk4K3Kh40
+q3oXeWDM6qpODLV5YwIYjVkPUXDkK7jMgQ9djWkGB1gFUO8apzQLMvvfVqrCYaK
Fyd5IJQ+E92TUQJWk4hqu16RH2MDDiDoLwhV8hw9rUQdQ3n68RYIYKtclh96BN1r
jwRJ7RS5PrR4KcOTipjafv8YzFOgIX72n5ILss0uPhMdUySAiPwaHV6pqbsraKtK
K3HkYXtOTcjjjvw/jyxDKse2qeK0gfCFFcjDhQgXWaafzeFS0FQ1gOhMcve+YF9E
wVzEauM059n92yL4WQ0yF3uZFGOi/jrm+WnBBcueAiKQQBPEddiruTF7k/RS/5O3
udnxRjakfowDVH/CclvXST1vmpHGhwaCWCJjePjx5wClMjNZtPk1hOYrF5kpU/X8
nWExB5mPUgNGLqz2W5a0UC05QzBxqY7XSXsOqjlz2/FFmAEe4Ritap32E2cD3M6r
ZX9xvPVp/1nHnGy0zViW7k1SSUrP/ExznW9PbLCufLvJFT1uoIeVp+pOKVHTfJGX
siDxrtozsFv+EB9xbjMDHfP10zPVvNajGcSUcGtFzFODRsy+E4fNZsxExuDGgOBR
eFi9Y2sSYJ4C/eE6Kmkqzu08d+eW7l3zTkSmcaCRV3o=
`protect END_PROTECTED
