`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gvp0Svt+OCVXyDQFdGz8tq1vsnIeGg/FsyCJ9ucE+v1tQiyICudOtP2JUbk1gNM/
00DxIxzhKqon3yj6CV0bpGXGMWrh4BKGkR/gc7sBIrVvuV0CHu4kWujMRUatFeU0
VvjxE56CYWUkq6HIQmC0c6PgGvRbTFdHaJTjWPk28RNMVN3lGXPCNJz2G2aoPlYa
/5uN8mPcbc13b+hCEPK0GtrqsyGmJohDburBHk5CBGIL0/IMUMBAllLIK3vUwR2a
sWlLbjZw0RhaQ+trYe2LdgH1mU1xPK9Skz/HgYVbP7Fd5bAk8R0K5RCMSFK0TJZK
Kv51If1+3kOSg14oA7Zd7yYg+MVr3H1I4/EAUG/WBNt+g7SWmr9oPI6D2qfZc4eg
Atz4NuH60rqPMpW2+ZEolVaog9fqvNnqpPj9b3W201iCjXH1l/X0ZPzA5ZKDm50U
UZRjK4hZe9pY5vMhVqIT4VAtZo612wmdP3PNupBNH5V80JhtRv2Dz4/D/+2qE6ke
LsegmiRW5t7It0pC2+8jgBa7ODTwWHt8lZjCxrr1XPU6qlscPB7UgMgeW5s9W4wK
KsCQLZtUxaengAdAmbK5Wc4ix8BQPsM53GkRb3sPwqVC0pQhOnehpx1Y4cxV6fC4
rlun1FESDSggA2wIpMX9beL2Fex8koz/i1YekGA4Lv6l7Y6sxcAxW2iSwGZClmvm
tcZ2BGgcGYkzp7tc+tIsy/t5E8SKTUsm+UKjGZyWx1UQ449DxtRr7X0F3ZK0p0AT
LasbkLOszWEy9TxDmHLdJ8mNpEnJnirU16bZWCwrPh1BUeabkcmB5gEWXGBrhq6X
gkXLWfmngn1yRu5wjBZBzaUOyzkWEAW/10UQiPSLF42mtuKUDXjhwZKrjFQ9zaI4
AXhTLkJUDbj50F2LsBOJXcdUIjT6Qy32D0uV+jWmFHXK63iTr5kj48AVMumPSsJx
xJeUsQg+w96w8/YdXO9zcyVoIlyee1vLiwQbhIKwmiMgCgqninretX3Z8FgjlVWm
ZzyCxuLorETQDeJiWPk7mfskCuMdeNgPwCnCBsIGgLSuYTYcSpOh3gSHbRr+dZnD
`protect END_PROTECTED
