`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JE87UVxsSfTwXy+eynPSZzLMrPbCTwvibXP6eE3KrOSEnYZnNZoXlBxv5xjwyD81
U1Obg/FKWgY9e6dmSxht1PkUltITI7Rrs3LVdHcKlLPOvLqOc8P/c+sovsPgC5AT
YkgLX5G6PaV/3xM0q+izWkOUThdL2l/ISYKB+sdxFfb8rtTtlIf2w33VdGEwkRv6
7kK3LwR4AlghVw0KVA976DHbrGQHo3pibdOwMOAf+hldttuFpo/3UiAq5gqnievM
ixgVKKLFPQ7iFed1BRaYIcIK0XtwwknrYj9Bt4wFc7d37Bumtfa/UU7I2Vzj6PmF
Ai1g5fYF2t8ZeFrXpdQiJo05o530qqweFiiCv9xI40DnxykmQvdldzYBXaWCVWGf
6fTnjTto5JaaWfWpqFkPYgeLNVJQ0sN65m5CARqgbrp3JjnLdvENKIbEPZbsVtB/
yoxcKHc1mE1b0ciNlfz4WIl9AJtDE9JaaQ6PXkCmCU6DHghhxEk27rY3qlVPcmZr
sBW2Tr/vT9/5jL8VlBBim6u/h6VXbHwurqG93Q1mQM/x1egeETPrN2eHge7Htv8G
ZwJIC9iUqM1lpQ94ijYX4w==
`protect END_PROTECTED
