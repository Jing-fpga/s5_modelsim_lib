`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
khSE1JnnoI2Z8lokUgLFm8z8Uj2FS75xztyuf0ceicinAbcLdr7pSE0tdhdHlrm8
Z8cwvvBG0ClKUUSROtB34Ng9eVRSYRJhvhLPdyq5axE7vc5LLeYhcXf2GtGSvvPH
udfcyCEUS+ndlxvYE1u/tGBowU6ykbcDUmCtA8qG5dgUckFXXyOZMWoa4g6lgO62
2YZBFe66rdNKYev3mr5mTsDgsDoBhoyzIbU1dVC4KrH4U5uaHucCIVjZQOvZPN7T
bBTGDKpRHRh/rDlcxehOr/3nbG5Z4Zjg9ONQYu/acz2ZH6GB1hpqqE5vwt83BMaW
Obdygbqfu1Eewz0KsOPQx7yFGMAzvFlspUzfGrhWXbE8CilAITfIRZPgUvDCp4m1
yTjrAJJeut6gYkoBuJDhp57oS2a10jfRGrMbnKp3vbSym+bph4EIsYpxTA+iqHHa
uDD02/M4fLLX44CK6tWjbRTuVsg+q0aRJpPYhCx5oXm1NOz8/ClDbO9PuOJkfmT+
ij7/DVOFoxqJuB1HzCyaYiQSNM1QEdDRAqbP3dvtW8HLVF+jeRCL2IUxGNRdXsna
V3eCbmrczjmW020fHFyPGnhEQQKbFEQfozWc69zxqPiNBhMaFRw7FahFisxEDeeP
Ns4BcOXKX5feBgvCxdfs0g==
`protect END_PROTECTED
