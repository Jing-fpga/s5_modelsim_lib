`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KYX+8xcWSL9xJg7ksuLiiX/RWGHHoOC3D9cHTp89yiWfbpUI4qwzL0Ed9JfC2MN4
nzIW4M4VhxIl/nQbHsqB076/onWEd3CaOn7AY6wY7eCt0fvmofgXyGQApuJyhiaj
zfdnTAonNgDKE/QQNurIPeeMVmXnk+2KKKbCNUEyPftyMxxZFkV0g3Bv2LqAiSi/
bE6ytzawWcrmPq2Jz8bNcF2+t+HiLXSFEcd9g+pNnR83mKuJYHcMgNn7yjNbKXOD
agFdMFY/zBDt3kvXOFmdAf93WfDyUbMoVxvWNyVUVj9CJ/Yp1XzXslm9xMx8dI0E
v2Z4d0yku0UHB10CItUaI4y2z+yG79loOzxhvs2AZLtscfYzIPTs38hAllfediKz
7+icmSWbbrSwOo3t6Ucra1aeI9hwRaGcYI63Rd47oqs1Z4sXjPZwzx3GX5vyXBaf
wy6of80m/yyNpFwsQtJDZVRzuIOfjhvjGxUhiSh1QmrOsiB6KvfcFWTu7ygwDpd4
Zrj/a+fpoK9RVKQL9nN8U9ROeBkcK3azQ/RTp8RID/ywXPAnSIIs2oxooNH5MtSq
y21xhABUYS7WXqIUA12qLCurE+2rzmKbyFpHAF3fbC6QBdWJZ8doW32gEKqC1Omw
GPhu3bTpKiXGa31fPLy0EqiVpIHuPj6jhrAtEiq3T1G7dHZXBphFUd/IA9wmiRq3
PegmJ2wriw/wkXlFJ3YVwFhHF8FivhLYoo0LetB0/fruU2ef/R99aepopmRli3Qi
NoNpQUgSJXkHgC1DCnlHZxGZTwfhW25OuFfN2g50pYk=
`protect END_PROTECTED
