`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QiDy7y5MhFCe1oprRyoN22CVdOFoUtc+jeFcIltatHiv6VYg/2/xpWq7e5f0fqSg
68y+ZJglAodxvMCrSnWtQjrK5yiOm1T7GBxrg6gWHQsCw7fhW7sR58oQJTkDaSPc
I8RV+sD7uSYnFwudbA7PLMGzVo1MZphSqkbTRwwGH5BtnDZ0bhMRz+ynemHBqpGO
9GggrjehHYBKgkKQ7thVLQBZlJ2PMpd/5Fj2d3gG9Are1o4DEcuaiZbsAV2VXUb/
s6jrTQFAkBzXKf+IK4R6T1e685+S6lm1YrUz6JzxUlyLLb42SalsZPUeKz9ltlAn
+Ge0+7ySf1lDH6CEOaEEC1aQAR9sw80vN3jt4sIrxXYCXFZclUqTO1zQRRm5a8oO
EiZWIGTENyy4eirQ7JqqvDtuiKva8xy4AY7uSrwRzZjZCphNuLoc556yc3XUclpI
XlKM7wodR6ZWTyWW9fmZ7C5MeEyyEQtTTjDWGJOGv2WeuDt946/E7fa+R1ORpVad
ETCuIZPuV+YD/PvZZRkvdgAvSsz35ynHbKWhcfNqpcpH9ZmrqKBdKLI0zoeqPyfT
g9oAog/BThYhpKNLeiT4qj0qg4KCf5oIxZRaaaBJnNsbAORYCUyyy3+Tn5CtCzkD
egjzf3P1Be1u9k6xP9XX49Zt3MY+RA0wbitgfl1B/96DvZ+QV3dBYfDncoZRJ6mX
EZc9cdOANcN/yPkjRI1FuD/X6NCY12SvyqVD1G0nrpNK4GFQtgNwnunn4E02+2KL
plUqetfSB3ySvgKQ6SI/vD5tZXbXfY5Osg5C37Iukw43ILkTDHAaI/m8WAAH/imf
p5Dnpq68cL0qlrQwTWYThmi6QMbhczCbeATgjcWp0CKGWfvJLTvj5T0hkEo7h9/1
RuhSpuC0F+TUVrF7stCj4rK+BJUa2mtEti32pJ83yw8/hNiU6CIIvoyBkf27iQnC
/y03wUsYBhNmHziRfcGPE+IylypNVYvr+SRrsL6FXsFnin742h943fsLp/Z0X6K6
NXtL0JSixfDwlyVSrhRhWpQlYUKjCg+IxsBwy2PE+0Gyaip3849L+Kk5MVWG+bWN
nNq+KwOwTHcZoNAEr+omsE7I8yTMwwDiUmfOj0d2V04ugInZqKX4CkK4thGCCRZL
sHtFss/rV/nif0vjnLx1Vtl66t/cjwR7gHBewfRDbuXCpdKAba5iA0nM1nPzGGRw
daFEDcw63LEOoUOVeLDaQNFNXnEW+4gBYswIuebSTm17MReFu/79au4lCgV7AOZN
ueevHJ4i1zF9thPHaEDDvOgW34O7tVg35kxdN16gNwbl6ZDJ29G2zfbV9tr+qo4B
hp1qZ+CoQpJXxNE+HjkssZe/usU6oFuVAfD3vGmB8V1bquRZPvJgZdaD7QeP/Wd7
1pLCOdgk/pVvm/8AdFzZy61AUeiUDzTaryY1186txjtNIpGd8BUNrRv8l8vBbfGE
ht8j6rJ12E1JfZRPDUzgpCLHcQ/jifM6T0ruluCRJQ5n5YjVR9hnHW4aD4WfzefM
clYT8CISAkrZUxLspyAIPnaiSH/D+FljjONe7nzoXiW5asyPf63GMnlE8IX5rl2F
`protect END_PROTECTED
