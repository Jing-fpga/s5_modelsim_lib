`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eHuhoGB0XVX5egwvpeyqt8en9j6kFZyQUAMUy2DhYzGhN+y+0y1HsbE5UF9ZVDFf
vOaEKtOib+i1DzCNj/o2vdqfGFFCpVLq6/+v/WarxJRuRaP+qi5sGMRfDYm4FxAl
UJldbpwLl3haYIO2nygKyahE7udCJlOEBDIa0kgmzYDRXoxNCF25Qy0DBeZ09V9C
r8t50+QTWfUwEQWbJKhCFSLnbELNbhTZVzJ88OkE6sXmsIn/N0CvWsH84Bnxr8Lm
lITtc+Xlb9Fl5/rFJaOgP183oURqJQNFwtrppj6bImCzLGdNN73+6lBgUEdcYKI2
HXY34/M5ipFQMy8z0N5SkRfIzgn/XHEXHexX0r15Slx4IN+9F/EivHzVQnXuwfmQ
2goDEVk8JF249BAGrn2uSeiKfcIGvoVWbPw3zV7fuSF2svwYR6VMGeIGXwlS2q+Z
NHQzv6m7Bv1FmAZftVLB+nl20zhqTV+Mo5eBxMM1RL+/oZqLAHgGDqzulBgdkS0c
legk1pV42kvrWk8bVXBfQAsYHvDKdojGsaAG0s4bVlLKyAiON/7oLmrDceukR6DE
iC0bZErtjQ80l4lXwKb+bP7oZY5ribW+QdCFY8p6Rf++gXTWaVyQqYyoPPXA5a0i
XO0NyL+J06YlQ2YlTuCSXaJZluPVzusKiUUBjSYvCEfKuW0wQOcGTdPsW/VY9mmF
zZRgzodMeLbLBO0v8IsmVGti9/ROs1AafjqicWl2hqlcNT3ET4mwgZzWxGJL2VFX
wDUuHnCw1TrNa/0XqHDxXEjroPjENfITy2zH2kb4zzEH3e9v63SZB4v9rjB4a0Wh
Nz5kMPVCKdz49E1DI+iLv7KzH9C4VWEFKei1C/wdVTheB1S2vQnVtawu6eSd5IGn
ecppzPiUdWv+rL4GdW+OM0WboAohR1PBq3am8NpHznKVvp0ugizP66RyKybCvvPE
C2PrQid7YrcgvUeyCW9TVlcrEjcibUc8H8FajG0KdIHhDGNmf7cKMjWsCuP50Lur
TO1sJHD2C/j2Bt5tiOqPCd0ViEq2SH+BSQMalhgrX20XsSO+m8GWqcw0ckAh3ocz
Ogk5N0/cYu2EHR1jVTs9YwNl7/FuLlNrhfTOg8zhvQ7FBt5ckgd4LW1AKNXhjdxU
YWMD+DK5najGz7d847gQC7VuABAGUYyQN1q2wThJZdIib0dJMOe3qeJNIINBXi+G
lVoAV5FdpnZ+1NLgk8gnr/jtzFUgZIQS/fMeopNNNIWaBxKrDViOL1ws9voL0D3S
QfcoAbPau+xFbRwVlki4TfSdUu0eEjKVrTLTNXthDserzfq3wZqhEXcl5dYXs/iy
hpZwR3vkjqmGL9sy+JLGwQ==
`protect END_PROTECTED
