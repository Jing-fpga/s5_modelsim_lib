`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qVYQxaotnaAxrpUIzhCxij5eYC8Mpvtbe6jCJSe27yXCtDuSfKU61AJ8rqNU3NHz
8ZMizHNE4RU8QSb1HLF/mde1ER4CrmgkVz1SYpIj6FqeBuVzhOJMob/EwVJu+6oN
SGg6QbeuGUpyTlsahsQ25VWrvPgIo0rd8JafxoF7CRswv1eHL6zHYpeNzXcTEdyQ
NGN9XpfuBi24/zILImMMbuexYemtxpBENM7NuEXQ5NOjbsOm3bYiFUTKECN0JtjL
FgYwjrMx7LrPGUhsC6Nm3kZhfC8Of2HMMv890ts5O76j70Ys/yZFYxvw3/vhAko9
yPyQk9xfZYu5VZz85LsFise5Xt3XPbrSrenXgaJUo/tpQCWj92XnyvyeWQF/+dRV
idiK6bNY/5mSmw+2hHXgBdyyA62sf20LS06zj0icm7sX2NZ9mi4blXVPGKQZj/pb
dNkWVXAyXHHGNY4NarW3jhUxu+w7JvIlbIC4OhEldW4MgKYXtzrY0H+hH4thmG6L
+dnauLyUqkWP8Rv2T5fQx77GbHJv3P1uutYY6v1MVseGufRR+411nNmnA9Mtx3fY
1ZUP2KmUVsXGJKJaXmgmq6/lSk1vUDoGknIQlBy35RXWX9keSHbqhbcPF+/V+ZYF
3gWScvwVuW1gICAo4kYjawkveeErgz5IipVph/TYkAEvX53BO0Rn3WyzJO4wmfHQ
j7x3arO0fBKZgCBi/0QJid6xR8+eoHaw97Vum1Ce4lEowR/z+4hoVEGlVIwVf6ZO
5m6l4wfMhprDp5nVfLOtRDfVbIB74sMmmwLQF2rnrDLe46cCGJ2Z0rK6IL91f0/X
5IwRzG/ImwtQH1/4HOLjWkbVtHZeHfsIDB4UJzjho1tgGZV06OKKhN0QpgWwTp0P
NSkw8fK+sIl3JaRaFrC7VPGX7Q/eB9kscXVf8O3nh7pPS4zpf7KD3YkqwAzlESeS
lQacP6c6td7ui9RFMrvTix1xawJCEhtOwNlGCnWNryinfTDckSV/IATwRhQHp93j
pnIgBIBKXWfo24dioXukFX/bClvll3RR1hYWjX2op4lq3EIzU+4Nh1pk+qzLXUpn
nLonf7rnf5dYnvTRhuQoPIZdqXPxNyzrs6ZLctWGcjKZRiINbYoRWNGnjzUtVg8/
+WKBDhLpjS5YgSI7ZLD1172vFHa9MKUR9fAOi6FrKyoxr3wvILGwfTPEh5iIqAIE
bW0X74oZ74c8wE/P4msNEQkIoykGRhBmmpyZA/iYAQPHlbtRg3alA7/0+no3+Q2K
YfKafAdYh1ZgiovFXOpoigin1vbjGNbO2/U6YdmRCBnpoM/lP+0r+8Isb553xjCz
Q2siE7A/dbp0BE5z42goIENkvtYmX4ijQXDS7zT6iSOKcKWttDL8Rx5eSt9rHl7U
yTfkcw+eIznWQ6LVF+hHTuwtt91Z+jM4pTvyp6h5fV3k5jDjQqCox98B3ggPrAdR
M4nPMWyuViSMkJ3j07/NUqGSCDkONzzMANn4UuFnzIoJ37fmilXhP/P0Z48bFZq3
FjK85h36gMvJxLZgd8UXsvqC0/y1EmRsSXwqZvowWqA3IAsImCLEcu5+FqY9+hrl
`protect END_PROTECTED
