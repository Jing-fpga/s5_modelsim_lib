`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZJlryKapyjrOH84UR5gZ/6tQEX0ha3dJ+AuOShzSsVndHSMa7zh2gYrjTwIXDFPJ
zONdyrpmcVvL53f05B3c0AXoPtXOk1Zv7KX1q5NvRDPjxUvImfkD/lh0IHn1KY5O
7PqYFqTMcfXCl0xpk7cD7URkfF+bv40R/g+fCh6dXpIK3B6NBhecho7yVIRM13/I
HJKxtrIs6ohDKqY/m2t8hsjuwAWqj2XVQb89IWVBgfwLIkVQM/7TxeAGjrSj9mOG
ucyVDrX62p1fv1f7KnNBT19Pmz8/r0Vsp9PnPJPXjU5Tws7NuNQAwZCVT3tRpusH
8XRc2uVqE0OAVFVKGTBUHjLI3TXR54q2BJIuPnobT5DhHkf2pF57kqgM/BazTP8a
k+QVr6c7XJMmZtdigRbNPYlJ2kqEe0Gv/2OSji0i/EZ2ATwz7DD+/AOnOvuJnyt8
i0mnJDoCn+m1mPbC0SZ8VLqNRIqccCp5HmAlQivNgqSYyq/wcS4zK0Hg0jTk9zZE
/xNT0NTFnJy5kBFCiWk2TmOm9Qm7H1xT6A2EDEMf+WAjE7ZtoTCCQWefCg9hT1yN
P3vaQTtAmjWx9ndnO3QFKMjZUbB3b3l6Ss6M3EVH9je8/2jqQ/5RTslRZTFOXfU+
QB1sIDeKq7U2PcMBCAy6DuUvx3OhC+nhYklwLeC232hVV+4gsxvfOV3tCgiZQPVz
n7oJ10mjGnmhmzAkmSJ7NNsmAi2CeUWNUhsQXufHCYChHdVG/ToYPnip9nMdotSM
l45a6EmfWyJ1JRwGBELg+3QaDRFLeptpOwAJoco6ainJT3zlCc9ahq5GplxI/Y1k
68JZrfkgrUgBUEhgnZu7AlcfzZ+Zm3L5PfOn87L+gOBoSn8TI/44WgT0Pg7cQ7Lw
Qi0/PabAxRsKomK1B2k+dhTyGghWELVjW9fKyFDUnVqcsJWZwL7CM6wc5i6Yp39n
glmOri6i3rram1NqqQJRfVdz2R5FDKUGUEfaxMNMIyxcbia2dK8j0mcYIEE/BeAH
nooka4s4h0A9HDJ4KIQ9TkDZob6Xf0qCx1qdSKX9WaS/jv5Eydt4aMerdjB89ZFd
RHIBnXaxo6l0vKYxzNm0Hgcx5LFfKSkp8yeMdHAxlSBPgkLJ2O4i9iEJawEhHY/K
SV+H+329WCqCif0wPc6ZN34S0LTfYqOV7b+CgtSmH6m2PdqlOKxGjaFmpgAZALea
U+P1VoAFT7ZxRP0PqdhB7YHk7YSSqUBWEXO7lLr91W1R4maL65CFNUhoD/m+zvx6
WeIgpYqOcsQz8DrM/DzB2kmhU5H+Su2f7BQTFqIhYc5YajbmfNrh8XhsogBRVXWc
42+j97d6IW5Ja21BD9rNdF7HU1Gg7yi0FJtI4tiS6t5nGdWb0Jgag7HUdHAPKeYZ
RbjarMnXDYXgVq7tplhXQFzp+LWHv2zneBws/mqvQ1mk6EoJzR0ivWQ/4gwU8Mdr
BuNLd1lrbtT2kLTJWEysbsvygt87WD4xy5fa6yi5mFnyQaZB5Xk87QNZ/HAs+1bS
qsqPRRj8cbKsb7SZxjTzqsFK4CrgUdIVIi16XxmwwtKRmcSFlxtWQTA9sNpmDDqT
bFh4jvI1SwPI0HTM9OtG5jTYMVRgA2+rKXXTxuogaqAfn5w3jlqSacDESuYZfVn4
Yvg5DyW6mOhkOFgDfqOUxQX4A7TSeKiYOl2XxB+yDvslPucdOATcUvgbZoi4AdV5
g3CN6AxRA43Wu9a9vrM/m7eeamfKYgTG5H8RH62Kdva3Zj6VbL8iaeysp67fO9uE
kaS6yk9aBBWBqyLoPUh0+eTYVQCVLZ85Iul44+81AwcowcwMZX5jg0B+WE4zLCUT
PSoGTExPU1VtaaMfH2/YGIRjZPoyV7vBFrTg0ryhTuMyBr/BrQxchRY5W0b7nLsl
yZ1PRYflkvopBVCuNeSGx0IkotCzmZJr7BDUpZlYAngnULhTHs3BFyuCpQ/W8TTc
IzTBLqoxSFWfyTNhBr1dvlVMFyXyzM688RUPvFNJAjFfCSDgZf6aPBvw2mv54QQq
Is7qjIW45v40hHCvKmaMM+vX7ljzgNPlDmAgU3vQXcT9Wvw5WDqhrJ2SgAXwBACD
lWX8ysiohVgJOhGaRl5/Yynh6+E9nMbTmWA3okosbTnsBR/29sC9gMEeXDXH2/Ub
wlfuQp0RPQurGqRNTRAci+EbfGFgyODvFv10g/ZYhPj3n8nUiTZfgvyV0dyf7to1
uXeu1bwWXAoWSIiKth76ha+dUFqsv+ErJRzA6tY6dQL0VmBiAQq3zdOak57gvRS5
eyH9N3D0PTMbagJEPnnTkMG4EbjlxLdo4YaxTUFOdGlq7E+iprFVLJnXs7I7+bhI
6GFOaQvSnZFhjJaibWqBL0Dm1T1xDTHXojuk12MAPHSlEUqB/L9AT8hNk21B7UKW
ik+CT3OfFvAXL9oJjLglUTvTwyE5tKFMBLuIfSYKM5l4RpCTTOVZgkbEySYoydJP
EUju7yqgn/Hjk3CBWLZgwPqhpFqsK39c5BUgWaZIe21aKdjhC3osB5JMfch2ps8V
huZB7Lyc7QOuizYCp18+LSr5W8q2y7mf2R4Td7Z5Tzwm6XyQO0e3GGyeO1JUM8nD
93onS7ZfDw9FgwWgsFuuDwEGD/rBEeyqsf/zeUeThPtu9DiBFlNTpHy4Z7ant+VD
T53PqNeiEpNb7k4ap1G1K+XfdVGYso3hblyTf5O6buzjIfP5CEc9jL34Ivqnw5aH
SzBZblD/c3oa3Bnr+GBZEwLdnfDmj6a+NSUP4iPE6nWmSQ926byY5D8gtK6K3aAN
MIrLJZ6qmOyThd0DGkr1ICVXirttNRmJL0oryhC/6fGXLTezHfQZNY9iekexqTH3
NSF+CIBRDHrIRlrFrqFPRsSeyv0VUdQ2m8WIqZKNuiH1o09O9iQjMtkERqpdypWU
imrDBNZgpQU0ERrG7X+dyt+vsg0HNo9esJA4LVjjzjNAVjZxdWa15ck9Ubhb08OM
O5eP5HVUL8OW1OrEQ29fZ3BUryzsK4NkG/i+ngttEapjxsbfr+9iVaOr57UpHwjS
DEn7AhNybbkHFU+c1LDBycgpxDtRpczl6B1TtZWkQWOk7kON6PhjRY5LxElHMoEK
8S+lgXt/e7Iga1ODDj/vnEdaYZw5S6rWBSHydiWCC21mY2xZg+TDRbjVre4PP2te
/uzDK+STHFk2oW7Pb8wy46HskgTiNI65PNhdQU1zBbHW09fTXyE1s38ysu23R6bW
JOst6Q8nTrDJAX9SqRDKZ7KICP+BgrvASNLxeEL4KI/48ORqj62hTng9KxlWzNvF
MJuK8zShuMKpq86znazvnclp5bvMOU8XCvOBTKrmTq/exKbRRHI6Fp19TQAO5wvT
iRCctH6mRZKNll76f+51yuOoGDxPgcEbC2PJJsLaJOq740qvsRJXBNtssb6VDshJ
WE+nJiYs2YrlIY/AlflN4b+9SmvoPa4d5k+zFGGjYPLqFL/BEzeh6TcuN/sB59VT
YX5D519RmJY+OXarutED16r+wWvqIBb3F0NG+sqU2DZ2/FFMzSASaXPlhN1F/TkT
ZAoU95fMf8JOgaJAS9rySz9/sXqfHgLnayz4L898eyKq3GC8v40JEVYnXWUYny+7
QEFa1rVfVLIKdzg7+jobN7xLypbx9+YyYzL9+COBramaB1+uH6jBXI9P1mJnpjLA
rlZv0yIrjHn3yy/uuFT8SAvXGJrBfFtGJ8YjCecYX2AAhELFUoBmsyBT5MwoJMTo
Hj1H65IzufCEv1tc6GfchbMRCkbkqgdwNeK29drySdoZRlznu8SilwJ2cFKcXibQ
m6vd2vKBuLbYRAv3HGzxqCfoLmfKhgujdnM2480cRTB7QodcPRqp3ppWGQQSYcfz
zoJeo1jKo/rbjU28r9AyvTmOf0l9JtSvtEs6RZCQDeo9aC/q7zfJai7HIv+/lEsy
wJ50IANlc7GT9jvmMeI1qid3bWPEmGEmuXYh/zH/4dJ4hav1HLli1iYD7tvJNsGn
45y3ZICDqNOrU2Vi4wXZitNYSp6mpv/a5WE72QsP+K1Kl47JXmXSXRoe3ENuBwBA
+tSE4KNpdF9Qae9ayVFQKx1J5QvEToahZdOiz0HehW43Juh0znJN/LNA7Y5j6eB4
kitBwrt0X8DGLonvmVha9bcSjrds2vJR1LH1nUtOcD6NGW9wkykRBg3hOAeKKndl
Tyj4O9CON/BwqnyOAhatTOhxi4hh4X7wu+2+7VQFdfWWBrlpdtJHFHvm0HgibzII
sEfIv8ZNJ5xRf62znDc/cAHLzlxloVJ1aJU2ucvgS28wlCSqveUHZpcL/a9OKeqy
kz3+PZgj5il59jP0uA/VumeVyAT/IbNZtxt6fNWB4mPx7shEjnkIumg3tvPcsrZj
q3gjzR2Yd3ZNhGGqhGZ8PTXzoi3AHJBfSTj8R3J3WkjHD2xkwR3o7EDHCk3KwE3c
TA5glo3+KiBVJbx5grh/VqXv3FPQHObklUp/8qfE/a/8bgMW0mZZNwG7BDlK/jjt
2tjeNKTZ4GdDpeT/pADIwO1VxYqKTCGHpyaWlj7AwZ7Hw3Yr5p+/+W6KDRoiS2LV
b5WlE/YbXFu2I8hkeY23VL4K/1JIWm+74NRTP+Qpl16eyFFEQDCBpIkV7GG/O+Qq
iY9FRMaG+XGeGsITG5k0S6Hb0fsAnU7209WQGCL+q3VArtaEz+NViUj2iyeMxFG/
qKArcG4IPwyZsT8jH4TAdg==
`protect END_PROTECTED
