`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X0zIRdlSG/QxzvpcN4fU+jpDpYeKQu8tyc7X+32gZGn5dn+HQb24cKeklEkHrRKb
riw7o+Gpp6jILdim6neFC8kMyC5o2bXeZNkdui27naroHrR5HFLDivr4ZfzPouRw
XM2T6K23x/whNWqsVAZuPo/usM9azg/cmkZD4v6HhL6WGCiZsdXSZhQ1DPxXZVDa
w2JdXKs/5tQ707f0+WG6hqkkVjRWapvRGUfsXbeIkmNWPPJm5y1Wwr5sl5+nocTP
3ofsuGsjL5o4OuNvdmGlocIPksY3q3braIdu4EQ1+WhavlPq7hUwS+4406CDolYG
751ytN6S8gXxhgS5FlItkA5tOiUTusAD9fZSkIAl8Aa55PPUwtueertNANdcyy/m
oEKf7atnZPrU7JRtHwnAbUVxAdkCOGrqQQ7hwTxDRqdTdPWz6gjkfOS+6JYyhkbb
6YB0v50bfVZWZGNG6zz/jsrmaCGdt8n7Qz2H18erKk0=
`protect END_PROTECTED
