`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C/lcqynobWXJZaftYdQTq7DPugt3P7bGl8GS4z1B01Yr6hTT4KVKlEEQgoQoW6UB
KptHB/L+c/mMO1ruX3kLmPrZ0f3gVNwjnMpxHskhSUdO69nMQZ81d+45+j8UlgX0
4hmY0XWhn3uo/tkA7Egcm2RyGsFctJ00G/kDIeR3KXIN7dyNWTosag/ryo0mLQzw
AA8BtQkrLMN12+pIPx8BgbZ998+w7TGZ90EpqzpjO75D8EI8ibjbAog8ZIu2Ke99
JyX0qdZyzcTM7fCDNy5CNUoe6tADjuIsvYio18wOb0EMuW4Oo1ntXhyibmuGWSb5
8IvchDLSs76W+2gyu1nlHo+gjfQLorRJEAFJkZMZn1uUD+qRNI4iL87cfMhBJieB
da66zkWt7nHsQmc548iciQ0hmm5Gv2vHKVeb94t4xUa9b6fb45LLTy4AtmlvONG7
tCUOc7n+vzzP87wWAauOhWMelrRBXiNTdgriYoUayzTcbZjAgZ84RdbwpIm8wucS
NjAfbC1il2m72TeWkp/5w+TmDG6g/7ze5QHFFJuZv6ZKidOpF6S30EmvyrMRKevn
KvR7NenP3BmRa8N0TDAqC++oleK6R2AvbRU6Xxu95uQHY9IN+R/OcvIxFw36aAwC
G47UroNNr3XWd0ZqS2BF2coXmhoja7m405ST0kAtoYeavnExu1OQQ9iUMxRbcFzq
+wXxzq79l60WPdbr/zEBJBHU6MeR1iha0pOSTTP33m63uFW8NVf+6cV1GUcYGu4A
tC0dmb8lxCOsZlsueTIZEHDekoXCqy5DQ1HAc5GZz8MYR46rJv2kJxztxmv8ezS8
YOXY331JZ1hSadeh0GdnRdfzVkk06Hj4WoLJJbSZqiytMukHlKMzdWJw6rXdPeU4
oakOH7AmzxXM1FZlWNdFbvlLwDm9dprTpeh1vtvOm66j3L/RJq/gPYg0i86JBY0d
g8sQP/Jkalm/ISikOVeuN/ovUpPb4pAosY2zBDTmQDbv/15zal5KK5MUWDEoQZC/
yaq8OBZIpE4QE0AAnrsiv4gtzgh9fiBp9XF3JRFMYgyaiKZ7rtBs03UfCAoXWpi/
Y/dlI5GwRHAYSlRIBz0fV68rmfE9qPpuhArgc9WE8Eb0i68Y+TQByhI339n7VxZR
ke7mq7PpHhiTXsSq4dGVn1gX+clM8un6DKfQUVnflglovpeefEAARx04Vuy6UEBc
3Q2MIX+hq9ytV1NfJkoMNmG42sbr+5adpHSswy36RkW5Pz5YzA9SDXFaxzcq+UXy
nkEkayNzKV5TanowrSihRTQ0ht7lkiVhkXtS724Bza3HFR5/1CYMtR2OWKUAAATv
dAxOpsncUokV7SWAxTYSaRwZQY/SGF+iMb3W7s7LgRW1Ifok9lBwrWtAKpDRxsxX
enMXdbNNRBTP7rhRMNmeLmb6rUQAPdDB14R9T2/BUEqRuPaaeXeln7awyRBwOSgv
tTAnvBhnZkUmwPUoD0szupiz0YuB9IBajg06eldly+9KiJ4YWOTz057L3OGI70O7
+YBEP+1Mmbaefm1yNWfVh3hdv48EjQzpBqHmpf5j0jF/OEsgsHqcq9sqOQ2a3GXm
iT26M0aU4hwg1Abh3VUxoHl8lFtlFtEU/QRU7Mk0GSo3kyVeIhwObcAUi0H3GY3r
ZhSDYvWpfM6nA9K8b1MwJJpxPmlZQeeULntgZZhvL9UgKBtVGjQ2BP1XpSEbCEWn
Q7nc2E5mUhywSkC4t97LU39GyXIwN1qo9D1Wg2p3ltW149FbDKgMjvPhGbajERRy
FOoecHYWriqjyC4+oZw3c/sBp3i0nvAYhc9pj4FzdUmmMG2oxRVMt1dh+01K6DxG
cQehUGsalri2WjjUdmSvig==
`protect END_PROTECTED
