`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p0cFgNGpnxAMy+y7fylvO6RUPw8/C6QB0Sz6lF5gxmQShSF10bEXNznx72O778fM
qwxEbrtM2chU7hxnD1UAsBHV8CC6CutBsicY2DNA4qW4EGMM4Q8l25wSCAMoXV2J
OpVmGywKIQBV/F+8CNroh1CZJ82D99tswzJlx2v5f8hl+Qs9pyWFJe2bsyCVL+ek
049RcDVtD5xNmvvF5YSZ3aLCZ9kbdXth88t2vDSZpeRSi5QE7epFfxZod2FBnbS2
j8t2UDz0DcWWhTBI0hMaFHD//hgp9Jd72B3LEsEMHIpse6MFvtx+mW8/kGXnH7LE
7poRN9XbWJb2vBEr2wmc+KYip3GHa+LUhzNtiMHmEo70f/LJ8F6cBO7oGHxbkS83
ciBH5JyYrxXJlep+6GqjvU+xOmP5V8KbUF0SHHHQxXphxQrYDB20mE1zyiKo09IG
KQdJmHpAw+qfQYSb28DQlzP/Qm81MfaOxphBaHUa1suxu+kKht31FzCBIb5n5v0K
8kA0mhjIuYEiaR3f5chz8RTCa2IuswR3FjtiWEGqDpdjkPfXBewBlgTttLtTeh1/
/1WbZ5mGNO2S9c1bPiJGIA==
`protect END_PROTECTED
