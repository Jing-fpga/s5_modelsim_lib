`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xUFdnPxUK2YAfFlWGloUzy7/qY8PIVWfYvpjREGHJ3SCy2y85HF4Dhb+psO+EnQe
1mw5tX9LYi4LQz6k4Km0in+TuuVIpnXA8gkhrkreGH2WskhGJdbdzu8erU8rzPKp
Bg2Z4oaaDLwhf0VjHlCEPIncmmuKy6xX32gyrNZeEZMEw4z5itviClmG+ChMxknb
/w4OtIbuF31Gu4vwICGQcwXF0y1Bma+D+hbEe1Q4NZPfL0JOvE/UN7w+6ljb+sZD
//H4DPJpb2noPglS4EhGV5oFLvs/VpRtiiYxR+V73E/x126LkFk2/22J4zwXOkqe
owwT8glGY8X5aU1zgwICcvDWICL929GLGISlmmmAIjUzDOeEDbDFWas7M7bExlYN
ia1xKjPQTs1DspXUMIGuAGazztigJ/BIOD5SXPGQS+Q7gcP0QF3DenaTP1MTdiTD
+E9NLYrNi71bYUXR0PZSXbNugx+Mp94bB1f2G2PrEedrHFIGqy1OUVvnlovVO+2y
t9HTDXdJF+8Ngl4RuMX3d0tFE91OB5aZqUos0Vf5ALpw1pMYqSkLMHRlMsCfEDvS
JKUXPA1U1bSanGTPTNSHU10GGBYZT+ussO0jLbPEy5Eo611s/njmNBRSqNDb69Op
CEpM4v4D6pO+arrA4ZWeSmVgXYJ8Sxax3u3Jk50lLNm+064OD2U11PMhg8phbe7p
5U86htKBVxabIAxDTXvMpb8Irlcszv7GZMeAPXLNmp8jtCOiSnBgbbFxNSNbIDft
eJdtMtAWp0TsIpCeEjAi9ZbrxQBSI2WrobMeStcTEq1RfJMd/xnnJyqeZEKGtVf8
7yZlB6Za9hpFD0jVn7AovrdcmiA4nEFXKBPDtLZjiCfDpVwfIajbgucWCLFDS6Z4
tUT6IresXh1C4MuzCsQigwKT0ZBssGP4drJN8gbn49iDK3VA0nuUpNayOag0ved2
NyDxgmtUkD+/YkBkMSIy9NdHPJzmZWHsZJcVAb6YkEb/+v1LJ21Ew95hCfWscwbw
YOGbbJ2lFA0Ydd2LZQSNXVeLpHMnJqMggEf2y3oEprchAL2VN1d3nLLZIbNdDAK1
toyxJwDkttllzntYGwcoC6p6DmNoebyDaD4BR0yroAFgk54ujfUwOSjfMgeyieJ0
RFysQAY/Dm8W6NLW+LXZilXqoSuh3vW4GHoU4wpKRAn7ZAzP8Xj5PMaqT3NXsXg+
73pZm3M4UkzHdAR1aDm58BzLPEQjozL77fCVsWFd/IzzZekZVsx5HhQMNhk4wAb2
vXPZ7ubKCXm9llTYKONA6lKa4yySQBEJvAO13dWItIKE9JDQwf6uzP6BsvccQodN
DOfp/FT0RH/Lvk6+XFQjv/171CgQV1LXJOOBSczEXMCCeystG7dCM+6M6p468iNN
6VhqFNVXcjECVtxfi5vf1/D7GMk9F0ft1dZHPNsM0Js39SVCZi7WRfKMerqAstp5
GmkxRy3nZHqQ+d8VHjtYwQk1tnYMvOrPdVH2+tekvBq0fYYickw/Yh7Y+JahV1+i
GdidsiR3dQe94O75ECbLL0RQYlw+Ntg79AsKhWmPwgViufEMgloUHeC2U6842QHY
iRuWhFuWIQz3fCV+8nkpXtOW9L4nWLXRqY5+kTUbx6yxi7MoThHGx4pD1IEcuegW
nibzNZ6fw0XbzWsFbYuwbQZBF9Ia6iWIe5gTP18EH4Hx4iNtT+T5aLFNnfEQuNtf
Df8erJV0Cmfx+JGd7WEnCcfCKKKq0pbRfm5cDhaYc4vObxzzp+Wyut1ISuqE3aGh
Uf1CP22I77kv09i+1q2UFj0MZzfsCEWkhBjHIVdPDUvoEpBE07HXlUCfyGq+PNyS
XagWAnX04Ap4B9SPCSEf88z0Fxup+n2LVMzoogt5B3QWaEY50NqH5wLJ0Eo7oM7g
DYF2+CA463xlki/iBYKkHOdupsepsNaULFz/Fe+/ZxZKokCXOHR5N3IKeHJ7syMF
rN4uweOQWPINQNEOPRXJvM2Z//wPByguYx9OnXUVXqv52bkUEjeBHluCBmpNOZQC
QFCJQ13gawGfOZPBAGTh54eD+WxgA1bd6qSSusASD10d7wGsIa1reI4btw5Y3bi3
qyRUBrXT/647Yivdczdi+0b9psExaIGWNCv0ebpSI/2qAKZCCAaTR4KruEKy6DUY
fbyfoz43oG5YaGYj4FnlKwRGV8y8X7c0kppQl0dgWOkgj4omyjJODCgtDoCEfJjf
RXg6cyLVayS9bF17ETqJdZwYJNf1m4Eep+a/nKIpXm+rSgNgRuzLX113PVbbn5NY
mfs5ZaEfP1tugODyi5aJsvsl6rZllQKdpADFOeWYcLJb78A4pO2UK1H6CDGcCmKG
btO2tLsLfEPav3VGbdxWOjd4Rg4760WXs7qPZGbLsOlMJJ9y08LbVG6MNS910zxb
0KxLQwx2hUaDkLYXmQlasy0p6+IuIi/ohX0bZEc4tU2WkvSy3Jq8Hk3Zm14njOYB
VaDFW7vHFcINQOAN0iY9sDf/Ha8k27KQ6oqmL2ycBiRCA9FXrymQMufbj+YXxxeL
gdXjCRpUr09eNIez1BO6ANTuHx5BhgiqCAt9tzH7BzZC/CZFGmqJFz/ehLEPdxsn
GR4fvkxVM0vsDzA6cJ6fUO9YcoSZjmvrkI/QJZtApk8F1B/EQD85KqzGKbncXRQP
cq8VRXDHPiz9EcqwMX1zlu10hswhIt5phpQnONEkj9gV/7aqMlGxYB8nEjcOyMMk
WvTeJLgLFL8nJneNnTNQV+TkPzFw8waG8ftfcRWIOK/ImLvYLWaSos8dSquS5ptm
9CLbfJy+4g/+hkuJy1zEwfQv47GpxDZlFqwgKgrsWxybp1guIWHCMkvVdRJ8G9Gr
ZDfNiC1idb2RKONMXrQ3QtAB+um/ujvP7B+fPZ1U0u+vQm0uGUCz07RcCT3/cqYI
+kGgvHeirSKmeamOtx7A1gMfUgpSUdlKMSVyxeo4yButxQCcbZ9DKK6mwhEFmgMz
lIRplA0buaxrNx87kHSuDzn/Bpgl/qbpo25Kv5iQ2D/BJoLSCDsPeWOTrV4pg8xi
jZU3CywoC04EvZB3x8nbxbn7pgshkuAv4X9+VldNy1e9vvJJwDsQhpwbapsQ4jSk
GP3lCbjW6a08Ey6XClvVxu5OXV66M2hpqlNcwBSsD7PNksNutYGXENHbCrXSPVbx
Ry6di9XASyvawpJzyY8zsXRr5X7wfN/MsJfZ1rZ0n0njNlznuLR82MLnmiu+xbnI
pIh1DrqbuB4+eID17zP+d/W0PZF1zExwc7Y6fwFLCX1vgCHUjNpelH2kN+nMVnwp
OZvzush1YBiEkjjaq5Sen2FmSPR9/6Q3xlZ7vtyYMrbRhh9rRoSnivYHGZqTSI/F
oN0bMvJv7aCqK3fe7MTBusrLASCFXqau+R6QyGMBz7t+HR5dnbA1Gy1Ht0E1jhYz
b4PytUlR4e5e7dGlJb4R217k0j4CQebshR8gAv+FtU/0RtukPsJs9KwU9tBoKqJw
gYVSlDc7oGhB0WRFS1njGBABe/UmzIN7ypNZQchg/DZ/I9oi6kyDEFcUalqCRqCM
F/jHEsGbafdxsUtr579VdZjDVSzycK2yGdltc2h8uqbJyN7j04aJmKkSmKUH0dsL
8DB5b7ra+xiEtihHwlcDCF7cauWCcyQ1+Qa/OOXaHfRZ7i+atYMuG9dnn5fMEnck
Tq8h07V8deHYSSYrOTS3SEjl4JWE+FPm7bfbGFihpTa5/GDyulx3TEykAY/53wn5
IHXhIRb7lUafxCXoVw2roEt9jPCdywutbDW+td6giqI22dxRPrsUhFadXDeFJkZM
D5jl+J0Iu0ZcLOqx4tL36UGn33oiu5jcjt382yxVB2PYIB9CUcTInaQlL/JGSUx9
pAe3kk+r4ZtayUrO8+Ac77kSC7dbpbymz0w8b3/dyNv4V3v3pEZbrldHWcyk69ey
MjDYWB64V4QqECKcrv8lxo6A2iX3hWnBKAuxuRjdyWpowGyx+O302Y/2XW4Oodv6
Bdw1GsYVULBeMYkXHvSEap33qfN0BA5nPmuvDDb8YLormuc7jzMXatZKdroJTG11
S1tidZmRMvyw8BVGCj5Gh2TIsUj0+qOnHEE9Jg7Dg2YyFLQlD8Z393n++hWqXDzT
iJRzIPDrZ1AREVOu7EQi6MeOJlDAcgsONSjNeL+yyyQmCRs6tvQpg09WX0KC57Ms
Zu3M7d0j2V586lqaLC2SjhXABSFQ71piQTDqQCDWjXgei+5g0VpQ+M9NPHVVy5bU
bx2/7YMDO2CRHQ769OmC47pL2+kTosnq7pCz7ofvVhL0ZtFdutXQlPg2ooEvHvge
sWq6BTsUGZ1n5k1akjgV88MRZzAFYaHVzTdrGm0oECuKE6L1JSitXSmm4MIvxF09
IZzSHj/Ngl9KVb5ExP1dVVx582Aw7IF/1fIC1KPQeA8XDwbIz0Ncsq+3fpLyNT7S
6Zy+7kL3gpNaopq9BzQOAPiDqduNQq3rIw2LVJTsTnt9zHElKPR27cREf4D1hAdx
dX93Lj396aIVg4gzXEeTYk2LMouYfjjTT6jjlBP5w7cOGm9n1wc3G397swwlpZYT
cYJg4i5uH5iGzHouTWW5aoOmj0wutDPD6d0+xzMI/k7QPJcX+qbdv34JmT1M7H47
/TdHeQZCmml/NLeDu327iNTrHWBjYV+6oJotY3cZmXK+AhMgb9I1oFVR81ix7Owm
qmYhg9PWWKy1mOBfnvNvFBCBJ9yDQi56MDO5vKLg5YIbqrpcf7xTkJlI3QOwUbXO
YHIwr2fWxrubIamIUu4Xp/YwSBFsWNo/wTmse3Hu1MbiLl+ZseOL4nIlgnHdEs7I
g5PS7rOnQFFSboc9EMszZ1g88Rtz67rvaO/6iNzqdzzM7aJ93cml+0UV44DvLXr4
Xf279XRFW/56YUo4Ar32udpcLwEy3aDeNCOLOFvKm9EyMYneN3RqWCTAgE46brtE
GWVClv5Lz/8ULYamJ8P12HgTYm6IWtZsWwsNevuVyyW9DZegHoR2nJpDa2XvBfUj
6d/nDX8XI/D9CABFaJIY31/UGkH+qQwGtasQRJBiy9xLF6tuhjIMJohaa9PSKV9W
aGJFd8A8u1AUci/Eg9l71yIj8xCqrVbAohS/qNAQq9ECwWpSC1YlzIlPPKeSkg15
LoWacKACEnnXBEkSKckE6lixM2idTzsSwzyORZ0xCa3si8IHgNY3pudJvrzqhQzo
qgpa4Syj7Jr+vZqPqFc59xznID09wZwp37CCkhYEcK9HTZW/iT/hMOk1CMfYQ3z8
VhhFgSv1jqBAtxdUZM1MWFypZKxPF5QTnPNuzPbd0M3SlaR/1q34ITtlj6xCt86B
8ASGgckKIpjI/02ePnx1WTnmbrNXiFN9q5j681P3lMDygAFpHKGy2YJyt/h2W3VA
Q9KXvgbNszMZkiG/N0JocaQTeP98uUQDYxNRMKwGTAUjSj9p2WwugbgzzHs2RvY1
4iv+Q+Irxy8rQgFszRhtYH4lkZnNkPQk6rpoXuMst/86pJNKq6BzXQABhiMDfkRr
aMFbQHsv2LHoVVwJnZkTlsbLWLZyXKLsSjx2BjEOAULHUQdUVuAcQRKyVUPN3Jcr
GHNmr/Rjy7U4arkDev4UExDnNJlMidbXFrFALa3poLpLRSerG+hcX7t1QV7jxf7J
jLtM+XMOo614+kkEmOEg5OzjHi9+KLOMbbXbrqPqW+vzE7BbwhdYFT+IMrY0flLj
HtCQO1SVOik8wAKEHWywi9bjJzbDpGkCg4Kl9k9qCzXlv+OcquHj3kENy8Xrs9+G
F5rViKt9JviiVuP0GFMVq5BUHPG8aVkNeU66PbCa6kNekf9Vr1ezbYBHl0Y2+4DU
xA/CZZ+hrUS+IV0FVdukED7BjBZQtf4hekrzNDIBhJNvoKtTQWllcUBCPkfQMQyt
HLRBoG1sKEu81fFuAfQY8q5AB9BEi/Z528G/jMzF2SbjxBOZgh/YWrR+sOaAhHrE
Hsu7dxBT+lRkM0o45ZRh7Ap3EwQ8Yw3tI1blg1QD/STAgl0TnuMq6DoeUX/aU8QZ
N/ImxKUH5CGTo9LieKtJqYtQfslqUV3DS5f+Qgfd1XuGGS7JVnVpLRBJiYNU7Asb
oC+oAM/RiGiGjDOAlJOjVkl3RNQWeCd83cpkGOGRRGj+dHte0hm8ADmXNpG8io+s
lFuK2EfEbjg67+Ia9trLzp3+Fc3tOBlMszUqf3AhxiQ8bXsxVpuLICmJbx9B2lNl
zz0KFObFQA4lcJfHVXagsZOgYjpvRMefQCSlIPtHEUI8HzjFs37ezwzgK/lKTLmc
mKwgl3TxsO+LJfAMQsDcHNCRuYDLTahMzCt8W6/+zp/qG59JJUOOhzczDomcFlZ9
o/A8RmWOBegvEAtRDghusumhV6lv+BkGr0fGMEBgTfuRgksC15T0aaWh7xlpXT42
n5LfbFBKgD1bp4jsc1VphIXr0L2or7tSMWRZszj4oCfF9Kjoj+FZNsbZl3/AYDSz
ydnp0SUf3UKUrJeVY0xAhu7vWJ4T4nc3Li/0AbqVCY21tXZxdNEvd0MExb4+LL/d
bCeQ+yFRDEPjSIwGOqY1S2zZcrG46XaC41n7Sno+/+CeaeknaJvCcWrjctwRE2Ew
/mlhT2GL39r+A5dDTP0CIY8KT/Z06jzufs8bzAOxma6dJrnYrnGV2/rnRDvOqzKw
YJ3Vo7W7SzIA68YetJLsPikUh/F4vx3K87tqIC8RZttSKWfumZsn8LZl57hDO5Kr
E8TKP/a5ldquGJLQGx2KDGhqdFomcQJA4/L4IJhZZwPLKaJVLQbN5lnHaYXKgqPu
jneHhJmSXOxvWyANIuxatOqRfmYZ8GiHWbMSw55zmL/ppDxjQClAZzYM5jlgOM2w
oj2wUPR4uPFxWofRXfhMWN3v8EucwuAiO8z3BequhCMRt1d48YJ+voandhFWf3Tu
bkKMWs5y9jfu2L7/qlEjrrvUTizIVL5iYrFoUn/pucnk7NXr45TvH1bgsCUULF4E
qr45hexSFqm/5CUAT1l3mlJ8t6JLxCqhWkeGWVIras2rqWWOpON2aIPQAw0uzbUM
depthBPjnUPG5Xd4jE2aQWiXg9YiTTnTQELPMzaDjAHhkjdvVr71r3phCTxHLCpc
sXs9JFVcVnGMYL/Bnb6oYh5ldwyRicZN8/R9bTxCM3JIApps/nQEuS/2NrOBSHxH
34IsrvgANjgjjk7eB0GafqsWTNF5QKA4iA+VjunBBHvGt/xaCoXtexbB9aqH4baY
Y+gi4nPaF1vBkYdTnZoktBYhLBssoWT9gdgVvL8T8NLwz0RLLSArHWx3capzPEZt
8TjOKA5mESqbP1tZzD632Fe3Rh7979iqtU5GIQhulR+dJHnwZoMqVsnpuhdJTVYx
EYu10PRK024MIrSxiBgjRbnRqUojPGZ342OoMJfsPLfEYbyqQd7/sqwVIg9t9uBQ
3XyVoVT/Mrnfi/I9IyQlzbP8dYnRF/FnzgEL0EPlHW/r6KzWpDv+wmFCCaIjLtm0
qk/eL1+3HcfJ+QuL4m2qOd/yEoYt2xRnFc/auF6NeoiWhlFv/rpdX+14KVevwfJe
Enn4I4pI2aulBVjPszUI/x9WbqX0XtHA4wcvcJ28t0XLiMcru8rH2YDP2XDGCTDb
f6wnziI4DCIqW6hESAyHdqh1fOGan1UZJ0oDieTbjo4TLbId79hG3R31pgSoqrL5
8pgnerx2NtRJr97oi/FO1jjtUKoIgc2V5tgXkafElpWZV8kH1KYezelcNXQmmSaq
woNBfJkMMn1LCVfSyzHuOOy4KVUZPvBAQ+5nMhvV8P4eCleIB+XfGdwLUwb/WKia
EXmckcIJIE0vnlrhU6/w+NfPneZU1sXLuD28ngOgNR0i9n4blCoG2R+INNvYWdSM
qPttnB4Jw3pqMTCLuQMM3cpqhyfnRfsptdorWZmtK/M4L2a1YaCEcDl9swZ5L9JA
oHI0pYFRCDt0ZtYRTQNBgCsovMziNrNsk3kxi7XiTkC1fXXqtZqq2w0ezQ2KE0tx
nsVyv46KEg7xSnol43RB2+1ocTnWZafQY2t9acGi5QHqFCeTBKyzPfpF5SegXzL+
fMMcCDj1zokFBqrDzuM+F2iJfUhW83LJeopLAaZn4CI+gU9wm19H9bOUvdT02+wt
4qBnNKBk6DDUxO0tQnYmDYGGOBZWXoTmTHYk8x+yRCH2ilQmYw/p0kdZ5qp8C+7b
JxaLfc3sNd8xAAAswJShFnwryZZX0PmINZqNt2440SS+4mKRpGsGHBgsBB44E0cz
uA1xSHewZ7G8vdSTy739moH/8sg9LhbcVI3LJxqOL3iVVNEXmgX8i/s1TjrXATxq
1yrpcrx17DLeaZVyuDQJYvB9ucV0DRTVMX0outpQNUcz9BmEFf1mPC0yv5O1SWLh
4H8eQ0hn44AUmPuLHLl9xd2hg8Orvp4NbeNUO5VInxBYzhVI8/vqs2xlz1MWzQ82
bkPVTAkJTGZtawr/ZvR8uw9X8ywI70KbJRyzEUkfJte2iTJ+cr9mfh1o+CggQJfn
mM726Ua58beTNIyq9fHCeK2X/FxKaeGEx4pTOD1Q+00o/O4fJo6G/ytBaA+q0oee
SKWcELN2QcfOXBZBW+WsynDQTDdCJVK0A0fV6azMwcO7XcL9lEZL288TEhoKz/vl
TpMb0a/VQ+LVHl/OuPpW5eUvYvicxgv/e66eAXJgMWuMW+Nd6IpUOuEGQwa94ljh
UA5e90OvWlsCTQjHLNBqIQHX/z/F8eGn9diy+CxWs4VpK38IIh3H7qlUjnG2cTVw
aY+2MNe6QR/ooZdv8ioa+UPbJZrH5DmgjnkatwraWFw30ad/KG8BFG3uABPtqRPZ
WYtN+5FUrfBNRkNIHvJbaNgOpi06O8puUm+12Go0XDCu+oTxRdE+DtWCKY5s2LmR
T/77fWg0zINYFfHvuDPplshSKgjM0ZGMqMM9aA5n5ylH1uA70Jg48EURaRyGT0Di
1zwaJNfsdAz2WbPgTTWMOQazTYIC6CwWi3jViREpXVZnUqdTQP1tAZnO9O49ffC9
rAcDfP1oDgtXeQle5QJFILwUfaUNJ1U+CPmLUCh+AcCJkIhF9WX94iumdf/m7soK
OY1F4gGAx7zZ3o5yazrPUq5mzUePIZz/UMGJFpABQBdiQpdgvFIjwkIB38wGXam/
5SNEDwLcUAsys6zKIzktPiYQUvxR0sq3sBaJcR6CtpFpIuw6dfLs1z5JXh3a68uN
361G6M+C20FOiszSc/daJc1CwytYFfbBWCtcC8Gkwnu/rUERk4MTNBJiH5FNTCIH
Y7IG98hmJrjNSe4K4FjZvy9802yvgnbQ50hR0iiYdmMrMbCbg3o5LX+e8z/mSsAu
+LI1Rx6fCZltJ/Ot4y71sBzyXdnV2XXqsgSaNkizCAUcPMv4SQTYe8wxp9NghnKy
Ea8d8ToFeroNLppwC8iZG1+P8Afe7/DMmKr6QdCQN1n4X88jSZwxJDvH4RhL0rG0
1mn/cZ43zYakx9bx6BP0AwHE8Wsj9Bt5lntAMy6JTT0N0dEwqR6yefcIESvAU6o1
Rx6jcqnmqiJqVclJevCe9cqrokOWoKgZm6T1jMuFRRiiQgRp6Mlutlujd4px8G10
0RSe26+46380IbrXK6OdkXR29KMpG6VwXDO/B7BF36CtbRYzrkdZT1MhxQgJcXBH
VgAZTASj82P7cb4iYyi8tbGg4su58IBQFcwwxzJGg+GfQI9jSDKxQeUfq28uA8ou
P26ctFS3jznXc9WytRXPOGnUHGzetutRI7sCbYWrkZxiwdtXn7XC2H6t78k2GdwU
u2IvTlBtSBTqGUYQGqRJIVajV/YAqpDeJpj5KyGXoztr4uEVDkwPAEcaYcvXONFQ
eNQpRpZcTrXVKDiZeVHE/7EagiGXDXZAppzmAuhy2DS6VBNmzXYytQt6QhqyVUoT
c4/DvRxqmthQ0GIjzIbY8z3gkvDKIGJPbeIF7Vt9NWC5R4z9m5AjamfvkOQ98HnH
sC0GuG6hI2VDt4RtTQoamLk/Q9Jl4wJG2KGK05gVMOIY6N2hI6Xcmwbvzhp9dvaL
70Av7k8XVj3OQ8HFA0FlgtluwyajOLM65oRqltvY13/5nu0zLqkurgHTrnzIMQa8
Xug8zLtwu0SPAjZCbhFYdA6YyRciroDvUtNKyMEap2XFqAGcvSYNN1pnT8IicgNZ
MzNjRgvqXmbKVmburpczcV9r0todbQRB1vfyS87og34Xl6HXIE/07xyRk7zulSka
zLyBe42bPbX1CvygYRX6eoRi0vT/79ieTQiso/lS/AdyslnbHzlfvXqAxqnu/F+T
ioSOTJuMXbxaetHMiVPyQEnuhGzhdpFpsSaH/rFOTggZlhPUYnsIRYmo3FAx8GPp
UcS8kWrNBll3qxqB1gmplTAIM955rXoz5FD3bOkCd3fRxebaWal1XshkZWWG4rnu
B/8OycePsgT1Iyr5eJC6vi7eEt9OAT+KnaK2Zpzkt2me8vnfTg0Hw0seuBw4UleR
vFBWCP7dN4MLJSlyKh4aRZA33CI+mmE3ZirqmeuqfVj8fSNwGXaqQGCKgsZIgk4h
Fdpxm0CVbGN0gGafmZjdSiMs1WMDzvI2nkGElNzP2g06XOEN9shyh8P8R8gSNESY
cCkNaP21fVY0CsOEMAY9Oizv4EbczN06ZCYx7aRUz3NdQLTRA0nKgBIf74NurfCP
gvzl58ZJamaeLBU3+2YL8nc0znvcpx9i+CqXgqP6T1JpLWR74gLAfJvc8a2L3FA8
fLXLDL3tLlfkfKZQjKEtQkI4BCyT15HJQ2AsgrumHGRprn2+lAb2lT8eyWe33eb5
bUYiExskdvPeAXZBYO5d27FL5m5v9E2F5TbeW/E1PneAJbmKCrlNeb4BHsIVZ5Q9
3s9wHWabgDVOcZIzT/hRmt78GqH0QHMw2nDuut7DIsZtozh0UQMcjszot2KSwNmF
PtTuRjdOUdmg5cS5rY67Xrp942k8wl40aP3+jneFkWl365LqFHZcWzYAImYwmsn9
8XuuubyZQuZI4uwjWe7JOP6ujgnegQvNLSzvmaitA0l6plPTf9AaVAboOs9J0Ssb
jW8o/LRvwzemYL5c4l5WCPM3Xav6uxT1RSPbLOBQj3NHXGS5WAH86+v9FJTjkpPQ
1H9IN20tqNTh4neMetmb351H1vi7IBqzjO9em01QOFVi72xbP7k5MY83KCkVj+4U
stLF6NuKprydRdTOmqfU4U3vGV1X8+l6zNxLOZ84nmIpc+sDRJerVbk3NAdOoHZn
t7e9CrrPrjPXZVewepGS0oA48FpfqxQWbf3E4sl4FQbVVjd9igyw8AwHBUfIl/Ja
0U5Wnti9j5qooDbIwHu3PixwRiLD/kE7ElAVp/ZR44i4cZDZa3xK1Fl3DKI6ttoI
GQlUtVKUmVFGAlYmxeDRKvAwKeM7ymYm1iwDZI52B1kdRLMu9A2ZgcWyrSOGiWWR
pit74+r1M8Wq35IaVvZIJJbdWB2YPq4fDjERK4xNUEPtN4TwgpQIeMUYX3DbOHyU
Q8dbK9l81G1WZv0OZcR/er5JpyMYPEuNG426SEKCeDrCf5xwcG+0pYy7Avpr71rX
/LOB6NUnXcinH5BCudVdahhxLczpRujEgfb8S0LODoVdBHOYWlyn7oBOaRDK8eqe
eBUbcO7QYZtRagbZnW8gcUlNarWO7KKv9P/8hKrn49R5tbJ8NPYErB8MEzNOyoBk
nwEYsZ4iFA1wLPW/6X7liMyaLKv4AvVqsc8HVomJvaXcnzSg1mSv/sWHqx2Hq/lJ
JFncFfPQoFGFoMYVjLeT7jcAnnPqI1aF/BoXOLcAS/eIR2t95IU63ED45VPl5sjX
mlvEXALq7QtSBzuX8If3d1iJLjuXkZNUgcGG2wmXUEEAIcSt3gU+yTFj8O8XPvcA
2IrrJNFMKyGRDlN063lLl3CE9mMgPTh1Fmp7jY5NOpfhskKOwHpBuYXYY9V0psCd
jsrVYs11MkQm7zMwfEa9Q25Pa7Y6EAddcrbeOBO8w8i0tHIzQfBicqJoHlebKKhO
2koRYlkvkePLS3S061r97rFl0cFGxp7jnKtcr+TcwWVr9gGXb5QtUxx8Jb5ALk/k
Iln+h8+4rl38SlDAA6rNd1AusOAVaMe6XV6cqWC+5vePMr+4KMyqZ/XrK8CUWQgJ
aH6hEvjga2Zc3ARRZd1GkS8eseGb42z4yVnke5e7erWDJhKnb6KlQn6FDx6dSxDQ
e4JYBJzTWLcOW5kQVWz8Fofct1tTLB38/ieEO6d3N1rAVnUpucQ3kpl8mIb16vbO
sNQ9d+tqJeysOiGN6tOwW/nrHA7ODggaZCjtafvRo1XAcvkp7gzfvoRGW73IFrd3
Pn9itE+RwRcYTfg6Ejy4MwyV2GPzflYlcZyHUlK4KAbzv4sjI3XLClxtd1mN4zxr
yYkaj4khqoy6rVktLt6N4Wq1A8zuNx9fEq3xIZ9TlEiGYNHD9WMm6J4bvLWjNZev
aY2Lf/R9eWTJjJ9DUq2JUM65fqpO0HhZVlt4caAXlYwI3CjDV+rxBZrG2K4rv3+i
5Sx7Bxofb4/GwUYk+pUcK0eCum0ng3nu4g5zJrqb9BaLQpXBO1K0QVrm/dZKYTXq
101j8yEUTpwN62XOWBB1jxcIM4q0yrPF859piMTCfFUahUlhBViVVnkb7lPjdmAu
6mfuDCPYfNreasOGIterpHbn6PdIBFcXlPWg91LQclc0QfeNrokeiNR0xRfVYmF3
3j2tmJV7v/lsxhy41oG/MuFBCGfYmH4/dSb5wOtoVdGfgTJoXGA79bjKhrv7jGab
o8AHISA9R/XfgNUMG8Xqh/C3fZvu0dbTlB9KU5py4McS/9sM142HV7Wm+gFxXnPP
NcZ/ETMEMtoxPCx6I7F4Vr8EzhXOhKhBaHqeVRPb1dtBv+hPpSPrTn65Y639T02A
7e8vj4OE+kWndXrfZmPsgNgQrxRB1HGbu8xCZ9RMl1TkAFSWhGQ9MSUBQLv3/3/3
TAgmHvHu7uqsZ56UzRNvARy7ogLYHOcYnN0xfe8qkhUj2z9QE0RglMuPid0C+KxT
5OqLULYZNXe4XToPGKXC0Y/KGZL+/eSUz5MpwVt/ip6Ti0FxTA6V5INbS6ywI3C8
M5/W0DbUVT9oX+UZ90+tl3OMT7K/yWSm4yNYfUxtqaMOhJMZpmhFOWXk0bQqthp2
EL9UIyvkNKek3pavN2WtzBR/9bg3jWIPux7gZ9ij0/9aY3ajW51z0+lbvWxi9Pu2
Se8SRa2xPP+SmdBvYtPSxSliOP7OBmB3g2zStY3yg5FJygXL8XY+NiYq+L/WmJIp
rP8eRSfTKxkTGVjjteWvMti+G2YslC+L55si7ZAilxyhVRzC17B5V1on9V9ouZGy
0BjhvO3vjcLJHxRVqPazXL+02rBAr4r9ZXPegCznZCzBepy662x0wXnao0wRUW24
jxVd/bQgIubgmHF9DQAA+tm2Oj21pKalZ7vqh0MRZG+Hu6HUyGIYRKaXEYrdK9mS
YFwAIc3GeSEdVRGhDkiXQ28zyqndmhuV4PWaLDS2Yu9KUE78RqDL0jQ/o/pvn95O
f7qgkVr0P4A9snWvukmvEYwkM+ZXco/DHabZ4eP+O4aeywq5ickgLA96a9mh2b9S
lDTHld8o2/Ndn+YntY5rUae/aQnqI7YV794RvURMCkzlJURTYBgsaU6gKceBYDU+
2Q6eT/a8IkbRRcrSGSFv8y1YJhFJh1Nq4w9FwOgJxczJr64c6/w2K+7kU9XPTSWA
6nC05rT4FxBuUc3hOhEvEYJu/Bs8wAi87EKjyWQ4D3s7WT4dJX11WIbv2Mc3H0K2
8vxYnBc6Z0avdgbXPPwek2CbJE4QjidRdb2xR46HS3Ek22q6YUkgYWMVVcc2TdTj
lK5+6SqzLlMkR2Rqi2BMHGw/yJ+3ddTe/3YtxFDhVA74586/5Vvs549Xh3w3Fq57
1JqXBL8L/7pRvb/CMug8uyh6vV+rYlLZIsAxzzoo1xg/mH/78b61q+Tfqfv8Wqzu
tm1sT4HEsiT0YA4mu0diuj0iU/f9DjPL0xAKdGeYM7sVcnTK7oOZy6H8roKj11SI
VYypMqocVzQlqfTPJSHWBVAvgw2xXaf2zIdXivxtcqbYpN+rRyvFQD5RQdSGxJpD
I8ss850NLd818tYRQVVxj4/2tX+LqZSbxG6sYopj3MXuZ6O2SXOEbNrlXPzlSKN2
16Zf18FkFSJtDHzNqPhNJul2VfcCahrVpXIFm0wgM650HWF4LEKcv2YGY1gSPXOc
ZygiX8KNeTrDmmH8OdhHzDKPUXohMl5bVMPOI8Fpwe6ZUmWgcpBv5UBmRBtI055x
7E6wrzPoAd1qTLKrI819C1MlJm3cdfea3eRiBFdraEblKTyJ6fvCHqlK1RvX4hwD
rVerl7vox1L9Yt633LtzUkEWkE7y7dcYVG/TvZw+SwczOLAm3/IEGctuu37XKaz9
ld/yuJE1+nbUWyEaDX3keZph9gHcQQtqA33v8MZvx6gbskx8sEL4Ss8hjx1V+QVJ
alv1U2HNdmbQjLLSgZhHabWdyPwjCkMp25nzQzf2tGZ0AuzEEoaGqJS1385kkVh9
PPj+3h5scjTaeMva3z9NdLhEGsQ8ejyjym4mEWCIoIFdLxtfiL8ndABwIbD7W1tG
DuraTW3LsiaqCTa0AVRzynmazZ/S3iGTZA8Xbhg1IF9hV70M0PWGqrwpZ1X+cTyc
D4QW1JhUiXpJj+6WYKJR0aVP6DhWkLmR3opUHzJSd7JDGj90ULyO98D5aRjARvN5
mkeKuEHDUeKzF1O5gzxQhc4XB6FnvRMGCG8zqLykkKz3ej655BbBtL0oTEPdTA15
a2g8u79j7fVHzHFt/hg/X4CwIeb1iM/ogxbBpR1wqbMPY67W4vRMy6zlBs3Lh9jK
z3TEn7tvyDcVLdr2FR8GLrPMgVfyxaCFjHnvGyDSRpRv/6L1YURShLeoM29L0ZIP
6Mhzo9If5shLGB1/+f/kcuLVSWaZWnv3g1ubbjFaY/X3eGLtgiWHJNsLj1ALYyq/
KmtWakMoLXaaPFE331LBwlQwammTtI/s8V9WQkUtXaGklHUZX7rHduNjlYQ9trow
5P2aKg0nJ266Qt3yyd3pFVREJncoV/WewkJiRg7v0z409FVBklqK8hKUscma6SA/
Amx9GYlS7Gae8dPXgKTwJlDQ2Sid1ZpGN+thWY0ZmkSYUfnzfyB5V8r18i4dNg3X
WAWRLrnK7MbFan1b8OIqW2aEna0VcCs9VLTYMLZaSB7HczaAPkAe73vJjdbtYm/A
+BxKa3tQjVtLxeqaoWV3HvYipBGQtLuA/UJD+TKAEHwf9tKJj/La7vnEuMrIbZj0
7CjhIhFvS0bwbfCCKY2KOI9dkgwTb5s8CUP9dM5PBLRR9zZkjwGcCzftUdS7DCPY
zYP/IiQuO+t++X98NMt9W7oc4KKuw+qwIvnv1RXISMLGLyy12AR2QTZe0nZiMCPI
0wtv+qef0aT/C1/0K2T5FLDbvx640qeX0o8dKQ0ZQ5ScOYg8u3S+Z2ev2D0bKa7V
wv1HEHGsHJ6KzOlpGVCdDgYvElkoYb1Cz6XJPt1tvSjN2koUVn8SYY8buX+j3cZ+
bjeoyqs/z4Fd+67Jg4dcKAOS6v80aFAF9bW0HQAkbRQ8TEJ4+DMSxk6+dHtqPc0n
PbCcWzj+RuD7MioW8hbB6ol/pLIb83NrpfNPG2H5LbughynrCjNPlEasO45EMUyu
I22GbKEMOGQJ1T0JjMPRbDcsln1RXFkJNacz2acM2MDH1jmfMdtuYCThWXW4MV4P
/Naj6xEro5EP4bmuC0Txy5NvNh25eQuMwwLDFCr9M506adtojkxcdO+x9rJlzoGp
U+OrMGl3MYKRSZHACOd9H9SKcMPnQSc+X+pqy+KsBaJLY8kvlv+ByxaTrLsIaaoe
d9UoUsebawBEY4zFEd274I3gkEt5ZwUc0o5wg/h/2poOx0wPkhHswJGMvnX7udGn
s8XBlmnTKckLtz+T4CcbySlB3GeEZzdiMIVWeXsDHAxW2fz1UAWzCFy7kRnn/ptN
oCOkENqVS+mNV6VeWLzZ4boFOF4FxLbaClHdihd8WNLgc8cQzOemajtV4NwDVqSU
f86MKVbMo/7Lmi6aKGj+RBMfV1yVPAdp2OCF/oN0gff5ZCc7fYc/ObKKrjlAjI8H
0XvQwCZ8s869LgJ93bCNLQrsk4hwN1dqxVS6EBQhKahKdhSDR/MfB8FHPztS1pDA
15fAaCtvEjLiDTcd9adUK+6Um3XBoG6bvIJ6/ObjKre04nXSyENG4K+GTVSEwJQm
GwkUkQlo8ec6kLIY7QqnG/w3ivXuB6BAfpnhi+TsucsPNIQ0Uy5sJprT+e8a72Rv
QRcJdMN8aVnM2JPu8OB4D+Jo2PDkC8IlyMYVe0ugJvkhFvsfpyG8+XxgwNgN73Af
HaMILoO+ec2bLF3Kk5qLb0lDFsacpplE5ro5ly1TpjoMc0BuD0Vf+TahM+zyYVVC
dO9PrmdrboIZr0Q8BTTI9vL3HEVet7o/FtP26mMoUDALocNN0jqMJ/qpb4xWj8XX
+hU48qFnMdle45t1/tTz+iZh8z+wRUQYbG5yuv+a2KVQW/7FahGZ3bEXskbbURgc
09clYgiSEL85kKnTQ3YFciooSclEQ0EvELlUkxDMNrhNZ+3ilH/k/f/nqLTfbupJ
8WOlaXLlPICTFl9IO3XGdDBJBnWBtBd0lOT+lNJBf0xTH98MNWDgiwuAYH3KdFZC
+shVvRTJpwZt7jO6ZQnWf+fsGKLAyha9xD/gMb7LQqsTlQ8vH6QSkXhrgHhIl/ns
AEcgQV2OHMUlb+1ZvQ38gu2B/5FTS0KrUW/LC3mPYgzZZkwTKcjSC4bmUZyu9kW6
PcA9KY7x/XzMVN9RZMMT5BOQJyTlSjxudoEDFGNPERu2nJEt5gy0puHAv0l7kGsg
mH58uFR4fu+fy1jr77nvKwrITAHnHQEVUTmSgmPmiR80TWdmXymh0qpsRJfPOpN+
Hh06SHZukGikiO4izPv0fXn++qd2aoWFbzWwNiPGNNOl6D9Pb6ayjLzoZvWHD5kb
519QXuyzm2cm9zQlQA0NSKEBlaqohlBxVay4SGzXmds4jA24f/wo7sX7G9hDWLkJ
YXlxOBHE1hm1JXxFkT1eVi/tZEjA2xzqcowxCegnHOxvDf/an0+AnhhF1VOwFBQs
zLZUE7W7kwS4mFhhjCvpQzNd3IgdICl7DhPzYaNLdCU5NW/jM1Ocuh1W6clJ3P5b
5S1FdMaaRxrYCHzrazhRtsOvDgJXIb3Hu/KlkxhIdecGdopk0TDy6nUcz5vm8bRy
HRwgoEYV/dC88GtLv0elgzCTu1nGom6/eND21VezhnVVh30f9+rBNqxr47QJO45z
zfCW/EZGN3L/NBHzFYmycJSB9CtHRT9paJ3M5ZsTeWQetIbWGf/w1AD5zsW9HMAg
gFUI99Dly3JoOhTdvrx/s0qGhgvlzttiYZN9M4V55oSKFUlR4d/XDiSYP6vpckIv
4BGzWwXVIgaBeIrnUzBTOwFFj8OOLKmpu6bqVwLVpzC6fcg0cFNAEz6YBJInTyAF
t9IEqOmozxy0E+/alK3n2WdWgqq6GevsHvzUCGRA/syojWJPt2u5qlOh1HfravLv
Mxknou1PQjBVBztEbB81bLqHPQ5i0Zu+TPW+tvRYTfu9oWFzgVi1NVUVsbdZ4kkY
t3v/GMPFaOMx7a/b+AUKV20STU6VuIH2X0BWoBBlpPN2zs803N8o2sgHY6IJj83F
0HjL1+Sr42KmcZaEGxAzfS5iI+GPFAQUGvva5Lns6HF6uRzn5ToPc/6vr6A1vYqz
Bh7asoM1l7sTHM8RjQuf7+2CnbzlryreMCAi3JZkNl6S7f44s+F4vDOgwd4aJXmm
2+EbSWsaRIaIzMPIpvNxoafKX/UHzr45WjokAemQE26Fi0nuD95+405cSgwoHtop
jIdQx2oJ2jEChHho8JvlARuCwCjsL6McWR78X2WJNnN/8y99xyPwFiBoAyf/qVWo
k50Nxfoq1jKFkjkt3BmOVTgE3B8eBENBeb1/OFU/NsLK6FNDLDOZUNwNp8MyPjPy
o+2Vdce0Sw2IFs287o0NDjQrK8RMCgSMt/B1EUkzjfvV496grEm+1vR6289rrjqr
sSG2P7SAKZrWXXiZSxhAnvuSIPfQPLRgEaQhge9pCmw7UFzZ8cOGPUHY4yt5X6xZ
SJYzhW2aYIbu5BoiN+DwWY8M2u7y5S5Xgx7V0c/yAYrQFrJ9MYUW9iHub5l/HbJ6
57f66+ryKPMCO0SzC3OVEm05gMYqlKhLpCtyo4Zqg2j8PJkBHz5Nz7JRtaSAyFvN
5zgD3/WVivyoQIxKWcP0y3+7ssMemAy2RRvqx02LZXMry1pZk7ndTIzqSiEc6VxS
AGaWV0bE7tDa7KPe4ng82AhMTY3u9CL1VVRNaQALSXkgGXSafX4fFthwKqgIgit/
OnPJfcINEa/NIQq7RV1fE+t2jSpuZmHeKzKjmizqlS3Tg2Yux7AChzomY5OEUK4S
Cp/q+CNWUFJNFlgM3W6CzihstpmeWeXsnkcf0v7pAWIn/WJdm3MrBnOTJ5y4W6p7
7vFNrYU/APFD54hO45ojEasDlnBDiFHta4Yulu6FKJAJYxX8djRVXa1OSRC20knF
f27wcCytX0mSsdFuGA6VPfaGqTmgQZsISIpPdPlJIMwe6V0XuoOm/r1p5uGYjsiY
o7hlVM59lQK8OCo+YNSfvtQQMluvHC5zwhhiw+ae836V/uJacEXSNjjis+RMz7jO
yZDPKIGJ0kP9aq3Z9WcP3jBQZZXwNVmYg0I/1Dh7rTxViHnTTqxq76oWjTI3YrUh
FA+z6zZ5p930IfpbAEaueQ11DuLNPVVt+DEiFXpMqlMwFdoRGyIDChxbjVQPVjpT
TqLMHs6pZWazbQwBoWVcHRbbxz25/iTagqbeMoz3djSLD21/QZxjz2RPNcJ5in+f
aFuQgYqgBXBfgunWPwDNGzDL9iz1rIFxi6J65sfugLW+1tdtiy0TK4cxXhcCkgYv
/CDvrXXd0PfPhbcSi1qdVM6objC9z85gGGUitgHtWxpGRyIJ3WCITvo5B4XDdzJi
ahSWADXc24PvwA+Z2rTpyLcImOy8WSsjVG9+Dn8SpfdqbIGirlOPOkBe85afKIKk
4tfibKAVkwhbkkTTqbWku1sYeSv4WepNN0YUP0WxTbv9wHRAv8KJ/cfFQhKmFL7f
RP4/tgPtJ77Vz4M5sJ0io+jWYFSactbfEHGmcMAnuIyQR5oitSLIn598C+KIZWjI
TRRXbdaR8UvcLCQKIlDWp/b88NqkWIVFM9nQj99knxH2c7jFDUd7CRCdMblt7YlE
73JS3lg93u/rFno8XwjNXkjuNftzdMLEtU5HUZ4bnYQ7mdKjlw64W709oN/Ch4V0
agfX2C+CmI7XjoE/vrvbAU3+OuI+f6UIe7ong0kHlncHXwRN1+2xdYItG+INOxoG
p/GoWXTqBPU09C1jTG6v0tNqygRM7S07DIHI40gR5fyu/Aiu7z5SuEnEYEo/zSr2
l5pSHezMDA9jUi+P3hh7H6vGpFFf7flWMvxYeDepSMMshv9hjhaL3uq0AQTtwK4O
38u4vHURl8LexQn/nJQoSc3Mr3c8zRGbciCNRudJnUOWmo/yLY4JrT8dJPIt8dPy
L0215bg65Rk8OP+zEsTU0UtYoajt3ih2UD75ptw9SaXHZOP5AUEy2ALHWYLa4f7y
RTC6qqr2YjhtbzfC4xvgv+sppekwxhGmm0bcQeT8wyNpeSIns6QkRJzfV7KlXLDs
AXTyLIgL1OfuZqfKCJrRObQe1iJ5uh9P0U+vddiGFefAk5BF8NgMKXT5wN3m3jkN
BJgONWo5IfDLPrxyDyD3dC+gv7bMeUiLwgcEHm0e7wtkQyfRZHSVA9JloE/b29Y3
waMCTDV32AebP3rxBgNQbRrVxnytjymXtJUZK7VFBw41qPbrNW63N2xzQANPz00Q
otkCJmlBbzBLt/5zbjEA8RjeViSO14sQEfZeuRSC9/cQkQn3EjPbi50P7zH7HwMv
bS1HwHOfQXWxIc/W8tjREIgPLLG7kd4VeDpIg69m4SIs37Jhq7mZdstIX6pFbQfQ
6k30kSF7xmbgLt87bzLyAJwG9wktfrpPJ+mpYkoJ5Jvba6zzZYTUOxVL9xd39FbV
38snmisBujsOOJDCgoXDux5j5/4AjiRuSj6DnBp4gUkdrTmhmYqddtNUdrA28mSF
HiQxq0GRpGnqJGZYlUU40eiTHE7y+WB+F4KPbkeWUpKHkexQvaq/K6ydk0MgeMZt
25BbOsXZazsDGWSJfUdr1rDJ1Xjn+CT6JYsDitVTpMDzWo+7ik6tOc01P7WXc+ED
31OfVlJwn0mbvIP2hfHU5B9sdrmkXCdh1BrqFPD7F0SrHJlHuzDJnyAeOIZtcH7u
JibsmmnO9ysOLXVebmd4dS3YJzEwNRfn/0yJkpc/m1ArCfi6h2mPLW9VvecZ3w57
hWPKNu/ZTwWCQuEsmAwPgqIR1OJJZdRiXGLdn9W+k+4xwW4KVnNVYeukjCkpyWbi
HaWohJ9rC7Mqf5F5UKQdBSBTCw9kJbTzCrLt5OTtfqZdFloZ7Y3kDCLBuGO9pTEE
kd5jM2ATW5kK34uRd8gmI4AjfpzBOFQTM2npnbsnHmd3E/7aeYEeG8BjheML5hWp
VQRNOZaaDSFedCQK8Rj+zEcjuolA3BHVtMYNAtLNcWfvrw8HI2OjIZbut04EWCpr
rTEnoM1n+qFfeWEirGHUN+efl2Guiq2ClqPVJf9u1YzAWyOU3sKcrteACPAHSvk+
rS7kDbqSozmnVueaaj5o70czUo3l/gR4ADfBWHKDheBmm2HJ3tv9gfystQlpRdfU
bHTf/gVy8C8KlJN9klJC92Lv7uWqukElG2selSPXtt8ZD7LvAiW5ow1PWwH0lxh0
Gh8MuCBxDIeniM4PtKOk1Ov1BToJPfCjLBl/ZzHdkVf/jMM2aNbWUSd5Oio+R2Rr
qbnrIbnaSbXMIzBK4dIvXw1ZEhigUTmKvsDjvobO6OEkDoU2oXGseIJXtPkO4FKj
T6SPaD9buyk6UrYVDHoQ3y7DC7VVP96mFARRF3yPAB9xPZUG9TAR6nVEezhhisBM
g45V9+rxC6cMSu4PhZDmpS8mbdtD9GAok8ZMNBV4wTa6uY4IlfPrnD4thVDoXXiS
avA+QftFxuiOrP7I4VyFRuFedzofP7FffBreSZ4oMJGwa/J+s3DUbww2ZO8ikrEy
zDClwbs5iRNjNauKnRn2Vf0CPESRT6Gg6+Z7I2zY/SYxk2bVLJ/CcfUdEvJRRdSm
ShbbeU8NadbrRN6dSjqf3+WnNdPlV8CwNkb62qS6SAUDT0/o9LXWaqa/bGmwL/OH
KMRRIejfhUks/9X15nwklFX0dWpzDseGEfrbWOIeox+TPAx3Hn4MsDzfKf+TMTo/
xG0iHBqdlBEDg8u4YDwyLyadtIQ5gyAsbuzZdUavdljVBYVbxZeQfXp0TBu1vSVO
s47aAdMrxXsfTKNK3wBODGgXbA/rREddFOICuGkFRscm4WFGxq7WhRp1jfmvf3e5
5inJRlIfISkOtZ+ysrzAmTaj+9XH9stBl2f3S0Dpfmm5jzIiEUhwF3hClrURAnlM
0MiPfDCQbhj8LNcGK7+HiiAVGJ3E3rhhZysR6FwOTE7XPZUmtjtoaha3OjWUhXgs
Rx856e6gJAtxKinZfkUJE3CT0+WqKnOQDCdH5eetpSK2azJX1Krmx7BumSPVvNcf
wkvNR35BXwWctsy0TYVVLrX0FihIo2tDmvwbKl9pQ3Majb7CijHlpvViAIFED21H
jdoKe16oeaVPTfGA7FHIXUzz4dgPVIUxQp+C2FOY1x669NucyYtRkANQub7UJAsj
IdqTke/8zqB7UcGr7lTENvrm2yx2E/3cx8wu+Qb05to6s7G0WkB/9gj/3Rk3EUeu
iHbRgksnWjUDFFn2s/S0bG7YiChqM9t5+BnJw3ZhfRT/6Z6AeJyuoOsdCopO2PvL
iCsHBKK4h7IiYsuPtc541ztcLSvuWUkAmiPCXyJ+eOCW2/rJ1GDtqFTnHToNHgRw
+7uxa3p+bA461p5Xext22wRuDwb6e2dPy4YPcHC0FU8hpuLZBLhAeAF1oPxI5mWf
Dv5EWzAqLnscETp/sfWKYP9veUgzJvgmVzrpOTK1WvNNR3VWMrYWCnZHzGQLbEcw
BqV1PUuCC9FSgSfJ+OCPRUTDWu3mCV2o/eRFAVll0AJd+yzLSubu2X2ubPsxhwTg
cjhTMjUpZsVlWq+LbdMm1aQnryeXa4pbqN6vv8POKD/wot70dIdNNUkjr3LcFFkQ
eeprcil3zYpd4i+A2WrnJPPuiZy/9ehNdX2hUYMC82b89wj5wGS/wq3YItW8iSRK
x6kuDZDh13YN+9v/L1aGju/OGM/mgc72SL/udlBq+fWNTLGQJPf4HPBJNmM2/Ybc
cLgor8mpbu4Ppn84aZjeHfGfIBehZ48hlG/bRAxWuZOFUrK1aFbMp/IukRvZin6B
kAqVDWj/aPqawt2wR+NxsZQ7veIsVFHWf6Y9yTnkY6WuqHmbd9wB1NelyasNN2mT
TVrA92bnNd+4vIMzSfofKfnAtszaeixuk98fTM+1uwS9IqlhcbnoOYo+fdBMhq22
dcgGmKXJqoE4XUr2GPgWIn8vsD6UAN5pVLtERAINppnK2Wx/6BLAqrscv3HKrA9B
Eo94AhJc7+ETpNFx6xU/1NRxJuFPEfJNTUvaJnU0xlIKJNg/9mQSAKoS+iB/R08o
YVykO0zGd4yVsw8Namz13VRR4qGW9mnaoapLIidIkdG4j2huDlTziH7eOTd3TSpK
4RrhPbKhGpCit0Sj/d1Md9zCuC4o6+uVpZWcvrpLdrcCObeb9nKIyl7Wsk+rfmii
qiUMHcybg9SmmMEGSBr7MKHSENTy+J1IOLrRHJtZP0JY/LC8tii9kdYoyzhjmJ32
c7x7sejXlulJFASukRQKuTLDzeB9Sbk/Rmr4e/2DUc1/3eVnPmH86rOegEiXobyr
+NQ/NkcGxPyqeAYM5xPxdMYydEdlpNvIlfN6yWG1nsA+nNP+Vk1hXZffJyzFgKoB
fsUc5f6hCzouPi7gSxjuvNa0tuzucW7wfQ6fCXnGN38ASs7d3LKaNCHwyh2f84oB
7wCEVCB5v9kvNLCOxY/9FVa1C5/hvGnF0i3+wCqfkgpwcng0Ta38MK0yTHM2mW3t
6FV9oqEe3xv35Nqzf11f/brQidSdqJF3/Pm5W2eFgOey+ICDYkpDzM/IMQs5ekBA
dmSIoi4vIudd2HeUlXAwScTkTxCuhV3U1ziMeBMQ7NaFz1/9zyQmM92SvKXr3IkE
eQUYljG3KTCGeDvwM90P53Q7q0d4Gy9oqZuZ4gVyU+GaA9NrT3xkNSWzThn0BCHF
sQ3wbbrrR3TDI3CusfshHetSOIuJg1qqfvCI9AQymQJDn6tqnJB9QFURsWYTPtM9
jF5dXdotIVcauN/QY0VXteepjvSG0umhhOIF0tPwnEGz3EpzYY9RORDeF26J0dc/
6uX6GUR1J5XKJD9/ZxjoKfgojeC3HtrNFsRfvuEnEMbtXF1PEKl2sFioAlemJK2O
4F6uYXuwnwP5BC4g3Oe41YbYw6kymNYMgwg2/+LqIoySQ28HJWxf69MaUpTw3R1r
9R157IlQxA1DiJqjKnziJoup5i285TYqu95B01HryLcxRNAk5Y9zIU3B+N+Dkvcu
I8n2eeP7Uuqur42TYITnjQ3PgrJjK9EdSzAE+hWDEdkzwcSsdO2mZqDCCSugPu7/
bLtk+X9xrZZO7NyFUlz0+KNwBc6PWRe3u1Dh8Q2b1Zt/J1PIm70Oni2C1e/QrBgD
/ZB4qsZzJlfuMyU761in+7eO9GgmYCC9aNrV6hW8TB3EWUCeWXp3bQZMomxGnIKl
gpwhl/kecXawUEYyndjMeVAaW1JqxeGRTE4XhvaFILATtGFn4YAiFO2grKlWtGmQ
z5SSc7cfwI/L6gr0hYxhP5IQX2hwobUk6CM/5qBvfIx9E1zXtRTxJ/BpBS4nqLbB
8VJjjXTomxG+JtY/2A2vfwsXtBKvo/ts9MAl5UJenhXj9e3opFi2MLRpihpTYMKd
C+qOwVY83MyLkZhRu8dTQRy6388R0zGuAm3tHKjrsiDLMA9tO4yrPhQ5HeMm7mHx
VHCoC2o9hQfR2Y//hky81tCi1mzCSHBFZffc1cIRMBIA5zfv8PM0djYjTRJRZ8W2
8c3I2HzzvAYhH2IvpUOpQ+S4xfpXSH93ocJHkS6mx/sySExYqoZB57Mb42WjE89r
hlWAKnLMN+YSoZpeis/uEPeCSIcFIi8dhA282u5ANjFsdyy+RCHqwveNDSTGIq2t
euapmDx0Q5bYY/T9m6Q114udq8+45uZDXYQg6r1Lh0DFa1exSzJfxn7Y0RUzAJSt
a1rfNlFAfukcl5NhHh2/YZ0ep7rIUvUtFZbk2bhNFsuMsHrMCAqLQm+/Tf/gt4ub
Csd78FXrU8SsynwW4UV8DzkpxJ5RGbOkTGcrZPzvDH5mLH2OkbCuHYXwy7Tzb460
QycD6P+jNfQX82ppR1nbWh7HHDvlUdL7b8MF9YEt6y5Uh9w7bZlEL8HV9B0Sj5Rj
L6nclUDqW8IY0PHmQodzs9hu9bfTHbAFDzFHzyo12fELbJ781WTYbwhn+/b6+cYM
yQmUUmKLR6DuT9MoT50YuggFc9C7BrhDE8EzSPiHRUXrWt78qqJ1tnd/7PARAxLk
aYxs2QA42kv1Er0V62H3v0T9YXju2PKEGoM1QTymiIr+hA68glF0T1WReKU8QnBF
+T4nCmH8Azle+g+j4iwgLqK67lmRXZQXuCnARZrIQ9OYfZx3h1yM6Zqewa4FbaVM
SEiBuTMUyB2d5AGNAsHxisJS6B5OcF56F/30t4p3UufSkoB48Ucw+OPCHKa6EuM0
7ZzANEUXofREjnJ3+uFf3Bcadwfd0i1zCBlE+a9OG8Xa2joAZcwFrMPQuGpAeaic
MQM/rkbJwy2hFcPGNgEBZ2itd2LvEO8XDAyS/dWswzxQLLlOLKZhH191+aOnYm2C
B6KS0AKFvuNuUI+qnuYgng7TdTi9l2VRE7L6SFcG1RTTwGspBiZxUPN/cilMb8Vh
S3sxoaVM46rwfXMtYzWEkfK2tTJ/68Pcv9qtJ9C9Mie25MmwHe1nTy1b5wGBFL8Y
nUETnIpRgNB+zILT4r107jN3UXZrRmlFm385XnptWqFP9snXbeiSRrc2SF9V7LHS
GllyRDm5SqDV9q5sngpO65y7yyXW1cxtlxpRUBI7ycErWgo+DvX15q405+feHvtI
kz3SEvdAkf2xAw6jejAd1khJuuzxc6a9kWDl27wmlVcn4ima3nz+wiTC4TWV3pUE
ZjwaBlsuJCza0xIqGrZWP9AJdBZ4u24JaJm4SGcUga0TjZaX/kMMRnwuo2gnfUNk
AIOoKxNm0FHCWA7lFH1clmNDwdAqsvIGM0fh71REHlZ+DjPlwYPAXbadua0OkZgR
2YLME3tZllyx0NKdn0thqFZveIBVqmobP+HxMYKNvzagDDFV3FFjpUBR02u7fWNo
meuonuQa79jfQOafMWEZ6d6xZedjPpMtNGDCvSJG8pDjDDp2pT/LGVw2jTzQlSRO
90/alUx68JZW8I8i6KTEJKGS7ZHHys4uOFmqD0jBKxzoN2eCvjpQLCYMJDkCuyjo
jgKe3huhhbl8Kkiz/HDC7xOc99xVAv+TqppgseKoAlLZHzPbAcgwxmfybU8mGkOL
0ilZeWpVmMVF6Lz8BKx57yaXfljcEUr7d4poG4F4SkhPJOrtheyqWz8cz8xKb8UO
sDSUc4iD9HH0TkPsyF1c9zgrcKKH3FBPR2YfNEGU4EYdf5m7D/Sfl8jcyb+002xY
YeGnZiJKAKiHWjkIygnoGTwK5jeYg7wGZ1IZ50NJ48NJ1ccXoDGvLiAd3GINclLj
nsTjeAO4Ex+8rjF0VbhLmEFjPCjJWU5zaxmwfr7bDSTP1iTbRpaZ5VrNkYLK0uPk
m6x3f+FOBBk68ZqlExdF9975ruLrk5/uYd+XGpr8HUpecnRHwxo7UgbqUv5A9xWW
uN4pqMR384YfBH4TGIeT2RM6ek1hisqoxtUgoSlo1pMcr7W5LKYbUdxbbL/lgMS/
yuM9HsEHBkBub0YFmuNeIgYukFF1z0QFtRTRm0S2mc2oyr0CZoNM/tvLgUug6+wx
hcodGnu5c7SwD4me+/CBPtgyBFAh0WUB3N0FB2976PjX/lTfeNWW/VbzEkHLVxSs
IkoBILuu9vmLsE6JgjCUO2JzzJg8JPv/8UEBAUW7EUgK/KX0EGwAkmxlLIu+ZXxe
iNEhL0AOKLibExI/fqpPcJHM+qzVMLxST8oPocSs/2NtXj4masXbJ6kXNzFZQFaJ
at649ffjHzjsjcsmsFG6zmZwWX3DNeR5VQIClhkWx8ZTI9hzjFwzUQ8UKOSvulmB
NVLv3YTWKvViRXi88lBFuI8QMGN2Kgu8IdzlRYRU9NcVkBXEONyhndR+0J4dza+9
5qgOQKXvibYrixLGvZnpOe+rZMowejI78fGPXbL4LGD1gnqfmapPmBXbnOCuVG9Z
NgM6CeO3d+rF+X7M+evZUDjHS7U+z5lEWc9tq+LHJYhFUgQs9t0Ix0iS0uPXkEUm
HJ1L1fn38lR8m+cescfrKirhJ1ucJFJFGD1ZFCo5DYn93/KvyJgXW+4chB2iSSab
0HbK4k9Fr1RzCo55jeJ0CGYBYHwAdLz/D3xozpC47WHqOWMtZPNvVHT817whDk5C
7KNS/zBk3xxnirmJ8Nb1X/mOyHhozFud3CBpQXrQrJuzcluJtsgJ1JTYZ4UR2ab4
gpBTjB4MH+0YtzeTsjtjL+ejngN8hkPJXilLvz3D82Gk33uPCqTUo8iZH/XCX1Cf
ZLiSsgegMWbUYbQStG4+8I/5b0o9ubuPOJMELQOQfXY0YnZpKpq0thn7YAn5ZOTh
yhiXT99PZUTPXldLCoBO3VmdE5REtZh9I9ZEnKZ3ZBADwWCRI6M0c20tDTNJeiNN
jvFQUh7FJDwPoHj12Cw+/1Rq+em6pb2G6RfWp29zVs8LUMg/+RI19SXbstblt0rx
p9vlJhuxx63pS7qqxUvaF/7jlZaq24l4iy8SjYJ66sGPc7uz/eKb+j/fp8gwq2tD
PiOj4E6uFrfpQL0OljMJ2UL4czhpK1/Yu0NGDYXfuQP7VR6MldLbXreYIbKqx4va
YPqwzhCClwWpNqkDeb0YGKuSCyTgoViSQM7Q9ySOsTgKKLeIjPIbf+kUV+I1HBsX
fpMzPf6trKIkrCll84LesaNgIoJ2QPt7QziHe/wkkggwBN5yXYfUkmyuS3fl2/BY
AJMhbUbI1QbLNr4S1rpUoUHzc+S1wQOw+ajEn9pLyEGJ3YYEpg5Xkgd9tTaIPYXt
L7z/LB7T74EbMlSeyGCqk57qWLu5MfrcfJGMVOZq0HZ38NhK3ZPXr5MbLM1R//9Q
ykPMMnjhoIZyg0lrO4WHXr3GfmPbA1zgGv/gnbVRNRPiubf6bgn3NK1cwzZHqhBr
vjbYYdNaP5GR4IOAevY8XQ3bA0kTe0gIVYURHoPgJp/BUCgDVtmbCn/LProOqYGo
+QlXZ7bP7ayXwevkGr/8dpxe3KzLJ/ZQCo+OFMIR05YCYaCvJKAg3iSTt+etJNv6
7cUxY5XvR6VY/T7lAl75bET9vx+NiFiXwr5EcRLx8guh+1vWADRVe6Q6NpffVVUH
jRqeKCGkl1/Sn5PWKmVF5FqADpf/k22O+G0sh6S7SOOUBH/u4FUQSiuQbSsG5MkN
ssuUjcMYLu8Ee5DtzyPOeAqYuQrilQysHJaPnJZXHhucqE1tbXmS5uYsAVkXS7uI
VSEaqto+6fTY9Iy+Eg3lPDrFhSNnlDXzmhbTHZILjdjVEFv0gFcfUh6c/LI+371t
mwqQ0zR2pU66CR8g29pp1XKqH6Z/7NZVBZzh7DLPBElzXDQDI0LyLlWyfRlA80WX
Xav0/zyb0aJQduU8NOo+vrTgbQqTGIGoXi5uKKu1qcncNBEZxPs57fmk+ekEgowV
ceIrnTLYbHXGs47L3I3epeDYZsETxuKDQVG6KoC9aM0ykrdBqq9+8D7u52vodC9o
qQ4dhH/uV/YmHxoxcbLuuh4P88pLxWqljkvXc9ii749hK6i8a/Nv4Vr8lD+jFKnn
Q1qWJI3jfsriqXtVaOy3Ff9ItrYhQtvYXhYZ6B5VjjDJwJgqclFMgmSJJsXeWuQl
HsIQuSSFgQqaR6RC1+h0f42f1Oha5ffDQhaQvh+eeo1dzV4c1wPNQwudIVw8bM/E
M2wCOijP3NL6PsPQpmsjBZriHjRF4fSQVrxDdOiNMkNNikSdpyjVbq8bVW7/6Z/G
PPNas4uip93xwwVRvZP+Oh+aRhFR7ldBaaWMYPCdLBc70aURWl1hfH+xkQHGObc7
+c0VAEK/cXlKjdjLqVMPIQ==
`protect END_PROTECTED
