`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Grf4lGNRRx1s6Pbb9SVn8ODokQFQ/2//GoFl1QU9FXQFU13gHp9We1mpXrkOgnF
8nMHZsfUllcSFbHuigokoALtYB8xXSXVMnZu1OVeVf5uzptPTVdinPc9p0KXyDJI
jwDqxfgxdLCreuOJSPlpAgXUESy5RTWHhLebxE3Q1pmvfxNPpAi2CKzja7BKkdj1
4s6Vnb7obAmoKsgtzR1xqVcim3JnQDiNpxCQtweiEzvC+T2DPsOiBJ0TlfKK1zTb
5PZ29ZyRezb29iD6Aa1iI6Jogetz+YYN0gtaBl9kVrRiKkedk3I2uiwBFpQk11CJ
W82VleBFfhTfWlJDj0SI+Qr5yeub5g0Gm56YMIuj/TAHO8JDkVdoXKP26XZ/u+7f
tAqZreuH8DbRl16ms9nLgTEM7ooJTNDdz4UiC75AdGwcFRSwoLtDS9v150Zowz/M
fUMNatvB7QIX5s9Uf+kE+BOQILLnzo9CV9HQ1orJ654JlT6XF4WsuYTn6aiAN6w2
bx4W5jPqVhfI8ldTE9SHm/4QrwCgnsB1UkoCF6iCMhkKuJrW+BIrJCkMIPFdQLB3
D+rLBqk7VyKnmBzqlK6s+B+T9wYGwAm0N4V99wTOWYUutcJ8qvKyby71jZ1vWQcT
LzPZmE065P5zxJHOz+HBMN1j3LQnklIcPbPU1bZi63jY3QFtssXlN7E2W3sKywzY
vWabePWiQfe0LCng9zpwakgENsslyUzR5rjNjETAAVFBaq8szbrYNjkYn3iapmUA
VVSIR8ePQ0wqX7rNSKixojWYpI7MvBhczKwQCyEfWi6R0fUuikZJ7S9MMScUEfGo
Sr9bqKUZokGWOK39Hu4vdO7wPyg30AG5X9AomqVAFdXBbrjpefBM8niL++S/ujBe
yMlLkBZLfGVP1hzfdb7h4SlGejtZX8kmnp8WeLs1/NwWwqffXMT3yKlz76Brx1HS
OCqIB97kdJqAhw6H7xsYOO2OBAooblwpJCINxeTMelJlcfztyVVqPzWkmapOYiQ4
uXQPgX/5WjmOQPCvPVFPTRimbxwc/n2pAme1MLqwVoxyHHFlay53G4xM3zfzmyjc
DR22DqgwYio5577mDGSlk0d43Hb+If0EDpcIt5pMBIIaM1tWx8KL0rfVpv4qn3RM
TJq6qOtvwd1r1C3YlqsC/XBHkfQZqC+KHkexYU++Hch5QtrgGu9etGjUf8UjLI0z
Yfg6wBhrDeX6tV1GtLjrenk3tARyotPUXOjgvSvxO0Tkqo1wF3K4SzbCOgZX+IXI
tnfZqvYZT/NuNMZrz2VVQVsLZbU8y9hiuNkSpqCkX5RUeu61dW6oIevGK1KIm+tL
zYJtgST/kHQ7nQJhcXyD7COMWLNixcBLPa/a8A92cF3yBxzAg+5zNN5WPzdxYINj
NPFIO2T3C1W6S5ocnNuTM8fZFaZvxcZQbEJAeg3XvIKciX7IJMjizROciXpG1wM/
sO9gBNM/O5Rg+JLKsBQtE/8tgW2DuQE6zwQ+C4HPWuSMHNTrS+0s1LXc8LI7nW8v
qEIzhnE1HJfgI9Ww9GTxxDIHwphz96DvUEBV623QlKynlbo1d4DOvFo0MhG9si3o
7y1CxDjmGvOoRx9UsOv9slRYHwfm3R/+24zzQKH8hx7xgu5P8Afh6UfA/pNDhU81
bbgzU7UNbGunZA+WgJMA58RpSpVHyLpJjDCh/s9cpfhSrwwHvgNLpM8zrqD8R/OG
cJkUAN5MGy5Oc4bRHwEartfvJ8avFUHRKpAOFewIxP/s7adMILa4IECeXR0dyb5q
0wgiAMqGBiwCDgrJ3NvQN089M+MUWZ574tluxYHsB181evVmKc51y7nEx63Vwzmx
mik35woGWLiLCD+LIYIYyiSRnjJeOsEbP5z/o+x0vIuWrdkUB6BiYy1MEteeEy/Z
hfzTIfpjAdWaum3pqSMbJm3EArA01XEW7qk+zOyg0qikIsWLgFlrWVU2DI/720Bp
GooMQyrSDZikCvYSXsFn+HtN0uw4S2TlMU+XF6B7z5PpCvQVQxlSp0jK4dfJZl6h
WPH/VXKCx9cdVy5WllB2TW+dSvqyTFke02pG8vjo/fynFTuGkDz0mZiMzbQvszzy
bWrwvsKdc2xYrxdh7Al0ZA==
`protect END_PROTECTED
