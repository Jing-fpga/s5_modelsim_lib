`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gcVrF3KF2cZbhFxb4w+M+59Px8yLyUwTUYx9g/W3Fe2GuF+Fncs6WXG0abOnpGRL
49WirJoE37NF0NvPN6LuZv+YZxa9vuPJGMbx7v/+HvgHTcfphuw2cmH4oivzJigD
IXEcvsL07WCCjGtZHjhgRrTWpz6yKm8CUqC7DOKoBvjN64nZ7E7/sM6hTCTpZeYX
fI5pitNkUolEVACkq3c636e+mFiyW/Qdz4nQm5bvpRM0cuhzkaZkpVlm+wiCvolY
SXzbBB05WchOEuddJnNxNSZud2GC+rEf/ueYqgvQ52z2QgJM4xU7sx5s4zPLJTX+
cy7fkvTI4kabEASOjFMXGdhxhYYYOugl43qE3AdR5lG5rrM0Bpzt+Ngg+zZtCAdt
2kLyB9HbB5qGrTi4w52MCCeFAnEytvXnr713MMFrZuwQ3bhN3+UFz0TEhvEUftGc
W/9KBm+O2ihvnBqm8vt64Ww2rBNowhLwXh3DsPs+edLozk7iS7WQpoHzUapzE7DO
ujHfJ2Z/4KQi4yBwiFc6eOSlSsc/i9beXhq9bkFKV/8SJNFrP+06bGuTUCSTRr3V
h/SMIl1h8BbVsJibLTVXmKdlB7AfbldMoXi/8IIUey+ZFiPzGyGPvAzVCPu/rEjU
87rlyTMI09exWx9KkwG4zjcmSSDIulUllDzqev9YG/NnOMyXM2ixpu6DFAK1JIM5
Jy7j0QhLOOg3fxR26po+XirIvRiFLckA9qDJOZ8KFe+9NmaOh/Cr1ICjexXrBgY7
kRlNUUwxNLj06nc8wq2EUTR1n+T1IktkE2GdM3rI6SIR/b9p5t/ghppwFfd6A6Sd
LYLE+SgZRc8juOsUntoVNjvvV4qeuvN++cUL9nMNViM9cRdEFbjgC9s93Io/pXa9
LV/df5AIoOa5gBWFrq2NFSq9xo8HauJi5648QvAhM1GeHbPAQl3rT3YePyy4ulWt
tsH7xsEMED8AYv1YUohdGEwWdnNZwvyE60OGfV4az+RgoKC9Ky1jMk/EFQ+K5dRV
2Z11j5h6GzKPgZaPuCShS/Nty+hf8PXLW+t9IXhTugmWylNih3mgLGakj0hSVh6A
/ShNSpIrNuqgAMjsmqbNI91KAIDZNxNx5cAeF90tSxZIo9/eHg/xFJnXrxEvY4y1
CWxFslJHqGck17uPMrpwRWymVQ3H2RGslmyObnzh1IzTZfGj+hMZTaiZYOe2nyCW
1fod7U8xsmwdGk0c/oU8HNsV4VJtImSV+belWorf93iWsjzfYxfivyCASDfRqk7z
5tvErcXnCjBgigZA/pHFR/I5Eyo5pu1q+aBYwihrhYoeU4MSEEZ+WgceagSxqS48
1op1tDRTBd/ahAR7Kt2xF+uhyuyppLCYiobBAE/NkZ8oZH7d0MNrOajhhqChi5mK
XKt7n4LtB8bEeXxOBRs/H6bXiUwGANYOmPnYa8esD9WCvWq6QLWN/yaDMQcK9wev
D0iAu4AccEAX7nDRujl/Jrid6SifSkQhhP/aUXugeYfH5n4ehmMOLtc+8hGfM06L
tGdLLWaHKQ2zGvc5+LjW3XThjvUL/Pjo/QsVV8lAgBba74c5ySLYodzfEKpIW2hP
TEXVFVe0n1MtO5OnZqfSDOSee2D+GmkGHhvfHA34lV+g2SahSr66SLEZebOfYR8/
+UynPQolj4vJSD+921PT0PXy3wuL4aQ0E2BojKmOM4tWjFUSuUKbZr2LcuDLG3S5
qYbc1zKVXGPKHIpBe3rJc5KGEZpf09cHOfc4YgGiVWd3D/NlsIt69RuDbk7hez7d
I2LzVs7SgzyR0QebzdX0Pi/gF3nMbRAC74PcHsoSm2QKF6OBT5RbCOO44v9e9pjB
zHHKKAFYEz9aDHrKDOnlimttbXtF6AE+AmxvJtnbnlcpee+q2RZDkkY5PgQjqDJ2
HrwMzqMSz3lQ3goddIhl36KRmMZAY/5Ri0Ni2klaZp+DjRA82THPR4nP3gc0Mh3v
sHViiTi9UmuWv2Iu1q6DMbqPi1kYjsU5ZtIBlg5yyp8XEBUIZMjOS6dyXN7+4YWT
4mPAuCfx+Nlhn/sDPaNxGTyyHxu8Ee5Qpd4LU7Mes6jjlSv6k8GtwnN1cqyil7hA
CWcUI/EWzAsANqbP7F91wu52Fm/UPcRCYlSEnj1h6rtTS0E817hWaAW/JI5g6zvM
cIZmHdV2jGqViUvjQk2tiyziqClwi170jfsBvE3hjOxXEZrJEEJtfoLHFTfin246
2QCkN3jbcBermDS+cm6gKf4dSLFnP18TnsYRAdOBlzH2LLQcixdL5yHctNfgXUB+
EpzcdVXREiFcEXlg4CMc0iN9vORnMMbm2p+pgXqGd4PS1EZodY7WVif0y30EWQBS
cZ+UFfAYTvFwvCX27V94mEmyt+xZP35qIyXlQp854rI=
`protect END_PROTECTED
