`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tTmenmztpoI8ZJ3+K63aiJM9vjNsAY8n7W/vHLPeCz4iLqCJSX2j6olSc0kMEKTh
hTveOvFOfx75oQHO6CnbOB2TsC/3yYmrDUGcM5GquoXNMLlSt5dgl9HoZksLCIw1
per/xDGCv/oiYaKNgVOjTbl3lzLVUN8i5s8M3Pp4bez8JoAPoSqOcJocgboCZTP0
m5P9NN/sfNBJu764f76QZ8an9z22PO/5FWB7tbS5I1zzgcwvdD8tRlyFomro3EPX
yPn61AoQKLuai9dm1WEN5zd8LNLAJiHnNA1bar3l5wunLijCrZxQfem0WUGpqDh+
RRvmE9aXHKhMC4ZoB0iwYDlEAKFX8Wy3Q0Q4ek/cRU+FGpmOK+Ae1uI84YAt/t0Q
/jCks6OK6vps9A5vEt0Erdj+BKh7M9fM5iKAKR+sXAPZaa9D8vvw4PSIzKzDmYNs
dlfhEvwYC1Xhu83GJ9yypxMj87c8e/y75PcU0fLDlUvm1+TWTqup8bdQwlEm+vuf
KVnBOQW+yTsiv6rUHCxtOaaaH6H2LOBZJHMfayhUxkGO3aG1K7EE2hvAnCMtD7ef
OiQipiRYrnEUDUdUVQfKNTKoAV3bvrRFJF0klDWacAw=
`protect END_PROTECTED
