`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h2Q/Os/nt/7nB/npsVGJ/feAb2qzJDcfeSMq02RKCa5R05gPLeTJ1U6JaGARpKvz
S/VrTB9iVa7OlhEtK2VLmR94KbPxzV1HrpPgZYKl+D3Iz426Z8xVuFstH1j/KkAs
fYBGOAcx/ZQ3klarzED7Sw7tpOjGYTdANbxigtvLZgdhm34pv+bEB+lxidPU3YXy
EiCFbObGRYJVxXvEnWHPfPCSjoglnGG7XNTveAMyDaOkmkHZI4d3QHaWqZ03F46N
SF8d8o4/X5XzUIyKd4cAi4nGnD1AeJLqkk5hHmkPPh940KRzQxoKxmS/IzV2banb
YqQIKYV0XrgbG7afHV01D9RdppWNGNZu6O1hQ0mr/jDrNDCZ1pmZzVFZd0/PBJuZ
JIQ0V10tpwYHBlgh44rgESL7Y5H0Q/3hIJWjAFKYedIncUNIvB3Rm6x8r2ooT1WD
VuJg+7D5+7SDEx0ucqFfYZcyLohnoQ/Ru/9TZLMmB3r6b80xT+vAEhyJxKrrLPnZ
lMMlwEOsP9kQ72nlmEVGG2e3VF5vZrdIjx1anCDZRVktDRzZAHCdH9x7l1PpnHpP
KeJ6Y1n/Fq145GUK2Zo5ZUTcQLG9KEhuWPTq9r3gSYElsZ/PTiV2XLDU/y3u26t6
IcBzvUvbk7tp4ZpJ1DM7Cjq4A0OF5ZfsbJcM0dx/pBIhcPq5bwJzlOMFaEroKccO
xA89e/JjEJLfInaYu99iRXUBvcHuLrMtUyUvgnP8Te4HC2SccM0r2LVCYH5aJf2C
QkoIG1cBsbCFJjFDzxrOaVdrjKdf2BaXiNE1HW88N94F2o2X8NX8X8GWZl9UliJQ
dzFirnuUn5g51Fq5ixGPe0fnyNZJ65u1iGAOrP51X/6uO4Vg1u05R1B75sNRUS3N
Gxp5hg9k8YUDJq8Ve3WN5XDlNNHTuo2dY6tzbG8ZG41ASU0cJiKtFcA5dkTvetec
8wFXBoCJNSC9HDDg9M1ViJDtwNFMev5xlwbkUY5MCuy4m5cWnObOI4BP8ddzPWJF
x1LWVz/oVy0i7jikjEnEjV/d08blXvRUw9SOUWgFRag=
`protect END_PROTECTED
