`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x5tRa0ktWjZSNTY1AtwW9u1XsJKoy/09grNHbiaGKKgHj04Cmwv2/FHno+OZPcaZ
aDR194bQwd4hmqObty542CWGQTVx8I1uVZggl6WNFGYBod2hT8+suKJldY2cs+yf
M5kEx90fOTOT//i1qrIX3gQQT3AlJlB0yYN1GFr2jaWEpqXKZxQMWA7CMbRA3n7M
uHMXlUqkoDg+J2vlDCqz4Fla2ZKHeyEFqMSm0v1YdpOk41u/VHQZul9a6WGqs5Uw
lYI0joxyzlvsYhAMT6TJPqoXkXUqwQQjbSKnBK4EXlwPBMWKY1YWK4GNIeyVnL7S
mSU2jtI9m140vzhcoKgAy0wsARMVTdz2cy8umL+BLVB/zSs+Kh2+/ICCF5Uw17CZ
0bihgQJVfHga8Rn7jbuq31Zc+3WQcXOjJBixitVR7nORi67xV3PPpdu05LuSCpyW
8j3cZrsgVWSoFAc8jtPfCZFrjpzgIoOorBEj49EGJiAeuoVlxHpduz9IEYGt33hZ
j+cFJaVQKkd/PObjOpU3l44ZmMxY2tmOs07/Tb0TI5412M0oenix4jroZ+x07Ghr
d39x2b3CWEHuJJ6bWr7/Ix3E6v46ZT2ltA8c0g+3NsZzKMCXH4Ot9LRaeFgy4S2P
hJQZ454voDQW4Nb2C3A0kGzPDfVl5FXiLpLDeXAvf0HNo2GhqEFgsW7Qp+2jtxMr
ihEpN4t9CHB3niyPIfLef/rrbJiEAtygglAMRAEEkaqvTo4akmT5oFqOQ98yQI+v
qOhDNSXO1YpuCiagB0n2RUesOGSS5tP0bz0ujiZm3TecuYLRpl25TCKofzIE37ee
rGqQuw+DyzmZGG+A3EOk9dOUhdEXD6/JLvPiSpdLwG1FjdpduhkUcy7lwrKvBPzB
19bt3dnD27xwXnLxwIVH0fq7Fw45HOjjaLizDay0PwdlA44GoR7MTQRk8xrqFgPM
tUBhzx6EHIbgKhdOwRaGeKcFJkNakO0qsK61DOXZa8NiBRNC/4pzSA6/K5xtLsPQ
piLdl/VNXf7AHp0Ueh5TkRhOJlWfBnOEW6itunrOOwDN2NW31kupWPXbno9eFECB
nbPdjCVedPdEHy/93+7BvoDVzRMWP7CILYbdym+8UptpwAb762P+ZvL6chCKJ0ZJ
xBQWb9qxPTJ6Tf3eeSS905RwKhtDr3Rk0efS2teZZOfF33kEDpFnQsQeZHxdYBoh
XBQMEYZgtaVgzIAm+13QpTgUc1rPTapE1RgOOOE7g4p7m45CFtVE+Eul9W17A/fg
`protect END_PROTECTED
