`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q4hKpgv+tAA2w2ZK/zDbmKtcG+QHnu3c1ZTpwGtfw123naF/eRZY4Kg9alzbNIZw
Q5PVpJgfzcLON07MMLBEbVU3n1OTS8p+4x5n/wCByz5fq5mihdDWWzP81Ri+YN9D
YIzQ8Q5Vfvab38UHNpij7YFYWIyqtsMhVfgbtQi2bZ52xTfDvL/kAUW2npBeyVJY
mNh9au8M7NWjbgZcuiFuEv48amEeD/zSoNd8B5HTYqpUE2zcOd9kKRxGyS6mR1YP
MSGK8b96BWGpsCIx4dZqKcyxRUgclDBCyCH7EwPSx7V9N4ydlll/82BGEpcHqvD6
BMH1bI/AbXe0C7NZBoHaQneZf7v4WT5C6WpfeqtGgqeLB+MFOsjD7YC6UjFXn/6f
xCgPPLgfbH9j5x67oUvcL/OkYRnesH4Uq9nllX/krnc25LkPNe+74IQRRlJpFb+A
0fRsAc4OxjoN2iiiZTKpxg7ycDL0G6wEM56XFd5HOPi4avs+Z18y7N2oTIa3Iq2Q
yXpq/uHRVBC54MYy0uuDYWoj+6FXmgBX/8z9AmgiWlnhLuOnaXiBqzoovAEmHtRq
8dO7DzT0mHVUiyeD7wOWCFwtpfnFYI3RrwHKamOjR9z7nL7zVnRM+/6DD/26fk1D
L6rMC1gzNWfQlwoU2Db0xGWdbBoYb1BJuYKm3cKZCjM0r4NAbSE+0LGv4WS4pQsW
AU6889lhSPBH3r7DehKnukoTGBT74c/OmLCpLDKCb9rifJmWpiWDwJohVIRZjVeR
thdX1GitnjtZj4hmQwnOZz2EvZ4emGBUFVZSSdqC1IBTYWZ/jUmybX2ibFsWCgmX
DF8Lv1NKSTyVs0INqzNd27f3GPm98+osn/bAtfWSPLVZWOgJERZvmdihAn1WB/2w
ryzbbc0JciMWEa8r5o2yzfN9qo6rzFmP1YJyzkwbCJ/NiKgF/OHaG6PdDPuX6eN7
iAwNFq6+weJaigYOkS0kxR1cYhmujj93D1I7eHQub6BymteWU5Fky38arshBOsVL
vamwbh4+OW75G72wMr4DHuHZ8lLNG9CrKxk0ThlXF0uOWUik/y/qAPd6KDnfs/5u
Px5vaBwfoL2TvPqMLCQK+NkKSs0dxLkgxIhlPS0W0W7xHlInoKOA1l6sePXTv3Ey
ViK9yb8sa1nl+piIb6MiG2q3hXcUv1mmalHiVeipR5dW08AWZhz2+vV1Qqs0dZHU
7oxNtLVqHAGfG4G5nufcLTKkaWMV7rOf8n0aGUFTqFcYgKZqGiXQtvZq/EbSozci
1gSzEZizoaxNmGPCtHG9u/gMNHynn7JwxXQTTRHAwl/6X335UYvEMvKRLu2hg4uH
/MGMj41UVwK/VeoOsFz/2tswRhA+vesHRusQwEmc7Ezvwd7AK4e0tDWtnnCsktRy
d+IBkbz08fN5318g/989fE9KUH4fTsIZM5Pr8dUwYVsMHLFzSLwdmEDTWXtuRr2o
+O2o0Q/3SfL2GCA7r115EiG/fn+tLANWz3At04KJlZm3pRgPZm/MaSBxUz+X3yrg
6ZMOqB4zv7F41/PHeRLfYNF9ETAE4yer4582LdWLfVbMcFwF7LH4rd8Ks3wt3b8p
XIO35f80+lclxO0YA93yyHuweQJj+5hR32xZ+MGE7L4TBwUFVvTM9vxhIsPeEwOg
o0HrMxMWu7ujbpLEvaSpeAqgHgDpcfddkvtDK4lRAWPLGAL3amyVS8PLYW6HT7sy
zItviuU2ht92UC8kCvwEEW09T4V1hklYNroRNFoiQZ7/WkeJ9WsaNyDce6q3F0ht
l0pt7u+toetBy9/eydxkVWz7Y3UyGyrVugPQpNZolq6tG3vDvYnub4zD+rcqUTAM
1lGXMzU9MEkgkpdpgLrqw3zKDBZIzXjQ0yBNS8vo6wCqEJSn+wv8pi7MwWTF9gU0
hZcytGWURVTBND2x7uTUhTw9X+5WAt7Jcx28//r5ZxIaG/nxPMl5WEJQmHmPxxGA
Iw4bNBRJBZMae4qnhnbbAaZh45dLs883hY7umgVPilr8w0RUH/H+LQw+HKCdMUgP
SLCAWbIohhBgyAHSZqddrOgjuzVbKr8cDhkWWWurB+MXb8xGXAzFrB06yb1eE8Fm
`protect END_PROTECTED
