`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/JjWNrdOArgjCxKW/W7KkIgh/5zBOUze/FDCWbiVSRfWcfoJXzZbz8TfIYumSiOK
856kxe/eKfrqlN6KnvLC9RAv2xlFYxs0/dQ0EjCTdbEjREyslWrRSKiKv6Tz8DBd
YB609phK+JqatWNTpqfh9DiedPLoktMc12YqWdSheK+B8FlwppRQrbwybseK5MDE
/69xA3T/cqvG07hWgJPB3B/B0ed5vU5fdIk7exH5wgOdn0Am1SUIbSxnGoK32JeC
GydAuPgkCrSGwbdsjd0I3Xh+DiLciVMGH+sz/i+y06gzJ7QRtZg19t9OlPUYKQgt
ytpZz7T4EI0Tmh/bN1z9fA1ycgfEJ7Ic8yserriNn/hp20EjWU3x60jBu+e03RCi
aBzluSSbd1FTazuhHTfGzRzaoWOlTq+4xA4gfReEb7mzDQF2DnLje7gNCel7Mh/A
k4f6IfH5VHUj7NDUxCKUalc1ltFqT+MGN6q7vWzFnda46KEQe+d+pStpKxSELEkr
7tmiOcI34VebOobxw3fTgN6HDeJReiI3e95SQah3HPvMq3y9cOhJJ+cCkZrjuk8N
GJoArHdJSqVfFss5mhdNHKj9mwYTRmL2rF+7zxca6h14NwjzXJydFvagaQRuQclT
`protect END_PROTECTED
