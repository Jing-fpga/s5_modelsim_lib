`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Seu2X0W+u7BIHEbG6n/OQ9WNFT6dzK9NqVbtTGjmm+bCS9eyu9Q5yoQUzOqLwe0w
9TLWiAxKcP9/Ej40cgBTI78BAa25Faq/wBDzboPAOzXIBpyINLt4KTF1bt6Ixa4V
xhaOfbBuKHlB3E8udYPm2y7G1Y0VdJJms/wfAgfV58Gf4/OfmG04tg7OnrxJ898+
KPS7rb+9+grBPhdLL8rMiddnJUZSXL9AJ4CDfcAmVqEhB2uqx5IM3r7Le0hLMMcO
VL7WKYQNh81rnUabRfOVb/Q/nOEh69Iw23yH9YEoetNVFfIHk+fOks9pYyGRpRZr
rpGTrFxB+ijiIrDzCXKCKu0KQIGC3quIjZSYyNMYe9j+N+70Dm68xltDRAXaU0zt
cjWPFjaMTkXutwvqJUQv2K3KGVNqdNqOgd6wgCmClCxi1fc7S+tSjCTUn1hrB0Eo
4oms5p+qlSawEVEkIHcUnMFvcBghcxTaFHYFamn6DyVS6k7MDhfKoZzpJlWDAN2a
NTF2caAI4MGyo3PicD4d2/yGwhED5PD7+v8WaeYoAqGipCilnTfST9nSXYKbzQoB
mjrFoX/fZlW6kBuzkj4n+uXxKeAYW6YXIbdV/ViPHz/UoGrqxkUmp/MYMEwS5NvI
46NgQeMC9sXfYXCmxDwrXlaRgF36fK4Kr10+vXPwXAtwrqH2fO5IsEpDMq40daDu
sO6OIKFx5AsJc1Y3zUTakadf/dnpKcKJEHE4/oC+k3Bj6Gh/ASHB45w6DRid8W6h
9rAVD9gPJtZp4oWPs0syxQYnCwc6+dgylKGjJkpefxNa2hJ4zml2IDJdLIlNcxVP
xaanfr2lhPZ1ZFvNm3Z4Q/t+SD1xrd7z9h7n1589PZpAyuM0lf136/BRZO0CDKnX
SFquT/H6LkEnqyveoxg+a1ToV+SSfgQSaR9nnHHmNyx3ExqH33VzjHsEWsBjudzM
QClPOBXyTYiEoBEgwdz9WiTfequcp6DC9EV4nXa5oq909GBTsHCOsmMnk49/UHeR
ZFXDqgjp7S6hOKYjtMmvdA7KRC0Yy3r38Fn0iWoaP0mAYBxHvFzKAhYNGQxvYw3A
+UsMKTMfUciP9tSDNmhnDnSUXbzT+7SE9axesAnStDkBNvwlmO1P3OuG6E37ri/9
m6BkulBH/ICggRhAO88aGztZBC1CMQufFqlmV2XimOHj9y8nWL1sYHofev7dawO6
ZrWDOX3cfYBcCx5uzuvIK9bpwu0hm97qUq5jEbp/rH76BYUDUWZaMgGQQKReI2p8
5Lv9HJckpnc//+/FXF0zE2gCURxVlQRLUCrsakg+/340EbNM+huVuZ3im1qVhtoL
vz8+XUeoEwP4+YAjkMYxWlvT0zlhtYOjcrK+NjODqL8Rgz+KJr8qzvdF26qMNmzF
jr7h7yRBI8kZA6OgEckAMdjZBPyTPFqsOCFZAFHcPp0vbjpk1XERswKif2ffRSCZ
XInzbcA+IBBITZe82r31UTW19xrjaXHHH8v3CI5qboWv85yUqMDje6uCvx8BKeXJ
S3kt6E7zLHObH9pB0L/uRbNeaeECuRB3MFjzNzRKDBvmD+77DDuIh92reQIrDN+Y
jglYsbiTINoiSkC54ag1QjAo/knSp2uld9orcC82jKnc9KB/9YrK5f8JwQor6sbn
r0EqR1axZ678ukSjJrhFtpoALKQT/k/cqQOd+X39hMfBlb8u2rf0csYRC2mDW6Ma
d3Iy5MKazo0xGm9iee+5OCQ9oN/NjaIOVcV+9x3hubmVRB6H1FO13l5Pc/XF9vm4
H8ts6KN+AqffkWdThmwOuiD8E7EvcWObBxHvOLekyOyOUjGdn2h0ueoT9QLXQGuE
2e2WzgMC401mrTF8u7NOqDvGSnhPTewCAwgQCzsPZhL3Dlmv8i3Dlre+07Bd6wEd
DvQNuPz9CWpySZiHwQClbBTHLG0nvqr4DY3kKbfgOibBSYcA6W8szHFdGIKK9MdB
wBSYtiruAJGm5I1e8nMmtgoJ06alv37ymDCyyUwGFn82PVpiDEUGTPJuua/CTq16
zydkOy2z1DnBF/MjD987m/0bvkw/ql2iMhTH4dJ1EcaMTn9nql+dvcJ+8pdG2UkQ
eNZXK0sB9c3DO9gFI6XtMf3J++1uUgs3p06tE7QaKqIZL4P/oI9RaONTedzdlGgc
`protect END_PROTECTED
