`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VzKz3oIvi+pQtU5IkH0MXg4Z112+ngksArXxxj0awibyBeYCB6ZSencr7hVgdDS6
1L8o22+RO41bOvH9P8z9l/Yn+UhPWLrNE2o9Obiy9mdykYAK3xvsNEfs7/F1h9en
3QtX1haEXiinfEgcMgig1qV8i4+/o0hqwO4ZneskEQlGFyRSP9fSAX5mQpl2a2NO
OpP57Euo/RdXSEItJ9jtegcjrNeWjCphALjJhXkEE7WeSpBpWg2V8e7G+E+w7ogt
btsVTuo9WQNMnrx0Rtv/szFnXv3OABk+mCh/isZVxorgNB2c/ptM6mu2qqLiqkjq
Kz4cn6TLA1MGLR15iqQeDSBTqoVgUViunVW+ny/vWjaBw7WS/Qy21DBz+OfVTwUd
bLGseFvNsaWDH3+/U588PzmiiafzdjL6tz90u3mcKDwvVozOZn0hO4FQivVoHJja
gUYmjpSAznGPGC2i7P1wxSlHx8dBH6dllm4QAbhwjuhYm6rqfZF1lvBn4EMXQCor
5NFC/HkhY4P2oIfyrtC0bAT+eYJnXh7vsZ/rawt4Wolka9iDKoNZfPdakNIlyn+f
Obs/lin4eB/dgCSY1eI5a3MR57hpILay13DM6EWl/KA=
`protect END_PROTECTED
