`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cXGFClvJPSHitD5l7iW1NKRo6GfUJcraxeTgj1vSgKDFCzA4QFzEKbF8MYEP4Vsf
G5dVv/ulIhtKngxKUUKMR0q5Sg/LMQGvPUp6gSmLVshJFuyjogjx1Kis9FQfyotG
8hA6p8ayg/5hQRue+MlVzMRKGd+iBD++0JJRH390nDRfkJKFinCz+EEDaZbslBYF
3FMjdKME5mrAzR3dQSwlEH/+i2WyMywlbwuUxF6hdfLoYMkFnga9Xps+8pOTJR/Q
Qh0uzW+a50DzPz9VbXlyikAghzMD/izKnnOoH9uS1TgZPIBktqBcOlhUuvgQqij3
PWBsrfBh67N6wjwLDH3GyPM6nRuCyun8OSpggXlrFEIt0F7rTM3w3VHz1j/JLdo0
F6lj/BztzEkENseNOrSXbaYv7yziRHCGgU/cYY16a1qdCRM335EL0jFNTy2qmv+2
vxQqkNishwDSmmtBwq8EcnbbLLmeffVYwuXi0YJI6Ig3HFj/9gaDFZHAekBiHhir
TS3nIZ0oLSCvRUReNMuOdfr8NvRiNq+Cno5nLxky4R55AAmSzB2sLdaqIt111Fla
AZI2w3HbF2ootCPgjV9XzuDJouxrZBwBHwlwuLmDfMRW/ZoUwPYTA3GFYJPKf42E
`protect END_PROTECTED
