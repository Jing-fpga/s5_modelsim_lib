`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
24XKisY1lT/vLaTtlS0x4f6SjeLu9DO+ElMkpH3REOO/GvWzK4NUD/+pGkbO1F1B
75ibGpng53HIV7kwSRLfGaPtG0q+UwXChbCqHxVghohqyZ0XmkkV34lML8ZCpE1r
1Y/sTuaHkcQRm/RDnPHc3w/aCmNpPK87Bj9PALEksx6sfxf/6/lZogh+ds1iFhfI
8aoVQLI8XU1G+A0sYwLm2ZRObuRqkY4uBA8Yh5ySxOW7yYegk2NmG/+633g7kFN+
f0rbNwA0EgVU6MiA9+hNAIiSbR/R/tmIDhKJbBiaBFSyveuaLtJLS+TNm/bZqJ9A
IDzdeUY8nj7qzfxBUfCNTfMPLPIOKXSrM+z2OaXf0RkiwX76LzCfGikN5nKLpkx/
SetLlCSRpv794AqI0E8xPLy7gXm7jRcOuXZIglKcp+D+0KrkP1o9FI/mec8kQYsz
1tXSDcVHQH1KoBuj+mqsQop1Gf0W1vpDoRJ+4zCl8VOZhqIiA++6OOkL5ptcRzqR
R9ZkP8LVic48v4TBk5YLq9pxH3b10KYhfkFzx1XkKmv/jp/d20qWm2mSx6vwilYf
3iLOPTzvmWKl6NeK6+ejQ0mgEYraB2wC5l3dlwBCWTp4uIgyhqajD5/m5W7z8quf
ttPNSTkvXS40GPKeZUECUg==
`protect END_PROTECTED
