`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SZAzwyObqjqnHSYkUYM15HTscGgZJqPYR6IzlB2XvqVYDpyMxaawlj1c9VKrjtci
MrN5rxTsqCVz8W8uMoB5opcHgAuJlvJUIfjA6dvwo33zd1gsfTYcImwPdyRB/dUn
Cpu74RUgsD7zj45JoHjPoa/1iOvsAA+9yS9NhyDl+v6PSvI2i99tGAtN2cFfZxg6
Uv8ZdLKnqY/QM/xPNMcE3So+zPCp8u8qKpVdbndDgxUGvYXpgmu/DzVKrNyGvCGf
0ftqPyia6Sf7C7CzwKHrdv+yhAZuDb7mnM8DPDX2M9Nx8/GjlCcQBog/jx0b2KIF
HbvEsemW8JYPAhu4nmPIW82F7Bmz7I9A1HX4rrv3jJRlTRNVdue0ojVD7Jl+E/db
NBP05mIsv5lS0F/GHqq/5dCx838KfHhil2ijfrRAp1CLd8PRmaQGhWWPNKTBnAND
j+MD9S9AtYBmIaMNCfUf5p41h3iAIWNq8tr3BESdLJbkCNC42LnJtv75Mrz4gHQL
BFQlnSNJJdOJjqeUMLW+dABM+m6vCccqTcS5GYARqL16pf2KeXECYKx3h4WYq9D6
TxRhidvL7cb+8TpQSTPonBrApyIMwNOANFXufc3Fs5+uhbiJsy1eRy6rxTiW/rxv
HuFOfFXoSRXpt1zF5FAa6XUrCW8OZm7X0RTy6Lbb0AmK7XKGrKMQPrUIHRCrfHBK
kIxj0lxeTkF15SeLhlCAGwvdLApggIc5zBxeIuQwPSXvRda0zk/NEbhvfwwbjyHg
vDe/cefKKFZKx4dAxRvWLIOXCGaFpqlAC7iC33e9Wmps61VCq6eg2tMH6SmqlMLa
WU9bAWUVwsz+/jvqS3bUPpGLTQBdBDgLqeC2atM74urA62Vu2z3dYHBs4KBh5yA1
SqpMNLjSOqP5nKXPlGrWK0UwXRstpZHMKWdp1AUdAceND0F+1BtWQnQMa+wl2QC+
RuOWEMRmO7UzSHdD/I0KyCHSFzl5l/xo4c4YyObrCqBliSBcYMhlqvNB3QSY/ucR
5j2HtjoHUST5POWFygKmRX3KtAx4+vZ7Ryjo3nNyG3lXFKw1p/xIPQhcfNqQrB6m
/WPWzm8ao9G8ZQnWwf31ghxgM8cpFLQ1PLt6BoLRTw7c+XP1AxB36iZ9PeKLaAPz
pFTPMA2l+vz8GOPJFbI+vkohEXaHHkrfMEGEVjXzRgto8NGkwK44+sT3CqIOF8Mz
MZCpULoStu4FNa7renhA1dImI4xtg8LbtyeGyjjzPv1tESoxvZ2RAUCiP+ECkrPJ
xggLkc3K084RmL8gjTFN9ATnqTBxx95c72dVTf3m+FxeWnijipa9QBau58c7v+qw
//JLiWDceQm/vJqh33MSudCyWYFlk6bBXT9i5EfXR1mQPpHyT8fWY4nIexHizygC
9huTfA9aLP4N6xGECJtdNKBDoJIc41B4mzaxLMCMIZufaULMIjY2c5et5xzb/g1S
T7H5yeWqRYve5194Aljib6fYQjC4CG8SUUgp5odOQvIewHcKRHXX+9BvC9I5QTMk
CnM4up8VDb78rsEP21J/+gh7yeHN5A4Jm8y28EYsXrKsmxUZgoe649f5OAvCvbex
buBTrxmO3oI8mOI6twhbQp+69exueEL+U+6uHgBRY7GoN7ZsCKlyHvSs/T8X76Yn
4Nk50Y0GLJxBgRcxp+WsiCoclzvDTjk+mX6I9nvdegfmZzrxKCQj4jXnVwRMEzSB
1rJTfvgKJa+IBaZmtt8yris2gBS3ayxm4Sn2y50jzee+Acab52XBgHi4tw4bxc2Q
4cJCBImQCrpU2eRcE9RRPg==
`protect END_PROTECTED
