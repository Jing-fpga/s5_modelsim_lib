`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zUweKlnmwboaNHOJMsSnqGwOnAaAR9URzD+z4r/h/hE7wvqtF3zX1FbPPR789jVP
n7xwaXky7wth+qaiDCliGIuhmKgn2gPvIQuIGDIFByHgSuj0ITshcFp0D85bsBXw
a7ed9eo/lxTBZ4dyrgZ7AQ1S9hltzriEuMvEULIOyTvrWnnjwAiPXhySO6HIkuCP
XB33ZLZlFv68tnCogR9WrQ2CI26OXXhSrQZi9hx/TtHbLxhtqECbiNcMLKHz8Apq
t+alaCypxgcCKELhhVDtu74MNUmLRNkh/CWj7zjwJgiK72QIQd82NJWUFzDrdoK+
EXR7oy874lTEaDwbdSJUAiHZzU9Xy8ZKdZSgarLYHRst0ZwoNHgtpWgrZRcUIQcW
z++lgieb2YmxdPDocqrIwy72wItXSLVcfYl/wNhHcabivWTdtDi2y4kSCyj4ZsDM
P4Waq9rrcrwaLe4e+6QL+NQugKC6Slw+bqPzJVB70TCMoHZO0vSpU0MORPi5cHCt
pQ3Qe5QHYWJqQiY1iG91SMu399k5z4PZjcxVaVYb7q/4R9kO1CBKAbmk2A1rrw5m
La/cSh1plO+qjcOrcEhrBJutCNi0MYD6KlFyGYZanB5BNf2uSp5gDsFCQ9ncHpum
9jBTT0kTQeQBarcRkNSwfR7s2t59N+Jbm37lO0TH6PzNzDLJvi+ylHo1Jtq8bqLx
SHQRElK2cVeC6jXI2l7QZsy2B84GryZTBkhvH0zpJUsIlSO0pikmWQrXuhg3P9AA
qNV3yVKUFX8dL41F+GLAY9ruSIUAJ17r2vrAWezG4YqkhTLGqjn+9B0qRmTA+BLP
Er4XXTlwDarEAG2bZoGeA+UJo+gj4wSLKd3ainB06NcgUHgTakPuYBvXtNYF4FA/
+WKFxsr5VtPHYAZGR5jiQBaJLWaxuCvgJDuSRj1X4NtysutU84FpQYaYy2bz6fXP
i5o2tUlau4WabBX1IF5beseDr+3SKEbthkQZMK5xxbYjbI5rFakHJ8qH3pzVixeP
+W46NFo6dy+Yp6DY4FekdGx5fjGGZd/4R3BebL+DgxNc6LPtiV3Crv5pG5CvBGyo
bO8E49ko63d8w9jYmzQPPMAZP1QnmkeCLxGG4jMDc4YL85hnxlDMi+XQSyfRvS8B
64UARsa+5gFg6gOgoflvyXjCvNoM7C4BKtXwO7quduKrBRshD2+ekfBqZyBEZG5x
rX4WLdihhDrFsZTy1ewBmNEzyKGZOQL3f4mQHc0imNHwq+4ZhCGwrOICQzJn+O7q
LNvQRod+nCCMKUPbrcdwiNVgXXkpxbRWlk9v77AMflWikSgABDpTeib1PM6WBa5v
vLyArC/+o3AK10etHWnsChMMokEFSfBtDf0YE3b20J6zgq4uoU+9WsyoQ/n0qNR5
AzfHPim9A0dlW4pdWtrUHdq1Sda70OxCSO8q4+8e6TAaVtySvyO8De/xQWIzZ1hV
FfS9qf81Sk2V3Q1S4FDcEBED8ZoZ8j/zK7EZKZZUcZ0N7QRuEdssNIg37eTvah0t
iPApKjf6hCEM9Piy4YpQ/bs/BwepQXpsYoHJrnpDtqQ2beuAAgl+hviL4SemxgMN
y6Vf841BXdeIDRqNcUKDWAqml9MxpA7g07Dv/GOsZkr3absux/hL5bJvCD2E1isM
Jn+T86woCb5uuzraEEOK/DhMuNGWuRsiyTYBqXL5z77mWDGFh74d34RSig2oQCVn
gov8a/VO2Lc1tZ88bHWipO+xUb3oej+Sjme8/k1DI/73p/Cz+PELk6iKq+cYkOlY
5w+TZU/iK63vjiXjarReYuSAT6JrAKlLy//ZFR9P31Eowacm2qwq6QrrIPxw3Hg9
7UIZkuG1V9z6M2Omhp+x73i5iUzINeKL/uzZv4m5wwvkR+o3eDUu6oXUilAsbWCS
2XgzDpQU9BcP9piu6t56tv6gV5WQ4WWH0WBxbT88666qC61kFLvuLSq4Uxm33Poa
VFM/xvk+2/cjVtN0ScoBf97kvNAa8m0+UIbeTsfzvGO8haCfxoaWdVmVHPwdo9W2
RxnEeHZ7Pdn6D3+VG6+em7Ie3oWpH2Fi6CVsFS8oBeLAHvMGl5q3942B0q9Yf4RU
S5HyE6jGc0B5BSrck0l7amc8qPJRiHJdR/mCxrO1B4KL/63JmOo3MekfyZd38BP4
v5vI+TQuAKY0MAYQrznPxUpvxBJ9kc43OiybD8/IpDrrf8flREnxaxTJNC1arVjD
lXa8wQsG3LSK4M+hz95oTmkehqcDOfI1hYVw8khLXDPY92c53zvhrRVDE29e2j4H
tpFS5fvd8Jw8nW5W9b9HLZ/JQVxS578fvDhpI5BpibgnlrsbPiBQf5ZfvPlNRsR0
Hpsv5n3BeS8Vlpdas91iqBX+m1NDYh/KHmAUfNvrl9n3uSh22G/8H0ny3glRA4Rr
/+v1jDeWw+MH1BMFKBnlD3hIBUulzX+XpIDbjaR69BpgAW5WJ4woHnLzBarfnUEz
WPtAmAf+Pgrkw+lhmkRGPFpLp98tPWetaSaCRnmFzSIFJF2jzYZmORP6CEH/y3JP
RtlatRH68ApCwB1LiNmQS2DMRJObroMWKJqUT1+zlYKIpA6cVztxt+8XKdSvZrrQ
S/c4H8YPi8I3+1giU7UuZfNLyk1Ud92U+fGghPVIEfBbhCJhsFl+Ypz3VB+iHlkE
dUZ2hOBOjwq9DOHXsxCzhSFMVsISrClV3iG3cL08XFjwE1fDsZNJiV+oI7c4BsC6
7EBNAeia8+JB+WnaWPSIUpADr7+89G4nzGuhNOhcy0DXYFI1hE5i6qjDkyP9JbZC
YY8M8v+FvG2oymCIzB2LgDWuzBrS4kRl/0ix+zhIIL15EnmxL/zI0lyFTWx3h4kr
pslSVXDsZ+TOpyVVxTUr229Ysed+1vGBilL5WXQQQktn8qZVBxuUr78dlDrelxNT
Fb/2F3lfDo6ehWyOqDCMcrHrKcPrNQ+t9YCUGdjBaLmc20ClknZhQLP3JYClJqEQ
e0fXfjY2i898+E8B+fzFv9l4eWFaUsxTFmzBE6piZv7/DXgE9U0Ht/MhaW/nJJ0B
Yt3j0q9ZyqClf7psKe8QMspzO9wPftc/x4Vn7TJAl1bQIaUubX06KTCe7Imm5S9b
gNlz06ZZquYxrmmFTEmLgwU335TKnBlrE996ZD1S9+z/+yrH+kinDgUg6fXmqV6Y
IF2Pmg/3NLffwGsJPhn6TAJpSpX6Iy8/h9ofWiDmw5GzgbFdC2CjhesiGYlq5WEo
VmmK56gLi5WYcv19uhGP/ZwDDQxmEzlYe+KAPzUIU7rIgtxrAN0SQRX+reAX21pl
bAEyWF+EUS2xnoj7z8vkUJ609KUa3u90cdv16AYCO+yzk5GuAMSOgs7S7zTrAJTV
lv/IfpIAQ+YAU+5Ss+wl8i7gYFRcdZ0qlxUpN9OIgJqLeXdlvC2bse9t2uMgw+vg
CV51+qV8Fkw/gCyFwBvwL49Xv471o6G+0ptyn3Ia6xHI97YW93okNefCfMSWWGvN
CkSZE6vYwE8wOLC9y3D1wad9X033V6Ev1KAzVpCV/f2PNiikDXUR51bDWYrq0h6O
3sJZCrKl1uAmdPYZ0Al7ZcBmPdEmB6Z/wu7hxYf7P/eJPFHVULXmOYEE1W8MVbJv
SYs33i1/FkiA/wzPCcuaN34HFwQ2SmMIgcYI2dp2rUGGcAYZu3SFG0PjLe8qH5A8
KUvWeeyj5f3a5EX1etg3InL/MSZjO+/K8HWWQKs5OLs+0pGhokDCDkPHFl435lfa
Piiyh1bJFZuiioO30fTDznQCOrvW8tDDzOcCO46TM1Ohyjh4yL5BuL623J/M5+Vv
QfLOYgZHt5z7E66fDCPw5P2UHKHSa9MSmuJRtGVLMHIHevfRyGxssankQ5ePJuFW
eFAea1unLT1n0/ZLjZB2DrYBInLbxZSGFUIuoFIAJi3QcfmGh+Vngza2L0Wqcs2G
RH7NCmK2oLlx2yfA4yGn01SnjiF9shmaduS+yJkhwp4i8bvF55HovFQp1U2oLOLO
fGMJPgq116zvv7cHCgnfBZ/GeVXwNnGHrMaeVX4D1nnZanXdevTA+pwu8qZbyRAK
Ll3z7KLi+kXM9+bdn989biYbOpd9r1veAQifYHd+UVBXpM4I/94s6XK/ckQAYD8h
8YTGgOEKcZBMFqgt9JURcjzlPo1YN9QNpAnnCnMfkgzQVKvuIjhuujLwp453NuIQ
MUyHwx70VG3AhT6tBIAsoII9+azqPkFO5QftLkX/t/kb5N4bE3C2au5L6L6Rdf2S
rU1gOQ5g8GSPscMibiqynVQWp/bFhKr+JLYgCiIAV2DfO75nrJ0AMAZhydD4xleJ
86m3fmKjiWKg72Q5VG8AX/5C+8KzH61gTPL8E5VEEpxdO4GEuQbk1QrTnoULqCdB
en5zkA9SFYZMX4LYdzPZ8LteAli/uwi038XrOiA6HiZXKGNX4+4MzPRWfwdRB2qy
VED3gwHU91uMBZGGpLMF/5so1KM6kz1PxEF3z5uYWJMT/3DguS8nFLchKahOjPXn
b94In6FI4TovQrWcvX8ClpwRsIbBx7QB56L5jVWcuwK8S45o+yQNbT51T5ffivU6
MBSqZCJTUSGJwme4FFG2i3cNdW9RB/8yptlfnr2LbEYoKstrXz1sKhcosmvPGM3n
jNtrJHDRs0/XCs2rbXy2G9dUvpTlWI+2VxEwnmGU4ptUsgeJJf049L5Xq5Od9MVk
ubtSeiDz/z3nYfDpOQXqFsMxhFWPLVEi5N667tXXaTh+CjUPDzcwzTL9DkF8CZky
YsbNtmMOTMqYiEBfiB5Qx8rLI4mc3RVOf84SWJN7l7um6Zd/boOu2DNV+udru7pz
BEmDPXniTM3nt5jGO0+RAyUB84mvThz4m7D1v519Dh19z7PlaobnWdRMRz7OlTJp
+68tTz2PVvUKgeSK7TsKjggIIRguPO2cim326rXgXx6NgsbUqbCrMbuhhDNmvMm8
7LYGiEhsgMYRZiMMrikWH6cCaRgwTUlNoquWnd5Hf+E+xdZeteIUwZEbxXEv4/wD
w/kGjGlLq8TBUrKsXQmZciGG47UfSJaO+17BQ1GT5B3R+8/loij8xKTZfDZC9bgL
Pliicq99kg3PloMxIInmhas6qZPnSiDtdsD7CQgGIRrLIx1hfByUAvxX4+kb63UI
T+g3BLoNhRsCTMyTB91jfyy8HxRb38qWOo5TJLk5lNMZNMJXv1quFJdNmEbMsBWL
JwmmeAHxcz/KbRgTBRyvp6IuHCTP06lBTfASUKOajQqRXFdVV8RWiuMvgFAhIeau
lViZF+kzP0907442jCZrpQwZLswGN2unZ6UU4Ezu7SRwYVMfUW1ZoHfvwzJ+/aiw
kEAyogy3v3PIFyMnLbi2jaOvOQkZv7zNmIh1JxIbPusS8Vjjd3CxXCyOLmU1a8Bb
nxlfuCr2bpzzfjoO5BleW1z406F7mRc0taP5mWNJVQsI3mg0LAUc5axIwg6d6xrD
rYn0zi7yQrp1HEk9O+j5qkWpQt2XUs+P9V+4l7BxOdtzwhBaVc9NoFDWxV6s9nMI
7mW2IHEdcztzZio2EahfxY7lverJ+NlA901fT42/cN10vAgEMsGV12mHi2QZ/1qA
T7Lu7HKTDPnGjnqGfZL+ZU8zb1cpq35211yYaoSSgR3Vz1iA1dO00NPzssfei1B1
eKce1C1yL8sENFGjJX3GosZ9wpsi1kRO+YuK1zFzEJEIdDJOXOFmjfCVxNTR5DcD
bJqc5fTHArjKbBSviJRUkFpaso/ZRA8sBaY2mTt+h5z74pdk981l7CeLhGFRmL1x
4GmHDAjXk6rql+H5R/y542HyLThQwOOghxQ2MaBOV4bt8W74H/RqJJn4xvo41IY/
KGqczyZt6ueXjYDE39xL1FbyrVWDwTxYQ/MHSZXeUMEBcOYq12KgurRygetmT3tq
WuVPagz25fW7wTgmTS9RJSA1YkghbmeUo2JMVsrDK+W40knV5HeKeBIru3m26dT7
WRE67X3RCEXoyuVZe2ldt/cMPD0r0q8TtyoxxJWEiznF+X3qSRQV6Qw9am4D5WQw
lCnDmtjhWKAZCgTXQY8GLtKQc8J4WzSSVdKf858AdJRazdc3Hxkgw/irobelruob
QxfmA1xH1mbROGtpPk5LEXDY+l1yCg7Mfdan9dpCELypP0XWWXiw7nHkQNsSpsUq
uenC0JoSs/g1sDAmRhdvZZ7ktRbFM+srncT+b7QB7jI19lPsfnoVHudamEdgr9Z6
zE0/6/OfrU/iHr1Y/RfpPv/Qe//M/0w3jgoFIBSjox48USSJ/AOxtkAFaszBHSs3
/NDejnIf84QA43R1spxMYy2Hk1nmhJxMOhXCdb8exqIKNyVsWLMMVBw5GjIDzGsT
E2b26nvvSHfFwMV0K6fQbH7NNvCAG8RGi6197GJ5vv7kl42dr2DJ0CPXECLV7n5k
V4E5MSDNfOY6W3yT5PH8HtI6GB0QG7ym8eEznIblq0yg+jpsP0YnVyxSlrkm/ehS
zC/BEPAlgOsn97BJhKHQ5mnwrDa8m26BuskFKgvADJL2gk7MsAXq+Eugv/2zdOwP
wk0CQZ676alJKu6RK76r2uZI5EAR6qNodeoO41iJRX4xX2uegpZ2vfm02gF1raeh
KSoKGTYj+UeRcGovPs4SQtd2Qa6Ik030eYDe3MKJSK97gsHTeKUkJHG65wZlgEQV
Uz95s9RbH1YcaFYre3pBbI6LwVBoz9IXzvNenQdpFl4BBVjigG2Fv5POsP7Hki4b
KAV3aXVtaqOLmfEWHrgg016JHC2NRVeOokmU3r1EsH3JatggyUui7c8YYaiYnCSS
JAA8utWWn8r0m1MJCe2OVoksDtqdX1LqeVmXlNp5ncU=
`protect END_PROTECTED
