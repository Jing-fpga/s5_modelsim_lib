`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
16S9/nNaes15w6SuwZbuZzwdtKnfiov7CzqADPZt3lsevZbBbWyLK3j5hhRBkZ+i
jC7Qbeb1jVGbUdYiYsWCQq9k8eGsf3zEph4+VESgOXceJOw+K9u8UPpkB61asYqU
FZ8eXScvRxywwzS94pwSm93JCxvGEinbp8AqqXuB8w/CHKd1+V3EQxkfJ9UTW1ME
cD5GVjx01mMxLe54vkiE2u2KkbyDVgNoRJfYLGz8YvyELokOHsi/LyDaXGiaXV7E
mpqhGq4SE/l3+0WsPH/HdcCkVjpI0Lybj0Lca+oBH1BtnIqjoOVHW3kacKeG1OcT
EtB/dip4pHF5y3SPh0hLnxtD0Sy1/aX56wMXySHzgF1wLCrPcfRW0fYKPn25XYAd
+Buiw8uuy0PO3RjJpwrNQ7Fj0PM5QycyqIwxfZIO9tNHBMMyzLkgOI4nGc4+/f4J
i8JBScEQD6lfxSon53f2d4dYyi906EvUBpHHT8KVFhL1OA5y1JE7ufNY9ZxlbF1o
KimJSsyZ5u/zO93Z0XEaH8XyeSKyIfLfpWqavsecRTlyuovju0LkVhmcylWdmsdA
RcqFBraE2mj11yqVvI+cegudymgjzpvlrAI5suS0zgT0qI2jQqbeYdcheflgTbyF
um2SK0Xb/HWf/FRgtjGpsCI9MYgSbAZJDj1r4DC1aMkDUz7Ky+AX4b2iu0DLf/k2
03RwnpjWvvXoCeDFpyGSS0tgyR3QQ3RIDaKbLJX0jzpaB93J5npniYEEfgMd1YmZ
oeNd5usJrp5EfohnHNT+Qcz9vBmrzUlGj8p2mExjdxp512L7xqSnPi4EIXQl7ZKA
EviKx7lW/lmjQC857zx7SotDBwLi/zi/4UUxfHQGPERep0FNoDydz7CYJ83ICFT2
dI771AFH6cnDLazFgpv0B/h7aNA0+LMMjMDWYIeGJs0Yy3xRMZSYpzZePPBrQHFw
GcAQFAhNzkeNRjVRz4h/PDIujS+A2xFTSsotocu4711tFh79FtDiIWsRMr82KFZM
qOMlgLXDpmdnxh85u7d2qidpLa4JK1qYCwiH0TVhyO8e+TTRk8yRaXhbWSJiy0f4
hTV4gs5JRvADuVNX7SI5J5/aMHo1Al3DDd8swlZcRnNYfm4+RfkE6bmOGQ7K1fZS
F8HvrddntN+ZWzsiSJVa5K/4aMGZ3druVoS6EirSQ2cKcdAxR/GiRHOw69k8mYlk
ZSDrOuiu4wooEdKQPLI8VeXMLOfomHRsVUnJEhrEMbSbrMOaEcppwCLz+3nr0ku+
nFKx9rKIcbUdOV+u1B9DrR/STLaXRh1Fae6aWVogQwWfYeKcchqdhQH9yhB4+7wE
hFTLiVRa9mpcFKHD2eVbTM8IPazgumLrfBwtwpobQWEBDzf798QCFHY4NOgo0Y2g
7+TgldHUty1jg1BgkYyhmDMRjEPUJeCz1rrMNBuP0h/PM8Hpe5Wzu07xu9CAfDkN
/2BnjpU2ZptuSIKJNoUrjgQqAGJfee7gfE8xz5443zP/Pjb1tz4MI2Hdbsjts8eC
Jn5KpVacp+oYp61gibaVbiA7Rc0oGgUhpZTPD1TpaFbsru/TVY6tUzv8SLDeHZXB
`protect END_PROTECTED
