`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wiSBJi9dzmGmTqkhpR4OlFRH4bBkBE+gqy6muFAszIpx0mjtcgWhtHktQX5J+a4n
jbGfIQ3rzD94CIDQ0alH1AhjAqO4IhBDczE5dWBD99rq3avtwrG/iVk81OEhg/qI
FDDAqCgxUWtdc7WwdGDSExWZXPpSezyBkEr1NGX8yv9jMuHqMiJU64801SGe3P9g
AQKQYRlGOKGRvEQfbbsO5JSqwk3+0oquUDizDZPgJA6Poycgc+yb+txedgSp633M
RvuyudvfF2hqB97uVD0XHJCPJ5LriF/FTkCQKMHxFE0PzjzE5YTQuLn0egQizzgd
T+vidaQE/7lbw+xHnjTR5quFVnPDk8gXKaTu+WoOucpRjOsBT7T2Nhp5D749/Oml
KUQnQvxePD5HDMFtR+qqxHfLOuciA9SmWtwqAvDKhGbm9ikwz7BXOkFaImF/+qWF
FIDw+hQhml2+uav0UH+wK6jFkOkc9IySkO//TmGXcb5bErHg4qq6jyIclwL9b409
WHRDjldb0qqh0vl8Bt0mldcV3ncdM5uWlLzG0rg4US11tKGIeyIXWt3kEW+tByqg
Dh7a9zUcXAkdVo+ipcrKnV67vQ9MLW1ab5Kq4/S9LqdczEVoX7yVmkAVPPIopcav
uw7iDGD5X/dEXlmfb6dywEZVKac94vC9OPLTMyscqF8lo6A5Zjhn1uChGTTeax6q
Qq9QXGMh9beBKI/I3StrKFi20JcCY8feY3vgjyxF5Zx7YjLTRGLlATwcZIaq6yLe
kUePeJ+E9Ui67j/LCWPQb9h6AO+oGHp6iAP1dEn5PFJjcAayZRvSFcNkIG7LgZEX
B2k0l71O66oqWXRn83CSF1so8BCiNcfy3HfpFGiKz7+hYCMDFWEbeWUGmZyYl/G2
Rhx6m2QR7xdiU9pU2diOB0L3Zm0t37mLmC8hztXpvIO2sHvPoLPW9D2YLi7z3225
TlU+32g1Ib9XIM8aL50LN1yqTABhkZcU96bw5UdYHDw/v50nNOJjYtCWyAWDrL+J
ni83tb2ZncHzQTPTmnWVVb+RxEstbxc6S0oIp6MG0L9GswGcebbmC1w0T4DBedIH
uifVmcnj8RWzlM+Mg49oUIJXmRDvlweAL2epXbkOCUk2OfDdWJs8OdYdu2gN2Ya0
3arEvKGVnNGIw3gKRm/68CJ5NPZ89FiDu7fLPTqsSa+9ObSKIQdr6LZrBmoMXwTo
uM8mQdbykYkTpgRc7zOGRilzRC92GgtbrIekbKaRQFnOW9wBc3xjI1eHHY/WFoxw
t949hlhoiBWb40JNjMzrn0iwZ7Iv2wVP5R6IZvldR/hXYihRCVX3qKN9B1vh7yiJ
RM4LXjurs1fVJ/407iOJi+hieRXcnqEl96yrWYEYF3+sljo2ghbLPPmCm0003Js1
2FT0ZPcgUZocI7plRBV62rCRSZV+ZYhZ4cZHV22iHIieS51Zy41pH21WwAZXdboe
H9BoRu/pZfwtc4qCpmT7BHptEPJwkl5+m8pekDrjmyWEwwUpyYpxeMtpQw4udnrw
vFw8nOsxEm/zyPCjsfNN525fP1OcQKdVTYVwnSouNV2m8d+xT9YUCuJ1YZ3KfMNI
xR+MSvHC6pWPBVoz65mNn5CEHhU2Te/RI3vVqem3XIiGskVBbVnuSvwkjdL0T/eg
tLoXin9NyE1NLzDn3CGlU+uCjZG27X5UYNrI/O13QZaX43FMZe3zegOZ04uOpSyU
Bl/RRCQ+mIEDhmPNVbXHIy3Mq+gtlJLlKbXvjF3Uyagio/RJm45rSV8hdacKoLZY
47XQONeuqabbelYsct99NK88cnnJNUNMUyLmGr5s3kN1kB1pA8Jv/0F4hAmWCzpT
i5vSp9gOQVWBM/sl0ouRI6LixDhgXSGnY2cvWRtU8Y/FgL0WmxTAKK79Y0ZD/l8h
Eqtcgg3EELicP37qdmtKOMmqPtEIaqI7vi8kPwjCgRA=
`protect END_PROTECTED
