`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
exkFWqEO76QpaVwpOwgBq625JPdK/uxIymLNYucrX3cQXxcu6fP85FhFLgKYGV7F
BvsuTXcFTNFds0b/z4n1bZbj35OEkr9CwfPeh+w6TDu7ll0M+rZvnj7JWtuWf/GK
cOkU91jJzF+Qu3trQM3idKnGZJNh0SN9ULJJ3QogRiuY1XXu0pWFwn4RCJJ+ofUF
sX+IdG1sArE4rtbQZ7zqzsFLF8UXaqs0pu3cRuOU6XnK8wDItaHjxqAThSzX4AkX
BnkxtD5lmNECWpxqfJjBopCtomVJLAA7XLxHW2Ob9wzhciFuLRf8uCu5M69vT0oc
KQYrLOcX2aD49MZX8YTIOspJW3v97Wk+skAgq+WS1q9mNL+f8uhGVuK78J86gkzn
UM9SfUHhqNwMEZSYVoYn6ILCPW5PI19T+O9GX2UO6OxnaR913lAWH9UPuMKsqLA9
W/JVVXiwp9m4frssdZpbSrDlUs+1lsrApcga4bIauVcie54gDALcnC4acsbsqYo/
hGtT37eU+dx2H7xgvgKBeqJuGfys09BeO6W/UPrRg4Y0E4FE3wz4ZCYhTnGk6hIQ
MkHFvORY9pezdvX8moffVXnYnslFrceGIAxo4n8UAm/nFbMMq8oCy0gLumJ1q5a8
cLGWb/zqKCRdCAlK/5pJf14Gd/LH/bvMdbH1Tidlm8Nsj2FCQbRzo4f54IpmgiSz
fmrDra00HzZU5LaJt0nRjXUMa8Z8Kn1IQYD3t3zd8ftYs2oN9QFNS6UKJC/Te1xt
vkVWNvoUf94dNgZaJCyhPxPGbpmTlqCBdMHXcmVglCu0ja6ch5mEe9lTfNRRyc5m
fjDdgZ//Slj4hxnRUYPn/8BY3Ozs7dKaRRsVpj6jS/uQjEn2kWwoGZlRFnHkMBDS
OLKia0E9LH59zkNB6zX06EctlP1DhUkcz4//+yNQlAGwEY/N6PKhDrxaqgPyBZE+
yopcixzwt9p+ORIcp1hbTJBcp3ZX6tAu5sxV5JX9RTfeM720xQ5bd0cKiviy0i74
7hiCZuCitG7r/pUBikXE3jkS+ra8dgaCu5ICIVy2JpHFGBbiswODoGxsr6vFasoP
N9PKmMS29F5SjUbUlMUGblXVHiiHbLe6GisHS5JbM2eRn4wQHbQnI8chAggTLcr/
JsBStycUodRLWqvJ1xsRJvemtQJzRu3DpikEPH7V1yPf/l1jtLQ9dOT6HTu9uaJ1
FmoTiWDBuu6/A28vi7xTuyUbNW2GsqpkrLwDlA2IoLv9dGd9dlrDeAXm3DsZ614i
q8p45yrsykyy3zIP/gFtfpKZezt3IwqKrz+dMIKeMx9MAhAoVff91Dv/ohv/Jjmm
nh/dycBASgjK8Py47A8K60d+oTmMVS+lGqmrvI3bmCC2WNssLhe+au+lUen7HCI5
WOMoRJ7Jk9lTKGmLZBE6TmA9+JWo23kUDSiHQN7o+tJgY7lrPL5zpUktQk2fkM8B
/een/iXFqDfKMInEBZTxdFq6DMHCTjWE46YCs5cU5jcsW1fL7RJwgU1X2DR05FFU
AH8uNe8f+F9iKITog4y5PHPgNj/Z9XJ60w0u7rwsG5tDBJBtTmCpxUBCrn3kj0e8
3fkfcAL9scD9qLwZVFTZscNjwKRYMGdq0o6qVhNF/vFRcMxbqz2+nMB2mweAZ5uR
ZpNL6CTfsoZH5+g3n2Ka8vCztLlfLrGqZEmVkrNx8rGcukDjDfdfM5gHUlc++bBV
5caTn5PIuDvJ748RSfTHDEfJGOHKc2XUEnqQRsG4ft520oKQHIOIcbdX2liazfmU
+pIHKuTKrAenGFCncAyMC5s4gu3k/vqJgSNhGITn2V1ugIUaIDjd0H4UiZ8HbdGY
GX9yVZAxaIP+jOw2crBKiY7RYB38qT+IQ+R95gBzn3uOLpm+/DxaoVE4uoQHEmqj
vuElA2/mx0wSbMj+9Q9Zb5glv64FhJJPE0DFKdpq1gWP7UZd4cOQzNxtaovg5aQ1
iIYAcvY2EpKRnF2Sg548AsaJ4MZbiXy2VCYrxvvt8OLtMWQN5fXlCsqR+IMuCx+L
WDXK4EwiU6Ts+0VCIUyYYibw0a7/t6iQJxvtXtAKCznQCsmLbw++RtzTPGZam3Eu
wwoF9X0FWat79z4uFeT/x/ZUbKy9On4KNrutDJk/Vw3dFJgxqLKblTqS047wDHkx
`protect END_PROTECTED
