`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BfyjKc6IXvvXwhgMY7IzxwFmyvaxz9TpU7cB/yvrIIb+pfhw47T2/1YrnqhR0dV/
I6re037zxjjlVVpitezaaXxzsPa6XuAEAJrp6Itp480V8f8pLm+6ypcIGwts+8RF
0lRg550hRVWnXL6VLG39DHsyDrhVjA3J6pTdLHsinFmp6jUcRrjHHZkrt6wUReJq
s+kKuUm8QELf6+GhOA0bl3aQMyYNdpW85T0BWOseiCxyRiy2HIPNSmP6T2+Ul0s1
A4siz30ooZeAQ8+XTm5eOGrWdHRS9m+jtq+MX0NvyWQ7qyO5dW9Z9n8tRkPNaPf+
UhnH84U8Os/9Gpdj9pv7IFpThM3Rt9V1KssZjPGu5QUMrRtfQ1NPB4GY3/y89TPF
Lh6SU9sKAaPajCwnpByl33ko3nEa6XOmHq5zBNgi1qnpvehyJo/2+YrCELcH7CWS
qY6NORfE4ENTfOoxcPNxlLJWgL+X0mWNRyArFG9RzKf/PDaeHkUGew5N6cgsB8DG
6TA98YYF7iBJP5j1/Th8TR8mRrLOsWmhLgNTJhxXn8bDFqc47qpKKvY2dUsnqp0f
B7ILDJHy/fHcWlwh3SZs2wBOcVu++Hj2S9lzWIHGo2Rw6EvT/2wvhOGv8vmNlnYs
n8zk/cyVu6CovLBsFDlvRuEzmuH89xAIXtY7FXImusjhd3hGlurtASRBkFrRPFQC
2MuBFDQ5RS3AFtGB2/V8d6vmNQ31Qv7rTrrNtSszpzHIdX1xkTULLaOUmkNFTSp4
cp5NPhSGW9MQVIeVmUHc2StsaoI//IQ2yhDvoOq1CUBIwiN2Wk9P0hd3KW9xgy0w
vQI86rVS5ioRDzjGLt6gpvQpTZezvDJcLhlqBaijY+ydqiBu/JfO6tix6/5Lzw8c
3Dqm+1OHYJfC0B85aPchz/4IkgULBN9DgWpaXuBsvdsokU9od6HYSN/stpRAg4pW
hg2IgPY62VP6dLCY2o3EfScl2sbsPAQibow+rnLgC92z/6+V5BPFlwpvTGSa9aKT
RPAl9MJDhCFKkX1emihxLa/i887eyGlwc/3vu3hU3eI/C6uZfCl4xFvLdtNKqIhc
KUvBngMZZw6i52DDqTou3omA20Hf5jHWKXEbsyPgtPr5tLaLYk90Gg/t10ePKTfQ
ZVqnCAku4YjDzK1pveyqVHtfT7yEVlGbHxsECacw4uE1WWorC8pkYms1ToDGnhOF
xpOGSwQnCJP20KneCHeoCJBLewzY/yeIhFfrgtfgASaM5YaamDgnKqEDlQxmNKxv
6ZFBrA5tnOWN6wmY1g0GO1CPu9QWXWR2PYDdAgl5QbZ7ofa319xJfqsye1DeYypB
e2dNFcJjODRi1ULkvWw6moB/c50KR3/3zpU3ApChJNwGH7q+/7Jmv8L0qbrJHFwk
QlEbAInf9TPwmjK6oqdj6pufSH+9Y4+1rCV023xn5H/StiuwlGdwdaQD3RL46/CO
W9fFvz+IEu18Ed7iZbHldrnslpImNZ9h+KVkZboLEXWhZcV/T8ECB3efHUPmVOze
R5mbdktYIkdxaZPjH6Y1+6IR/m1OS33oOvIAkfayKVVNsoLX0BGg7E9iNWTikQ+q
3+l6/epniJW09/MFnTcZbeh2eESFGngNmhvLLYfN/9aX2ZUpvYZeb1mmUIPMzR3E
K1D9N6LFIM+xi1gOUTikIjo06lS+okdO/lCME0aZri09Y4P3251t6+EoUHVJxe1F
DrtLXEZsHqhDjkN9mn0IM2ZlZ8zs+/sgawM/e3vKDHoS9X7QO1aMJamssfm2mA3g
XDkT1kt1I4SFiDQQcVAujfqqjewYWilphgArqUYb4gbKOolvSnL4qzQezwyXkLUQ
8t1gyls9XYxhw1aNUMUF9C+D5oskDMpkiTouC1htu86GoY103s0ba/JKL/JWgro4
JbRFgofGK4WBMJZ4mJMhZHIttWOwAbFZZ9IvRSIaoyjZ5baMBA/GQqmbOaXd6DJc
xufUu+uwMeebWMNU0n/CpoU/jSHr8r2zNU1oo+6HITrVACYoV7D3Ac+fxfRbpg61
a20v+cxIjcW1HEKI9M8+dTddi9hhqGsk8zPh+g3cy3C+/nQWYWyrglabvwIOorIc
v/y7vrVIIkrqv++xDc270WjNbiWVCcSaNMW5bsgo0HEpfT+MPtU7y9bzEP60T/w6
P41VNMmr/YVUt7h68qW4zuYp9pWz9gSbXPXIQmORlwZSuUo92WbMfKzlKpiUTYvc
JGWxwVPfl/Ra/fq9b0xuJrO5ZunqVHAeaTck8eHJXqp7Ne2i+O+JWK0DH+AG+5lT
RK9I5wavZNpOV6HDovOwOlyQQgRhss8fh0ip5aeyNgJO4/IJM7Pg21Qr2+jQik2I
D2RehRsRvnivA/tzQPSQpEkY5jZdfWgHha9yuSXNtJJD2w8oQqc4n/QzkywSVSXC
4lfffFp9hC1G620+InOGVbXfhzry/VbphpksaFsN3SMNmTw2f5BBt5LqD/5gjqgw
OH1onjvw/644FHG+vZqCdXyH3kmsWFxtwpxvy0fEnKMJKbTfWn99n/7Enyn8MNnc
YswtwQp8wmqd5nQ25kC7gPKvB7bdgsjoAK5icpyWqcRgkv8oNUGC1dVI+bmlbL8Z
IPvJFpBwKjdvUSxw12DVNR23D5vIxTd8vWHrM8mNtSZ1qC387OqWnnQPclOV6s9M
OncJjttAxmJD9gMqhIWpV8oVgfj8PB5PCyj8vQsQTTwO11czk5biDkQ1FhW8/3mH
jj3bm+G69vTPA7vx9mqXc77DsI31/DB1X+/oEneaZT7PHt4SEM17Scr21G2akJF5
voHozJKcgbmlsb0BpX+U/CiikzsR0VGBPXP7lZsV8HjNdnTk0LMYPXu7Adx2AHAy
VLA8L6907ABZOgzRmqwPbBPqdhZzceQjKuYYv9Zoy3e1y8A0ylk/LN1Vcl5/BUzj
CJKmrm1WdEAMawdaQzi5/fMv4VvLXmb8hUhtXpxTmD/NU85L1FBLftNfVpCiwD8Y
owjrJxlyRfh/AyHdp9EpA95twIC4FvElqgMb94E+8gkm44m7PfDMJsxkNKxNJKGV
2/VH7qKpFSD0q5mh4oDMxtcztP4CtYJDVQnL4qIXdDLJSrPOiOfi78+uS4HdV8A8
XBLqXVVM0p07rw3fdvQSHPUOgPPChald9/1VNHHr8H9XgNNScy5meEfmA9LOpMUn
kFvzE5fnI+jKHrmv4Yhz+Mmlf7PnjSW9ZgNvSXP7Hn1z4cUdI5O1bmxzxi1ySOGT
hm0Y1lT7Dwk6vaXtUrNfzGhivN2dadxrb2hzBGPQTR03oSMSrNnmcXeErY1X3YKp
Bu33RWEF8dJ+2jxE1miGTiWad6POp5XUUP8II1hUtDOjb2yOqL+IxrRBvvgRIAXN
PJtE7fS2gni4FYKc7Glu3vRxjW+vf8PCsyauD3uZpS6YQDeXAchz1h5Sx/Kiyy8S
Zg/jtPSALfPFzohQIVK2MaHJwnP4KNg7JY/uf5fHb3QvvJP61AXMrf1vRW4VZdOV
VJykbiMKaBg5SXeTUNHOK7bL3z7dVm2t8fwbm9eckInE3R1gwWCteg0Q5+zlpDfO
WUUNNg7+XmFDKoqnDuSrIOMkTx4UmbTLPnI2caytWQYF7FKmo97qEfEuNc+W8VAq
5aFTMkp8tBRY9EgwTtwLwesVAZVKGOqoL3KctDohi1ZpHzuHkLiib43BPmcPsjMo
h9bgHe3kB+f/iNlp5JAv63InL70ZQzT/qEvxhQfCtCXD6GQPDd+hTrGnoIgXKvUj
aZAAwcBhI30d4bXliJ7nIWVI9RaydUdAEorlQfT4fI1pswWgR7lW0h06L4Cx467f
e8sr6RzQ6O1NbOxMGGe15kYnszYeWoEoWwqDiQEZlakRVPtVglrzthYVwk2Bmn3q
47oksJhT8xaekXBmgL3HwVxiSeUPGPnDC8Ra2uzqZDsPRfmGzchll2JgkmUgWt6i
qXiaIKGPwJ4wZe7H/AampBAOOAI/kqokp7qW6GVEp4KQZwwBJy9IajHiZJpPTH/X
vqw0xf+CTXVAnlScAd1DJa0I/eAuhVVySBvRodLCF6xE6xKqVfa03TKN1TApZmxu
yV0u5KHAe5wpEJJDUHd+8Ke7zfhDJDeY/LiVrpxx9uj84YdNFLBkbCji00i1EPZG
cmkLA1RTrIezh3oNbM2MJbibSM7wELXmI+e/b9o9CGJalXicMPKyzAIl0r6EW2GL
ZgX3W3wL1AufH4tT8hIHbC7S/mRT9h1Mi0/Ke2X/kthYkFxgSOD7sUCSyIQD+C5c
zQxGuI9mJ88IxDoLiMpFRFYUkTvTYkqQDSjs02ELjKhUXv364j2J7HkVK7kxgMF+
kEjZxjCAYDzBdfhb11mSJ8WzWnOfLa206laPDBh3lBV/2hEk/A/rYpLft4cB2iNG
Aqc6y+BWDipB0KMz7OfaNFm+hCHmrrhcZPiEQgcyAkg1x1NgLaX53uh7l4fAyFu0
aqnDhjoH8ec42TJbEWWU5HdGZZUnotKZww1c5Ew/GWrW1eJGQ83jBCrZ2mglnROW
/2qt9OxYQ80mTSOHuK/8u6olUHM/BWL3iOpzHwS6S/ktHcMm+fBeRO0BefyY6P1p
cWz8llgz6mu6fS2FexxtWRlmsKOFFoQ/Dbl3lJGiq1IAXIXbAAXQ75GHminoG6eF
X3Q0SzRbDKgjdgwUoRuDeawpJprxnsBQTOXFBSvvgLwMvMS+CyrurnEzxoVRehZQ
+Xz4lOxyEE5WcKitcU1Oq3OjS06RZrKOWM5+i2bCm52OATXfv3zLijsKD/cESDho
pT0DkARgfYQTlMhAWUOpNh7qRU9ZjvG6Sn33yRcoPRgh09UHoB3jqeASMFLrq4tY
ZlTe2PVXEDb2+3zZjPtBtyL0BIoImGF5vaDTihF2eiL+qKyc9u7BiKUa6maI94Sh
QbZwAK04ctzaV7lUXZSQDPTZFBeL3A8GNsiIOljPMo5W3ev1K65WAl7ltTzYcVti
CTgo9+lxIpyEiIJP/lJDerGWB4ff0IiMkau9dI0wfhH3Aq6O6dKPbDOwwT/rGUku
pNEOlpbbzF168et3eJVtTCuU3dQI2lhEmEBP7GnpYDOJfyq+wRVgrhewXRVVaYl5
NlJGG8jPwIwmWaZRwjwDW04Wf5G+Pg6Pb9zMRxpoQakLZ0sqAfX5CacodbNwDNuZ
voQ+AtoVsxbnFRYwF5m0qMz5l/uGRjkiFzTmc26+ER4cAEW6vb1SCzUKSiSUSBPK
iIbhs3s1euiBLEe3iaLd/Hek5JoaG9YSdULgoQ/GziOxZRoh9tTKn8VBgUm/aM4V
pvI0Pga7BGDDOf3FjwBrfSk81kCNVrG2arcOm2wgLHaH8XbhjL5ReyPpnM/fmqJY
BGW10pGhZL2b1mtE6g14g4raM27frX/04dizqIPOIPCydxmyygxrwnkkKi4jVR02
1gRW3HKrynw4BNPfxycRKQftmvXnLrznjFO+SNph4xzbJlsHOflNAQUxe7J+tOSV
TkyJK0xhz3QhC/A6yqy2h5hw8Ff5jdEGVgDToDLHKGPFcOs+qpMW89+kYFRYqDhf
E2I7D/8oxUS6xJqJH6fZGxlpxsIV6FFh+u7/fSXe3eNZt1ChS5m4i9foX3C2CHIv
j/4HLZUDfJHq0ggkL12pRv/HYengncrXE3wCvgiMUsIS1cTl7bQP76ZK6RXmNDFA
QAHVcopuJhsrIWfbC+eyn5QxzOybh6EEu3LWcnvTeOVbJWBwLMf9xqpcQYkVzBMj
cY6dX7NgvzSGl/3IxhI21n8gZRB/TtsV2HBvscInGeQg4KDRT0v38FTr9RZYmFYf
a4BWK7saAHhjAjEwdyCmBzr+HhUgwRsGUZacQPuviSpdxXCpziDG/DPEZtyj0lIO
uEmJFwVRgZ75EdvgSglPZJ/K0ulSdLe0dsMeyP09hGiDW6l+Ol7zuIY7IJ7fuOp7
cjafgsIps0oqDKd+/xbG6yLxJhUz/AP62x5yvGVL94Jg49Li6lqSbjTAYyHANwrf
wFQWP7SsaGEL8D66EXM41ZAfK7CA5B2fTxRuXhJLuJgoIacq80NyaIS2GFy77+tw
7CY+yVGDaPlr0UYns4U39snzQtohaFHF1Wo7sBW6KJ36Zddo+K9voIJySMXauB3e
P1cwL/nAup5BMahdGIRWsMlSjYcBuJH3SEjcsNTQKcn1A4EcuCClaRI5xWjo4/Ag
oJy1KNaNbMl0scPdR02FY9oRX9UN2F8GJlowO3pn3cI=
`protect END_PROTECTED
