`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q0/Nr8ahNlNWt4rw7jiR+W0gFz4LOh/PvyAqhtEhmhmKDMkcw6NbiU+QNEcjPaYq
b/s+ZqPmTZoKKLFlljDzwI/dFeeDIdvtmrquod1aEfWZipqf6/g30xJ9XYIMJjMa
e4kJlArRFbbUDyXV67H2NqyoaecJmm91tEYMWQeJWjzaKbd8PoRlCNAnQGSiV8A+
gNY+FdeLwq9MGgXfeLVN6Zw0yU6yUFRy3R56iKYpyKBc8ijsdQGCMqRKMslL9ePr
jR9JTXfTQhSTTfxMrnHkAXR7x4MuDfXRwsvUpK68ASNR6IUgbzGroQR6hNkop+cL
vwvGIoG//+NW93GbuGpnIaj0lsWBzfUpG6VJrSTvZ3syzKZ7mBIHDoVgz0GxRjYp
/owkrzEusvsWNyM5nxZScaso0irEXcN5ezabLZIp3cDf03gS6AOkU8OPIy0nQfnE
JTmBAQmhjnVM/R5U1VGHeNezy91KraN5EOF5YfDVU1dT4qMhrVq08FwZq83OOFbU
YYdxtsLZLixcWS4iP6aKT6K9GiMjHlqVDG5rutHbWmPHI/a3+xp3k/azLlqFiMpp
tN9zOIujmVf/ifXpXKFoBwB4t3PIzNg0EGJ+OsW/sD250eKeewhiqeWm1WRZ83Ef
WcIiq1uqMqF1bXEUDeO79jiDJkBuFeaA7poTYF5prfHgqapFGP+cXqzsbM4c3LuL
yn9eUYyTQXv84gPqUTC/vgXtyKH/rGqmjLBKdA2exPVBxfVO88hgWvMOXF3mRaGr
pVip9KC1I8IU8kK16NNpHjA4yGYZMNAsHdoHzlcbqz37v9k0HGtvhTQD5gRE6ZiB
BU7RrnCab57NvLPnagkYMHavpvz9kCfG6ca1U1prE+oUVYNpgsgEg20i+09UJiJZ
RDlkIUbukejMsmDbCteNelAVNbvt8+ccMHwGwb1zrQJkNEaTeXXaW4o2nmWNCbP7
ZaBsBzb5duWjHhREpE8ia/vULCbMdZkEv41KlCOHGK8WUH6wCSJ78dLARV8OaDyX
0PBh+5pSknsmk9nPAWL3Tfs0YD+AuZYgCxHXMYMCfKViRXiAuwu/1Z+vPmeS/Hj2
eArGIST/RzoTudk+H7cHImWWsjavEiNDU0xwHSIiQpSrfolZqS86rRtvYkebErVI
CvGWSSJqCtkpYO7dFFrU2ZWzAnPyx0z+i/TeZh7M7CXu3O4PATb1I4QHl2EvI6F8
TjFRMs+7sRtq4LY1LhPO2XMaAdi81eMvoB0Gwxq9m49wL2GBrqLfnHZ5Ky5bOumP
nBCM0ylTHsQokAp8nJV7GdjF5dk4stto6egni/RYjuvC+FerGg/i8jfitaJGrRXh
fCA6Yw/QaKImPCCqo1pDSAvtja2juEg4Gio+8BOLec0q94TmmSjpwdT0d2Ey8ZFC
1yh6lJ9rSYdITN4M9XCRGVDdPqdqoXGe0Zqj4dD5p7rTHRQ94q1wZF4AGXDtMwoj
vNhKvLgFgJhmrgF6kQtZMQ==
`protect END_PROTECTED
