`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MhcZkXoBysRlhYZjIhOAgwdLwD17xaaeedqxLqq+S9aS5XBdfPJc13w5dY3Kbk6B
Iv8gimJ67MaI/8ECUNTolmV3ABg3lXRO0pfpApLsIRVqp8J7pgJaLS6YNcqUKWdo
R3oCz0l+X1vNwI3k1t+EHJGgpHFo5GVciCHmQ9z17Ge1DAHvu+rlLujf7ZjPe8Bg
9aZlfqDXJsiE0f9w9BRrykv4uJtnokue9Tl6ip1I8xWhCSuTzhcD9S0EcKbrQgAd
7SmBze5yVknqmN9qVJE6eafGXbVNaRLLCxe9RruXRsMa/buJVRpsEHQHjKWgz7kg
9FGzT2uBPShxLKL+Jv5XvLLYSlmRV6lqs3WShsAxgy82vn4IPk2ROrn/l/tzC/Wi
C/P+JdKLWzLFYWjvNxAnbkKjOV63u2vmx6a1pIc8WRia1fMRsY6/w1KkfojNBbPQ
BfhxwlF63wh6PUjHq7gDUoB2FxQJyh3NU/Xpufp9Jj++eSLaCWzeedIGvxmLxKnj
Xy8S299gghbWXjk4bbfXZXF3zRAtmIeYqs0wqIddx/uTju4fBbK8tGRZ0Zzn6MMP
HYEnlp3lAe6INtyD+UxDhNT+6rDmU9t8WBY9SOxnpJt6U0Zj+JI66On/zliDMoUS
FidMkXCR2DNWUmhekbwRaxFAv7DOj3Oa5uPPGM2yoSvRzr7LZlcwUya/cXL6rjQ0
DqxNbZ2gV8slb5Wls7eEHQvtHoV8QNLzmlQTZzGRlBior3fsTZ0oY9Haqrxz17im
0gJn0d8QmVhtHZfSkHX9jgU9j8to4B5XKrzrdCwhFe5X4ViHGgNewDdN4eJEJgRb
To/WxeTkXW/wv3CkLPSfmAeBrq+QGBWOXv3KzFkAOm79hP9uWUBYnwX1AdIoUsjE
`protect END_PROTECTED
