`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+v0g1DgLTwDz3iXtEGbq8D+enF2Bx5Zc1n4XTfo92D1mWEQK2zdeU8503EypKtM0
Lb/kpIvLIrTwypZvLPTjDtrwc8afZaVXaGyt9eGtY+UI0GP6adx8E1s4glo3H1XH
vXMoh+ZsuxaAne9luxwL1x7PlJSNKRBguW4XheMzG4v7Pko2yFUpGbKqyoWpYK2G
0YU6BrY+abeGVp0jxesuDtGfI186DHr9x21to7cNgSiLEPXzdQ5BuDeU/1TzWAP8
oX2FVbeaWtPLDP8NMnkR/yrwRbI4pUJRoM/Kf2EfrJ2b72l/S5A/k/Ziz0ZuyIJI
nKJWzWjHC90I36xUMxjjmGAvXUWnbZWXzKNVwuWO7RBdu0ELdbGjUtkIDJ0CWL9A
ABtL67BSRlRHHLJba22hNwl6VYEEJNMc9GJGjPSDS44w9G7ZAEHrlZceOgcuuJIW
W3QsB8xRol/2bGu497uqqwg6JHB1dG7dAnI7SfLffi6U5MDUAgfmApbq/J8yhdsl
xIkFrgbsXRnZLwdlE3c0dEibDj6MZHX49RIGZSnhxnSyYwg+TyHi+jdKZ9td9ArT
nR5u6CyfktsJw+77TxJLctfYpAoq3CxqX9OARirFzmww5k0gg9Kx8Ow6SURh5gG6
RY2xq+XGuQ5tKGx2V88lL2L8rX86YsXhCSq6/MCu9uadG9lEn8Tz/xp6IwZ0pbuJ
JGOBlLvmb1/ToMK5vlBAQVPisOTuHaT/XfVsb846AGDKaM0trsLrKyMd2SIiyHHg
P9cxpP0Xo1DEEg6oU5BlcVDNAdpmRgiW3AjmUHk2/4LteFnzW9pPcOtlaxlB4LTQ
w1T0rM9epyRL72xV8PMcfDmEXlLXwyaYc593k81YYTKLJHVnLFUc+XjNWSpgl367
a+T5SlWg+FSx+TgQgV1U6Xc5W3lciZBtrHXMVCXQz9DHaAC/IeQFQJwLEpjFj1xY
ow+9ovlcvEmn0pUYlHM+ANTLMD3dcnz5uvOA6vHc7kgfiJq+kQbSvfEbtzCEebQu
o5IyjUOlKZFve9+78RQxPCTWvItHnMVhYBzxrTrxyEbphFpqgTBMq7LDUUh5qrTe
DveOdopERvKf0V7CguqjE+9FBUQj9mSOxxg6hL4T95tECoLTMTG5anh1Zy+SpU3U
MsvBx1LGE4t29MbGBWmYAFczbMs7fmUK0jwh81KF/VGYSGaz8s90BGc0Fw0qEhhW
AJtVVwPw67J31YE+ff48UzOg1pg/8WSl1CDNVEU6wPHJ7rxP4q6+MYxlXiMN+vQZ
qA38g3dc1vNN/NdPZunYJYy60KjUOcJ3WR6grD3Eg4nqH3baBT1Jps8ioVqDDuWi
sce8phiHSwXqYOVD+w6TuBZ8ynlMyFY45c468LM9NuglFdI4PPKJ2IQMhaNlu4TU
aoTRMXTsipes6eYU4Bpud3EOnhiqRQIvw5KBqcrsx9boYPf2+uHnfWAiAejp2nz/
Gmr6kRdFngzDCwfQQpJHMSPxvukzZJB6EjvWmfG8n5ELobvEHzFSqyhn+VFIQGOB
MVrXhlPo31qWmoSXc52cX/38XOSOEK+7ygqvd6YIkKCGHLqsboOb3ostHTpZFvIS
4nPMYvnXv3+G+d0mJlcKU7CxMkvcM7xLQNkdRLWC8rmyTgQpt2zGAArofoL7NqgP
/BZvFNS3kl7lCg4/YOE1Hst78FGF4FYlacWc+vk3OXBSqqFsxHDy+V1XVq184gHz
VLLGQ7o833ViLTebaOHfgE8uQvvihL2DRxz1mtizKLwDhHZBXZQF49v1Gg5fXnzu
O3pwtw7nDSBX2kGKIAe1eq3cARAQLxgB+tVVK5D+qXQSyZTabGlhMTZZS2s1PaUI
yRs9rHFpIEsvpHvc0hXxgfNmOhdSOXJnpLHOO79VzW1wZ3utCmOZfZS8+n0YO4pA
nwF8uTkGwyqZA1QzoF3qGpp/IZv7v3nnVRpU0lmI+yX9fB0V82wS53Qjix0XD6SU
CkRIBGb0bfruU9mIBrWe8sdz9FauHmSpwP2bOJEQGS+XSfnMgNJlmIIfZ1AOLYAb
ukG+2iYC/CSLpcasLUUSbNGL5CBO4JGEajSF4L5ZElR30A0XuK1M27bB/aBFJpFm
7tgVaXE8XwR5o/JFlo01wVRja9AohrX/kvVx7CWjJw4WAE2dMTDO7WR834TWTn7O
cEYG6/44fnHR9L6wX4OmTr0MHiJsCMyRd3EEo8SbLgTFwrI/2i9QLamD3kqZZ8S5
BFk2tp7kcI9YfW2RwPjKsv88I6+g7i89BZBz0QyvpyDPAuOfiNAvhF7FYe5WtyIt
HAXOfogZG+Si0oXljRGPbgNZokYtRB2ayjiWhVtF0shAxDvnWLmhavQdMwjOFGS2
yfozutHFnKR05WUa1CI9mJcL+Vx4k3w4LHM4S2OBxS6B1UHZOGsTCndo5o49xWlD
jFqdjP8YbruL1eOktA/KtSpm2RCAOS+B3zxMnuODAwy6Jc9y7mvZlelO0tjBRbht
DJ+f/YMuYk+b+62L6GdVkEejWByfEYJMpChbxWbB15Nsb4nNv2xVJ2LJCo+R33Ti
w3bb9qQAcHfWz9o/8/XBb74rNrOY4obz1IrKbBBuZbMVHf27e8269n0plVFv27s3
1L3dKatKufvUXg28A65XoE6MG6Osslg1ObOnJqAi/tsHVo3lW+utgrYwH9uA0THT
2v6eOAFC42QQpPDom+OStG1nJK+rypzO5xZZET/S3jNJk8wNfQ3D1Bu9aZ/qIPSe
Emae5giY5Aa/jPGLsbZ95neh5XzoTDbbRsMnQUbu7QVHFTSNFyhXOF/lbFkDHMWH
0VrOCOHONSwu9hTQ0KMOPVGV4zvyLK4xodzMxYuHfvpcV32nRJXfr/eD4OLY7Vrb
XrdJJEAn/8+rTkPLdMzQ3U0ym70o5xBx1imrjfBfkswIMlumN7DlTQ3cxQCa/IGM
9Saoa33WwnrqQzOQwT/2ZxrYyCu0JuClGN8ve+lgGxV6Ch1m2rW7g+X5q3u9qq+s
mmRTvIbJUqFR505/SRWQ+p1aOBIswhOjKcI8xxHUVke3ZDue0F8ikDxksSTrdWPv
pme65hLD1EUtRe39jGewlYsKVQPppy/nMH0QnG353ulls79HlaGapEhyi/xJWOuh
v5aEJdtc4sCVR8lHfAB5ZlBOygyLnF5UhzmNBOGQH92qn/o4IJaHyHqOz8jbVqS5
yuVMhQTXCp2KsEA4lbVFGz3sBiubwpqEGMqjop9dNjB9w2E/3if9oYOzeWcxyQA4
oDiINr+CtnCqAvtn3dOP93PJ43W58XnoTXJv6p61T4LJA14LsSTQg31dpKkeR9Wc
oUkXxeSBNQbWbF1nDTufrqHi50UCgV9vNO/Y0QcTx5lXa7snYY4dkAQX6fRrfQN4
0FPeWl6DlxrxxfxNKgi/ac7aLqpGjehKjjnssDvjLe8TLHKaGl4AAhp9ScarGWTF
k2z532QWEJUHt1SLdCBV1HF8CKe8fKaCF1tcEarB9pxVbWyxs7s17uTVeOc+vzyV
TlWyBeT02GAW4indRVUSvVQItgwtk5xBx9sdn6yFlTY9TyZsmV/qEz521H2q0RPa
secrzxAQzAes7U1B9mkvsCCw7RaSJ/f3guOr57Msj+QnYr8pzSLpXdA3AUBCOgNr
7XLQTFLTSEY9hFDJosfUmknvcbSZw4UiBE5lEfst+q9gtWOk2aPmsSnIvu/UrF7I
T00dKP5FvOoSeoW2cNdXGa8Q0yK78ai3xAuzz6pmqer3zHFLrovqw8YG5yukHunh
CRCtIOBofz7D8vQhjrGA3n1YDIvAP+rPAmcWCCIY81jiYUjAoeKPO/RgK+tK8I4o
zaoSG9gsTQN3j1+WsrWJP70WYWPhh9/H3nALTDSXGeqjK8Ag/3XXk3VT7AUxBKUI
8uy9vF4U09wlt25NvavChTdEeMWjGNz2ftn4GxPsEybYwBZ6Dr4UMqRp4lJ3YbCk
NSSnZzYboQlftD7+Ls9P8YZylipAMr96wVln275HVYMlh4vej+oc1kaydEAEZTpS
7M33ehvgyr6w5M42lqs+aJSKawbKB9D2acx4rQle80nwM6I/jQLhc+xrHjiGMXQX
RtX74sucmshlyqZyZFfAIhlqq5PoHhC6UHXK1nfZkyioJjjuKBhmCgNL5Fy+txWm
1WHRdPcQjqQnujBkQNVNxEkYHJZhOZFj94icu6fh6iWSfMg4NFNvxfQ/QaMU5WEV
UdB3IgB7RlGC4MS8B+yj0GY1959VydTN/nW5yCMfH1lrOGtJWtA7LEFZ+TmSzYz9
/8nYGFXH/QNEFbEmqJwH9qI3ntFZv9EegA2yUdvSOP8KxiyQV5lKK8FBkih7iQ+u
1rHsQcPA3sU4BFYrmOZvMkReLsCjl+1jfAVni0CobhkIZPh5qQhfKec60CdrAwOu
8LvAzJ+jyT4E1NKWyKKaHKOnArmoIgwxApgUQAPZ+d+6HCCzBiyox/5nzvRMCw7+
mUebxFCEsEDuvoYdygeIraTbkvIBDeivr3ajWIxY/SoaQAnW42KB3dAciElvLJju
8hrFQ+nzsp6w9KH5Yg/T6FwYcwN7/+2MzDgpH6GmirFr4/+aEL62xOzUiHPRDolH
bTn20yJw9NMVBng360X02G3NjlcR68arfIadJM46fRAbva7yC0iR4T3vpHewRjb3
H5URBFBNW6/qbGTU1UmRh4Oi9r3gm9LmFYSOY8/bDqKZZCTjSSd8t6TB0fVpcQqG
/i+ukbyfY/RKb+KsNNY5TKlijfIsArI3fSWi/d8HOZwIkIuKmbltDx3ZsoLBYIYl
C0OXySxgrOa3FWjgeY7Fs/acxn5+Do8HRZAPaqEIU/BdiFaarTkXh49dB8ZnPNFa
NdctoESb6bKJ0FpTa/u7/1XSI9hxGU1Mn3eCIt5MiQCh6cAEKaOxlNa6kJmbJMlA
8F+cVi7uwhrtGgSUPmNeYN3MkMdgZR1ChX+q6lAzJlDNKnYHtX4VLN2Ft5NCrSSx
q0xNwqQn+YEaDXdNJ2/5Boo33mUoKk2vInHU/f84fPIBxBTCmOFhwR6gK9Plu5pK
lPj/4WYev0l7VElxojx50hQSnHbrDYU5gfHtWJVqfM1xQsihxjuPXrtN4uTDA6xz
BaXaopEejuTacInKmQ5BxSm2Xm/hVKX1+W2MJ38z2LiZK8cvpiPZs1vnGgsj9UX2
1pUUIf4hDlsv+sz1NrwXBLUB+LTWE6unC5GR5i7A42/43QYCqYs6BKE1uGz+i9ig
/zSqIRf1/HATlSLquZwccwzKrKVdHeTAS3XhXwYxqFqxapKXhmQtWTkWgdNwARZU
gPe7ppCnsfpHqcEwmATVxJ/2hJkWnYg3L49OxnUumYTPt4kloRuRXXssO3YnGNWa
XHAFyATugA+CrVnCzYgoGnvG5DwAo6rtzKLzazRajjjZfQAQsX13EaTIJ7Yd/RFX
JwgUsps1D74jZypj93h83OixST2YhmCOOLLtmt8qejg6T6sBO4F4y2WN7Aestdfx
dK2l34A/7CR35k7udcTzlkhk6LLpHevkROoH3DMBzFTw9lq5rULcIA2mdZn5M/4B
KLAaqMtSvY8e37E+kzEKuH3mXZVVW01bcjuOrO9VQCmhbAPtkvfo0tw4DFEh7ino
1vZce7iC0iNbi4RNsw5KJH+tXfSg18JVunSi6NnNsSscqxjFEuxMKUycFH/8Vy+L
CmuBweAa6TfTwuwatXQ8Wd3kouwjw9bbKBH8IwsVjT7RAVjINimzOVflSo3TbK2C
EsVWUz08bZJCZp69xmvvRxZRq0tFLZhP/mTkAnO5c6bCuPk1k49Fn3o5kZqbCNOA
Qgso4pVfGlkUxPSDcWFitbG4pxz8p983z3ymezX3ULetQuUeBxoFjLXRt6yzCIu7
4w35ay8ta3oMUXnskKY44o+0NV0yecFlaqsD7uV6SBqiE/KfHPy/ScsRsp4jJm9E
LieghrpZVfEjTF9KsFLPb9MVNlBM0SsPZYTuh+eKk+f1OY8nTEEfvuSNgaVNiy0a
2GdfC74A+NOI5XpBxPhmKhny6ur5RiY36xA0el7RYoojtfMhtyRcAZ7wKKrKsznn
t8EyG5H3Gxclf4QcXJr7byrNiiEVdQXNomNaK0IxgBreanxMDaR1ISLVGWhMXdz3
jZDJSnSzb8yqENch1pr7GJ+AqvSSsBxfYwaN7rNKUNtIuCVSL5XypiAyxFKUkb1u
2DBHjihJ+Y5/0yv9NTN903C5q4enuwmKQ2orISpK4L0bAzq+7bdgSHWoRcXU43Dq
Vf8k6gEFHxcSOSZd6VP2QbrlXhcugiqqunO/4a9jQMy/j+88AC0sAn7Mk9jzTSD7
POPBgAT8qYQ2cPQDs35IZPIc+qD4Ns7YB9ARdZe5qIOI90IX0pjgWcoUBLJIT2HE
3f+F4h3dJg3s96R5873jnjCaCoFcT92S/Mi8s6JXDKZ/0P4fKF2avpk4zrOrEpaP
jxWLoMUVPAi9ZD9bZccAsMjQM6461QC+X6v/a05OtAIPcwmxYLQdcjyK6TEAK3BE
e8D4yUmCUS113nKs+QylPMp3KhDHzR6KkkHGUUa10ZrJmarIj1PY4hFm6OjRzrpz
6JGF6xly6/Yedpof1WF5fGm08XLCzRJ4WjRGzTXbZhcOQNImjx8OJPBv8Fu2nKC3
h4syWknRvqCglKnC8aMPzZFpX5bUc8zlXv3SVlVqFRkUs5UCgjFg8nAce3vWIt86
HIoP74CUbrA3PYrElbvWNjrGzO14Vjs4nDb047Srdo1vYQ2VCIiRdkDLbHMzm0uS
WzRGgQal53x5L32QikHPd5Y0WyGMyptgjFxuCFHrH4KL1BJ0jUl1ptarwMIFe+3z
oveA/14F1oe70+1ZKIvf+WEESb/fQkCC5DSAlestdCKQU7Wd6QPLPn56+cjl638G
pnAXa3sMFW6nf2B57z+TzaWQySOvEjXx1qYiEAw+GDWtngF8TFsDypEe33gdpijM
hP0c/z5UsJjmW2cMrhUOtndWDLNjQ5nVZmegrbn7EN1CrjzlTTmybuxtgTgIMRUf
2p6kkar8kpqUUTCxe2ipH5mB32PuwALswW6FqVUHOdfCg4AIMv7LVlygKkY9q1hl
X/G/ncZoa8MWncCdzXbB8zIIH64qGKUpwr9zRyAYOE1iXkrWgC5d8gGMig9iZy5E
zAv4CkAy2aznm2lyretp87l3gunueIZ2W2WRW5qBHR4ea8w2KfTciUa5XpazOrU9
axv6ovYd3lKvNu3IedsTO1jhyVRs/pHGKy5HVotj2mwyEfm/UknTPgZzbgwAjjCY
DigFxV2teTsq/rLsglybsyGJTeJ0c2FcSwPCtJsWw1oh+WcaBPyTk+yokyvzVImN
a2ntbGahUVedrQyATSOgoyz4abZNpjGjFWOpUPK+6iKdc20ZqeSnQULco7du9i1o
3hbyoJrgPb99jB8AhQgdtETiLyFnMOstPgfGbDfd6tT5ate91cpVI8nGyOSLjjgI
f0BS+R14A+ZAtpbONQaeJZD7HRzgJJhcZUuksr0KFftDgSa8n48aJnl8pvFDIb86
9o/WphyHC8jtMDd1TKfNW9Vxhz2qkqwQECy338ZutO9lj+qg1CihXwioIBti7Q0z
QX9Ldy5uham2A6Xn2y3SGGPYSwHEq4AMRXPyYgcDPlT29PhEtQ94SS3oLQV3ot8w
wvBwOqxFmOKvjzzBVcnzEl3oLxbCnCY1uAxZo4cAWFx71V2mgTAMSk5putlb/0VM
e7Um0sS8HJMTCjbN/NaYp6nlBU3sNCXgDVQyaeAHnIeSMgd9MtLo0Lu0+f4unGBa
PK5Fv4i9O8+vwNIPQdioI7k91KEi6RVOfIlgxemoINUHYlsviLEk0fU9ZQ07as5c
iVOmNHDpJjhl8vbl8IZg1t7EZ6jWjaQpzdzp/OLCGgHLiCU8O5DP15kVyILEZ6io
/RcnNIsbg85CbPBvqTwqikXfSvxevwircs8xCR+8osmmxEVebq+aGIG9vt348Wcv
JtRwDFDDn9Yg+9dI7hFzlWw6fyXW3+9BD4YAPBle0lGEF92YaouECsVKmS91ZPNL
LkwEWYwMzAFi1R6TzXSrBT2BxdMC1b+RO5LZIJh1dAoDsiDCjiVuYD+4IjKgAeZn
jLr6KbiSSeAlnXjTOTCV6HyUIVxb1FNx+VVpUPz42sxNimGVxdcJ0cNxBfAekBlN
rp274QBFDrvRTLGtLb3FIfJDsR0FN3AHkhl3OG6phrd81KJXjNz/cPtdhN4YnmQh
A7p7NDCgmlaYmBISO8av0CrMZrGT+MFVgL9an49gnzMW2MDwW+ChCS6jC4O+lcUq
YVUvY14QtG9DPNsg/44BY1ilRu/UWR46WgI0RJpzqUMBxXtal0cyPcnJqObD2hDB
8ojbkcYElHg8W9Wt2To6A+FFhOhZPGwT9U7krP+kCOokdz+g4+CYGm7K0TER890v
shyroU7ba2laGU6igOmcL6JkyTwkNrAnSpsqsYYsMa06S9qkf8SKk4JdySMIL6x3
W6PnC3Nv26Q/Usnyq7awZSmdVHY9vmqubjF+pjyNZvYTOEpMv7UCpuGDZjUwFpfk
7l+yHFRY1c0iJ4MU4mgyhGLjXrQsI0OWm1eFDIQG4cHhu3VJggUaQRbwD024lz+l
xzuiOic8I9h1Du1LLkCCAWpf0QNg3X+jtPs0+4YQPOXPN22NI4NjqVJO/HEGhOkE
RmZn7vmlGCPF+U63/aDobG8bp6O3ouO8f0Glbj5HVyV2Uev8PtoXXWKLD9Prhugf
fCtg27Xisd6kd2dQSfkmH5iPKD3qbBmlBNCzQPiZoMqGcNesRrMIIwY1tEgcjciF
NTMh9zJckwbUi1ba55dNnZGgt+XPSpRA86yApXmr0/4p5ir3/BZSUTUaQNHmk81b
egXjEeCKJ91LQtj7qIWDCj/9DF+7ISeVbZCNRdAuTgML2+2y1m4L6baq1pW/1IMZ
zfzpyKF3rx9Ak5FJsbSXQge1g8jLBZiP8dCicf8Gj+8+DyIRhjIENs4fqhU74qJR
O/SE7LRSx1ZZvR8LSbTx88gFtBmqRfMdDWVkGj2yFEDlM0G2v9ZGNVTFsqXxsauU
WiARlDhY48/5+PQiLMY9IwW3sP+D0Wle/5G7gd4mOCo/Z02k/DO9manV7kZ5XnPB
MPXFq295giPASAL2eYtpemnBK28pnPqwrezGEVG+xUoPl4Xouyk3KMUKw9UtPLQk
3jmHYsm22KJJAx25qBGEm2CcEIUKYSyB+g9YPdXHLYei9fFzg9BfaUtWZTsm8aIQ
4sa/rmH+nkm6/gpnLgmH984H0c7ZSAbBu8w77NCtE1cTs8ZGa/zEMU/5odfar0dP
HzDf0onwYjdteoQFiZFCfjXN6eUppBsQxK0Ui9CyW45hp3cQydKlXyaLlMEREyCv
cPImiuAZIL2CUWS5ceysywOMwDAl/4g0yX1mb+kTpMTr6Y8eX+SzPld/JrLtBXYB
/c6xIGs1/EjelY2akheYxRVeOdJioM77wCccDrlHVv7bT9J8T6E09bZc9uO8hNEh
a1aJh2FHr0BXvXvnKuNtMnrroLLyl2Ta36/+sYtq5/jand+KFCbCOA5brdfGzYzL
g9jiclO990YhOuhrp4et6zvX7J9atdMo7f6wwqC5H2tw92Zr2l16+TZiebmWj1zG
bs+VQhWh8xRx35gZf/Eso5RIsiESkuQqFOpEVqNhfpD8Nx/qsR7DN6A+dIs8V85P
AsbWCBklYCdKxJE9CR+FbdvR+pZKo9BdVZE1cThu/OxExd6C3RQmNbzLHe3PwggF
fDoWjMlLCfOa7+oyr3dN5SbW8a5Jogxsv4DBNe2Wj3GQeuxeUvku15wPELK1KaiX
FXp5tiwNG8WyKXzoBCODpdROubEC4OWGFTG1zcTAaV13a9ddzXdr72IMPqdVmAsw
dLzz0JRXYlmkd46DIANDsHVxxKPrhAxFjecgNZobHL04iDAgtnceBUudQPQl3JK9
PM08W4WNpvw++AyAIDAjdd61yoLW5gQ+Iu+aQwl36Ir4s4SLcCdFIhLIC+mJMGBY
ZRw4kVwzQ9juYlHj/lt7jMuUereoGHO0GyhzJrJu+Zd90W5LNWwANeD0GC8zbdhU
3swRrH3/4GeT0v3vVybh0D8CU58jfMl7Rz1ZcKZmQiTmIvB1oKl2jUKQj74tO8b3
W3dH6leowRNzsMnjHlVZM3mo1r4jTYoblJJ/xgIB0xeKGOKJnkpKK9cOmazyirBm
fSLj1xiL+sz9CEtjwe8ZwAXAI/3y2k1DKezXxJ47d6q0LjW+rgCYh4CGoxx65+yk
bYxkxcK/lbZLSoXP2ToHrBXyMLUpwOJ/ekSIxfnuta/I1N3aARS0dXwSpYtaP/SD
ePDa7bB2B+gGhcQ8YIbazG0FnDkFEmO8wrZG+bw73r/ctwCWlv4x31GSHj+0kqJP
LNHokZ8NkGn4504rh3d39W97d8w3tYkI0C9zs8m7dkk30FPxLvrd9jV6D37TTtu7
vBs/+wMBoO64E3L+YFylInU85HBX4Aawj9rvQu73Sbqu3/QNkx6m4vQnrXCuIdSN
lI2oHAfjcQ5H8yznezmk4VhFaKzm4evf4yGaS3z4Z/j6OoZY+LwdrOk4PRmv5tpv
VblwGghcyYzsy+4+l/4JG9MB1EqLtXyPDYe7q/SehmdHNMWc/T/iVtsFZKRDcIXu
/UqKSMYeHpVoCKhpq0P7yvRzmUDOAgCPJx4nYAI2QS1agGM9BPNpSieNKHHRkyo9
8ttVSuMdMqWxgafvmdgAGQ==
`protect END_PROTECTED
