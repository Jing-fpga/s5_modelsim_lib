`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o4kkeSJTUW6DXKxKN8iFGLH2AtGuM08iwBu8o3qVhnRyczYAnTYnsz4iHAN2OoJx
RxkV99HUmMCf2CKaMRg7ZwRylNaFWQRsniT35GgOIe8rGXvdcO52CxfyMEOl3vDn
U4BFcQQB71/s+aJ2ogvDBolveHm0aAhwxG3D1+VM3zk6Pkyhs+49GtsUc6Q+VnEo
NcmqmLSwbCMBluIMR2x26LRqPG3ZPwn+5BNSniSbwH8NdNd8rnri1toR4rJspP5W
mhRe3CftSs6HphLgRsaQhJapSO7dVU+pG1dMGmcinraw4v57gpcBanvajl+cQQGw
Xlsf850/L7RhjZLSoSSQ9uMseHngNa5HSuOG7X7rnp9eN+Cn7zMyymXJ7ePxqOzg
wJODUcNO8Ho0mJTp9Avr1hRkNhGsNdOP5VLFE+dWMNoWQFzSFuSYAdsWz8xkKXPO
dpNUDgFF1BMXbH/3PJR13pK7PhldZ2H86xYANeTKCo+/IseCdXnSOEK96CLFw0j7
aYRkDlAWmbG2M8/LnxW3mtwCkj0i7hDzz/z8cnrRYvfZS7Y8qqH0MaArEynRtMmh
m7nU2zDusjQ0XRLm+G3KcsEX+/Rg4/N8M4U4VvzYFkX23+adwiIq8EN6ZX3KzK0P
Jhqjfb3oH/Fon98qdoEMxo49pY2G2khCwwA3momPUlAVwYGeTgcm5KD1T+1hnEOK
WmYy1vcaG1F/IrMFcWXd4diHKXNLqlWffK2YhBDGgWw7JXsiIfFUj+xDc2v4Itpu
elFDA2nIk69iJ06AMKa4KQw/rtjcZAO1bv4xVvWOfoKHfb2n1njTHsViEzsJwOY2
ccEuJygxfglL0Uxt6vPKC1ZCdbLx6sKfun48CAfg8s68sQG2DrlzlkXGrA29iBeb
n8e3r5dlEzjaay/ObWdjxqAEw1CiSlggbGj7Pbv9W2QGls4mgD+zbqdxSNF/qY6t
t68lNgMwIISRLeeYqGNKkszsW03bWYfaIS/8GzSfG3ckeQkz2itG27XRlIZgcG+K
iCRfUO2LO9gQvgbsayZjiPUvz/4K/bSwJFrbZjKpeqZ2RrPrIghnUWuM+ZcMJtBQ
rRcohWR/m2LaUTpWTpVG1xQJAmjV1HxqxB0yN9q5PuF7v/1EWgyJIzUYmM0eHYOq
x3dnuPTANFZTjOrtgKRf/6OJj8/u6stGGOzsL9L1MzUGEjcdwOrgrSD6iKDU77ZO
gnLGltRsSIKani9WZol8nQ==
`protect END_PROTECTED
