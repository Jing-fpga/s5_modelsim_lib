`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bnUZE6HP1TNHWJFd3rI7YWjjRFpHY0orAdd6iPlhGjVxbWyp0dPkPji0NAajzGKE
nj5/jBIjB1g/h1dwDD+wGU28YMpoUV4+xp4njDDRMgW90SS/A7JrKGW4j4dXiYdf
3iSciQJIHYyhnHlQAORr8qS26yZHbazcyJCvrXn4yi0eProd7x8H1h7LwNenXsMR
hzr8rTKSpl7Lp8x0C0c/KrbKZxS3MrgmIBqk4jbtSC80CG3Nyd9ynsdlMPxrcjzz
4OsSBSRPb4cx0S8kp/EnIOdikJBUi+mnuK7ef0WsDFXFGelpGCoQ7xjImKSU8ie4
h2mPcWzSo6GCsHwtlcWDAkpqOWUpwvFPcYozd8tRAsDTsEKUNQK+85Ivqv7ztyAD
2w5Fi3wuy2mTnDi2bBt6M5x3gW3yYLtMMfY0LEODbckzAfzrRjBGMW7U6z0GNBzC
EQ7XJBW7ubaVKzp4FU/f4ceMMpxnSzrPL9T+ID4OiObNPS8iv6vk1CdQmNOKx7wc
ZBnFfsJHULztS3f89PWrdGNkqyKE61aBaSQfnmsKr4R5uJ1zmXbC5L2ThMCXYj0P
9AuTde/kpvgzOoRDgWqGGuS5/5jLt2Kj2lzE4wkTnb6fsayfdLEaUrbIadtYEZ9U
Y5mgIAKQuddpA9lcq10TgZEpFxoVVZHD0KCe3WLHF9ber7XKZJyT1xZqSW3/lEYm
nQ0Ox6lWLQjQU0KPf9GiKOU3xp4U61JnszVikZo28GGifUk3abSn1yl16pLOmLLt
h8KWNRZ8vND+raqB5GzaymK+OBzW7nuFuJ9TDvpepEwCGBjbs5JLWPmvI8+u6Aho
F3rplQW/LEB2Bn3UToIDukZXm965cPVdCw5ccEjshfg=
`protect END_PROTECTED
