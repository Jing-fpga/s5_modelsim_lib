`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iI+7MqTiqpc5KqBivV6URFAc1LUfwNpWtf+MmJEqtxGhZcN++X4kk/07MDEVcfJX
hPLMT2g2/HJEmWZhmwTQch/z0bKthHQtoBPBRpK7we9luM1JuLazXXWuJSNdiAzG
5ncBSI0tXz640WvuGKF1A2EmYiXyWEVyRU/lsdJLLzaKZuOMccVJMlcjdxzv28ld
eKPgTb4FsKOTOrHmnqyo7yrzUO35P4h2DvkUrVWppu0htTGN+vR5isa2qj9PstIb
+S+ZFnIOKq3sWWzLrnTKpADs7KAkEudzO4zCbHRhupvxmRjmkc+CYoAsfRw+alDz
mTwTYBT0l/JbKzW4N9noNLwE8L8HPiuBk/3fZqZdzvBO9KrW4fsWs0PxWunLz+u1
ijvT7sVbx4QWkDt8vEofAv56w8OK+BlLSroGtRVje7vllVcghy+VdN9bUQ079EgN
xZw4Qq9wNjYLtmjF+kIJkP/3xSsD/PT6G+fanDE4/shHGP/iiTU0/WGBqiC0S815
zIRgfxoifm5lM295qENlcXz75KaCuoX5jPJFtnRAw6LkOKgfSr1g5uVz8LnSbbSE
6kxBrScOTD79TtbvoyZ6HCx/4vyAjyJJXUfSiu7dZdM9KrRqdGBNDPGM/DmVgMt/
5bGVFrpnMhrCA2hVj0IvXLG0mTVkkmKFyH11H9uNsNWpt0a1fmxY0ruL2bxZv3z7
umT66C9mOTJu2LlULbJc4+0DqBFruJ4DR+wOEQDP79oSUxAgWJcOiPdhX/UQXDAN
Ke38NqacdvdfHiJoNPm+iUSYN6J2cfoyDGbSIVWgLXvjaO0YOI6SKsLxRRG/Izlr
yCob/TVvA6CAY4KPGimvr5lKfFj73VQHpAoQblsRl6mX5xSCGgc9l9kT7yHaIGJj
u0DBsXx2U2km3BJdHbGl1pGKgzsD1t0hln0ZULOE8+sGG7ZFzZMSJN9bGMzNCP5y
Ci6K35eDV0GetQj8kz566/DQ/K+4+EYrRMMig0YkAiq9PrextK6ddpIjbV8ck0O/
cRmfnqLZZFN7UkiH57kKVT7wqhNvzjLkP8ZUOhN9QaEeZdK33xoWQfwgHe6YX5Ia
`protect END_PROTECTED
