`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ORDh0y7By2pVGa1FiIpyaw3iCFk33i8suUEJyT/k7wAVZibHU3md+lzDw12ergYU
j1bzr626S+Nvzy11BLR3S/LRC8SQ4/wHvjitqxFfE8J30vUEHpagscejXeQAi7wo
lzlbE2EwF8N1eZ/0RDJtCGpf4X8j470sZPYOYqiI7oFoZEvhekYTa5qFfpYQ+k27
uNuTPLsnTBI1wwm0+WdZdFWCVHijE7p/y4Ew+gOTgt845hectxG/EADxpQMhBKIh
yKss7T5eo7LK6QZLnHVALXUdZ11HlaGg/WsnUAZDOAT5ayLjRd5jT/7BjZuFKUCh
AmZHa6A2VENSJMU64oC2qCfnIHCib/Di/JmhWfmGmpUMIyBS6I3ahljbr/i49OtA
Z5n7L5spvXoPv8afZDThHWVm9vICIdQsqhXHah7irEoqE//Z2V7ih9AnXQMW8sf4
A8bRjuCzxeFA924XQsULKpA2BHOmD2n19NeLHA6z4ixt8BzG6q0VlmvzD+4EAKHB
PtCCbYz/S7v8w8VuvS15qAfAyMuvNANI09BPhLDmS2NI8BX6s/1d8jqwyQ5RdJWQ
G6mtwtIxdgluJZT6odMqNYIlxutA4TFIVAcyTvDHk/Z1tS9tonnwsorclhL6ZL8j
I/1rFGHWb2SFb2UDT1MdRyVk1CQWygZ+q/uBciz7EZWME9SZmDl+ko4cJ1IIPNgX
BZZsUO0lYKVxsadKxHQil7TYjLPC6y0Z2GSCAijDfKGqcVKtDZUxO8Kbnfj84/6N
9NNTu/V6jIhf/abdRe/xBxj5bqHF0vaNP61LgzFgKHy/rNgQHYiXKRyNpsE8eR/K
PzBQRTVL+LENRETwgag0xm+DUgZqEJjP1UVpJrynQFNbyeuU8ySkTuK4L6GeJwtG
9ANfWZQ7O0Cn6Pd9DdA1P4YsohogkImSMnmFKbTOa1dQcnORAG4BWkPLmnBoOT0A
+QWg4/fc6lnZqIauy+4Qx3l7r2p1UI96Go4RDCHiQxiRyjITV0qj02oYuHhG+i3b
ziZY8owif6Ksssh6JGoL2DSKru3sUexyZVKqIl8r2cfGoslxGZn7L1/1gykKWcp0
HfbFLPsCTVMl/a77QJ9LXnn6vRnCYKEvG76VJR1iqdA=
`protect END_PROTECTED
