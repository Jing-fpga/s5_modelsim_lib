`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rS9Ie2Nk27a+G735r7awbjKWrioawMTMuu+vQKGjcwCRW0n2jjvjoinCwV+K9yHs
N3ZuKAfuGuH3UWR6YLdcbfnEdly0gu8DeqcVwdZY+6/DnTHBXV7yN3H9rfd3lMU2
yTDAY6xX4blcLU3wBkkJGYIhXDYcGouStgHynvFeAgHK5u3mS5HlRov/66n8L3AE
GRgC8jvT2w+rDHx6xSqXPM80gbsBXuQ1yHru3cZQSZoB3Y/WafzTkRPZFZXcIuFs
fWRLJL1yw5+Ccg72hry0VV5FQL2JPeNnYL24rfup7za1nuMDVe4hXyLcM4HRAatG
AL5WIheEUTu099pjfc5sPRr0vGTY0rub4FuHRnZsAkKdESrGEvS4LfvTUCFQSTj9
F28GIIKHENLK6Vk+v2VIHNK0H0h8y1T1l0XH6HH/megMOVTrITnvAz6mse6wyNYT
Qea9hLAKnaH6CSZaQIIpMFeapp16PrIBc2PKveAYkZrF1QrgmpJQVYybHAFZgigE
8gd66RCTQkDSJckL+jq0tE/Fas1pkNyssbXOwGP4R/M=
`protect END_PROTECTED
