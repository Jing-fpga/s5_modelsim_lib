`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H9rBTAMUh2bGGG02n4ZpbCDbYuBfE/JDp/zTTbR0REEAbewCorb4ULdgkQgfQwij
Osjnfy8gGj6TzRHT8ls/5Ph3SLjC6zQQMAWGrgSFO8NbUueFIzh7WWonzlMjJGE+
nbotQ02pwVE7W2wKLVFtIQn7hkm5oak/dPGecfYfAakjYMmoDXcMAI5VCXITd+0H
9dSLfNuH0Oaz+vBdUZ5qgjF9PzMWJ4qseYd2IT7gyKf8du4k+cf7TpCdcGvqkRbM
EtRJxZh1bEcCY2QFcPhw/+uawp9y/YpSISekdaq2ZGAiA8e1NIL9HvP5/KItlORs
UNi6xIl1+dT/USYvDmHfwK6VZSAZDCabVzL2pw8W7NNYmr5XlKwEnibEzh++DshU
eQ17MTSOI53yo97j9JWmv9/8f+op2RKO+dIjbCMjkV1d6rcLgtfkOVf18nMd/roR
mUA7JIzy9qUCvsFkzD7SeC0SIKpSduUd0HrG/D0JCPEg8b6Utbuk64TcdSSRKb9P
M1olnZYA7xlV3s7lushSayrMTdBgSrigzKNAY5NDzzMFntCacsdsgRfCCk8lX/hH
/1fC2FX+qwIsNMhb1Qj5J3dn1fXr6DDiFeNMFhbsGd8oB2FxqpiKZgC2pb3ARDJ7
nSOALE/bqHdbamJ+8dSBr5EfiTQksVEW2OkUW+8CBJ/LA9ZVMF3BeqcL0pl1vafX
LjBjm/pIkh7DekutHVHHRmRa3LrZDTAFZmZpQinu0Gt4xmziM5+P1FVitj47UYhp
T1cgSdki+HPhv49EZyvbDeJcJzIWLiB39gv5lu6oVJPhc/eEVUj8HGKiPmwsrrrH
CAKOTHK8aX2kKSENO3tRb0I4RS5lZHt5MQtGy/gJ3oY7d4fUGtf1byZdz39idwtU
MBicRDgp2lFyAUIjxg0cmApMm8QfDespLkGDYdRZG/BFOwtBtommQUPPxMoJmSuq
VCI+bYdsqFD1j6uBzCkCpwRHZxLOIB8pvjO20332uKT5WsfND5diKXoU2+r3xtBc
67BrmRwFV4vAuNOID6dasSOUM8VfxCx9F+ogRZrM0VfIagxOt1p9DfMWcJBMngmX
Adxa+QETsMOTkqBQ8OLTzJorte/idaPxJzAZ+cEjI8SO1Er6a2c1JErpokvhLBW4
AiF0hCGMfYbsOsxWXX6lquCPFEK8nNRpCzmKhZTWIbbuGMVcy4rQKhisx/mPkCuj
0SZa/YzaSqMF+9WFdFT9F8uWaHqW9MXr0roUs9zzhkg2IY4tsCB0L9S40t/dwpBz
CBr5mXlMYqRpIlg4KwRL594oULRwXns12vUtunlHXdqD9t9iCxkVvqngvUUl+Tml
v4+MxvsjGxDo5I7RD+6RZP6Z51unpiJ/JvG3jhQy5KHk4bvWtFaVPgvUw2BimkFu
wYv/5a/lO7RkTl6hMEBPHYBNVoQzeQL0s/Bzh+NUPXZot65wbom8lW2VWiUmqx+m
9rfGxQGg8ThCQFc2GxSbymn3mCB8uD5gVU415nDN95/1NMFs4anSab3kKRCNXUuv
`protect END_PROTECTED
