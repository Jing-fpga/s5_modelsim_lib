`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NyUwQ/1j0qNHIHCR3mcUkTxLTHdfi5+erkMToLmNrXglnHXqvAYscjm1+Jwnse/u
+JpkEsg/QNuCrYZy9wGSargA8P0iix9jdCCo+tvL9ZOrfnHbyS5PwkkOzaN+lYSe
3bGEM/Wp2qFSALhY8kkl4428KR/gcmYtQMMG6Vcx2wmsr/TmrWpW8hac2usKV06K
cCMaRZnGFdb9GgcY5wWoJUvPzOGXQ0oTbpqq0dX0syrWyS+SzE/2+zMHZf4kayuy
2UhFN8zarHb+oLGd7hQ4vN2nF0vdGJRSIn0g7lpAqJIlxChOwkr5cBNGvbFZEZe6
MjpNF/InH7K04l2hf93x/tWE06x3OQyfi5DW5P9M8pDXwNlAPjsGDWfLQjRQVH9s
B0iqU/Xz1DO7N47AsBOZl/QBX/C8y/aOHJ/XkJgNgc5MTGd50T9wj9zBZEx980e9
DsZHjPI5lii0FiLZOHP/Drs71xNi0J8fvlmqg4J4elm1nyrCSSY6F8JRn3XRshoC
aWi6tJBfhg+LbkRIore8uaglx/NGRUdp1LCFuqD8rLSp2Ef85EPN9cm2JRLec/BR
IUNQdzCIz77fCwDzPq2c9sVp4q3q8EcBjAJJ0LqNS7YKMHvNxfk/WAkJxhxZ+xUs
1WBHC7WVyXi386TvCNmpXMQEZcfpuHgrzWIssDncB/GD3aQjBBPIIM/Xs9jmchM2
kxTR89taN1WeGTe7YQXCe5sYmbRm3knLKPp2zHOsGcRHr5bbEjd18xvxMJvkOPYY
354o/BGFDLUd5JZP6mN1gJBiS3C8fTpnAugcBmMrvljxyslvlYFcXLOvaKIO8mVM
AjmWZ9zUUrWiJ5A2I3EvosFT3sh8b8FxENcHk6BtcfJcHwrr+8rwpe/M8So2a2qC
0kwVbWSixV2Xo4bdOpMFn1fwiVEpATiGBHH7UwUk4dxvf7SgifAZEUitIrkSSsfy
/QgNZyhfnY3FraBwzOgzvNWQrzknPeikx0VZjaYjLvYB3l1FDZq1kAyHZJaAoHbK
2C9fVc74wVoTJNJq1d79126f1+Yzv9vjJ1dtqGpbts7RXTAvPn0mD3wb/R0Rw3Bn
dAHa4bRP8uHhqkfUj8Gv4AM2khUmCxTrS1LXGq8G7oS1PyQES6WYUX7B0vnKtw7d
zi9Ucu6lM3UDSXrimazNKtv37YyoQJGHjI2Jn42PnV4upGVCpJVZDis9o+Je3ogB
nE6h8o1xk5SeZU8fvfcLXugElmV51rZ/0TFNFmMSwbWQulsm3yZOPHB+Um4MTe7t
sQpHOJWfjsjeJKcXzI/ZcF0EB2qxfu+AmZXH2e6Uj97ZJz+Aot06lrQuFYojQqtT
G1/CtPe2rsJDxneYupb+34GCfJXyxdpyyXbBM2YaCxn2kFMxvVBSIdviHyJPP7cC
iNmeMuzBN9wZ4/oh/IlVtFgw8iaBkBtbXitznUdLHs39C56auUf24PMaSQbXEDUS
A5lKQkcij8nc+NQCQHlZ0utvtecfF9IaScj6v8LJiakz8LQtE0am/rkvz0cFMSG/
3mnTFux0z9BY7plsc6xvy0sDePs8zWzApJaD427VCKWnR6pQUrJHU0/HuVjH7Md4
vnWQKUDAsuglvpejAvL1Souh4HTRylzVvmq+tkY/ARrZsSawdub9Md+exDUIV7CP
jdpKe2MqU7JJyTy3i4MpPVsD1pxfMZosPGoLUyUUhOWTjX+8pJyhuLFLhzo217Uk
xvCcZhhtYDYkMrI84oIlOZgId7qmS0FX4SmKlWI79gzm1lQxN23Nn/0KcHdApx8t
oJTbSZ9M3Mx0Hz6l1UP8TQUFqQexX88jnaXl47jojdwusXcZgQstOoObBxI9npX1
8nwX8MEgavnzBeL11mWT5ah8ROBOECaiP3yT4fLhLnLc/4sbzfO5bWjZI9DyvKcL
HK8yG3247V8nmc13SCAriL4ZHabilnyeBXexwYtTSfuXE/eRtNt2rH45XiShxuYL
elddK2dfbvuFB3SxbER8J4hpuAsq4ihWpsF2O+y4RlM6TqM8s/E2FErEJFLr7sYt
nRYDCC7eMpc/AOxIUUDJ8XvqmqNq1ijrgXSWF6BsfQWj1X6eJsPST7gZiRc7liii
6ZIUDQmVUdaiQgQBnZXT9YO/LJjaXN5kuSyNGjCBVBxI2ZwIe+wiudgheX1iYUDm
O6qa7A2GAy0Q/X8dchOqsLA8LUnLwZggIsaVqavnlVh14vQxJUKRlCAp9RBxtAv5
2v6n/o1fKBzAGrB3RAvK0Q==
`protect END_PROTECTED
