`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8u0quPDy1bA/P/e4GJp+yi8IxG4/pJgLZdi0HmzW80eYiYpPqCi1GXqDiwaXhVn2
wfvFwbDV5XphQiswK6iY9tYD1+tfGfcLcE8JVi2d5jYjJKz2VQSMegRSUSFxAgL7
Dmx0gpHqqUVc0fh3oVSXAB7TeKVh6rUFGRFPOa4gMBPxAmvRctHebJkfsClFku9/
vnE/sgBiZIS1wH60vg2cu4vcAeSm4X5TLRLMqVYF1X7R/C8+D6/sUkyg7svsIRyf
Kv9BGzJ4+NS8jNTCU52Jbffo7PJiE9Iv9ZZ+JBTfgSTet3R27L/oVN0v1oor5r41
+/sS3FmsQ3mEsp0h/TndytVx3xG8K8hv76fzLSQowqKC0+pM9q6PLCKvsI7yKR3t
B58i+9J9qbcp/FbYAoAmc2mC6g3by20U/klB8MuZ6L7D2dAc9y/vguna38B/RoBg
HveSYqAzaTQTyX5ah2AsC3QXKpGHZ68yjlS1Iu1OguR8PkwHKGwzCdsHNxIZTFlJ
lpYninj4CsRYmIw3YjqpV+IvgeLTJtwvNU7Hi4BPzFTPkyETbxZd65lhj5EZD3e+
QqWMn5K06RDTXA9hDPFkIK5EzSmlIw7r3sMBqRvIfJB5p2zHoTAOK3Uh7/XTCbLZ
hjdEjAxh9SJcrC70HiZkXv2puSIpJffV6Ox6geX4jXddIvinO8/VWF5sMPlVn8oW
nB5KkVQbqAbZEWs9sww/JPHSHypGBJC1hn7IEqFCACh+laU3UI24MO1jan4Wiezf
qUutskRIy4a5+jkPepUKla+pHPZMkhWcHH6LZ9r04mJcUo4dDQp6HsDvt1to8uF6
PsEju1Yh0MOum+4efPTy9RXfmDdRSRrrVK+wAGEK5QsQS0vWVQCoxshwaqe9nGZi
Rg+Z5sttaJDSh6GC6w4Z0XLTIaqTNxXRru7m/rXDtN6imHz6TSbvRc/s1DYf7Ov5
yFcjgijePwIOWCko9Mip+DbB9MkkxgKxbVxaRWEXlfTqhAwM0ljap85elVCcdOr5
jmJ1VuikJKgTAPid9PQhANMXTfLOmzW9HhXWPFkblk4Vss3zuipgQQ8bAyixzl+M
Bw7Xy/5yo811aibGRIlLQF79ZfY3qPr9aeRR10GwgAot3amGi5ozof8s1iDOWKWy
9I9tuW0/OhfPZ0ICcML3t0gMwuPG0hm0mUX4mwETfHXqrDTy7OB82fYM5F58B0Sc
Jpuu0Fm8f8ZgS7C+1Idq3aM0e4dXi4CFOQVeN2f4PyWxq1G5ih06tmZtqPL9qJfz
3Z7YDeJnB7d1OLHJI11jetE+Q573Okt8v7foUbPhZ/tE2AaE3UGQEM2pMRfGBljU
4z+q5WlzSM+owIA4Xid4/Xo+fJTaunUJn+PiBOW7ughYaZ2Wh04Wmva8OyUJbC6X
DdBTbLNJZTT97zfJ0DtjTOVlfcW+FuPS+S35BOJkLtOZg0LVJHInqBbuNdoydXnx
ucU0mff8fjKBZriniVzDX9dO0sjIR/h/ZEx9vzrjqM0qlwAvv6Ejf+FkQpBMSLd7
yObMoq3eng8qHcKH+mG4dw==
`protect END_PROTECTED
