`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dOz14dKsE/izT3r0BheGDYsmeT/8CT/lpOf/nPmL/6CI+FF9qUQO1PO/bCM9PWbS
+RJbgGgWPo6tIHq7EGT0IH5/wOn8upLEo9gigNAw9tDBU8GX76GlF0xb6rP94OMS
gcTrD86TWX82nT9QfEpLzn1VMxxthUoCDYEwe510N1BOtUezOcqE6zag21d9ecif
qsg2KEMt1QdFgZ9qmPoxKz7iVUqaNZm0w5U663I5H1ZU/QmpAputJMVfhQCUSc13
ZLSexPMdlq8LlNbCcMn8S9xdsla1Bnk9M7h/q24S1dsUfyS6y/LCIx9XGoCuiWVg
T8u8bzjrjHkFAq6x06bXSvhOu5umx9yC2Yozs4jNFb8T7EUDVznHlEUVlRlheOXl
h+XCWdne4NV/OYdVOZeiODyt+jqVfUmhn3Mp1sWCxv9LxxU1FS7nKUMUnSvBhRcu
bBBFcdRilbvz/I4XvbmAE3aVrOBp4borCkWA3iRoXFUUiST+jJVNw/b8OPz0cSqq
gEbRStcAFuyx1IPyOFkW1yrYBPh8hc2LALheSUrUJ0DNz0WZ9pv7DSqpacutdwHk
qmxU/Ao+0Jfhpw/fAw8XSvyok0GknSHuSktukKcYmS3hFrGSVv9nwpYtgn7MAKM+
Zj2d9ZqCksBDGKf+wij4DEO0RPOyNItdko5x+dPpGDjbcFFddSgrIG3Edc9O7x+7
Do1PzaisnKIa85AWmw+zUzHCYgGD7dOOxPWLwOtVitV2uCyUKj1gzmoK/46GlEKD
h2WqHPLP5+lYRqeq+Uj33xIx+bjNC3VU4UKzVez5ToBBnr/G1+t5d0zAE26V+NSC
qnmWfjTP8uMOHRfoh1PIUos+0vEnPiwZ75L6GHP0QpaF7pEc9cpPURagsiMLYF1h
qGj0XHAVPLkzClzs4GdYL2TRaDKqI/tz2b5zH7iHys6EONWdb78xVPQ8nHBzytrw
2pv3QDpKWeAYjgZrYbCIRH82W7FNM3Oe1IXGP5hyfPwbQP+4pEfUcnM6x3hkjPuG
EXXJCbXor30bshcoNLF0n7B2cJk8/2m/Py6k/KFvT9efDRlRaoqszUvkznSdEnvy
hNTAAkBmBL3LeEOoSeRwvPxwrO6sRxNTT5rOnOMMSp+y4fSosv2dTmPWmkk3PLmS
SxbdPmEq5tJnqShgjyxF7+Sv64EH43tvZVgsfgPEZn1T7zoT9MAjSVh7F9+9sAce
NouBkQFiLP9rpu+Y3xuabKwYGSVZw0/UxzXgFwswcMu7QN0LkO7txIdlqjDOrbVg
dNNHaHH+t0KGS60LWijj311pfAwD6vuhH4+uRtWKOFSNcS84ZyEaBgEUi6cohhRi
5UiJYzC/OlaQ4cJRvSLYb58Br0ImuNkUnepZcsdyoGOSIXuM9F7ILtooMhdzUPsG
OcmIOqZH93tBV8aTNRIhrDMkSFqUG91JT1sSdk63AU3PocBUOEiNEbQPqj+dplA1
UCXNdXiFvpUaACxnve/K2g==
`protect END_PROTECTED
