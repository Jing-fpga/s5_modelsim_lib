`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HbUjh+oJ+3NQdBzyPnXjpHI9yUUp9PXOef9qU+omRkeMekUq7f49w4EKqkjUSqJL
8cadYXYEBaPwaWz0sfFqdIMbCF2thyabd06tkaOHh2Zj6LBRFbwb9DcwrJyWfyEr
z+chcRdMOZLvBQPtsCtqPyMxAnylDcHrgqU425uDfaQ5Zitxeva8CS18xbBTtbT6
P2Po0noh8etj9XVnIEu+hqJdt5p2poXQnJ7XtZkgpWGtk1Z95agYCFZoKtacUYx8
aJDy2SBuRwyQ1v1QqO20yayvDj4s7JfBOaQNymHbpdKUg7sje0pWJGG3e2PKXOWp
/CQAVQVHeZWKaM7r0Un4IzkFgvFCUR6Vvg532VTuCZeDTXORBPj2tER07BTyz0TI
GuLRPeqZgsZUwNtII/eyofANH4i2jNj+QeN6qqlXvSjdNkR4rJC2W7RyGkTuxIVI
nFzS1eAe3Zl52Ch/htVuiaUeAv5RSHHyhcKzxld3qPGmfG/OQ/S9GdxnWrbGcci9
pReekc0oTEbmVDRF0OrjypddVxc4AxEtdJEmI4nAgTq4xFH/s9UccpdKzo8WKaJ7
9NZuyx03tjPkRcWW+oynTYF+ChKL7vRnetIGLxeoqgJPdzFuUla6tCWql0fvzKpH
YZJ9W6M7VLd0/HJ3kqwzGHy4HlOT6Zf62eVdSDJevhhV73v2ezSYqXhDJSkoM07T
XbLVnulCtk7zXPexaHGFC16CBgNEoN9xncJt8NUozJbumMrq7gryVPeemgRxojfm
Ew2XWJQ/HC4s1iFNIjC6y26fToWqF6DZZMuSvzPRh2QKv0TD3JRcSDyhHGgUcPcx
`protect END_PROTECTED
