`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NRSGEH3MNAGmGRTNtOgida+Lpc/d26v7ZXCy25Kxh4lk4Xp2+ksRMu6QGoL/0QpH
rRycb2/ytbxD+cSUt0Sb92zRL9UPd4OJ31V8qaH9Sf+uAWhy4qBqrkaet3djo7zD
iRT3WBpGyFuYhqWvGWe6GJVutpzWkd/SghFgKQttyouE3bnW7OHmeLnk37WRZGTo
8aGz8CzgxvSHcD71NW8tgsWGTjHFQLg/LvdYzQju4V4+4Xlu9t3fuetbrdNmLkSV
IPA2c1mCT2yNjJJjFR//flU+aE1uaabpjDoZMLXtFgHeOMuIcENX2AZPWv3i531u
qxTxKUwQ1ufnjQrr6v4fwLCOJbMq377FRZKMpmpr1R+syvgRFV/vPJRcyfFzVUaN
wk5pzNOCnSodPxAiMqOTYgOz5T1oFNdhmi/F+o0ezoK0Nwtip5RgDbYtzf2qgm1Q
iVeOb79eRnR6M95szt/L9Mzkx0DDJ28wuV3Jq5j71pp5rMyILfFDWpHlDxDe0LMQ
Mo1F+Vgf7RX/S/P7WeNRACRyUwLH5CyBqcxWE2n7rxv88xBs34fQR7bpVV6RdOqF
FwKtrhQUymkBrt8K6OfB53XIcHlps96cSP8YTCIoB6FcRljSkdnX4kVfxdP3mUtr
+gqeFyCWNg4pdtaPxcDaak14RX02UHqRgevgchN++704kiXv79V42dQ5bjzrlF7E
P8q37I5krXh1KE/OLQCsXCSBzQsTuSSy+7QY+EBaxzW6pA+OxOwj42V8Lp8McYp1
VfpFJFbxb+rVhlTfhogR1goEBZqMB3tTEjeb0AutfyVK/aP5kmQs225751Vd6Tdu
e6bEWHmcswjopyLfh3/OcULYS7oz4qcSkuUknhysdb6HETOsDWR0HOeVJdR9q9CI
QrZ+o4fYsBrkWLk7QJYaFbI2xLG8RfKsVHk5+d3gcyODvpXMAwlrHHMfpBrEEJJV
`protect END_PROTECTED
