`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pkeHPtlvrDITsUjnQDKrp3vv5OU/XPi9DNA6yXikSmB/N86dLEKfc0bOgr3Rjmov
kOFA/h0+GtZFIIp5oWAFsvcP85tpYMCL5Ovuyj7Ovj/C173gEnJlC4Sj3rw3nmJH
Um1oi9RMErnQPJGnHDQzLr55VozF0HgwSQRm86PO+BDqmWbWrCzy8hzvVhvOmjRV
GQGFoUbSrmQDfTAwn/DHfM+Tpq6b5C4dNFsFfKdGE8/I7aNRC+C2Xe7MsQjsRVQL
Y1NSgp5Z+6YctxVFpGRaXfVapXuIV3n2w8iwQ1a4O0frtiz7gu8HYpLj05nzRvMi
EjNky3dXVfORbUfTAbhzSXYuVD9Yb6c/NNS9fWhWaSlcjIcZOHiJwP8C2F+LMQLo
5JNaXiELHXP95r7xhYYYlvA23HcAjDLDmSlXbe2YLT/bndaN+NQNniIsToNQTpsG
oAHTz/S/QCYK9zahR75DDS4jRbJ6tyYhtJxTmXNmTMy2hwUbiY32q1/lGdqIKSH5
MImmxYe8AsCi3e6JDxDyy+wGryReV+UIKnUo7m8UWbee5VusqD/YmBhHj7+t6VSe
U5i1GECzWkymkD8ZDXLV8UwqKN5FEMWsvfT0AGn8FTI7UMgkd3tnbus8I+lavTBL
uVl3y8HD1dvDAHGilQLtzOP7N4+qetlxtm2/khPDN84=
`protect END_PROTECTED
