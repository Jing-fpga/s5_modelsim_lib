`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QelNe/TREqU55XTxnZxcuqWNAPDxMLOfPrH52pnOMh1La7Y3GZOm1nK1moueuLvg
OXzDb51JXNJpjlR8R0MSLOFquZovtXIIS885OtVLWLMV20dr4TawNFzhISebCtvq
j7ji6ZLOZkPwBpfO+hVr+yWL7ipHDEKNtBDsvxE1s24LGcuhWpj93ggRJwtA61PG
CagmMzMmNg5ILfPanMTHPAo8fp/A9EiTT+ktdW6mRL0qipcaFlTuSSA52aWtgEEZ
9MZvUxt1PsnJK/wboYqmNgZo4qE1JhOAbcSwttrZjswlUMrcHcSk7PeB+k/PwIkl
V7kTBRkUooUWEdbjqXfUNQwG+jK35FQAq0tvixOtvkwQac8BYmhvYHG/t1umgX/V
`protect END_PROTECTED
