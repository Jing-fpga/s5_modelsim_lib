`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L+Mzst+RKJcIAK6I3VWOkNbGuHRBKJNG/VfIhC/2XyfoEQwDC4SbuYgq3xDt9nBJ
ywFEYNFCOEusNKECPXoOLJxnQ3QoI4yEI1vuB0nptlrq/mQYmkZiIt34dNA1fi6s
CfycaNz+E0ku1d55pqsDK3BRHf44kP0ZhTC/0ihQMcVd2X/EK9MASq93INqbyzaL
C6mWwAzCHqWHWvm4yjxTz25dtcoTvySQQi/Kr09lwK1dhd1X6Ei9NWHlNEwAsQw5
oT0sDZCgS+EHaV4L/pZmjDOq5mrkcF2+3MXdybY9y+SGtaWoN9qozAESAHccOQCD
SdRCHLqkpdi45PFYgeH4va83hwX6sCSnFFLcvwq5JvvWKogzCjLNRQVck/rod9oK
7K59Tu5XL4izUdfm2NKlriFc7Qmne3cuXdxpwpmj8HDGBKd2s5RllBS0iuDNsNG/
7Qjfer0xtwYs/UystAG5Zzt89MhU8CIYGieHka2L2IbjNsq46b7cbeidxz6SVXIO
GJ0jpx93mUQI/bnv9Ww8v9qbhl63KgX9bWiNqFX6KOYyNvkDyNi1ouFAGt+STZ5s
4COWlaUBmr5QgXcxyeKl4NKVo3OzR8qKLFkO6IKhYQRAPzDPSVJvrL6J+i7sGR+V
6UHdD5aFeTvOpRih4jM3hgxCRphyCotT8ozDHKeQRaAncVjWrA9OV06VUhEmFutn
`protect END_PROTECTED
