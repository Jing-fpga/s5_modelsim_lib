`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/XFv9r0ads8JqOx8qCQVeaUzLR2ZUnHs0lNmTTeZsJkr/7UM2/0KqLlvF/iMQtfm
6nRSgzqn93pcADvaRey+aoTozrELygTtMDfOmwHHh80wLATl+2AYKSiJTz7aGHyc
IXbcFrhdc0QwutSWnmQU81uZY0xba3/udCU0cKjrW3mnAWrvamhS/7P9Rn3vGfri
if9aHLEEBeA2JkVKuiuYmwpyimlMTPeOQ9h9qhpFBr3zLL6AksU07JxU/wI3vR2L
WzCP0KgL9wrWBMu7ZG84ayRW3ZO2oWU+FCk9dPTG7EQX9ijHgVdcxzdH/5NJ8JGP
wr3fty52qtyBmwkK/N9ABDGZdbdsohSHOjE4mtp0ZCKMSE5WqGj3XQ23WD57guml
UpHxU7hj1w0NryQdTExTb2XbphXUUdVTfglbcB1fJMspnIsCR+/OpzB6Tm+IQ0Fm
Hf/HdrLNoSfcFqDFa7JGJQB7Y++R/M/MDypPpn/LhStix4seHL4mdYQKHtqYVxHk
PtumbM8x+8raurAsodgiBg==
`protect END_PROTECTED
