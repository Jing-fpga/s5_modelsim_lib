`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K1vBEhU/zzVXyYeW/8uHQ8lAl+qBSzCPYa4WNU4pSwMCJDbZ4yzr2lseVzJBpFza
Nu7XznYbQuIUqjKFk76zf/aCf4Mv/Uk/Pnzq81fg3KLObjLu47P869xeWduCf/OU
ZSXsmwQTEtBsPkt41OAEkrec6X2fMkaznuLKwsyoURGNQPag0RfyslBow8rsJay+
UYqD/Z7HR9lGYjV1c7edunTT6OblN11kexthAnfudB9bJ0iuloMluQPGgaw4GTm0
mIIPPCbD2PJzcPEkHXOygOC3j9wr+k649gzIHsgh4f4LMppMwDOa/Pn/UG8o/NUV
D2EyuKyTKidIIerBfXqdB+IR5IO1OUSCyfrCfi3C51lT7b+Sq3ntou3aIFLBj6xB
Fm/0Q4QyTJ1b8x+oSZPScOakbxRh2/vGYIyD3PcrymRziUE+0Gag2ZECjhusYcRS
XEBBdUX81etFctDXbPot3W6mSkn9ErOaadJ3qsM+RsX9JEhAL5bzAjxdDkdR7eu/
Js5l6O5FstMnTeyp/brgvISvAXjNg1csPV5qUu7Tc6ADIN1eIs1LFAwlkf+khVCR
5eyESVOyeuf5KmpczjiylouABev3nSZeypdJkHVHhtZaZul+RK4fv82Hb979yDdD
H0fk44hOF3HpuND5/8mMQNq2XzN3HqTtcGz+pOpnbG3c3sQYT99zh6tKuO1uky+X
8lEWVJyNftOfeZWTJ9qmfSjic/KxPMnrsW+IDhsCwkfS/tqwCWQ4GZonUO0L0/pE
Hcac/a5x7Qvqw7SvSx57XzMe0T9bMb+DYPkLT4LJ76ccTCWE97rHMeIZUoNZ5nkx
QQ0i/Tpl0rSimcnDl1GdNia9T7dyZtJUde4fAOxz/FYrQxoB050tcYm5yGAjflzb
T1++XWFAqwWwggiuNQdJ3wHtIroVruRez47dE48cGPrWbrpkL91rnWSoOZFPbkFr
uo4Kb4/Aat7Wk/fbdr5SI5tHEYTUDePmRE8H0Y/Ax3CahfNoApf5zgudJQHapvcM
uGo/39YVGEOoohaNlxLg/BW6ePDBJAbzOxkYfhmqJYbrTuriWQXcGVpDoTMVGeFn
9BGGkRoMkgSDuJn423CUPqDiGJpUCeXCM58l56Avu0sD3Y6jCgrYGkrV9C4Jvs0v
+HhajU6y0L+2JTq6G8fxrWBkJG1hZP7VRqX+01tA3ugozAxKCs4ZemMwYuwhU1tr
uxxipwHpZtWSHLmAzsEy9piaCmDY3Ep2qsM6lZYcZ4yVbszwRS+pEuDMz3hT4R83
BkkF7hfX8s2/L6+i/5H5HvMjztdjMUNi1b3ITPCv7Y/cdbWqyeIFoF+MFKqZ8v7k
VU/ugBeBPQsrn47pGugmv/iOMwcp8kt99RgFrY82Lwyh8+EHylXfZ984J93I8cJd
eVL5t6IFLEk+2N5ZMpRg63fSi50Eb36GUeQt4RqnJjHkynfqGPfxI23A5h/EE67o
LYpBYJn7Nb0owbN+E6C4ETyFd0cpoQL0sHq9uubOgqWbyV2G179kEKCgCKLFZfd9
3qMJ/Lqamby3w2ir4X+nzZi7BtIkTwoPj7U+YurP7J3nPkT4iWXvzS9IWCx1kCWr
DHHMfo9+MCOhI6m/t+xvwPcBxScBX7slGEa11yMtx/CBGhsa36voZUaFJLDG9DU2
1MpkFn/orLmY/tqZOHW63CEqprf/KBR8rbfGfEKkfRcCOEj33WO5A5xHH39R2Gle
`protect END_PROTECTED
