`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8CVZf2+jn/aFBbwRTC9pf/PZpPPCt1IZ6hPbTpaGw2b5j55NmfTRROxytcpvZnQf
meCp4zTxR9ePaBdPmv4kolxT6QemRtu9NfdlcOhY9I0TPEtWeLHu/oTYDJucn6Kk
f2dDLZVliR0bTiIaQ6tzLiduvqBZafOQ7rRLoAoJ4S09/c4K9Fk2HTbrNx+j/HWO
uNdtywwfqoPmmSZW2ZPDn+Kz3cW2dUZBQH9QwJEIFuETivanHRFu0o0U4arfPF5h
8erUqr7PZ63L5YEFBWb7vbKTNyXdVGj/2Ehg4hfek0ccHMN398jH17eMcK5VfA11
I4QtB6AXPMB7ejl8/p99saetybAXhf7OBz2K0tP9G/67eVALXpjPhzN5POgaQNmN
zvyYqDTEZWnHShDiYMU4ooNFs9P7BOwRJcBaY3PvLYTuTWEZV65moUTyGPU89YQV
KOcRFkcqizbm2RYXCvgBx3gcvDgfCfD6e9PappSVqox5T7PL8oUzDi7CrA3KjEI3
fecPmyPPLOXnOEf6n9/JEQVAMQyfyPYtjnYcWuU8ueac/KFR+fVMJMiq3x/NyfuW
1+5eg0CcnWnP/x+53DYJgLkeOX93sTnTFx39zujf58eUhrBfownE3hYCbr0Cz89l
SKLUpaFqUh4kBCA7WkIsmo9S7Zn5pilE9zI+BVc0/kW2xjMG7omKuVNM4LyIoHiy
NWCHnk8BPcUMhlBfZwTcUD76QDhaSiBTuJ2PHCp0gs2OYyE97aIFADID+9xqHz/c
FcAgmRHqeSsSSY4N3hCCGI8EbgI032/F7SXg7oIPd214SQms9Y/MGH3RPqyOlYzK
9qUpG1YpFpQQG8tnNA9CJKE+IL3XenbdghQ5b17jI8bFHi93+Y0U969LiI9bNSpy
upnk7D1jsQhlMgV/cyVdoTyzdgokzz95PloxlBqzvmwBBkZ+gIogg2p7b1XStGx3
Xtep6PKjNC+e0ofs1UaMay2V6+6To5UINwNSoFBK40SDFU8JeFLOiQ8bI+wc53Dh
4IWnD8xMJJACNWWsZadBd24xzi/jYFVmZHqhk33Urw/chFk9JHWGln+KM4VJ0QSJ
0k6wWRZH4Oh1uHNaTo0yCCEt8U9o2R9b++CRzzBnkThxIpqYqQDyaXWbESLZq8jg
OoB0LSjOSRmii5BsJkSXXNJLjt9cWPHnCQV/mktExH79FijM7E8EzfdrHqyNNVq+
A4k0wDmXvP9fQ8C4yW5Lk28CFsYrp15ly39FTsmFM9ATMmoK1BEuaPuTyKQY9RJQ
+/wmP4i3e0H+0l9zo0DC/E/xbtR85EI15FgSI2/AmDitSWOHq27xRurelhgBtIuY
sdE6UPOCPkg1CJrRuSiIJv9vM0V0wpvXBTBzH1GicMKIIVxz4pJL7myaZW2VWdQT
YP3FTkQjIDBcUJoKhk0yWM7/uvDqQkBLOdbmMvjc7TFZj6ab0YLuLYQ+7gZ5QSjJ
s80myss7iKGpuPK8/FQoxzZliQQVM69Fy92HQfVn0b7SDDHv+bUgF7lG4uI9ls03
zbPG9NZ+ieuMQ8VCYBBCaDqd8NGpLrowmzHF7BXUObCKFygZpMvMLI65M+Mz6wLA
SlMg0kvCbnxkp7bMcXctH7RCCqVx0gZofJoc5yt2RCgPnezdJI+F7h9AY6X3Sn0p
WdYKhJSYlAhqtMtl3dpJLSKqmpqidIuS4ssaEsEicJKSQKLkoWuUiVqK3+zwprBS
/M6Rr2BiJ4AQp8+5q3+XqlZAYSjDfoX0kv7OLB7nxDh2IA5p+skS/idWpGWS8APh
d2g77teh3b8myYbjUVRy2c+8LFnUMXMO+N67jEVV3iuLaSk6kD6E/dBDHleCYcij
iJPCRpGB8g/xlCOfGyZLrzAOqIAaqg9LoE54gqjpY93bIeW9BkSYtVIlluIYPyum
xPauTL95lR0j6foEUJkJueSI4mbTOBV0tHGg7QpX/uwyD/ZvY57bsv+lQLTJwitY
UG9H8/IitiHSiNmB0FcwuAQT6NVoqPOL+QsdA4lSFzV+rySfBZSo8RZ8kZ6x9TH+
ODzYkE2IcoFfOjwOD7Hs7lyb/APLAL4sTo2qDgNCG+1NIk978N1vg+tdDPfUEUrr
JwmOFxyeJtInSAppk7+z/DdFJ5G4rdZ/nWgik7QLeC0F9EoaAcOBS/KMPZz91TkH
Zj8pE4lDJkOBi5HGFjkaMV351LA55UeRE7vY8S+RAwTS2o1Mx99Xm6eJxbqvGbIY
WMD7ZbcyWU1zjRwFf+fEIF9vEX0Ysg4LsQlc6oEHMaB/fpvHvHzG+D5pjzqB0sPG
J/b7INPo1Og9pvCBHiIt92ZK9o6pDdd6aUhMl/dh+anhP5XHCyfa1i+lzlbL9UHP
oGV+FmBER0KkS3z8ER8C0w==
`protect END_PROTECTED
