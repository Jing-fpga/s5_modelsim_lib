`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N9Clba2Oju5VykiMZEud8vZDC/Ql/SvpARGxVESVuNUPikjZUYrqQ5royzaU4DTV
8UyGMVoe4wZjTaCmalTcF1q4q9tCVZX/XHYJjz4kiaeM8C3y/2bOypDQ9WNKmCBu
8ye+Z/vJbeXYEj41Ei8gmyP80ZrZoHkqa/CrBi+DGUqmg158qFZTeEq7E/1irkaY
YuPICykJSsqRTUWd5aNHVVB51go55vtuHfcJx3c0/RPvalPRcW7uHuQBz3sz17ML
5LEQHQX/rf0ftNbIFC2B4Ttw+KdRjcXkN2ufHtB8I7VrSV9leUPi1xGXh6XUl8S7
Lbz/v9oo6LXcpNccCAXngt3MNYf1mz5NLguN9UTjIgP+YNOwXmX0mfTAKBFeHwCp
8jFPlZuDQOxsfgyn2pl6FzG/xDxErMakmvMyGc9aitQODZ0GIy9ixqndscLk+HKq
DTvVS6XeLiclIdvHTx426j3X9d/xE1bkop86bzRGv5RBgcrvI2xjqSBm7enIOLBT
aBzIBjHYKQpcFRUAYkfZR4urus4nR1qUG4un0YxgiiOamgrQxfT2TCp3rFMo3HAM
kGwx4AihI/5eOxETdeDG8+JpQjBI+z9ohkyC2wRrjbsX00oddYMpFjFnk89cRGtL
KFF9BrE5BSXS4KJFJDAA+tLbFObE14e75fOIqWd0lwGkxvmEGqyeuW2fHAF1JOuu
YpFKdL2pFJbfOzg793gcbQiS6dIjeYjj/A090fRORY8+zCcBOOQfr5L2JbBHzunr
DLDhCD49Bo7Ltyo3QqASPAsMi4LEAyfKZeZjMDg3CRU=
`protect END_PROTECTED
