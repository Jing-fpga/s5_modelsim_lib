`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4h2aTGceWOmW1DQyha1InHFgnF45LUbKDh7vlYY3HL7ktq4qva3qT+Db0a1kUDWY
F+zJgn5Na96X2oENCoWPEvMlzWB5XH0d5vxhCHPEhymCNhGkQuqBUNOtYlcSPsaO
tjzgISwNUuqI6/Ryj3Nw1bbOrDkhdVzLwcz7iGXgbVKFPEFnIub6ufA8IuJg/Ucs
EO7kQcvHHMW8YozqtUUzu7RMLxR6WwvudYx/65N61/6cGfEAchW4qyD8mkJIyHyC
bZIG/GLC0+It0tcV/HKnpBVbl2ONZ3H5j/gL3ammHVKKSpGrpA9oKnc305v6H0g4
IRtzHUiN80bBAAzKso1iGo9bEwhiuF2k/V9EAh42X+bBgZ8N531watnP4TH7QZaL
e77eJD71hd8HECD2mRKjaVKxFsnTOdQc4vXlkpDQSkKa/HPah/jGIx/AyvW4HqLy
+oOMIcsSRixHSEyK/S4Bh6Y9lxBdZlTs6BdR3YzxMmknEFRjkqng7GLE8a+mSGrz
Mq3WMsgHTLIX75nuTLLgJlnrAqgvh2gtuBKl+oRBApeK2U1UUokqS7tZWAqVup88
hI+d61wK3u4bbQdiPQwkb7YN9t0j/sM8xe1p5macJ8M+6dIm8Kc8dERY2QSNhlKd
2K6k9di4vLQYy6Wup7UoQJCESrqXo3ElqdcwSrXzyx0U7HdNoOZK980wvjS77qWS
vOW6AZnKkDMw/8pLGJxquvbN6ES+tVRPRGLvcKKM3oH2ZP2F/MjfqHaEfHQFd5lv
mgayj3EaRZAWEzl+xzJP0MPAA2hYeP2D7xuHNxWXtLIye9JkH2XmxMSoi2cfS9XY
i7ZDgVZRD/yXBZpjHpg10L15Sh5hlNaUgL6QBTe19QMkkgNidrj6o6GxlEutEopg
U9WGbTWvrWzPs98k/ZDCJQlTU+qE7uQ0XGmt5XZStLhg2lTToSFX3jHhQL/6SPeo
FRjcFXnswky5r8nL7alYjdZcDS/vuNnVKVbfa5bkP1wk8aL8ejhfDC8l0rWrTmJJ
Ig0FtwqugEU/PZHwdSqygX8ohYEdkj1PswOUDQ8xGLlPfURYqaFwDFMVBV6D0nIg
fjyJNIGiLdLy5hn4QXhqCJrGCM5c3DqR1hl5NseAgbpKUrqWjTovrtjCU2B298kf
NX8nuqqN+DDO5lkYAaF58gp/aUuxxk/zkJdaYzNqj61HMZIjqgQze+VHVNliLNwf
XQFNYfE10bS6Ls4eFtLObx1EGTh3Mj5GuWHRYUoMkF0iapbb4VUXFRYmLfy1QOWH
Jg6QlrQmusb+o7JWB9Vjqm2vn24wangP/2gr12kTLSSnksvvumky1ZiOmdjMYr7w
FvRXBdaOzJuqXJcLGslkR+50iHjGsi7eBrd+60jqtuBR4wUVM3vn8RI+T2GZw3ei
ARvxTWUrmBQ9029NPOfGpYdIMe6VoIfQaBSD9rQksgfvhraQMRzVeUBdri/hLbMM
DRe5pIG/ApNwL7z4ksDCMyujw5Sl1VbvTBjyxbwJ4pe2N5cLU4cXIE5d4sBWAULn
LazXRHo4capipEY3RhOPW86aCmEUfiDL2/2Jo0nx/eten5nyxxcxd0dOOD6E3Zu0
HK9Fpu/1npzwCZIio9tYCkqsyZNowiktZoztoanENEvk+HuZMXNO3n4KAYQAmajV
VqIjkx/7tGiYo2ygazxWrmXJ0v4U8qqc/fmjJEh90dvuYzSZRaDa+mlAqkVIKKyL
b9uOEC7UCPioeRVjZX+OH+Uyesrzzyf9hDeXaXH9d/uYQMKmP0zpeN5aFapVx8VQ
XeSI6QyHhkbfZzGYUYs82Ypre1o1ptdliX9bIOqbstM+PfINmhfSHshCW6oHJkRj
jGQxZFqb+lqz5Q2QTyC7eNKwrVYEsaGCNbKvThr1JXpMLxNLA1CTgmAoy3cJIQQ+
Oq7LH0Iz5SZuXPwUm0xEoY+NzahfkymgNr4KfqpsG2pgSeLjWfiSq3qh3uJAik64
eminfD3bzTH3VhbCju457r7rYxN2kJrncNWxZBq1m8NcdX7qHk2KHRo1STFy62n5
cckdXCQ7UsApWRETuFawD68HCxdUtUNyhe9KEK0BOQIgK+Z1gHvaXYyxH1X21j85
Upzw5Kgp/Duoe+9Yo7vh7Vm6jgwfBCWeO6uttU+B4wTylFQX4jjyrtKPY84Ssqg4
ERpwWphAg99++FSe4qtRBYqwI9/hn3VAtg/B0fpmEfKI6BYODrhSpBq+75VXeX1Y
dySnj/RP3cUjLovOjQWveuFpsoDgpLOsGY0cw9yMw7zClHlOqunr9UcM+C8CrxBS
CMS1N8eD8G4AvNYApiF4A04y1HAvYApgRtORwM4RtSbAGBsR9szvWON3ScMbychl
itKQtggiCDCDwiEt6CHjq545+zQY+byGOR05FtCigr42sXDTL57pXbNLiKLvCDYI
dhS+ELMBeoJoE2FitmagN9CoxApeB8mUw/KzT16sumbKm6sQF9is2ng5NNB8Ytni
Ns91iN2a+cXenvULDQdbiVm5ZDY0uk5cylGDhltbt5s3R5EPLmwZZkEUw4CzE2cd
KLktYx8ynIU3zhNgnCKFW8u7QWGYraSxIl6b32imPW7BX1gJgAKeELfkJ4Qn3JnP
g480fS2k2Gwv/jscLwT34EETg/JwgNjnmDBYqOLxYaycIAWBx/QeHCSgOmqqdzDk
O0IaN6F+3RBLzAAD4DrXVDh3HanJInjTNbRRdvkAqXvo7UCoMR4jIKpVIqhI4maq
GfVVv1iSpnY6bVWLoCj6nZK+E3k4qBZ6ygfroTbyE0GIaxK4fWgpBeIEI4aO1yfW
4IG3Il9YmjJG0dhnwR7J/LVwjeq7n4s2ZIsRRYSVllxSawIdb82x87MZXptEvydU
vGbq7Zj+gfSuISEs+rKvr4XjxXlDODazMtfH5+3NTnjn2Qdaa655qsijntLaTpBm
XWshNT4O0H1mIp0LJ5V4hYpQGSErKFRZManl+fjwZXMUuu1TLgGt8diNtR3ingpP
wYhtN68FJ9i9EHcUGRWkdux17f3FaekrmW7ZLX1oEfJND9LCWee8B376cJINdnme
FwNAyyUZyPUiEJ/VguP1mXpAMP5FqswHzMTdnmR/oKx/EDzERIUgmb45Yz3K4aCy
HBj9WkAwtQixqOVauFnZAS518PPBPF3GXzJpw+pXlJiJKsoUv1ukIBSUakWkiajm
3ChAOrntKvPIzHj62UzRaiDrlLCE6ojvyRha7IBG/AO86aj0DB1ATJ6EjVF0lyeH
gXqm5R0jRiUZWr8RvTMMyjTXySCSlV9YuSZZH7F1CgzUz7NYQtc0tHb3XXnamcRV
BKAGb6OLWCQBScSVH+3pysQPkFpXnfxXRrif/iEUpriPxlC3RVigL6Cu7ul61X0S
69kL5RL+0D87ru2hohvbbJPoSWjgLXTrb1Hp4Wtn5GFIitiKs2ogADx+eebQpS+E
Ic57I8lz5SXYZ1fj7C4SyLvnK3G/i1rkK2y8VUlTF0SGoCS4TelZ0ECjP1lJGS3v
8P4yrvEQ8xq5bHB9zq/jwAULxcZrgQgDwTEf82I2+eumAd3L8ifERAqy5pfxU15v
t8Wyk19RVRgRNkjGaTbf5Idrt9OJSbPJIdQX13PUNrM3ofzX8eUeBfNfVhbWzrUK
FHT/12kYBOMwy2TCMKqR4BvwowRX9x3Ocha5y05zyvU=
`protect END_PROTECTED
