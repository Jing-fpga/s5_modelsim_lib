library verilog;
use verilog.vl_types.all;
entity stratixv_hssi_8g_rx_pcs is
    generic(
        enable_debug_info: string  := "false";
        fixed_pat_det   : string  := "dis_fixed_patdet";
        byte_deserializer: string  := "dis_bds";
        polinv_8b10b_dec: string  := "dis_polinv_8b10b_dec";
        clock_gate_bist : string  := "dis_bist_clk_gating";
        test_bus_sel    : string  := "prbs_bist_testbus";
        rx_clk2         : string  := "rcvd_clk_clk2";
        cdr_ctrl        : string  := "dis_cdr_ctrl";
        deskew_prog_pattern_only: string  := "en_deskew_prog_pat_only";
        wa_pld_controlled: string  := "dis_pld_ctrl";
        wa_rgnumber_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        eightb_tenb_decoder: string  := "dis_8b10b";
        wa_disp_err_flag: string  := "dis_disp_err_flag";
        re_bo_on_wa     : string  := "dis_re_bo_on_wa";
        wa_renumber_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ibm_invalid_code: string  := "dis_ibm_invalid_code";
        tx_rx_parallel_loopback: string  := "dis_plpbk";
        rate_match      : string  := "dis_rm";
        auto_error_replacement: string  := "dis_err_replace";
        wa_sync_sm_ctrl : string  := "gige_sync_sm";
        wa_rknumber_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hip_mode        : string  := "dis_hip";
        cdr_ctrl_rxvalid_mask: string  := "dis_rxvalid_mask";
        deskew_pattern  : vl_logic_vector(0 to 9) := (Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        symbol_swap     : string  := "dis_symbol_swap";
        wa_kchar        : string  := "dis_kchar";
        bypass_pipeline_reg: string  := "dis_bypass_pipeline";
        clock_gate_dw_wa: string  := "dis_dw_wa_clk_gating";
        clock_gate_dw_pc_wrclk: string  := "dis_dw_pc_wrclk_gating";
        pad_or_edb_error_replace: string  := "replace_edb";
        wa_rvnumber_data: vl_logic_vector(0 to 12) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        cid_pattern_len : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        deskew          : string  := "dis_deskew";
        eidle_entry_sd  : string  := "dis_eidle_sd";
        eightbtenb_decoder_output_sel: string  := "data_8b10b_decoder";
        sup_mode        : string  := "user_mode";
        rx_pcs_urst     : string  := "en_rx_pcs_urst";
        prbs_ver        : string  := "dis_prbs";
        agg_block_sel   : string  := "same_smrt_pack";
        rx_wr_clk       : string  := "rx_clk2_div_1_2_4";
        fixed_pat_num   : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        bo_pattern      : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        eidle_entry_iei : string  := "dis_eidle_iei";
        use_default_base_address: string  := "true";
        comp_fifo_rst_pld_ctrl: string  := "dis_comp_fifo_rst_pld_ctrl";
        wait_cnt        : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        clkcmp_pattern_n: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        force_signal_detect: string  := "en_force_signal_detect";
        clock_gate_dw_dskw_wr: string  := "dis_dw_dskw_wrclk_gating";
        rx_clk1         : string  := "rcvd_clk_clk1";
        pma_done_count  : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        invalid_code_flag_only: string  := "dis_invalid_code_only";
        clock_gate_cdr_eidle: string  := "dis_cdr_eidle_clk_gating";
        clock_gate_bds_dec_asn: string  := "dis_bds_dec_asn_clk_gating";
        wa_rosnumber_data: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        clock_gate_sw_rm_rd: string  := "dis_sw_rm_rdclk_gating";
        err_flags_sel   : string  := "err_flags_wa";
        ctrl_plane_bonding_compensation: string  := "dis_compensation";
        bist_ver_clr_flag: string  := "dis_bist_clr_flag";
        clock_gate_byteorder: string  := "dis_byteorder_clk_gating";
        clock_gate_sw_rm_wr: string  := "dis_sw_rm_wrclk_gating";
        rx_clk_free_running: string  := "en_rx_clk_free_run";
        polarity_inversion: string  := "dis_pol_inv";
        auto_deassert_pc_rst_cnt_data: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        user_base_address: integer := 0;
        bo_pad          : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        clkcmp_pattern_p: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        wa_clk_slip_spacing_data: vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        clock_gate_prbs : string  := "dis_prbs_clk_gating";
        clock_gate_sw_wa: string  := "dis_sw_wa_clk_gating";
        runlength_val   : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        wa_pd           : string  := "wa_pd_10";
        bit_reversal    : string  := "dis_bit_reversal";
        wa_pd_data      : vl_logic_vector(0 to 39) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pc_fifo_rst_pld_ctrl: string  := "dis_pc_fifo_rst_pld_ctrl";
        mask_cnt        : vl_logic_vector(0 to 9) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        ctrl_plane_bonding_distribution: string  := "not_master_chnl_distr";
        cid_pattern     : string  := "cid_pattern_0";
        wait_for_phfifo_cnt_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pma_dw          : string  := "eight_bit";
        byte_order      : string  := "dis_bo";
        wa_det_latency_sync_status_beh: string  := "assert_sync_status_non_imm";
        clock_gate_sw_pc_wrclk: string  := "dis_sw_pc_wrclk_gating";
        prbs_ver_clr_flag: string  := "dis_prbs_clr_flag";
        clock_gate_pc_rdclk: string  := "dis_pc_rdclk_gating";
        pcs_bypass      : string  := "dis_pcs_bypass";
        dw_one_or_two_symbol_bo: string  := "donot_care_one_two_bo";
        pipe_if_enable  : string  := "dis_pipe_rx";
        avmm_group_channel_index: integer := 0;
        phase_compensation_fifo: string  := "low_latency";
        clock_gate_dskw_rd: string  := "dis_dskw_rdclk_gating";
        rx_rcvd_clk     : string  := "rcvd_clk_rcvd_clk";
        rx_refclk       : string  := "dis_refclk_sel";
        channel_number  : integer := 0;
        clock_gate_dw_rm_rd: string  := "dis_dw_rm_rdclk_gating";
        clock_gate_sw_dskw_wr: string  := "dis_sw_dskw_wrclk_gating";
        auto_pc_en_cnt_data: vl_logic_vector(0 to 6) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        wa_pd_polarity  : string  := "dis_pd_both_pol";
        wa_clk_slip_spacing: string  := "min_clk_slip_spacing";
        test_mode       : string  := "prbs";
        wa_boundary_lock_ctrl: string  := "bit_slip";
        ctrl_plane_bonding_consumption: string  := "individual";
        prot_mode       : string  := "basic";
        rx_rd_clk       : string  := "pld_rx_clk";
        eidle_entry_eios: string  := "dis_eidle_eios";
        auto_speed_nego : string  := "dis_asn";
        bist_ver        : string  := "dis_bist";
        clock_gate_dw_rm_wr: string  := "dis_dw_rm_wrclk_gating";
        runlength_check : string  := "en_runlength_sw";
        silicon_rev     : string  := "reve"
    );
    port(
        a1a2k1k2flag    : out    vl_logic_vector(3 downto 0);
        a1a2size        : in     vl_logic_vector(0 downto 0);
        aggrxpcsrst     : out    vl_logic_vector(0 downto 0);
        aggtestbus      : in     vl_logic_vector(15 downto 0);
        aligndetsync    : out    vl_logic_vector(1 downto 0);
        alignstatus     : in     vl_logic_vector(0 downto 0);
        alignstatuspld  : out    vl_logic_vector(0 downto 0);
        alignstatussync : out    vl_logic_vector(0 downto 0);
        alignstatussync0: in     vl_logic_vector(0 downto 0);
        alignstatussync0toporbot: in     vl_logic_vector(0 downto 0);
        alignstatustoporbot: in     vl_logic_vector(0 downto 0);
        avmmaddress     : in     vl_logic_vector(10 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        bistdone        : out    vl_logic_vector(0 downto 0);
        bisterr         : out    vl_logic_vector(0 downto 0);
        bitreversalenable: in     vl_logic_vector(0 downto 0);
        bitslip         : in     vl_logic_vector(0 downto 0);
        blockselect     : out    vl_logic_vector(0 downto 0);
        byteorder       : in     vl_logic_vector(0 downto 0);
        byteordflag     : out    vl_logic_vector(0 downto 0);
        bytereversalenable: in     vl_logic_vector(0 downto 0);
        cgcomprddall    : in     vl_logic_vector(0 downto 0);
        cgcomprddalltoporbot: in     vl_logic_vector(0 downto 0);
        cgcomprddout    : out    vl_logic_vector(1 downto 0);
        cgcompwrall     : in     vl_logic_vector(0 downto 0);
        cgcompwralltoporbot: in     vl_logic_vector(0 downto 0);
        cgcompwrout     : out    vl_logic_vector(1 downto 0);
        channeltestbusout: out    vl_logic_vector(19 downto 0);
        clocktopld      : out    vl_logic_vector(0 downto 0);
        configselinchnldown: in     vl_logic_vector(0 downto 0);
        configselinchnlup: in     vl_logic_vector(0 downto 0);
        configseloutchnldown: out    vl_logic_vector(0 downto 0);
        configseloutchnlup: out    vl_logic_vector(0 downto 0);
        ctrlfromaggblock: in     vl_logic_vector(0 downto 0);
        datafrinaggblock: in     vl_logic_vector(7 downto 0);
        datain          : in     vl_logic_vector(19 downto 0);
        dataout         : out    vl_logic_vector(63 downto 0);
        decoderctrl     : out    vl_logic_vector(0 downto 0);
        decoderdata     : out    vl_logic_vector(7 downto 0);
        decoderdatavalid: out    vl_logic_vector(0 downto 0);
        delcondmet0     : in     vl_logic_vector(0 downto 0);
        delcondmet0toporbot: in     vl_logic_vector(0 downto 0);
        delcondmetout   : out    vl_logic_vector(0 downto 0);
        disablepcfifobyteserdes: out    vl_logic_vector(0 downto 0);
        dispcbytegen3   : in     vl_logic_vector(0 downto 0);
        dynclkswitchn   : in     vl_logic_vector(0 downto 0);
        earlyeios       : out    vl_logic_vector(0 downto 0);
        eidledetected   : out    vl_logic_vector(0 downto 0);
        eidleexit       : out    vl_logic_vector(0 downto 0);
        eidleinfersel   : in     vl_logic_vector(2 downto 0);
        enablecommadetect: in     vl_logic_vector(0 downto 0);
        endskwqd        : in     vl_logic_vector(0 downto 0);
        endskwqdtoporbot: in     vl_logic_vector(0 downto 0);
        endskwrdptrs    : in     vl_logic_vector(0 downto 0);
        endskwrdptrstoporbot: in     vl_logic_vector(0 downto 0);
        errctrl         : out    vl_logic_vector(1 downto 0);
        errdata         : out    vl_logic_vector(15 downto 0);
        fifoovr0        : in     vl_logic_vector(0 downto 0);
        fifoovr0toporbot: in     vl_logic_vector(0 downto 0);
        fifoovrout      : out    vl_logic_vector(0 downto 0);
        fifordincomp0toporbot: in     vl_logic_vector(0 downto 0);
        fifordoutcomp   : out    vl_logic_vector(0 downto 0);
        fiforstrdqd     : in     vl_logic_vector(0 downto 0);
        fiforstrdqdtoporbot: in     vl_logic_vector(0 downto 0);
        gen2ngen1       : in     vl_logic_vector(0 downto 0);
        hrdrst          : in     vl_logic_vector(0 downto 0);
        insertincomplete0: in     vl_logic_vector(0 downto 0);
        insertincomplete0toporbot: in     vl_logic_vector(0 downto 0);
        insertincompleteout: out    vl_logic_vector(0 downto 0);
        latencycomp0    : in     vl_logic_vector(0 downto 0);
        latencycomp0toporbot: in     vl_logic_vector(0 downto 0);
        latencycompout  : out    vl_logic_vector(0 downto 0);
        ltr             : out    vl_logic_vector(0 downto 0);
        observablebyteserdesclock: out    vl_logic_vector(0 downto 0);
        parallelloopback: in     vl_logic_vector(19 downto 0);
        parallelrevloopback: out    vl_logic_vector(19 downto 0);
        pcfifoempty     : out    vl_logic_vector(0 downto 0);
        pcfifofull      : out    vl_logic_vector(0 downto 0);
        pcfifordenable  : in     vl_logic_vector(0 downto 0);
        pcieswitch      : out    vl_logic_vector(0 downto 0);
        pcieswitchgen3  : in     vl_logic_vector(0 downto 0);
        phfifouserrst   : in     vl_logic_vector(0 downto 0);
        phystatus       : out    vl_logic_vector(0 downto 0);
        phystatusinternal: in     vl_logic_vector(0 downto 0);
        phystatuspcsgen3: in     vl_logic_vector(0 downto 0);
        pipedata        : out    vl_logic_vector(63 downto 0);
        pipeloopbk      : in     vl_logic_vector(0 downto 0);
        pldltr          : in     vl_logic_vector(0 downto 0);
        pldrxclk        : in     vl_logic_vector(0 downto 0);
        polinvrx        : in     vl_logic_vector(0 downto 0);
        prbscidenable   : in     vl_logic_vector(0 downto 0);
        prbsdone        : out    vl_logic_vector(0 downto 0);
        prbserrlt       : out    vl_logic_vector(0 downto 0);
        pxfifowrdisable : in     vl_logic_vector(0 downto 0);
        rateswitchcontrol: in     vl_logic_vector(0 downto 0);
        rcvdclkagg      : in     vl_logic_vector(0 downto 0);
        rcvdclkaggtoporbot: in     vl_logic_vector(0 downto 0);
        rcvdclkpma      : in     vl_logic_vector(0 downto 0);
        rdalign         : out    vl_logic_vector(1 downto 0);
        rdenableinchnldown: in     vl_logic_vector(0 downto 0);
        rdenableinchnlup: in     vl_logic_vector(0 downto 0);
        rdenableoutchnldown: out    vl_logic_vector(0 downto 0);
        rdenableoutchnlup: out    vl_logic_vector(0 downto 0);
        refclkdig       : in     vl_logic_vector(0 downto 0);
        refclkdig2      : in     vl_logic_vector(0 downto 0);
        resetpcptrs     : out    vl_logic_vector(0 downto 0);
        resetpcptrsgen3 : in     vl_logic_vector(0 downto 0);
        resetpcptrsinchnldown: in     vl_logic_vector(0 downto 0);
        resetpcptrsinchnldownpipe: out    vl_logic_vector(0 downto 0);
        resetpcptrsinchnlup: in     vl_logic_vector(0 downto 0);
        resetpcptrsinchnluppipe: out    vl_logic_vector(0 downto 0);
        resetpcptrsoutchnldown: out    vl_logic_vector(0 downto 0);
        resetpcptrsoutchnlup: out    vl_logic_vector(0 downto 0);
        resetppmcntrsgen3: in     vl_logic_vector(0 downto 0);
        resetppmcntrsinchnldown: in     vl_logic_vector(0 downto 0);
        resetppmcntrsinchnlup: in     vl_logic_vector(0 downto 0);
        resetppmcntrsoutchnldown: out    vl_logic_vector(0 downto 0);
        resetppmcntrsoutchnlup: out    vl_logic_vector(0 downto 0);
        resetppmcntrspcspma: out    vl_logic_vector(0 downto 0);
        rlvlt           : out    vl_logic_vector(0 downto 0);
        rmfifoempty     : out    vl_logic_vector(0 downto 0);
        rmfifofull      : out    vl_logic_vector(0 downto 0);
        rmfifopartialempty: out    vl_logic_vector(0 downto 0);
        rmfifopartialfull: out    vl_logic_vector(0 downto 0);
        rmfifordincomp0 : in     vl_logic_vector(0 downto 0);
        rmfiforeadenable: in     vl_logic_vector(0 downto 0);
        rmfifouserrst   : in     vl_logic_vector(0 downto 0);
        rmfifowriteenable: in     vl_logic_vector(0 downto 0);
        runlengthviolation: out    vl_logic_vector(0 downto 0);
        runningdisparity: out    vl_logic_vector(1 downto 0);
        rxblkstart      : out    vl_logic_vector(3 downto 0);
        rxblkstartpcsgen3: in     vl_logic_vector(3 downto 0);
        rxclkoutgen3    : out    vl_logic_vector(0 downto 0);
        rxclkslip       : out    vl_logic_vector(0 downto 0);
        rxcontrolrstoporbot: in     vl_logic_vector(0 downto 0);
        rxdatapcsgen3   : in     vl_logic_vector(63 downto 0);
        rxdatarstoporbot: in     vl_logic_vector(7 downto 0);
        rxdatavalid     : out    vl_logic_vector(3 downto 0);
        rxdatavalidpcsgen3: in     vl_logic_vector(3 downto 0);
        rxdivsyncinchnldown: in     vl_logic_vector(1 downto 0);
        rxdivsyncinchnlup: in     vl_logic_vector(1 downto 0);
        rxdivsyncoutchnldown: out    vl_logic_vector(1 downto 0);
        rxdivsyncoutchnlup: out    vl_logic_vector(1 downto 0);
        rxpcsrst        : in     vl_logic_vector(0 downto 0);
        rxpipeclk       : out    vl_logic_vector(0 downto 0);
        rxpipesoftreset : out    vl_logic_vector(0 downto 0);
        rxstatus        : out    vl_logic_vector(2 downto 0);
        rxstatusinternal: in     vl_logic_vector(2 downto 0);
        rxstatuspcsgen3 : in     vl_logic_vector(2 downto 0);
        rxsynchdr       : out    vl_logic_vector(1 downto 0);
        rxsynchdrpcsgen3: in     vl_logic_vector(1 downto 0);
        rxvalid         : out    vl_logic_vector(0 downto 0);
        rxvalidinternal : in     vl_logic_vector(0 downto 0);
        rxvalidpcsgen3  : in     vl_logic_vector(0 downto 0);
        rxweinchnldown  : in     vl_logic_vector(1 downto 0);
        rxweinchnlup    : in     vl_logic_vector(1 downto 0);
        rxweoutchnldown : out    vl_logic_vector(1 downto 0);
        rxweoutchnlup   : out    vl_logic_vector(1 downto 0);
        scanmode        : in     vl_logic_vector(0 downto 0);
        selftestdone    : out    vl_logic_vector(0 downto 0);
        selftesterr     : out    vl_logic_vector(0 downto 0);
        sigdetfrompma   : in     vl_logic_vector(0 downto 0);
        signaldetectout : out    vl_logic_vector(0 downto 0);
        speedchange     : out    vl_logic_vector(0 downto 0);
        speedchangeinchnldown: in     vl_logic_vector(0 downto 0);
        speedchangeinchnldownpipe: out    vl_logic_vector(0 downto 0);
        speedchangeinchnlup: in     vl_logic_vector(0 downto 0);
        speedchangeinchnluppipe: out    vl_logic_vector(0 downto 0);
        speedchangeoutchnldown: out    vl_logic_vector(0 downto 0);
        speedchangeoutchnlup: out    vl_logic_vector(0 downto 0);
        syncdatain      : out    vl_logic_vector(0 downto 0);
        syncsmen        : in     vl_logic_vector(0 downto 0);
        syncstatus      : out    vl_logic_vector(0 downto 0);
        txctrlplanetestbus: in     vl_logic_vector(19 downto 0);
        txdivsync       : in     vl_logic_vector(1 downto 0);
        txpmaclk        : in     vl_logic_vector(0 downto 0);
        txtestbus       : in     vl_logic_vector(19 downto 0);
        wordalignboundary: out    vl_logic_vector(4 downto 0);
        wrenableinchnldown: in     vl_logic_vector(0 downto 0);
        wrenableinchnlup: in     vl_logic_vector(0 downto 0);
        wrenableoutchnldown: out    vl_logic_vector(0 downto 0);
        wrenableoutchnlup: out    vl_logic_vector(0 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of fixed_pat_det : constant is 1;
    attribute mti_svvh_generic_type of byte_deserializer : constant is 1;
    attribute mti_svvh_generic_type of polinv_8b10b_dec : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_bist : constant is 1;
    attribute mti_svvh_generic_type of test_bus_sel : constant is 1;
    attribute mti_svvh_generic_type of rx_clk2 : constant is 1;
    attribute mti_svvh_generic_type of cdr_ctrl : constant is 1;
    attribute mti_svvh_generic_type of deskew_prog_pattern_only : constant is 1;
    attribute mti_svvh_generic_type of wa_pld_controlled : constant is 1;
    attribute mti_svvh_generic_type of wa_rgnumber_data : constant is 1;
    attribute mti_svvh_generic_type of eightb_tenb_decoder : constant is 1;
    attribute mti_svvh_generic_type of wa_disp_err_flag : constant is 1;
    attribute mti_svvh_generic_type of re_bo_on_wa : constant is 1;
    attribute mti_svvh_generic_type of wa_renumber_data : constant is 1;
    attribute mti_svvh_generic_type of ibm_invalid_code : constant is 1;
    attribute mti_svvh_generic_type of tx_rx_parallel_loopback : constant is 1;
    attribute mti_svvh_generic_type of rate_match : constant is 1;
    attribute mti_svvh_generic_type of auto_error_replacement : constant is 1;
    attribute mti_svvh_generic_type of wa_sync_sm_ctrl : constant is 1;
    attribute mti_svvh_generic_type of wa_rknumber_data : constant is 1;
    attribute mti_svvh_generic_type of hip_mode : constant is 1;
    attribute mti_svvh_generic_type of cdr_ctrl_rxvalid_mask : constant is 1;
    attribute mti_svvh_generic_type of deskew_pattern : constant is 1;
    attribute mti_svvh_generic_type of symbol_swap : constant is 1;
    attribute mti_svvh_generic_type of wa_kchar : constant is 1;
    attribute mti_svvh_generic_type of bypass_pipeline_reg : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_dw_wa : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_dw_pc_wrclk : constant is 1;
    attribute mti_svvh_generic_type of pad_or_edb_error_replace : constant is 1;
    attribute mti_svvh_generic_type of wa_rvnumber_data : constant is 1;
    attribute mti_svvh_generic_type of cid_pattern_len : constant is 1;
    attribute mti_svvh_generic_type of deskew : constant is 1;
    attribute mti_svvh_generic_type of eidle_entry_sd : constant is 1;
    attribute mti_svvh_generic_type of eightbtenb_decoder_output_sel : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of rx_pcs_urst : constant is 1;
    attribute mti_svvh_generic_type of prbs_ver : constant is 1;
    attribute mti_svvh_generic_type of agg_block_sel : constant is 1;
    attribute mti_svvh_generic_type of rx_wr_clk : constant is 1;
    attribute mti_svvh_generic_type of fixed_pat_num : constant is 1;
    attribute mti_svvh_generic_type of bo_pattern : constant is 1;
    attribute mti_svvh_generic_type of eidle_entry_iei : constant is 1;
    attribute mti_svvh_generic_type of use_default_base_address : constant is 1;
    attribute mti_svvh_generic_type of comp_fifo_rst_pld_ctrl : constant is 1;
    attribute mti_svvh_generic_type of wait_cnt : constant is 1;
    attribute mti_svvh_generic_type of clkcmp_pattern_n : constant is 1;
    attribute mti_svvh_generic_type of force_signal_detect : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_dw_dskw_wr : constant is 1;
    attribute mti_svvh_generic_type of rx_clk1 : constant is 1;
    attribute mti_svvh_generic_type of pma_done_count : constant is 1;
    attribute mti_svvh_generic_type of invalid_code_flag_only : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_cdr_eidle : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_bds_dec_asn : constant is 1;
    attribute mti_svvh_generic_type of wa_rosnumber_data : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_sw_rm_rd : constant is 1;
    attribute mti_svvh_generic_type of err_flags_sel : constant is 1;
    attribute mti_svvh_generic_type of ctrl_plane_bonding_compensation : constant is 1;
    attribute mti_svvh_generic_type of bist_ver_clr_flag : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_byteorder : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_sw_rm_wr : constant is 1;
    attribute mti_svvh_generic_type of rx_clk_free_running : constant is 1;
    attribute mti_svvh_generic_type of polarity_inversion : constant is 1;
    attribute mti_svvh_generic_type of auto_deassert_pc_rst_cnt_data : constant is 1;
    attribute mti_svvh_generic_type of user_base_address : constant is 1;
    attribute mti_svvh_generic_type of bo_pad : constant is 1;
    attribute mti_svvh_generic_type of clkcmp_pattern_p : constant is 1;
    attribute mti_svvh_generic_type of wa_clk_slip_spacing_data : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_prbs : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_sw_wa : constant is 1;
    attribute mti_svvh_generic_type of runlength_val : constant is 1;
    attribute mti_svvh_generic_type of wa_pd : constant is 1;
    attribute mti_svvh_generic_type of bit_reversal : constant is 1;
    attribute mti_svvh_generic_type of wa_pd_data : constant is 1;
    attribute mti_svvh_generic_type of pc_fifo_rst_pld_ctrl : constant is 1;
    attribute mti_svvh_generic_type of mask_cnt : constant is 1;
    attribute mti_svvh_generic_type of ctrl_plane_bonding_distribution : constant is 1;
    attribute mti_svvh_generic_type of cid_pattern : constant is 1;
    attribute mti_svvh_generic_type of wait_for_phfifo_cnt_data : constant is 1;
    attribute mti_svvh_generic_type of pma_dw : constant is 1;
    attribute mti_svvh_generic_type of byte_order : constant is 1;
    attribute mti_svvh_generic_type of wa_det_latency_sync_status_beh : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_sw_pc_wrclk : constant is 1;
    attribute mti_svvh_generic_type of prbs_ver_clr_flag : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_pc_rdclk : constant is 1;
    attribute mti_svvh_generic_type of pcs_bypass : constant is 1;
    attribute mti_svvh_generic_type of dw_one_or_two_symbol_bo : constant is 1;
    attribute mti_svvh_generic_type of pipe_if_enable : constant is 1;
    attribute mti_svvh_generic_type of avmm_group_channel_index : constant is 1;
    attribute mti_svvh_generic_type of phase_compensation_fifo : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_dskw_rd : constant is 1;
    attribute mti_svvh_generic_type of rx_rcvd_clk : constant is 1;
    attribute mti_svvh_generic_type of rx_refclk : constant is 1;
    attribute mti_svvh_generic_type of channel_number : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_dw_rm_rd : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_sw_dskw_wr : constant is 1;
    attribute mti_svvh_generic_type of auto_pc_en_cnt_data : constant is 1;
    attribute mti_svvh_generic_type of wa_pd_polarity : constant is 1;
    attribute mti_svvh_generic_type of wa_clk_slip_spacing : constant is 1;
    attribute mti_svvh_generic_type of test_mode : constant is 1;
    attribute mti_svvh_generic_type of wa_boundary_lock_ctrl : constant is 1;
    attribute mti_svvh_generic_type of ctrl_plane_bonding_consumption : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of rx_rd_clk : constant is 1;
    attribute mti_svvh_generic_type of eidle_entry_eios : constant is 1;
    attribute mti_svvh_generic_type of auto_speed_nego : constant is 1;
    attribute mti_svvh_generic_type of bist_ver : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_dw_rm_wr : constant is 1;
    attribute mti_svvh_generic_type of runlength_check : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
end stratixv_hssi_8g_rx_pcs;
