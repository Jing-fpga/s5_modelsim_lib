`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EBgLEwvZgvB8WqiE/awbsTXVAnb65TCMQqUtbtaZjMv/6rOonJ/vM50u57jRBHs8
4KItC+f175Kb7obPlNDhVfT2n9vVapL/U7MUeiryXP3xY2skRgzPqTsVcYoix8CG
JZl7XubvgW8kFz0k6n+/t85li/jLCLSZIrTN5z3CuQ+VzOosf7XqOxMcehmvtZuL
HfsNet1y+Lh59Jj38ZI0f5et/dRNj7b71zXibMyHAqoq4Gs57hHrEUcJj73JnLpg
kB4l1bgErO4AnfLQMykP2LRENgkCMIMg3dXOIXvjbhHTRGxULROVduVqORX6uiqT
5fTeOZ3hlwptqRPMf8pU7c7MUfuFRc41Lx39EqoCCMpv3curccenOPaw29B5rmnr
2tMRG8mBcGXrneDPSQa+zPijAEKR0f4SOQGoe82GlADw60q4xqnNsL2NtGt4H3lk
JXE5O5sea43vfR8ffbEXZgWYQfGVu6XXI+EEYb0jMpuNz4TEUDIxqy3LRwLni+4h
Tsi4Cp+9BQ9qQ2uZDWfayuU0OAqW/DsLI0fIK0xb8w5uk5xx1iQ64ZqdnZ5xwUoK
cgRfMowAEn8Llr5OCqX7ruYTR/SQxVyy74Fq365wDY6cGJ6/rOMD60MdQNCZkdWv
laWNK88FAJS43kGRtVObY2XyUEOGeymW+0kAuSJXSPyEd6Ir4QVhH3pJB9U/XuTm
UXN+Ext4MCIeUM/bu6mVbUh9oKWdLPTeQEoW4iZpK0chQP37Ioz7W8yqsT74oww4
sbBVPDbjUa/tLgjlx9plN8hHs1SlHwbKpTVm3JpJK0Sj6Sx5dYwp/TvkrFL+1AyM
Jx6M96ZPRxB/dNHs3MXLykYHCV9gkGuzYlsMtdBOjFDdDCWdkB9EY7QBGJ6605yU
CqO/2RODHv6C9Xjwublf2/wZW8Wjl0WgxsXNWoE+l+Q=
`protect END_PROTECTED
