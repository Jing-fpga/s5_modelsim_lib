`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CTf15N2Cz0N43miwrm8QKdqGHSCs+4PAe0YETz3RfpINuAxwkAFqZ+NN6LVLxVr1
i9MlHLmBIDTpdZx2N9AuodZRDKcjRRDk9s1bgSBtIWB/I7iR09XFFnPcwnl9FQpZ
Js/9Cm1sVcSat3291B8EJSxM2ppnHNLF40NYvzLBTjAf8VIJFhdsb38m42CFyn6V
XPUhvL2yDZv3c6gqAfPjyWTqGZI4hKum+xPPABcCZlgckKLuzpR/dV+X6GMlgiDP
B+5Lqk82uYvixMajM5BUoSUR60t1cprBLCN+y5G+vHywZoStY5Au0gHFI6d1xh4s
9Eif6iDaqxv/ftT+auRwXkECxCzbfKcEpB6KTqp++7t4O3wSepM8S0+A1byiU8qI
8xDk/BTu4jbjzOH7FR4R1fULb2Gn247iV3lybgWdbamD1L6cR/8HOK55v+6qOtWR
zJt/7bKARrqbXCBsLbni46dLnzudDoFDH6WXnLKR61WOXNYtYcvLRPiVNzuzivw4
ToDqgaFsAOCn+WAbTJBSLL5b8kFMa0PjBqkVC6HBLT9k4OVgElyaPtNuYLcBmOJ2
gjSuJOrDvZsc6QiKCVAEU4dJxeDYRw+uy2aDJAw+MADYnPbVPw0+kfxfXbzKTvXY
5J4biDE41Phsgb032Qf9xVqHuMG87cgVkRG7lseLXcAdAdi073mRtVUpQ+qcwWSK
Ia5syK26SJmBxH0ZpCXwXaIUHLU6uDP84bzYOdVUdOo2xkICTz18Z1GiWjfe2A4v
T6mRrlfIYX9eb4aeX2hzc+dJTQGWF/+bSZ4wc+9/palfK7VeE5WQNtN0DbmP2GsZ
INH8rYb6QOXCxqlpk/qRbuyIigHZCM+7/jQfO2KrdA0ckUmYS8LhSGHOCCek2Tu2
4alSUbUOFTlEU5eDIL+vWYF/PWjkdeEtT24rHuPmEAhl9VdNr/9+RV8QGOrq+W47
eKtP+D8Abie6pgUtB6bo7AZk6eYJ8MoY3ddn/MIFygyeFnzPEoOae5LrBo2cBm2v
oKktJTgXjIGmTHil4xi4lRKyuCPs/Xs9g93v7i9rx4mleANret9mNW7vRtid172C
97jLgLn47Sup5VVL5MCQInyLeGVQYhRU0D+FVWk1gtGts6WpPk+msgLytvFdXwLg
AMuPVn22p2Xz6qQk3zC/3+2aGqTzozFk9Y3rRaj/6gcoSTTGXk3UmtK7/CBY0CqG
dRPCLzZD9qPEz15DH7FUkcT4vTPMyvnXNabdEAKOG0kLzvWqBsWC06Y7GM/Oqka4
fb7kwsz3koi4OoZwfogWwPKPmthY6nUIrKmzI7i7RD10jSmsFZNDuqbq2vUO8Ijh
YlXGmAXCgnAm3RQzxoaPbXDOqFQl9HI6VEvpIHpRtXf1CwpjynENvbzP+PT1qAYt
t5H0zNficEVhV4NICy5JhOIaY/eoeAsZRS9sU54oQkdcwCfRue2AR5EcYcDSb1f9
qOSzsIGvgDigKDnCaawvu5MX5WCFhXtcu9ltExQAxdUIwZ7meWsCnqxIalJrWZ/G
68956ltsiWtn7w+xRr8k8pRlD+rhgsdtutKPlJTHLbnYkgXr+F7OdW+MrwgQQBpx
DOc3+b60Q00jIgSf7b2fPIc10+XbzhwTKDLMTlfIy2c8eaU0mspY6IZu3S2u0aFD
SCsKJe+8dtsy6D6bTwq7uw8uPEOrLGsPwEe5aQ3Sjcc0KlexoAeKEtBXVkLWVhY2
3i0MR6mxE3U9fbby69yppTaHtCoPg8jUd1FlKBuI69k=
`protect END_PROTECTED
