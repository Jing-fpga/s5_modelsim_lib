`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dwfnZgbVWkxfgTZgMwIKkpCFlVVu6GkA+/NhREvsw1gogcs7R4hK6IUi4JGlJtNV
dJbYl89MBVUJwIRhGhpX9fT9obz+vFCdJj3+rzYgQvJDdFyxjoDvwmXzSBhmR5V2
HHajUnYgDhtsmKa8lAQziahv7KIhHY2ISTMUk289q59VMPacqJpEN6f3XvFfUddG
0NgcSDJszAMf+Zp8422PPtdUi2ryTAtw6IfMjL9gxqELqlvpT5XbVoK+uK65nDm9
T97O27aNWkAI14GwrEzU3NjaAKl8aDbUZFklwIp14vOyb/T8MF3gRU03iVoeVRJI
ZpUqNlar6rvwu0QKf5iFlQKF0pJqXOSZerZIIMeD9P461rFzeVVcsTC2GzjRY4ke
ddvFavc6XH7i9uYLZ1mgh9ivtmANwQ3OBoMriC3jhyVmXM75oI2W05xS2TDR/S5H
TLl18IRokLYWPFPn5XgZreXo4mK7r2+tvSOyCYLqTREO3HTTrQPaa47Do2l4Cxv9
0vf7gb93M8v411O+stb/VhL5AxkodcUP0j55L+/TpJX3Hu9EW5dcQqMncnFqN4w9
0BKucLuL8JuCGpJF7hR5Ao5jVGWFrS2/qL9tVhn4HFkR5pLFbdtJ72THU/J5dGYl
147s2wG9UCUU+1MiOZYmM2kM1Fqe9Eu5CLLerXnkqjXLoXE8geIBL8lArKqG72m7
x+I95ZKNk26GvSpcJ9xa2JHBYvzCVGuVCXNJp4midzvv5ne4TnNJYeqORyuxfxVo
tTykIG6ahCE1uBP44Grx4F/rz9PPe+g6TWJ6fPUVN76DeusdIzpKlHkQVp4alZvi
KDdll6S/lbl7YyH6c3DBrdd8YD103J9kGVxfNuM3joE=
`protect END_PROTECTED
