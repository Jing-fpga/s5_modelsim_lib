`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BgJdo/G7q6PORW8DQyI4qe/bQN8btkPMG9Vr6T+y7Z0K/QfXXb1bE65Z7BVtEdeZ
ia01gsmsR1XZEZL54srqU+BBDNCc9RSeKUbdUfaUWDZrQ57wmUiLpYJIk0rhKc7i
BY79JKxOITe5QFqD6uOadyekJrBVuhXM8kTuJ9T71FV4p2VPueS60+IR9VHrphNz
gJyxaTc/eSJq5KNbVAyswVTpUYSdTNdx78fTWJ0fuOTbS8+XUvMRj9rXzGAoo353
WDg0DTkMHsuL5ZEr4NT6nkC4s3uU/uR3hZiG3/KywqmdIEQdNWs33iP7+lgtO2QW
r7yGqMolK1aNlZs9h4MBFtYYR/SdbSRXIIxPRwdBH9iEEUObellLb8lrScJJkKWa
GKeg3Y2Cr92yDl8bMOZdJg7D1nhV9u2UNr06IMUTS+XNptUn4c3WVCm9Ykjczxw9
RKZ68EVqgkIdLCRm7LI+/07I2jJWeFl/5o/gGK9wm+QLPIdLs58UoCQu0G55/TXF
QIWSBP5iDPspVestWEAyjIrXm104A7frW4JtayjzaLFYFTJBKeMJmGXGRnEo5b/t
UentyV6cOWJbFCYc0k28aZYBxXmcD5eAzVHmH47dynxeffwPdpW+RGmmkrl0GK8D
fy7pxQ+/EHtfVyt0PN0h/8CBzPwSEzwVOwc1iSopGJ0BRTi2pW6aGqZgAVgMZ6Ax
4JkabnkP0IGwF5Iceknky7uK4+pTdjEHepd5SXWUxGx8PgOlV0Y60Fsk8sMjaf3d
l4sPpHgv/N8/td723pW1N2Wi9L/Gz6cpAXhQvywpRdAW+fNUMDw2pWnqI6bJsvfb
yloUGwTh8KUehB4FaYPt3ycwQznbmdvZsR2kfLpcFV0PxVWXHyRNS7/YYX/GgMyu
XTHIlXKKPjs5YVxnRHHGRsPPOQEUgd6o2xOrP++2LwkOyzwlP8ThEjs4IcbFORQ+
2FrHZWLktVy/dtGodTTnBYHvfJAHscARw7EeUuE1RcRpExiMOH86BfiH3tUwk484
TMI1JzX+niDXQxjs0aEUK6CJ5f9AAOi2tNxgPUOEHvkm6RpN9TAcI+FgCJmUhMC6
VSRUrG/2HfrrXFSf82NTfgEdDGMYzudXrfHWEGH0WhZZXt2Q0WTwCg3BT1AFMVPP
zHH2TOHDDM4ZAA+cHbyMlN3DXdP21XFgdr83yleIcHvg7YsZ0Vye9YlIXK5OxBZz
n5DiLfThxTPdXkk7gENFbERkd0eNc9WEluIeAwQmy5Be9tq8M7/JrQf5zr3I64fx
sCtn1xCbYQSgXhlo0t0PBXPtZisNf0+ReEugsiBvFa5ztq20L9dx48e+OXaWCcgm
JKu0AG1QcUusH08OJAUvDx04E22yY5b/CwbMuZ/zBWuvoTqKs2HJHoRt9dnSpjCA
W8/DWP1h5KsJLHMrar6YGujPZxk31n/Lg5JmE+CeWPrmR0/TRz6j4z68OVrvsA2n
skKvZUdgptFA7BFwn1iKjWrvWn43Sp2bL1fcHWPK3bvnr0fjFB7Qh/x58v7sZ3gk
1G+BaIJSoPloMizR+JCKDn4oOrQLPVY5dr6XOnLJy30SKifWIqcWZUo8WoK0cJfo
t84XP/6jIWfUwPo/SYBKhYBxZIUQWL3rFaMuXa8VZYc1TyDkiBbFZKKhAy0OImod
J53jrNDM4SVmS5px0emt23DSW2ExM+g0D5A8ex9U4woRWLALq2PLmDaOn78ToR9b
B94H32l8x/9SOFYmcCMmQHbINie2F+/8nBBqGy1G5uvFsz9+ROuinhxMj/oZns9t
/IcOByb9RKd1HmHcn7e3jpQQLuqpM0t8A0Ba7wesRAzAYOtXCKcfGekVXidLIk9p
ucpZCmPfPbAq92Jh7JLuRVr4eylhwqsYIZayy6jyakftgIyycTntfgbdJHl8gLJW
4VPgfnyfblW62fyTrqMV/l8zX6s4i4Abc4vyySL9ZvzxEddNyvD/bAJBPmS0rJQ3
E0h+HJ7NYAEVUeZ1qRHO5MDQbwUjSj+6oEsdA4c99V9pH+bxpSA6KNK+t2jvoori
tFBekljTiwloNJ5ubF2AB/s82Zb1P3Xz59TcMJoANijhly4FqfiJ+l5eTmmrfRhz
19XlNFV+M8x71VFPPnd1LUeGu7D1VGLKFqr1ggS8e5M=
`protect END_PROTECTED
