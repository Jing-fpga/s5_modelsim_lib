`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yfqIEbu4WBc11+MgKnFZjFLh7ZnaK4H3kMxYHMgb7ARCj85LrQBsgdFADTCreO7z
PXHkh/E7d3geJxh2BvKxw0XDnFTUl+0RLnGvfrnuYoQnBCj6TIfEJscPTiOXSFVi
bDZFzbNL93b8waBE3G18xSa+dbBkA2fK/I0wpr6sB3ylpirDV5lrI8/1yEh61brc
OWMvMZoMwZlCtSCRWmgJAYd7wv8D1w+gLqgxyRafBrmcmmWduwfEdQl4UrcBq0ZO
2HMiBuNzdu9UjQmpXATtEbA66TM+hbuDPtTUYKMuN83HtHdvL077LLtszP6pOa58
NEmRJSN9vEWb23BSuZQtV0GJazkU1nIvQB/tJH3G7qXbCkDHBRkeruEB1VnJ50+X
giLzCVdhK0qlRsBLHsncglT8cxDIPN1rxYpO2kHwnAwA4wL521fKeDrLdvdv0MF4
X5+8pOslqttES9WI9UDYwrk6+3//U5xkvgQFZ5Sh4NFPOmNPt/auSXXMaNUV2x+I
z5cHr8+fmgtGAyNFz2MldCjXomPjE/gnd4ybfUU1AYNu4SEQ73F04oM3Uc8tVPCm
Zcgg2NpceQnshGnbzpNS+Qu5isCxkTCPcWkoDyFU+ecaFfzBrysWH/BdNL6v+6cc
vUzKRlrN6qwv/Vn7Ppzevc7ayD2qd/7pBTgzOAzW+7ecXJhW4A12EFPBccg6T73k
njGSFxywhkLsg40b9QhXRnxX9MPSb0gB8QaA6vBwbpighF/F1jNPzsB0dhJGzD89
yAehdUwy+bdFqd5zSImoOQz8vgEo8rYhS3O4oADLFpNvuE87bMUX5PnFE9j3PYQH
jE83KI8Ely0eP23O49hYn17ZJW0hK1RpSEW7g/qR/BMhgrUfn/8iJIYrN8OKtZK5
e89TIjWmk/TRXMjnq1DP2InDKOCIpwLI5LTOoCh3MJcBFmTMk8Ay/8ct6wDkYBGF
R3mzYUxc7pVVy1j6XHIkHg6Z0G7jxZxEYLrfVbkNlf4r/Pgd34Q8FBR4VDQ/Sbp0
3h8HJ3uD1GuL2MmAzI/GiaVZZxMoqS1f/JgImV9iapjeICIWANGUlo+iw/0YFCtL
ZoR1KIBaNrQdixwvr3rcwG0DCUyE0ggutAmC3VVJ5jPByqKSL3sK4LtzpHai5lDo
Xqyws0yiiiZBJXHtw4O1WItr0aHnY6nFZ1XRgiO3kftLJsmtEJE0O1HipCUn8NRg
+oXstsXe27uFPwDKRUSO4Mw15vudZewEUVa7x5ASmbrPLTdzF/UxLoVS+BZg4bnQ
1sNAibOLpEROv9CiLVXJ32shgxANw5TMo+FXGjEVXirwRj1Jria5mqHl0zKtVutq
ltkelP27N4A7INPLLquk+R1+3GvCQwcF0sCzQvZDGT2taL+4aO80QtyIDt67yDzQ
nkvguGNguDHMOQTv9qbaVPLKjueEMyv7ESH4LxCUQaNdWUbc6y0o2jqZyADeIT4s
7Y0e4rd/OeomRniV/d8t1t9wmUZ5ea+HJR7CWHopOmd6yETmpsjxg/UaJpMiB06b
ZTwAb7sHlrV4WZ47H8ZdEOAFT64l6kyC2J3Aw8VRWWeXgcT8DDiPTsHXG28NhlS2
hoqmeHNaB11IMJ4JegA71TJqcukgMzQhnGH973hpbNQ5zupam9C4cz6s+bIB1F/x
OmbpMdhKfQJVSJPDvHPmcqWxTO+HsWOXBu0EXon1h4Jer+/fM1QgKO4XeFQnKYps
9wStnlqs3CFFQnATQ7svUan1wwwZD6SKPKS8CHs7RD/C5vv1Ci2J1Z4aqFk0wStR
n8mE0E51NiHDNALq+dvVzgQAQf+AK91V5qtkKbwp+OVBMKJEdGuslQd64J1YDCl8
HbUcn28ks1OAwFk9GOqOApbLb/1lNYmCafo8Od6nCMG7nNH9HEkr4I6KiIwacJl5
w/kFvIBgxlA0kovn49g7QABTgUl7idnOCM8/LJd2oWUTJsVaZJgK9IDXAWGjA3CX
RUvKD5YcDOv00oc0p38otN4dCMsPZ+6taCUPXLZmcZ0wdYcpfoxKHuJQCT36It0K
yiOAM37PKUSU42cpvCF/eUvXpNMmUeGOEDbtvtNv5Ut2pGWXwHQ8fEwmRC1Gh7kz
oAEQ317w0g1oACGt+44XXFtOyETTq/wAg5LvM0rt2HIluEnXiIQwBLJQFGsdHEZY
W+oQpbS3ZbrxVZfrWSOt/neffQHsQCMK+PYZAq1fV0QVnSL4jxUH4aX00jlxHqPH
byxvpMzJiiqblGsaAb9Xqas5V3WIuUh4ae5qAgRvEw8/4sEwEnsUB8GrNi3z1yhG
jZ7wEBIDZpWp7ZCi62jiv/UD22RJVRKxLeyrW10sxHRWIj8oNA1rDggxYoTmCaNS
Xd1UcPCdWdy9HiZxaE3YrBSyH/91amB8LWVTQG4/+pWUitc6iK65gK8UcniSHp4/
XdblbpjtTQ5kcOHdlYogcRZQCNoFmGlyCE7ziUVVJcX6dnNgE9KbPXKVjYt+fHuf
LR7aa8IoYwrU3CcxfS/uIORms+SlhGRE3DNTVdFPGwKVYW1zS8hZgokDmqsqXHu3
zMpGxDiBFmdkN7g//7gENu0X8gK9A3pt/fqsmxHsTsLDT/Zc14eP73xXcWDFuMio
seHnWPQI5Ugbmip5yXmiErhERsas9awWPV96vho903PKEmvF9A+mCbuSQnZyu27D
qmwO5R/dRB3muWY0yFwnN3Eg+FLkg93uD1Xyzv7OBGgQlgM1GuwfI2UqdhuvD97a
Fx00x0eLbDurg+3ZgCHJOuRv2wPB7FlFI8+iu6c6cHkzBsZ2P9nw3VFugipaPL6T
T77SgsXRF1n7P3/Ay8H8yfupml/iZXXdUBc2BP8EvTbOpXVZSvpoJAsupWGvNFD4
MpqKr2PGQcprIIw8T3GtHS6P0bx0iD+lGJrOoAXjXcnaRXYrSA3Q3Q7zPsH76P4W
9tzmd3gHnOAliNfppk5HBjbKBOVpaIx13aTTOfMr+veqLF5sc/IZdFVd0wtK9bYk
GEM2Yjxq3EuSXBTuoAA+/Q3wkHFWJqVcoE6db+qPjo1AaIEfyu8aviL4r9kBBX+7
PSZwybWREOX+RBULS02Cj70In26s+szRaWuYNfGQUaY+2XH1aIxfscCXuftN9f2l
K80mq5Qdf8gCDyVwQR2ALJ7HqulrZxdAnvMApppC2s+O8DUIjVat9+iZ2CwPTGsP
AHTCXQVKr2Doq3Fg84NEPhz58KNkdxQO3CWrnT8tVQqkP4zH8jdH+elEGxEExqJx
C8vAqJI2cV8Ov1SV/9gqlKWIw/fDkL1KGasxxb4J6ZRsbgTYqLApdhqyA2Dy4QVj
t4rkqL7LKSve1OTofdkpJwcDifK1zvD5f/Rx8kys2vnttnM1mmQn6ThM/K3mgbnt
GCbqwl9kbRj2pw/M3pFrrmdzn5uJg+cfO8KZEppkMYe4dv8r3xz0JlA+chuAzstC
n/BcWb/jWGz4GiZhocFe8sNaQ2gT8o+qMkJM3t7g0MlcvRUyzmD/SkxGXV/18ZZO
rdVdwA18tqx32oMf79GrqEWqEiBuwyoXiGOVtL04OHqT/1pULIER5x4F7D7w/EPQ
FJbsPkaFs/3/KU13wmlUNamimyr6KVS6Mz23AYcnf/VfFMsT+ZFXCcFf5DB5ZQsy
Y6a1zY7MlTylOC5WOr+JOrwXptwYW+hSs1Iq1PdbsKaQ9frsc9C/6MJyp6GjJnNu
fniPYvYcB+YO4aZQblS7MMjYdNSTLHTM+KtVJBftu3kZXTDQjN7TbPZZev4rwgsZ
rx6W54HA7U/RTdm5NdtlKb5wscb+2kvf9jmdEdmSqumrNDkzq+g7rJZsQel0hWSc
6pvTKraN4R4w6A5rt3nIWO4aeMc5Rud0cRTU8J+u4DO8Xyn7qJBAquwiUgHY8VpX
C3ptz9TOPpW9V3fJFMqgNB/sOG/YBpvHL2o7Te15tNoydP6oNawy0Qc2lmCeovvm
I35WlTgQpS73Mg8Wbs5Cvq/eo8XKIbTMsHzYijlcv3do4aa3DD9lW8Ofnm5uNd2S
/CwQ2S0x0BXrNemRUUUm5uuIlqKYIEqgjHwaNMcPex7y54KQZBASmIJDL1Wu86Jp
nEb4WETq/ogdaoucv8z//aPVeJEdv0eoq9JJNSJ9H/4Okm25Qb+HW9fbDm5bG+y7
Z+CcZX354Z8TQrPawFqAyWOQ65kbZVV5qAkIwqqJb0ZcEdSqefaEbJmsgG/IxKk2
lzGN/77wQf/fmyW6ImoTh04JUGArOt3LGjp56lXlmC1O2bMSk6r1XDpxzQQf8Aez
aPc4yt4cOEfwLQllFs9c2tsDusqexr8u1v6U9x85qWj8yiF8mqulCfvF2plAGtM8
EgbplrzAgaZ0/E59aixp2angBghmRzzol5wG+v4a/TOXEUir9jJcYUflMWcWEYjd
/0leQA0ioo73A1gGmET7gySzpSyQr7KMAIE+Br10YpeB4tj8heGLkm6Xrz4JSWWg
biY9tAfpmEmwEesFiizVAgh3+Q84PGPPau4nWidS8Y34zxVnnpfwDg8v7Z0GHWKR
NlsaX4prktmsRInR4PjZY+8QnY26Yh/cgaZZ1uQk2ahgqy44EUvxQ682kkm7A2W7
UB5jlzE+SPjJVihdDCIn7tmJahXhr7EnT0VdlUNy0AtsckvRTW0+XNakGdgUYiwz
wd9Lw1OTceCXuu9fvscl9JZCinmN7o7zdfFA8NyTwu0JE7sJrwduq5cZaaHdaYbr
/pNzq+dlTFLcPtlgisLbRW7cu2Mzq+x9TOIWq/ETOibzUdqWUfHv263B97nod5v4
8FF4zJC34EslYl7hVzglSUCz4IrrhvD9mps6VfKousjAkd/ST4AhWIPNKSzPzp02
QfhSeNQjdD5OauJhRuQ9dRnu/Je3B+Uqvt9KO/etF3CGrClarPP/ITZCzZ+ZvECi
cNdsHn5a2kxn1etwuCE2z58IWbRRt9DOaiCAr15hS0fBNWtIMaaxm/ivEyVqkV/x
Ql+3nRBokRllrthXSiPL7rEHWNXbyxtf9fBZ/uS4OfN4cGqbcgjaBkpNELAN9l/E
lhlI4oBGwIJbfn6YPXM8jIoH34gwEzfZjJpgSBtnXZ59nJtnyrYSpA4B4M2fSMCK
fw/ZCl/bHQSTebwdP1cLgtx0UGrS1inkA1UqydR59Bc=
`protect END_PROTECTED
