`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0IBrZnaSy1KA1nYuObgjERbs0JY2OsWe67AbTp0/cRMRIkyc+buabYLA0eGokjOM
npUPitevdB2alm9apOzLPOUwXij2CNKwIiHhDMQnF243Rhj/4uPmuAOORfl4RFKZ
NdR1cwGW6OwFA9EO+Hpv6Y9/iPNiq02InsueO/ue7pwsDiGnwVjpPOW7TcDSkDHT
ebOQKum0cvfny7MnKSHr3/Fzo1DP+5yGDdM9xAXbDNgqj7m0omIHBMasKJBn/rpb
HmgM4xfoN4kV5AwqqZJrGhPYUfD8fIqNfilTKoNBXQLejf7CGv0r4FAaBh7ujrvA
6UuNOLf5FZMa4FLfnC4ptfxGSCVDMARUCWPn0O77hWieuoebaQ+9VYkKfPZI1GvW
LmJrkyKzf7IWwjYProWoNozclbyYbZeE3HzNVm+0Crv9ij9CzfHHx4gm6XRCC/z7
Ps/D5Nq8uFTJ9QJde9Ko57W/f8lbpI0OwbjI+69ayvSNDeGRk4qlxFVPfUcI3Mdj
VsgGc8iHgDnKmuFD+E5y3VNKKXsi4hmhL7xt9D8xrKewPya0zQykMaSNv8QPytzd
dBLyqBeJX7TGt/8ApThebew2IhxH+hliqRCtSEgSfzJcYO1g6rtYBSQQEsU2iUqZ
ZaI2aNNCaKwe+MGUtR7epObYjl0t/FzL0X76dDFRV+0UvF85+Tm59TBcnUZWdG1q
3RogoKdWy+JrdT4Oq8DyKsaQZVUTKM1q6h4MPeHheoxBlDghwwjN3FajDl4F+wm1
TsZ8dffBnGA85y4FiTryrRZf2RbMM6Con3YcmdGsoX+En0osVOQfeUTVbkgA7qLa
`protect END_PROTECTED
