`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mrKrwesyQlxy9qDHFWM+cyNaZ8WscB/ccs49zWubp1WAMuMCwFQLdzNeB7ClR9/C
SUwC3Xyc/HanlcKRzrgoNT6/AgbCeZF9eykpD6zqSEYc2d2tZ9Ov5TDFlxI63nDh
ozPV9q3JVlok8JbCEWZIiiZJYbBqVJalbHub2vKp4Gt3Uwl/SfZgcKepgESisUe9
dkGkKRA000WI/9nPrMOCmmv9XFmNQFgMsdFmzUWEDf/eiX1xCsAww8go192RQnJL
IOQjdeFZrIJipgJ+F7nMXcyXWA5Y07k2PeV6tZlzg/FZwslB1Dn5DY5N4e9hLJo/
bh8iHdbg4sTNzijhMwIxhQV6N2FDIcos1IBpu7WjwuE4WkZOrc/4ulkdQmkhhpK+
JQOOromcR8CM/mGhzX1AMzY95uu/FCrTb+J+/+uNAjmto7hKywXMUphkO/iUsN5E
9tB3yMEvU/TmrxYoyTtEGloRxfNFA+7cqBMIkcUKGMq3OfLX8PzridUEoS8LTnLo
YJqcL9HtmBwkAUkCLJGF052UN57RH38VWlCOoLc5og/vgvIYMFGLuKiMCJNg8CsD
DhuWNEqeVjducE7NkTzfDMCsc3svRZVUQuImnFPmKzxg1uYAgFxlQI99lInwgPEY
0XZaPSNSXXHmd1Zdxfj7EVzXXcumMgU5TpO4nV1kGC3u/mmZctpIHMG085+u7p/f
NyJfxrOrLc0tSmtc71s6B+Nb+tMqrk0fCYIXicrFTmvdn5BmeKIrb2TubSxP73F8
zboyRDGqQOu8HtnAFN9gpjg4lDFSQjuzbwUAckiQgCi3cnEzgXi2AI2pq7Zspm5L
`protect END_PROTECTED
