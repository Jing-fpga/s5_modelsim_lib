`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V7yVSlben25SqPuEOXoszYNYF4YthT+N9c1i4jj78RETRpwQLoRPsFiOmEFCE1hB
st6CVDrMqciBuqC/agzkiQcFBUedQqp+gF/sGD7qUOcIxhWqNkhnjjrdZUvUGO22
U96oHO0/I5FnKfqFevMaQCJxfJQ8lKXwy4j7qfYuCC36dmLbuKZK2SvcynZ5Xfqs
7M3zsclrb/wWnWEsdp/3ZAds4W6kSA7auQdQszfHb9JXCxuwH/siDdBf/Kb64EFP
vEaXZrflIbuveDSKYyyxBANo4m6V/Nz2gTeZ2vSiVkXxC6iNzoOKHu/LS9hIdkVO
jRfLcqq9Dft/qqkw7fOEbeAysd1QUsTvssH1lyim5J282KMf3vBQqeZFCbN/czNR
MlSrXIMvmLbHdaJryG2P+WxxwNjMQLORE4fHaZJBeGPqnLGSs7bLgGTBVGdzVm42
zgmv0Ydigrp4XzyyyVaxvD+McUHLJZmVHvxaHpxdszDC7JAeLufwkhrSZwYiB6lJ
vL4m+OIwz7GU3CG2yCF3Zsu4qNWzRd/BhdYvuK27G+U/8+PTLjCOjuvINTe7qbTR
qg+LJidDugtw73xmYJqj/AvweGDI3Y0ra9IjeoA0cwSKL+g97gLE5ui84YwneaGY
a3Nnjst9JJ0gDLjCIDFfiq8FLyJL+C6wJB4SYG/2jqD3DwoqMRl/NA0ekVJbbAUB
8lOkURe1n4CsaUEQ2A6cE99W+ipiGcKMvZvEuSJ/Pd32Gn3Lq5ETttN6QcFtmE5t
Q548XkHUUvdF3vJZxPSOVC2GISF7AUhT1D4g6mnpVvJuFh9/Wi7cv9Rsvlc20+eU
g31X8yxq8324i7WHBXcndSCq5OMYES4tgV6Mgp9xC0tIEWP5hRMSXeBV2H96XdY8
oSp3HDth6uXuwvVhZOZi9UKpQvh9/o+Pr1KAN3SrUt5j9a580DZgQtDEiRq8CTLP
oY6v6okI5FsRIA7bxsftFw0KC+P6PXldP6Z1aN54TXdJppq6dLXg+YadKjXeG22L
eCDEH7PMy07FFBudZDCAQjzuKVxzvRFcMEvQJ4fuNVqb+gXcMvmzpnRnxPvA2w39
JturKniiF9lwSTmInA8at9jwe/V2ADN8TrerNnw3bEj3QP2RZZLGFBqdfDhoPfFz
3ELvIzM0FBkC+e2Swu2vsy5yVq1BqiLZAB/ila6YrGdq1BdDrdC8QcEz7Hr7SywE
tZF9tE+rLF471ExBMviN4eRYCGs3GE4LQcFy+8qGMCQwtiOQ8nZMiRYd/4IeHpzg
QOolRa9bhsCREMIykTWTdwO+ffQ+OGrUMW3OAVwvCaqEuYgH3Ecm1kq30K2b2My4
AJmfvv6PjO1Z2lTu5nzrBlq0K8qcWzrK/7d8VnjrpIFBslvjt8lF67nUAQSEd19O
1C0NlHedSfBrE2O5dzMphgQ3FxDTCo40QFTuCD4PCgqVEexsbid40k9AdyZTN3qi
gQ3wyKGwawEV1TG0X8z4dMbBaI0NtME18HDd27ZMe2EEf3+HfxlLP15LAbM4vC8k
fZ/eZMR9Z6Zhbc/KxTecybcxg9PACoomIyB2BhCDn3jgVXJuYeDpnspchtbYQA6N
CcOwTaVYUc0jxfbdVA+dTush6/vt36Q3NlByhreOo0ur5vuqBWkQNh5gV7ZEHkCS
8+ZMgVZ+RKIRpc5Ns8OVftT9l0Yt3LFR3SbwJXdSaFXA8vC9PNIlY5N0fPdBYY5q
WfgLiPV+tlFghOgu5gOK7tcDHEFcz/4kx9+3qoEVBkHifFED5O9C8VxP/LpU0zpH
vDU/CKF98DdUR1BLxcVTC3+AkXK4IW3F1OHjEsu+jl/Lmyhw5pWPgh08nKOam9RW
fEK25aaE3vBjfYlyscsC8Mn9eFlmogjCKuNyng8ZcdZIFXz6UIL/QF7AKZ1Ub+ru
6BISqzpeN2sKLAuU2N+RJA==
`protect END_PROTECTED
