`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ndUigJ0cnFkjy+J7FFLJitSthKQ3lk3jzShJfYlbSn5vSWJVIyOXb9twnocZ96c6
7UYPVIP9e4lRDbQjR+vEZd50G9fFsTuM/z92sv8ZwJZDrUhXodisS71DovYbb8TI
7o/YzU99KKF4Ov6lA1ZPxGBidTxdJ05vXuM0ZA/WBi275wMcrUos47C2zk7O4tUy
fxC04wej4+ulvc0oPyB4UJ2XEU4DEGEc+m+72h9Q7S5lZ0d02uO+kFGiUoSaiVD5
T7tKoUgDZnNofn23gGWNbau02get3V1p3+KNVeRW03BTV3czZkIT77idndS9fNDl
Cr89k2HmyVH6zsPeK1wonMOzsBb+hx9FWFoenof+3ANiV+kQ/clVimtgpGAmFTE6
Qp80E9kh+BGLMeQ/XQKXkm67lmzHE/Tsfa+KnSi3HwNgt4adyxDo/tT0fw/gh4EZ
Ta1DxvytZbmvbHjIDubFs4Av7n73fdoniB/kz7BfG5Ldm0qy+r0UpTxBpAa+LHEd
8FjXkTOftfuTspXZsiGCchHlFQ2+zQQPydTtb4Z8JIAeBT4VKZblY/01Wls5Wymh
9NqyIVGMH++JJpSbFrpYTDUNAKSuxRMEPoUJ3Yexr8tb2BN1YIhHZknTmjgB10Z8
+jy8C73QlPpZ5TkDiLX6x0nCt3U/3bA5xtzAPVrX3FGsEK2R3Ea4y6OepKg+At0B
XiZXHvbQcHVWLe/tzKffXicTsRkfhgEaJ/l6MsSVsDKJgZKEkZojk5Snm4Yak45w
fxy0XiuBVJRBsjDgYlcn+a8qfcDswE6Xtm7vcoKi+l/fAd9tn9RpqBWNBS4MR71y
vZj1OSFRGBluID5B+Gro5u87vVCRQ+NX/Pwd2x+EkmZGPt6Hqfakh02Mtxx3Svpj
BRI91rtZAf5lxzJn1r2nP9TfASOKhq9j1wyul3PLwRaXk6xEiGoDij0UFg1FM5SS
wic+JM/4eJGi8C2R1VsxTtLj14QJFlIkoDpoDwCheKOrB/DOvUNnOhxKryeZ2R8K
ELiBt1SQSlkb2qkUP4bjW1SM6KOxQwtnPDqYvuT0aExMXvxUZKvI1XadrMRqwSKm
owc/CaT2/1c3trgcjmw+UhtCOQmNTgVBfiO49H9QT2D5C4/tTQddqeX3e78QuX5P
ayJbC1gLbPxVY8IbORpySHbPAriwooh9ggJATzMXpsGVRDny0hD6ReFaxwSHW+Qh
oO2AQYoJfAGhecWhWXgxRTnPz/J5z+j/HyJEUBQdcThftM0cmVY8eSonNyC+//+Z
qDWkBcB1BH60yXJ18r3o/lQJeaeK0/ZRxaEtPuG/FVdl85K1jvjsNaVGtd6sg1AV
Exe3D5mlhMWx1+3xhQ+kOTzB8GRfqdTJv/71JP0h5YBLFe6TWzj3KJtp742QG2mL
Q42WTqP7bm34FIXZI9R8SXSeXu8s1LvWKQRWZis9d1rhpjUS0IAeXwfmMDxHz3H2
3jZhzLUK1XTza8a//26skB8NwshrXz7/uFaf7fZpmx2sE6st2rxDJ7jXsjTmSmte
I3+xMaNN+iD8xa0LzJKkVujTPVo9DaDo7yIjsPOCjCpjItf4OLmr9Qw9Fcy+cfu6
EaRW9CAW7/ZCGua6eBA5V3Ii0y4iV5eggs0m1EXU5KA0pK+i5UdftFPjijn0HyYr
yfeajViDMfgjesq8junOP5NttGyDrM8Tl4MepTxp+3mg27mj/cA+xYrQS4q+JDxH
FDc22fdPHuP9fv8plG9ICKHW6nE4ptFFlku+Cjb/tTctHM5BFJnI2QekdbgemR6q
ZE/CGivVATigc2jrgu+yHK8rBABtluADl67lXZe2j1xzaokibipDtFGb6T7Tq6gr
4M7lOHlt1YhayhKr3QU0vpPMHi4kAgQOERz1w2HgptI=
`protect END_PROTECTED
