`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3cDWIrgjjCFIuwzRqU1CaBwakW3/s35AdNdW9EvPR/iKF9DmO/Tba0/VsF3mN9/w
0ju2niHRI7sr6qWZYGn5XmjHkQkc6viAFU1ciyeeBhb3jwDAa8I2ihF0BAHMkoIM
fq8QdGYRPke8WHqswVCMLG6oJUQ79lgdnrSgM3BjNMtBaJMEMlrDyiOKVo5q0Thz
IC38fBxr0lTG5A7UY+zZafMVKw92yJ/7awHD55IiUFYJ5aCog9O2SaLFmbGX9ySb
uk9PvznnGlesRpAx+OKNQ092LbhimOPWZbs2X4veFkUJxSU29MoCCjSVyk59j/P9
w+o2Z4enzgmTTYf+OzikClZNSJNmi5EsmjqCQNTgTYylSCnZdx3UsgZzhCtqFXPt
8xIYWiydCpByLw1euxxcH1CF9KRQlS1OVxbxyjDhyT3LcU0uWtMywOTPDKKFGEZ7
PdZ3vBRhp/B+zE4xTnXAl9MX7LftnEO1Dp7/iUOCUwpZkQvdka0cCg4VOuw1Vdn5
9RTTltzDBsv06JsQpcXYxhcf6hmCsRoYw9O0jEUS/cKLumEJrOWN7Oq3qf2AJ9DW
9q9h1eUhZE87SyP6PKz31yJtD+a43ot/WecRp39swOvN8Pp2RNB1xBT+QIFWfJCO
8a4HcmUZb5Y7F54MbJ7Oa++m7w155nfTzLdAp781qfTMEH2pu60OnIL8unk+sglN
ya/C72+PkLOr4NRF7gTZYO25W8PByYT3PM0ezs8urqlj4KqL/IytGme9/jxu51EJ
ObP2a6Jf8CMA2Ok8zemxriAazks8xuNIfu7B9CUOlE3ceHJNpzexjPyiDDLilpJa
nZsRf72XRgyzzBiZKLrVrsz4Twg2NBlauNhoeK9RhSvDeNnMNCd6CJAUywQH5dUW
GdAWk9gL0a3EyWFqsukOcaY7G0PEnbcJiBZukObSLsPwkHnmgio8+larDz+AsxAw
c9vGB1Wh8An7isj3XGF2fxMKj8Min0I/BunV/SJ9Ceu690otFQtHo0Ska8HKEaBd
0/84UhLxTHnMc5Je8C2jSg==
`protect END_PROTECTED
