`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1UT/6o/O8Lm5seCsrQ2674rn5QjpG6cf3x6hR+3fEIpNq/G7BbF/no8WNr+Ye6qE
hfWrhABr3CoD14zruZ1bBKuUyZrPsDQl2nYYE3F8/qmm/UhwHzBwgp2Qr3KIha8k
P7qIVo9aTrsILzAMl9rqICbXNTirK1GRCZIS5OnpLPlbaZb5fEQ1fM9a8fgibL5+
ZhnpUw2ehXR2XyiqCQFQSDABrLnv6kKWEHYd+4bLq53o5RxJ+fhVhgDD0Ev4+xU2
07iOthhO+pzEpfi8VOhehfWlrEhPoZBUZscdL72ICyz38Uq2U+09r+w9TlEjYWTv
sc9zkclhtsPMJsilR99ENpZA8421GnZwHY99/SJc65w8vWW2Z99pkbeoa8BSyUIi
KGVvk0u4FPZWMhTNc6MKQHYghstCFJzvpTYr4Gco4IQp0vbdO7FYCAigqvywBVlN
Lfjc7E09JXeyC/m2900KAzRiVtb+7jZX+k/X92YgDu8t3ZujL0aZEgjrvD++Svts
tzwcODAQtpgFjrcQzFX9O6j8jSzFL2jAA7HwoT0U+IBn338JuNNHyYPgbhXwaJEh
EOE7SvT1LkGKPW5DcQUbVbbJICd6qvfRRJMcVDPNBfL31jN8SY4qu7X9ygjSsHmi
+rQQlz7aPwLFDnnMyoJtKmjSCwT/7qBB+/jPvEeqROG7mYGZ4F7k6WhNCXrfkF8c
D5dVf1exc6C6JGbYuM/L7mfaXeqECUWs7S2CjGy4sWzZGJYyUvYbos+kEMoP6lcc
mgUuIO6MepOSIaiCHyrwaAfXsaQCY+5qT2/i5etI33gmBETw6y3qfoe7V4r/opAq
6Ptp11NaFk62EJ6h5fru+6eucu/hAytaslPBo2r8rTfG1ScFQ7jMF8yuh66UZGVp
dm2EthZ3/VToLWFXS+5OgIt+CuW2Cn+5/PdS8GSSh5/PLMpvtjnAYvMhoyLHkTkF
kUEznzUVDwcqCRG03fo10BhBwWV/iTN2ntizLApe5B5+aCVIKhEK67Ymx/N+eO/Z
DGeZURSxiq5KwPDQKew6+spJJ1Oe1nWzw4wqDW7c8b04sv7ZNG8xBgjN1fwTPjEB
QnQOTnKhluhdf/jMFvERnixRVqvdHNR+YUURDouhj1tMY9uI3al9i5aQRNPtI9oJ
BRtBAliFQTs5JxtASX+dJNjxhjAVT++SCeaGrE9GHX2ed71La+C/OxwbCVKKjmx1
jm4vt2LxHtTiXc215O6DeY7Ii3r9lo/ljmH2HMz7zvAi1auxIrFTcl37vwHOWwrn
qA0TV4MQIJi2AiHylCWG7V40ImRknd4dnh1l5iuz2sv/jTHViK19/6grJfTyMNgt
dx+xgLSw61h/pKoKNIQ4IOd8MLrjDAGxtyHP063R8puAjCHj3rq/KlMwGGvAgDZl
M3KHxPrphyQLXFBA/e2xN9eWIYYdnh9OsyKGQLdE2wiWah2Gs7mpJH0Lhsx1Kz2r
HoYI3ed6tnVHY8jgqTEwJhFeBHZcaLeGrTCQEc3CV4iLHJfW2Lr8DLXdxHSQyf12
jqBQ7xrfd+rjNcxvPhT7Lt1xlBCNvHj762OTV6DKucdTPlbqefoSSViSCDVixL8e
mPjq0SKUpTuSj0+QVG9RAiG1gWhAbyFPeeDsbfqDzvF5ucovVbLTtHlLebwsmeii
AOz+E2jLJBi6bipN2iAO12FettKIIBbG4YbNPM8kVy5jsfSK3LGT6dIN8oWXfI3v
wZlXCApO1JSsid21FOx3r/ea629Z2HWbOTXHYMvhIBzTQvs1fZue5lTBcskXdkG2
6ovYXhVXL5y25OrcD+995DtZNk8AkF9YXBFt7skFwJtpYgCnzPwg5KpO6ZthEwuY
8V+gg0UUXZfb+xVKHkyaoAn7yC/VOMngywhYtJWoU7WwEJAcUJ/1ziHyP0OPdDwk
DkUWHVdZ4EUhbpW6xSifQ1Sp8JUMq0KCs9oAefz6D0fDCUpu//4GKIigg2wtwVV2
zuw1Zrew1NpEzeoRirL0fsnZ9P7PpR/m342LDZkXOwBymamB1edvlZsJeOyIgQc9
GwxuEovl5Fmq64Nun7DNuOxacCVOh1ksVDR6DfpJHBQKhH/NJmysLvUR7SNA1DCB
GwgRVKoUYa64/u6YKlzqEzR8HBq95Tynjy2iW2cUScDxmOcwJ63i9DTYHQfppLgP
JauGlDdUp7vyRNqu/uME9etOU1ZpXC2HvI0ZfEFOmuRMb9E1z2p5RKOQFYR3Guto
z/vZ+Cozvty8myFAeU8mhFpx4zWQodPXgenbBkjKAbdjgeuyLrziFCjAVPZdl/rd
JQpZ1TmVIpYth9pbrVBat3zALgag8NXLM2FeUvCxFdS2DMnpfcr6NcmRNlXiwDYY
4P3uKPqjbDqkqgiEHA1cPYj7x+4wv+Od5mi/3ehe7QZFpwqmMZSocG3zhBGn7C1B
Aox2tP8mnGju4hCRvnT8XyxrgdFabjQJELga4H02KPqxgkH5+VRI8JGqMv9lcVUC
hQdc5sZcBGIwJDSaCJzMGeQb6oMCu3TAht+uBw6m5BBwZ0L1Bs21ooe/qXQhMobt
5slani/gAaEamY24O11I+um0N3eUXC+69Upa/RXvUF6mwM5Bt/WkH9XI/g6pXEvi
ZmSAk4gYhUaUNZC/1eGocKJ0yXXHDfQyGwQLm1vIIbHOE7gLqVTfWxA8oJd76RLz
T4D7DaZTnEukC3Vr7tu3VojLhnvgfFCwUoUJAhw/hb+4vnIAkEl6Z2PxUd+GoZeU
dgXPRQR5ToaBMs+v1DESO1D79K6N47llOLtfbVczxOY5HMGFRK3FHX91HbUAE0gN
3+xfEcUzPfMpS6TQqgZCEh49FdVlxQ/XKx0kqfmUiw6q/kRfUjuFu+/Vn1PVN0pw
CEYHULYcsJpdexB8QzGm3c6EjhIunsdrfH2+5RMRuZ0=
`protect END_PROTECTED
