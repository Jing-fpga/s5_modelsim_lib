`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l8bLebdVzLfWzP3iBQRLG+HwtB2X0kEtNvjeEQfu0RH3b0iRfXxr0kZ6JNbfrYc+
WXqO9PB1Y2y648wbuV2Y9d1ZLcAJP1pbYfOeclXzR69eIe6yPhzPIHrm/M2ILe99
tluPKtTL/w8HGj0UVLDhw67KsrDC38BaU8nebZo3b0MiKGg1IM9Uah0KA+4TDHWo
0hgd0wpjQe+lomeedkFAJ1ZY19g/FFE6Y3ybby6MPvCoqv1oa8Bk2FSwAPL/3Cl0
5jCMNx0o964VBHjtopGxTeFsordApLm6JnoERO4hlOFR2e8LKVOrgfRMHDIvJQBY
ko922OSOaIoldn8De522A3CNNInpSWxIUVSbxvbM0pzGP88fZU9POiS8t/Ghpn91
oKmr08NKux4PA/gLT7cAqwbq4ZXECsDgAkaw3rS5+OcEB5S0+fLKjrCLIjsAcjVW
fyiiMZwrtR51bp0xN6sT/NGe2p7weoe/0F97+lJxBJQbsDdKGXCe7LZFkyJQ4ji0
WrVBI3ig2IkO4y4l2sEQw7Ragc78k1SDofZmyekIMnDqW+nYFmfesGNX8YHxa5++
DbZ7RN6a6s5gqiurUp/pI0rUenxJxRmNnateaijN1DQxox+OAzGMFVesM8QsnBgG
34eMckwbKpSSeH/Ye0FQT8fCB0yvpjH4FPBoQZyXSfEX+FXrMdO3A11xaecgtrYa
VQFjZJO79qeio01T85Dmdc64WLMasH8Kv0Bkq1CVbNV/AjeDwZNHKBCud/4b/I+H
kfF970XEW+d2sz2gyeiPlMPTc8AP8dDmI9CAriZrjQeNfFfDF2FVe5f6b/9++CM+
11PgPbkwV6TrB+NB11zTtdZnNA6zxK1hvI8+FrdpBR+jxP5eG2dQkNVn51PWx0qj
AavhA2phV6AlM1QtQjCamZ+c5XOpcTSg0Ky+Q91xN9X3hslJq1f+LOBY1O94/C6I
CizbUxUaq3wjibFxoVKZdTQTNT+8sKOeS7WV/cWcI+j/l+4+a1XAlfwxqdGf7fbs
wEnuJzK4OeJnFoOuDRISzUIDYN5XjUEhE9WVNOAMoO7FDWQvuPkYJjM06I0SBvva
3gTd4mnJECmIwvh/M33KciOyPF1VM9OrMHHfTCoG4XRDqwDr/pUb4OZ//SP+0TnV
g7DjJwY2Plyj4rzhExcplhqdhc+4L/nJ/tsWZ2g45erbR0UjJWIy2K5z8RPV4bEF
yOhn9Hj7na7PZ3TXWJzun0LSDv5ffiHx/v2jycD7JlOMpBiWoV00lCbKifxUFDAv
8niLdolC+d1GMrMoRAK9wJIls1XKcIAKkFwupMv7qR0hQcdQd8Qmf0Lj5Un3lXT8
uKD5EcOu3ZbceeH0a25HDiEq6I/Wv6qfFz/oH6mDGFPgQyNAXl5FZ2Ak/nenY7Vh
zAMeVKkabe+Uhcp8BpKRvsPVDP4UI2QkkwyKczG2lAUCZHrOb/jYnilRx8J8rkjO
myPLeSSuD1L7wd55roW9+wWmfT+neN1929rN1/0/+sRQAxleaXBPduh+3CAkBssu
kkeifssmbrcbe/npim0o+rWoZ4iA+PfDqmHrSnvLBSx8rYK7MAVDcfzvA2pM1wHs
odfmKn60I+RQrVmqXUMvCy1TboYKy0nRapJ/N3ZcWiOZpNgXnrN8Cyr2egu3WMF7
an7dX4kNYpM3OrBuhsPrEsQs+nFx3UzQ+mTKNCadMVst2Opbvg7evdns+dt5SnWz
uN+67dzF2lPOSZeVo3iTfYNLXpp1CLXAqGNoy6oJJ0dWKpqeFEfcbvSyeBndh6kp
IEebGv2/1qFFE01rssJExw==
`protect END_PROTECTED
