`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/7PqL2ghCsFOT+i/Y8wgF31VgUjpDHkUypqTLQJA5mDIu86hhTXw9gsD9yGVclbc
5NtlVFUfE6ayNnxj0YY/rf7MMp9Hw1azrxIh0zM0dOemvJ6yZmAQyb+0PLgSPOLA
jFhfQoKBN8hz5TEECB7/LOwbuaJ4CkvOZ35xPCk+av13NmkUqQISl81OBDfHnqjJ
iuiTlYzyzlXE1Xx5uJFS05HLl5Pr0qGPHvUgn+zTQ0janXGCESQYMv6uF2B9ULfi
DYx4WH13dc1+FWZo3L4hHqd8rJ0vHZMAOj95XZ4zT6ChAdRL/xIFSmVdQ85dqreC
djs3K2ANHVBu5exmN5AanKPrcQ2HwbNTUJN9NoUseGiBb8P5+QzjcfrK8ZsheNwI
5MmxdGGp+Pv2m6D3WXFvDqR7DjJhn4XwnjEpgZLk9NENCNHYbgozvCV0Z+5VtyuC
ERDndTUhV+x6Krh1NWda27O8eLdj6VDuQ98W6bhTy78roy5YeVlkrhxvef4NvjC1
Eh6Fh3YookEt1o6RG5isVohqVB6F4zL+oGqC74EzI/9p8LzXTC+fztwmNK3tPfGT
DdgfyY5nWfgaeq+7szdkmLBcYYfo6v7Hd2fWzMywRlM1BKRoqUGsWKX7vXqJWxHC
I3iamdxAK1mGYfHDt5yQ60pfKC710RbYZVdYyzSAiw6kLL6YaUNDFIrxiQRAfV8l
AyxxHvuJPfOVgZpZDFw196HWQSXvWvOijgbcWXDsQX0YRU4TpPFUyW0FaHNva/sT
tGt+lQoEuMhaIRuFYNoiq1Nf90RGm00JFgWvgyB+qMm2Dk4E6oTe9+E4YKzXKJR2
KOCegVAFjagClVv/jrsCLUUf+2t2QHqYHJ0CfIAxhKAVx4WY3vjW1LZM30LXBupN
YNkd9+GjNVRuz/8+V+vd6jneOt3/3aUKCU/8MI4SKemWauZdrBhWRqH6k9dIOKo5
G0mCzpu8wb2LEPR2tvud9gsmt32yEpCioaoHoKa9NY9b1onWVNZGKkT7JWDge4P+
kmXgeDG0ZIjR+kzs52ND+XmVbAGYkIP3GWs/9b1lWmzL5YPr2FVMJYJI7XWDwbT2
2lExSQOtSVQYlnZRYsR1Now9WIe3ZKvZfDBZPVfAS3qrKaNrXfge/InUM+VE0HQw
jrIpF9knG67rBFIoAUrIPEGPu+rk0+myemgoK5Iz6Exedp1Ue6OULRxCEMyJlhUL
sndqMbbhf489iwq+02gUxNnMMeDYVkMGtP1oC5Va1lNqEW7xLk4NuE5o3hvefDCy
UyOo/Iq50Ls1/4saSGd9NKOJgsOVZVkmTbqmqoJdM4D0O4bPNNTY9CpqSzYQ4MKL
3wZH1lmXiba7i3QiNoofcyO7CrK+yNwIpnVZTHy+raQfa6w0v0dUqCzvLecP2cvk
TmODQboRoctc1b412JTd818kR4VP8EsaBuUI4VyCtRP4n1tI/d8Ewk25wvC5z8UH
VQnMWzIMUAZ02W0KhwQqFdfo00HDsM8E0yKtkibA3HTvzKucbuMVqaed6MkweS22
q9EmdCKEd2ZtTgXW4XSNs9dJWDZITkvBV9nQLQmKc7sS/GQvQXz1Ov0IaF8g4jhn
tI/xtpJryBl9RUG9cVO4w9ICf7u3E/FowhiprmFijP+NJElHfS8rF4kxVSQ151g2
/rHkHZba7wjwSzryy2v2y0erbPtzlxTQx5arkosSr5xRztDBByx9HceLQwCN+CMu
DojjPHY1Q77Mcfys7WsVXOecz1vgbpHBL60VgchSOtnoqPmizbntHuVBw0kuY2Yv
uXOM90VMLn+eAGN3foPln+nePYlgLd+mRkbhG8uXcTAE5+AMYuxoTX7GtNJw5Ffk
uKEmxcHO4lTaA1TwAGE62sr381R/o9SXhUYjCII/FBmmu4wWjkkRu1ZWicWDBJ8/
MrLE4SkHjvoxVH2hbTEjdsH4l3mjx9lBfaOrqyLi0TeyuG+uS6d7ACNe5NZvewHu
QXcPCKxJtVo+ASvClzccnS6iAeuzdMMa9PaHXpejMdQ7BBjCAGrOFkUkMtpJHKFf
ltcgBG0ZSHqLiK/hW9+FxIwZiMh9zCQzEVYt5Z0UH/ZNBjlVnDF/Xp2FXOr8FHos
8l6TiwuVAUPylbw3D3fsaWiAwejLeBBeExthm3HGzbtb37OvF/9jWgdgUiRrPcVQ
gVtFBCvLwFMnxlP4Ty6uGiRecFMLRuNDyLoJNg5TbSDeWzEJTBzDl9z/PZMixLxt
XHMsc+j7EQM2vtdMlIrT4cyIPFTEP6T9Rc+uKwj+H+ZnEFvwaHtNDVYgBZVaqJSR
pHt/ZdL7kE1UF60HHj0JZuzLO6+Ro5CXZHjsW0aExMGY3foXB/UkUK9qIIhGFxEz
oLz3DYXH0V4lAH1RLchyF+mgQ0+6zY34kQgsv+YJkXsw0lh1sB5oDbspweSfQQBw
UMzduhrmxudvUQPWpRIgX36fzmH7mtP+aT84hnSZzOdrQwalOajQAs3lsz+wOHYq
PjKmIHG83cBmvxRSCpX53yFRwlWmppKgsduZaEHySAS30TU7NLuWo8/PACHUPLq9
UklGthidt8A4nayuIkwKR4WKR37DaLEWV7Mq5Cxr1NAXk5HLkWzh8pLClbvTxv3m
/O0HWzpnDViiL/1fYiEnG3vN7sQLGALQhz3Gx80y2xxwf/6g5vX+3KCn9bX1Uh9+
OvM/4phXix1McXrSdNX3ZF0zUCE5hL9CzE9PwMxjl+2SYjYhrMP2wThe8zUyrWis
Adkjrto7eK52LprDegdB8MNT61jCvlSqHYkLfaC1iQYWYSMyOKmtY43ggdmG6kio
j2+5uzKMtKIJkMQsNFFLcIIUmg/mHgnMapXWQUMAJj3d27KB8fDkx30FBaf2jtV8
2GI/Av1GbwHRfw5RawaP94WrPOP8+Pbw2sOFlAPzPhSR5wiW+leaZc5Av6JVnDFl
sfG9F2iFhjKhljGTzWFx1AHWqmFrK/oXg3C3ShAkeNo5VImV6U9zvMsqRf2kltSu
mStsGCKwolUjyB8RRxV8fJUSLOc70pTCfEXfl7t3f+lffCLOiUNHC63imy0ri5kA
82ZFFnK1Plz4li5s0cvhGLXcveR8ziVxXVVd9sFMddCxJJopAW0YxRbLs0xngTsj
r5XSEvBjFPcs909hCqv2BPkrhrt7fCvLkVTbravGUc2pxz86aSqgaf8V5ytExGBb
weEL7Y8oVydvFqsb8V6117VT9C9MNGbjwAaSGTVjqqEggJ3/JOkXnQjS3kIi1d9f
E3kqEsejPHVMQYDDCRvXIja8hvX5ZY5nARdbYDlVbT1dCEC+7T1VeMOMRskMxXg1
6qqUGYNmZxt/+ZxSPFNGPqPkAzVQ2++a725jHC7SGNYk1IXNFHtauLrk9FNlv+0g
2CmYmPOahWlLTP6MztVpNP1Je5eGyzAPi4zDOrpr9KSVlL+P/+gr7q3uRfMQhPtf
xRVIsHN0M/rqTsRmLBZm3euGMgMEaN1ePYC4n/pPtcUaWMAmG9EHSWoSaoug1U+Y
pYjmmE1aoRUqTXvkvNwBmVl8jo+3ttnjOooFsbXjlMm6av48E5zEHnoVlKDcwuk+
0k96ylD3QOKHGY7U/NeWjHPsEt3HavZgd/d4frDuHsgMA3/QeS6cj2SfjTFteZ/1
tz5z/hUQ5dWIwUOWU64VxU8ljZwYs1TEFmekBavbboiWbf1j9iTFHyPv8Cq8nMX5
7JHHXUvB7YGz9MC56YpAHkmbFjizJD066YDr5TM1xiJyeAr6HwdO+VWo5NCoXFX6
VhSMcfVY6Rwm64bRtuBZUSG8z6is2qLfW/HYJKFiJoZ8nbGDLYkQ5AOdb3KjLlrQ
`protect END_PROTECTED
