`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3rhFMD8xzBfxNzmpHDRzlCKzMFa6cM5FMNhlISy1PcuKSO4JdWG6dmCgsOdXD34j
iT8ogF5q6FQZB+dx39mO/7mCQWHAiZTLBBVOwf5qWAkUtiC9MhF/03Nvem3ba6TF
MhC5ztnPxtRKA7oZRfLhctWH3ie/Um+WE5lNNUdfugQ1t+6p6eE222X6/xhOSHWI
J0pIx2rud/obhJoRySdQjV9QuYoAE1OwzHStXhW9icxvs5w+D6Ij7T4gpebfFG3Z
+fSesuDokqyc8I02S8+WtANdnPuVXTjYFJUVMMMN+AUapIp5fE8G1NeFfI9hFeap
JMuIKLYJeUDRqE4O0II7vaY/OE2hwJeLMB+xdZa94Q0UmV2VD1/D/gxWmK8l0/MM
fowYJRv9aaelrETr/UhOR9Yambwi850Mq42y+qsu2ae0bQzSbfNzxvj34RJyjEbM
k7G63hJmRU9XGxm2wc7NXLTcACHTf5Q84w4uHUo/Nbo77F6Czni2WoqZZnW9kItR
YgVzbPTWcaRNp/YFPbdDNZsBD2MMXMhbS5evjf34BI8bi8RYg1ZG72bIdnVSFQRU
SYAPmlMZUa6V9RXN9q8MhJzNbtBJF2qb8oUHXZx39UuE/StwN8ahS9iYHUp92Bnx
yVq5VziFtp3f0XjWxOnhUc7CihZ3HI7Npgb4vRMD0E8S9dY3KvILrEKf+nY6AdNy
vE9i3JBUHF82YZgV5HN6WxJHQVwBZmqlqXA922f/Ebzdw8Yk2Hj5OznX+bytiFZB
knd0SmKI/q7zDncHHzMSIX9LidvZOovfWI+kTMctWy2/MbKwFJX8CbihKfU4AlUR
OOM5w5jpMUy4fRIn5HEYXoZ85oDpne+1vjX34Y4lKh/N8cjLS1Deooz2woRbD1Lo
ijpsLprdR6toHaiQPDVWmcEMT6WD+NL7cLlrQbvwgtEbok4ZtnEJNvqiFM3lzrcA
IU5N0wNq4JlXLeDg6eS66ZvKQjMLEyc7YA+eeRJQ13Ay6+QB3XM9sTeeg51lik4o
x+AU4SZCyKuJUHjIOrLM5e8mAu6qVDuxStxgtTwGTMSHwjkqjoeLFQx4RmWfqYlq
4C/k1evuFoxKdrTvFSqJ6qchm3nusZM6Hl0YpfDop/Sa2VIVn0duDWXvYlf0+HkC
egbn+nRBoxCE4pD4ner6B1yxw8DhQREXzs0TKLE9n9TS+aHL1P08vcAXV1W8WR9p
7UVFgGB74NdfUuHl/3wJbtUq4G0VOGn4/S4bxfKNJUxFZ2753apvqTnBRi5jBYyI
XW+dU+SnYiMvvXgnEBbnYyK4BLHaT8I0fv08c35gGyTcQ2+MQZhNsMTA4GLnY6PQ
uCFi31DkoCyt4rQR3DnGgxmz0HzumVHl0bPcvDE55VNVt+BN9wsixNGD4a6AICKi
xCkGd7W/Jmb+BdumX4UPlXOsGLwQilt9yfWhJ0z393liuvmfEEYOS9o7oX+E06no
EIkrdpnba8sUgp+UoT0SdBOE9r1IJppWYlLhknPX2NGvjulKEH9FTcf/tjnWT2Hd
9rfcJGIgBueLkGaq5UVsDOuv1aa0PaeJF/6+lmdQCR5pr+8uzi1GNxfVghTWMSiG
pWdxkgey7SSYwajoPEpnDufFwMa/6r+XfxmKcQL3kmja0xAJB1c63aQgAfnxHAID
xVDfQUIrnWRwgxT4c8rG6yCHuYtkBuk/ewPThdDCFHVolviG/vknJFHBPJfAyWoA
2geyr5jKFdy+yf4GgZVRPjxmeqXp8RZoHuftDC8Lab15AzCUyJaeZ/pCYLjSk3rY
hfpJBVLJZHOWDwenfk5kNn+sLtKoNGpaS4PJU/stf49aSW6bJKQqbMnLPLHJFWXa
BJQozfa8IQwrN8XapiTYD1TTgDvkL3Y+RYxr3qg5X1RttTT59Mgnl0hSLEFZxAr2
l/JJUk9feoT+/uLIclybZ7URdmiRiVH+iRF0B1/OJePxXvCL8wdn2fbJXlTIU8nL
CTQ39UVYprsWxR5lQ2mj9kotSKgndIXQZCsOeboAP9DYqJdPdmcYbgHX3e/BSgx5
NnN6N71kEc1BwcT4fLOBDfcHHU+6H8QjWMOsog6OcXBWsiT3ZI5aaYClwQrMivbS
zTz2hVarah6xv9zDiNNh6lcHmTxeF6pCd9KHDgQyUTXXb0yFg9X1G1GqPq1yg4JD
K1DPnx715Vf8QRQbjw7lJ56OTE7VsirYEQ/h/XcWBmuQNa0LwE55vX9MujlO+xbw
Z3A1Ua/LVPv9zaOYFa6/Ol5yX6B7irvXbIDQNRXf0M9tjE+am0iDNyvDel01dy0m
bM0o0fBLeeE0S1Iy1+5Kwf3UhcIVndOsU8hE55uAGkWLhcfAe74jim1a9fA471Xd
Z141BlyJ6VezavXCisJXJnnKjnaE6usf5bGKKuUspwKuHd1Ue14ldz7ck240IM1Q
1hoZBJxIJiRlEWji24MzhBetOWgbDcQL7gJViLNMRB9fuH4JYzZ+Cj982XrpFATu
AhOtgnd2I6ZySTZwfwUbYDwwB17NcvvFY5bA0NWQfgVWEp6iSM5PONethT+kcRfS
Ho9FLa7vCi9pPJUGbnzd75rLlpF8ZOhX8OdAVCDcjqSY/1aBl3tVbjvi05oRMOYd
gpIJzOVO4VCKF1onWje1gvf/Vz4K7wd0ahEr4pHGbhp77ibV2FAAkocHPCOeJ7Wp
dG+5L0cEJb+EHKKz/QZxa1YZHBJs6xgNmDKvtuvb7zmeeYxaNiGODTpq9ya/ku0q
MAp6X0vWcu1IHfEkIQwZ/fwt2jm0dsnFoD6+1fbBdX+1cSzJXy7ZYM8QDi33hhAw
PdzbcM77Qi535w3k6R8p8S6qM/MG0f2jaBjupD9bxrVpIM4JBaw+VI1EHHy7zuYq
wcUQsPaManjXBQyddlmMCBwIZy5m/guZMIbfEUoVMzDRVeXEXozzoTzDxBHiwPNO
8SHItmbDFFcfW0buJ7bWISGVJe9ejgD0G94eIJVT2p6puYKsw6hl6cMpWsMbGY9l
axTqBBcjfmJUe1vlcFnAFMl0vjaKJnXmxbdbAJN+pG07+0j1Ik5jkDtznRqHPI3r
sQ/YaQW1HpQScbamfHEYnuZ8sHOM83WdYhhcthvWyQ2tJ1+8HDCw1WEmaYPgTb5n
ypRPN/xnwq6T5CMKpaVSaGhcS4YloxcYnDbF/kjtKX68uwCNRH5YqDmZBm4XLkDx
AJO5JSSVeSF9e63XhWEdPfRSQng5gXz2NmCUCaFCz+r6Ee97/uXpi46pawZRAgFx
bRdkYKQ4dRDgkRL+g28VVOoyYNWxAQ3N/y88Ac0Fv4xD817zE8+U0HZIHrzkPdmI
pJpRDFr9TtrJyf2tjv0GCGx5s5nawdvzs2MjMBMtPB3NpXizuBCCCVNDDSdvAjig
QyLUfD3prNUYYRdQJXJqRnYRV7GD1mUkdZ9Kh6/TzYplhLOoGCQ5IcUCEtH58Af+
5X25W0PrcCOYBsX1MEY+SDjpqJnKFMdRUG3aTj2QLUrcQ7vyAQKBz0qgl1no2O7q
ACR4sXvFdyAZN9VAoSW2vDd86u1AEIcBMCCc9jHu7CdjDPiqvM+mcCCSb55RCVRK
EiEzY32QfvlE0Qv4beoEiPiXeh4Mfwx1iAbBvLoST3rlqPrOnJRSCRU7WDnPMdtv
1ZfJZnip5+N6rKAJI7YYIT5SDEJkJB5DfouUDnQziJ9XVv7qBD8IJBije35O5Ag+
yn04Rbxr17yAeu68Ot3fMAUwomhjT2i0ED/hwC8qcmfNL1lQuSh3YKfj1g1IsmI2
bVdW+1tFmBPEB5HLb+LeIvoh36RQexqwro5UvngyMs3K37058AOv7pAWjcVD/zlo
s97SWfSCqhLRfseGbj/9Rxpy2l83nTDt3zpN+MKmvqNaR9LZlxZbYKMWpQ/CeuZd
/+xqNNvyA1fg5RmLtkdrdYkK3iziV/DKfUYE/pbExT1+wJ1eQfPk9JckD544UZPs
5UwKhcVfwoNE948oyvEcE+CgvFdQJDMBW3ycia27SG9qKa2z/lDLU68HQx7CYq/5
cVH6iuvcEbebGtz5R5JEgdtgbYL8WkIFYqD3OAa4s8IbhfxZW/Fqf/QwVT0neoQI
1fZMx5H3dpSMbqpVZhkqGDk3/aS1xAgKz3Js32H6VYG8MM+VtHjBdKb4shdymij3
oDX8LoMCwwgKusH6WE0GzmdC6AQVVh/1mHELU7FeKbPF2sMJvfQGhkBdcX0+fH25
aRPARmLyua76tf7YvgmEt81Z5CYMnIT3S6cHU+fssrnI5IVe8aKfkVaumQ9EfcBe
TIEtHWETNe61DsA4LIQrP1Glh+uGjnOhBLXyh8q8Qr+mb/Kwm0tlJ5WxcS6kd4NY
V3ItmkWpKOs2pEfTDBL+oF3b/RS06yXZMyn4uGqkMuysnQQzuG4Dwtl2Rxlc3Jmu
QdTBxBeX8thi39933xNlxZ7zxP5h8NmeMdtcj2GYQFX/FNOgJ6THXwQuyPpV06Nz
Eve9JJfWB40ZK7xcxvNNTH33QQQ2RdNIaCWDi/VjMJ77cvrmdq0Zlwe2klT0XUeI
WcgZPrKi2vMGWRfsR4hHtyEo+Uk7nAZRLm7kRtiHpue9XNanCwVwripKxNmgDQyg
v23tP6uMyhbzST79yf2OY7dPB4Au3h1FehJefRc5QdHAmAET9gKNA4Ph7MIyvoXi
0eOhycvBJubS4sOcIrwjffUQ7Bc3LSg457/dXd+0u0aS6Llw1XX9TXxNkUw6xYlJ
LiPoTf3jVY9RiqEELu6Z/Y7cXMKI8HrC96ceDWbqgDKnSFXBw+9gzyCQa9BqeM58
AMMOBSDA4t80Y2GLQ+EYYyVNUEtbapOCO7FvMdLs8ST3DQ2VjxKuFl3BPhB1Zj/S
mOxo389KqXVVVsuVRIQ+8gEU/MFjbui/QJpWWUgJ/fiWsxHdTX2P7Vj/n3II1Z8P
TXXhabEde3NpDt0ynWH+TCJJu+cXXRsmYmz3qL/nt4Nz/mITkLikj/pBhHt1K81L
enbmqSf5DF2A/rpiJ730dS7M6gCbrDbjDQFXLxfh+HW58vQ+tvyCy0vqkOKnXas4
UmWc0nZwEnNERjY1qZLWqn1w9vvjXyspDGKsqGkTKpiQOqTuSgWHfnZ377GyMePk
sO2IYsSJO55/XflyBTpddkC2SXQ1ZKVmq7QHO/FmQ/xxKGqXa7DB9bmHZD8DBEoI
aAgQ68N4xTAe8/Ent+mqOpn10RD6ljDxiGeM9eaTXOtUU5Bz+Lsky9FPeFNfXQDc
I6EO/gmGWDgy9/j5hXn9e5DcZJfiDrmq+DdjTBSB/wg3YThjr4phi68OeKM5MDSS
9jR/o91XlCFUOZBM3U4Q2RzOrzjMVbkdwBWhg3s1c1FeBWQgvpL3VXSHL+oT5Knt
xvNo2rTswb0DPa+4jayYll3RY47H6T182t02hsTyGVNVH40wLSDJ2MrtHlmAP7Gk
7I4dOdgT5b7d3D9BtidCv1JoIQhysU1W+Z8ZvJ3rlwygAmipUKhuYrlMgbcFR18x
FvwGLSvxz24cmLfKfHCA9tbvrwGCFnhxg1Ei+7VyvP9mZNxEDyybRHNkB9kaBkDK
etEzF+0PxqlJE3N0evLzPhtIxawZlZYs/CmMpQ9ibB09m+zw6iAFCTH07Lu4M+Lt
IinhATbVOFTmWNp+AcIAFH0fyzFpu+teAY/xqAW65NserVzs6FQOdstVM3A5SqH0
0SJnZx4no6w3aWO5C3K+lWnat1E4xcCXPGPEup0tEZo8GuKVyeh23z7p1BBq6CKZ
ApefUhyhI0Cgv37r3sC/b7nOXiO5U/jQlKEw7wqoX+JqthF1GJfs4I9qCzLMGlvU
S/JHaBwy5cG7bXRw8PhFk5y6V//H+Ofx/jKc+1RBoO4kJb2ZCbDDxZK/U7hmKzJW
7CDuy+hKNse9Juyddkc/wV2jqgdAOlVikK8G9uL6F6DPjBHxziNiO3rh4FQ9y9XJ
4bx8Rianyz6R13aT2mbPMUM/fTVmRfFzLsc58Raieb0vKDNvzx2x66ikAcvMYQSp
NExQd8BQu0SPHULtS9iUuw150UT6spRj6aQt3deGKkEHFrOl9seS3MODT33dryYY
d57lwGnfD4qTq3cM53Cbu03aXyURjBNqL1Q8bS6jWaZdwudcRQUR8LMEE0jZf2gX
oCANLlEA3u7oVK5fPVv5Md+Xn/jTtOdSqrNQixfurqSCJiYDybx1XPbaWje37ADV
0D+vCLNeX3RZ/vRQVILKcYwLWUfuZXV3dCunX/SA/ICHrkyUDaYWHLeVwbgSLUJJ
glk4NTVACmCIqCQeFzCkh5mVp2LtwHOh+rYKxg+w/hQZfb4eXkaGqnpOAFW7w15p
PduxfPcuqvU5RpwkSYuCTN5khDn9upVNn+9KUZfKlvKNreejsnZnagQla2ph6cBG
vcQxteA+viBNtysr8QkQetaULRjDZupc+43i6Jeg2yMnxc+vAbLuMbwbmhvqjBth
wESYMA8vlf3kPu3INfqz+rW8VQ2r0nlpWjLX2PWiQLWPiHPBDO+ohPXoFhTLRVwY
X/pudKmXne8nIanyNPsuxlyzVmyCoT7lQMt7lkKFQVPgTA/SmkBG1k0M8wFZl1jZ
ZDyPzLpbxbt1xK9spE9Dher62zPtUNCSuAt8OSx7ZefH3JFa2hM1OeyS1WgJShPb
7IS7hHc3eIctryKoX1Lec3sxjbzt7NTcsB2RSi97TVUrAd6Vd+fK7S4KRvHCMwMn
07Tcial5imbJ5BofyKoQsCCErSCn4pt/FSMERZGgoF/+5jiSPKl6AKz4ff5OOQe5
ite3wqioq6cMEMyZgcPbJisyI2+pbwXBXMHhIk8EqDbztfqQQRbBnQwFFXUJ6HVR
X8ZQNBv13pZNCyflAQOh7aK7SJLaKFIGe9j5YakvXpsWuiuehGYZtleXSP+mACrR
idbXeKwdzHeuo+82SONKOzWegD4BlBqgXMlMEX0DgmgE72dAjQUS4W1AyeQdDiCs
5eqms2oFvTXnHHZfwLpF7ADJYBnmVVcbmIP3mOeVhCflLlbBVLjSnuSfKx8FPoXz
td7u5e8Rpyynxti41WS2gmv3FeamJr+OYk56qS4oUW/M+Gxay2ySvVVx4JD5kgqz
UEHaw7eWOBne/AjzaJGSD5cxiP8KftIFpCOxd7Z+/UbeJ0uGSqOjcwFa1UfQCInQ
yhT1zi9wF4GbIB34ZIMLz7qooX+skLhE6zwERFd/2WZLJPEM1uEhTND1abVEhciG
nzDRw0x4w/INb6rhFZgf3aLpeRKiuS1TxhvwAc6vUrksnDpPA31i9hmGcx7TIk6C
Kvt0lFGCv74Hb4mAUdZEZcl1moBuVINVs8nv31ZuMd5ypCuFO8ZO3h3mm18XHv9y
mTPhFHdDC8/TwD3gZwMPQqEOag5PF4jtix8hvaWoDMOU113PtJECpJ42vx1FWbaF
Zde77yz18YXhqxBeF66LJnGBkBdbiJo9SOvBpLbzqC4j9hzPuEiW1vnhFCnGCDME
G4JKSOLQ2RXKgctDn52choH3IJmJRclF2hMmpWI11DuNjk/XUgRyCOstziUtGiq9
`protect END_PROTECTED
