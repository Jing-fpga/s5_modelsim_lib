`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
91PdRgNry5H9469gFR/bU3ww9VAJLqTleBjjP/vltFHkFwci0p51WcIhY9z0BdX7
MPopQzmsPT7THFjYewrqBq1ABsY8UIWRCtS6zPBTBOtPNuR+6GJP0ygoJfhsvXj9
Zrz65isT0Au2bz4KPJ6NIEgBF50TZ1qsKKRQw9IA0DBTG55W112JBH+C4v3srLxp
Mel5lyWVbLN/cz54VJ5KE0A1C8KIzogwG7CFZLLK1ggcrOGvmAlbFIgkFJWhUzt7
r7WBD+chk5/fa3/405zf1kGyYznp/ndtY5io/7YaYGeq68q3kwxXCLiMeND29rVq
1Yq5t60vonq500UoRn0sCobn5MNpsYEqRqvDRO1vmJLOZLJ2CHqdUO1ErvWXyd8l
XRaGuA3UopbfMKdBzFUvzFkDwIkAG9WJb8BVFNP7af+7Gb8ZAgIYck12dx7DEArk
rIgBBOzOKsGG9koZyM8fmiD7ROOcICfM1C/wlrt41jRgT49e6NlLKYqdhYmB3qlU
0jwmBv9DNCZ3p2NQDCNk36oQ01RWqvRnzsYQ8Q8MGLKqL20RnrvBal4Jij7pVwRA
i99+al8W/IHJnsKbXOQMkpVVZs35HfzLoPv8Vt1g3x9xe7UuTR9rmrFNrHniknl5
AnVj+A0YBLNzcHpTAqG6dOOjd1k507yXqfcO1lej7BT8V+TMqIXu49NlYZ1j2m8e
gry+tB228djIAePUyKy/7IAh46xX60ak/K2jYs0fScUUHSOTXAYs1U24i/uVnlUh
IRMaB35F7Lrt+4MP773UlvHa/1aiXCK1q/C8QzopTY2Xa/wiRGJlb00G/aa3xWdB
g6KIJNFaILj8bWOLXDJv22XbLM+HX9TDfrPmqZXpIsodY9mRZ83NycbuqYrrUUbC
1Ve4YwSb8UZByQJAGL4t4U0rHECItKutAQi2YeDalBsLz/dEhWQH3in5fyOis3YT
8KInXcUCbpGV4P6FVpX8hMM244Qkn7Nnq2PdxsK21zZiPTXxGN34LQ+0FVNGWth9
F4laDYp+faLUQ4MXtkypDWK3AUBJwT6pvsmSFrWJH0NIay+QjAkQv/vDmMUav/48
bVn9YayIZaPaAVrn5CTF7YgSIm3A3SGSPMRU49EgXtkNaW/vZLBv6Eh37cAmV3pF
Un4vOOC76rUFHxuo7v2+QgTqPupXLS+Cbrmj/OI+T6R5V3QPNE5a6ODHOjJ7hmuL
LdP0NRhQnfcIjE34m6PrxNcayzozvZZZJ+DHIOzeFk5LcpsJGSWwJGObdOuxnjT2
SAVeucpb3ZEUS9ghUNulJgYtfoUpuJzgeIq4pJKSFIhtyEM7zpbpDcX5iG+I3Zcm
SsCNuE3WKWhud5N3LKq2EbJpNXvIIvWxUeask68H/b5rj6nJyvEC1tqMQVW13Gt1
atM9JEfRx/JScbTzuEU6kYm2lMVFZpRymGdK2tqalcl3VCXgu861GHRlXl7xwQA9
sgMemxevsM7Ibwp/7rAU0DbKibzP93JVoghiZCIL+i7CiOcSpElzVMVHRasmvAMr
KPMwXpvVaEcmiHM+8kddEmepycyC1EyQhfP0Zjiq3dB7Vl+ggnh3sVXdtFDADcKr
dbaX5R8aAH/PqqsHk6/f8cIY3Y1EPlauh736b7AVSwYPo53VcvjPghQfEAjQNEFa
jhVgysjq5cKBbLvxoZfTRxRGkR2lxbK7joawxkZAoz7kDiCBcNIxNf6AWZUipaCy
oTzDWUA8kdccPMB8CaE/J/Fkpj6Z1SClZfuRzy/pNCHjfBIdDTFc2I4E97f8n0SM
aqSNf0fueQTbTUL3f3KTFOrx9TRCcRyKkF8GC5p1ks7GGteWZSbfHu7dpIgNuB22
qBejtlmWJlFO+egUjeldlc0jJ6T8Q0Dj21KhZCj2FQ9nGlRdMSkXE3MnpRi+ynut
RduKX9jftmrheaTPsDTb4ed6qbPMGmcjRiWJGtGs1fJev6uHz+j0rUK5+mzBNjtt
6sz2S8llGPJ8XX09acx8VFUq5aA8haGY4sh75bQlqA47HO6c26KKBQYWlmkmvfkn
+7oIJYUh8shE7D5avCWLGRyQiqNAjI4gZUofAtWt+fMErW0PbGFrfb7RPqV2O5Wv
4vUP7EVvnungWknp2Kl7+M3uAMCIRceChzAv2s0HWAAmU+poNs8dO5LRRdL1aCPm
BtdqlB0Pr3t4MKAkFm2boquLR4bYMQocA3pR6LxVeVgh1oo0TJvkcJDouZfa97Ak
4eV+/vYXftupf796KRDUHTu2SzaNckVe0ddr688u+ZfnmgN5dz70x08iZbrfr1AP
pnQRhCiL+XuG23oYxhpuiE7Lc4nCViR0hTFDMrOyKyKW0y90RicUULq0EdApKBFb
I3GsIsJhrX3EpBHbyF55/vdH8yGypeKcUrt4BV82MeP8bu2cyfw8w8fIsUcMMGDK
BK0KEuMgZM/O4PCsR+yVZD0olVVj0sfWonPKplYdppg3dpJ+RcnHwEFLVLSa0eB/
dMIeEbEr16Fcn2WwFGTt0X5arkihlXzpbHqAfldvBryVDuPQpfi5aebtMaMwemWA
EIwlKyD2hKrwA8soVzonnjE7T6KYx+s8Jfx6fncSlMQEuZuV8KKX5Tpc6wLxudzw
zb46TyryPMYHJW540D2ma/qGJLEF9HreD6CHffJ/g27YVm8aQOGqtmsbwoCmthOW
GgIe8I/1pj+ZQu/jjw935aSikzMujO3ariCT3FNSRJYlFqZAGPhCJO9fvo/RhSa2
2Jh7p0bysEnIh9G2iV9VSCuaSRw+1cQxRD1AmrXIIFCnYUCs/2CSbnadjc58HYz7
0zuFKOWGhX/b6AGLjDgDiiqGxp3i8QuUQ+8pTk5Djb79tOWtlk1+j307aBpRW8km
UD4YZjI2vR+8mY5SMRg7HJqQGcmhuhlIvnpUNm+GQ4wuqoea1euNLIVZHBrO2llh
qPRjuN28aBpsOfaorilmQ3h1Gh3O8SfefmhOV5PAR5V64NNHIfoI0/aTb4TYy1Se
F35ARbUXdhghbjfwB8qFAn2xWxQWHYY+GbTemfZHiPH5zI/hfzdKEe8EH3MJ6Cec
GwDH4pubw/KkYaLHeUoPkQG8UEXQcAIpqVsSpx7NSn7HQrLF+yg0qWQhCFM8mjx7
Gu3TNU0o+HexXc6mbKXvh5S5sDfWbzNXOPi3Al+b4GQRPlIiQ6yUecnqTJHY7Thl
Y1S5BJBWN/Kl8a464xxiXHbQSyiKzLJsHZX52pFL93pNuN8p+seKz4juhRQdTHO0
saa8NZLLIQg8+NJGkg1tyatTiXG1qUf+zUL0P6fY8LQ8k2FwfJMIvnkMfH20ZpGs
64gFROWMwYI+6mYWrYJiWQo/GkDlMvf5wP1dHQyLQwK22NbMgcxeDMKjPWhTZpbw
GYSZRqp6nTQ54mykjVzOtPrvOJo+BjVGT5WuUmMI6+nfzhWahlxRRIirx9r4ogPl
gcWIDTcf5FI01G9ElvablHdXsh3LZjhaRL6BQwowgWRl6beD5WBNlzX7Zscq/37C
peZytS5MVGHS9l4GbOSuGTtVg8jF+JGZSYpUHBSzQRsikV87wXCxRURpE8uzrukY
xtyktfJKxjjLuCb9iDuATn71APItkWeXJJrwKAE1Vozwide5m8gomvetU+n3H+z5
5qe0BJpQupJqoy4AgUX8B0ACwPU4Mta8n42d1W3G539pPt6zm5bEYGsHsWlmndLK
cs7b6tskBCkv6h89hmzD3Wt3Lg9kBlxX/6wB3iWgg03QTHQS7jxGH7m4LTMTF6k9
HGIiYpzYggtpBVga7lVAxuvwidG/sqxonNK9aQChpKohadlUmI8DZFLUDm4YUlOY
u2+zIm3KGv0mJqeXpNpx/HgZVy9VZOtyoo35YsEPDYIaWosxh9gxpjk1y0lmTKwC
Az2b42PtyzUux4p34wEVQ9DPfFY1fTzHtlggdfSb5ga6PnavTsswnS83YcuO8Mtg
sMgTn4wfOz01vftUR/ssQiyMLACw7W4hBTVRBOYn+YRS7GNq1+a286jKWKGzPLiF
e46yVf03tKSdPiY5AXCJXQGCZcH8gZ9A8YL7LeQPw5KVp2AYFhJHZVTvXKEdiziF
avsq6w/lWStFjehWNU+ZiNgxxQdbNMEs4wlFmsuvNE8xDx8NVrQ4gUPhe+b7rVVY
eV1OSeoms1pP0gPYU2dkfrso6XfTRZh3fgpgGiZXw8DZtvHft3SZ42nMFdT1+h5f
RzcRk/E7TCeZ74XDijkBSixRoc649aGv0728wncqPwKukS3Jn6GLbcgKJsjaZ639
E1d6CGDKAKeAXnUGw3CmlKdJU0fcSUR8Vb0FYA9EzalB11d7/dvveK9JeC4p4E9T
Uwj7F45fo8nS6ft/XsHoAzGbq+Z8F/ik43gCcnxFTG5LA9E23Ryr+MA+0C6gSqip
lVLJVqX4VR+PmDr9ZIijDQpwjqKBBLiG0lICt+KwsfjqEVvy8tny2kJM3Z3GTUyf
FmWVXprpLdWpZshYYjoLUpWCuagbPMhTlb2CK1d5UfcI6BFyK2sL6yTU7eODnuJ4
oWWbWU26z4ZJYCGq08DK43C24TOcUdi1+Krp0NJmaAIzgyltpttfRJQQcgmHSgvn
h1f9GuoVcnVRYEDvd4MbiTkVxNIgMPI2kXIFFwvKhaBDPbK+4PNvRCWxBJsdYpSx
69P8+xBN2ZkOUNdms4bbMnnSvUOYaCSKLO4t/edwg/4gXt4IE9Ol5bGIkxMRJUj4
Q419Bk+q5WrQM1c8JebK1l8H3tREQFTx0fDmhjBOhRaRjM3IOGIrhOeQUeQVPE4R
IdtamyXmrzSXkQrg/ro9sKGr9xUVV3rw/omcmm0vcSMGboWr9JbznawY3tiSnqkQ
cbkecTHme8VwWUOxJ3FuDLmtOMoXiLMBB1azeyq1P73e8ut8AQtsgByvimwHWbTX
bAzTgyomv36AHj0r0hyVELM+5cazFKFt/ttVUf7v7SCZz9lugcHwROSsl3eOG7Cr
0bgYgj/pWiRSQ5el7lmdQtVxjKILCm4w9NJMPjPE+FRykotnlVbmZFo1u3FLCNyh
14ZXyIxk+xvFO+KDdjCTZUkoDVUswJzL9OH985ddzLgnIrfnbuYz24VlK/xNrKA1
gpQLHNmVX6hnQZTSjABcpwz6ZvTO1QLnNOJRIUXvE+/qLsm/2XYzQuJK5e6C1CiL
kDjwUqbBC9OrEez/1TxmbR4CZvAC2n0Iy9DWM0lxhZBb6Xj0l1nhkQ0QTjmA4z4G
+etY8qcffnkIO4rwlL3AkVVbeydNTbblRb3ivUTV0WUS6OhjiQd22GFx+1uzJO9y
UGLLnnn2p9mqDBpJO8mNG/+JUtm4Kd7VoFuigM2yjJ0XWhf9hNzRjLEwDYRgu63M
11DBHEOKSHGsu0F9/MEOAIqn6AileBolPjPTxKZUvf94suKgayAp2y2ynaJAkyQE
huHmPUuXX2M2vvhUYSSm3BjGncXh+9YaV5iqLcCHCfYFzTG3aTZdmZyx5FD5gy+/
ahxJirKiyEP2Ud0czJFf+YUIuii8dCTP84w7dU/ZSAmLO8xUohlFK4XjTxtLjTS2
hg5HGSpqhDuz2sn9f2/5ZJaufDgBIaJ2CSASv15/OaSlouDHAKLDNFJuilDchhAQ
IqKv9MKrRGIoz1hWEBGMts1Yr8Mh+JZYEbQKcybDl2uooTxqxJ4k3qAjvSvPu64s
MLYDEuJD6mXYjVCNKirY8NXxlug1wUbrmtfcPNEDeSU3XP7sAiLbhfvqOcC/gAJL
v9fMrpHNUsyLKqw3h9aE19HqipW3v/FQ9CE48BWXtOQW7/ePkVO5kUXwxgyD1OMd
3+DL9kuJS8SfCRpqKsHXrSuec91SnBpAh/NWgC7yX9wWwAx84U/cZBUC7Xgm3l0l
fF7lzt/SCY795UXlo+gtRJNIx6IP3iywM0foFifsv44SAI9LTiYux8PGKW3r/fcD
8cCJzxfOjGf1aQW5hgaeBZ5HI8EkM2dRK9JwXpsAvWji3h+dZs+/Be6xulLWY+y2
kL+iYzS5qqK47dfPW1K+3FudWCHTtcQfUH2CJVCmWeEQTDWtmpBQrIN0oyXp6rLw
wiw0dQL5vrR5cGO0oVQE3hW867i1fx14LrLo2O044xfZlcmL5mDmCCgVXyXcr383
Y2Zm8X8Xcx8C4ROAiM4Gk2nRZ18/xiQG8U8egdBCbyk8thUNeG3CQ3yd/FvUTQl/
M25gtShG2igG/31HIUuLW2l09UEqYku6mu0Dc7EOsBhn3fucmOm3QweqRiOuYVQH
QbVpZCpwKwJ+GlwT0BoqlwZ7avIYvUD5/D8k9gvrr/M5Idc2ADPPqqmSPCWmHsJj
fn1qbdiYT02fcVeMIle+tGi40zHDYQelLGuxOqRR3cpis0njGlzN375oSPWgCsAK
eKFJfwEincYSQEXksxFHN3/VoxX14g20+ujZd/BWZ8cV/EVzS5SJCXzrVc/3fMvE
Swuy1jPAUDtqdSP+TWPutiUBbPYlHb3kk/21Uj+SDvy9+SrvuoK1NaFV3h1w1i5U
lowSLAwqjeoTHXimjWGO16I74X5wX714g6Muz9JqLmQxEq+E53pxgrE7SQ39HGBJ
qdCLPVGDTIiKTMU6TQmjwhqmQvgp5HH2EshuVaLyIgSCZbhNjEP87b5j9yZeAyTs
nbLBAdksonyzjWgF9TamZpLxGhhDbAI+YwN2wMW2Vu7ieigE0c60ixlHVbJKMaH2
PbiStkNJYkTzeIHBW/qNaFW8iu53hk2wLrN/HIwH8JeAh4DWd4kSzayCciL5uVex
Scyb/JWjCmmDUAQDMplDLq7Yy8fo3TNcHdYKh+eiXLinqs/BlWu7JdwFTzucUS8o
YJhBixlfuhuR53rpLoR6TR1Fyhcrjhez1yXSzs79OLxSvLAvWSKDzTEGtuzwotRE
sgawD67jRch+TIcBRNWhHrysuXcKTs+fcaD1iZ3BZq6zPIDPz+AkaGzFwAIfaRr5
s7ZrA//vwlZoad0P1cF5yejCfRj4128+nW+0Kl7O2sau6ZybNbm4yX94sazTO6go
RdN+3C7o0Tq8kJcD4h6vSZRlmWXwu+94JDnP6k9nM2Na5Td6l5s6yKbVxS50sMsg
Q7FFSiEMq6HQccmtK288uTaxCBMeIMx9dl/kTFr62k0PPeul391nqGPxr+pUNRwp
CC+ase0yYKSS+ArK5j64hdDa3FpXiIgBq4thPl92iFxiuyB1OHFzjOh++vgPubSC
83/4jm97iDBFBlyNaCstAHTukZmWkqmymQEVxhFt+PZwUM+hEL+ifQ/9R/K2Np/8
5nSroy5EwzgRIosytezAatKAsDgrx/hajqTOJH28bWsLl77XhU4PL1UpQ3Aywe7M
hpORfvDKzPbMVb4tArFjPK7VF6jBulh7rZIejj0LEGmbOV9giub436eQIjF65z5N
Mc/HqG54r0wxwXrjXAEdebw8saUswDTUhSwCuy8I+tXY3LCiz4LLlDsiLfgcFVFV
E12cSthPk2b4EgfJP66/8OK5dp2kREyjS4RDE5DjwEg4KCz193eR88OnL4xSzR02
z3JI6GMjuCn+tB8KlCX2/kv9Y/EiUh8aE8qn/OXLobv2h1jjN5PgUIbKjdgtodnq
gLbF/FQNwwctvI6qkdWEEAuidiAc53M3rQK/JJmzdGE7+CPqMZr9DQKwFhS9kM5O
+RTNipH3Ons9zs2g/sPAxxypBss/gjrZVs7s57Cc6ftOUGtZvpK6wOyk5EsvPBXm
zFPUsRC1EDsiY1qa/V4ehlg62Q7Le1CZ8iPm+DVkNKCndiZ6+PrSlF38gzuXWMo+
DUq7g+diedzP38q+nmjnveKK28a1OGmCB1pXdX7lWPITliZnx1Gn0INwiRYVRjmU
klj/Tfc913+NTs5InrGXN6fsO9wm0aSarX2q7NBwePuUeBbQ1TRe+Ehs4rhpk5Da
CNGxIrbl5ZfrAVP+SjA8G9jALpE6jRlqOjg8c/xRrVtos+SCfsHH641y3xQLKfQE
BmPcpe6v49WaN+v/gozelKTSYEspCOXa/UsXCVr4SU5sq4ITKi0sQUusQUY96rLG
8HHY0KkoHSZNedCGhEZwbTs3mVsuvfqmGx3YhVDObfu9gF/PQVLD3khAv+yNsts+
wDusupg63++7VNZewFSMRBYjKYWwQK6njVsx8q/jVfXU2wPdcnTXU4AqhBekGPW7
VdSjaUJM7200civnzUuWVH0ZN27k1uRySkSti6Ju74/TcXmcByacW/Ztwds8J9kr
2mshK37ZV8CAvE7+skNhPj/nHt4kt6mGYyxAmQzuEqzu0Kvdim2A2Ae7q5dmCeVi
KLt+AbINunsSDZkNC3X/TpnYyxK5N1azGgEsYdrfS20xvMn1YFH03OeJBt0N8TMV
RxbBO86UzoxDewds7Jb22s+9bybmvXhp053BRJAL3WWoeRQZLR3qHWSiXxwvJcOu
NbvCVb5Psmc5T53KHEs7TxPVg3XTdoImKjvhXWvFO75gRcLnRAdP0jxGt9drM4T0
dLWCHcQWoo3Q5MPZp2+ir/C5oveteYMvMfEFQiwztvzFdQkiDbOCaqSoYVUuKtSK
k8JGyETpGdaG1cXeGaQJZrI4btJGWeVZepjy18lhdijaseJRB3JTswki6mr/rAwZ
TzrFFU+H/GSJtQE7a6GyTqc0pqHg7uk17nVKUoq8tbtgXTRLEUdy1vOafGAJY/Wg
ovVGoPX3fyOWSdTQDkXQatLeBpUxcyXNPyphNreNCpopzz2k8s1Z2V7E3dxSs4yz
PEsRKogMXeipWB70GUAeNm5mnfeLZAQCEfINoJA4pcU8Oo85EJgMjPCRNtBi75xN
OhtmePT2NuzTFeMH2eY0XRh93RGYldoomdMqGBchX5y1NS7YK9op3pFAyQ2LCeW1
h6OiqZNd/sO7p+SDwQgjFfL9aG6V6eKFdhQ3rhKHu68exzov/L4L+yzJlZQYbw8o
4w1icSZ6LVAaGFt5G+i8061ryosoy4D//pxIonXne8zoKG2AtGyEei+aKV5ovGZR
uWCPwd5RGNsEs9CsfuE11x+/qyZzq43qeaAeDsknYLzEVZ0pUrlrUa7ebCGpR68S
LrnYmShIea7AtcXm/mRZYv+j79Wbt6HoLsH/zw+G/2tx+lCipMQ8HVUoJfTPbV3I
oqDlYy9N3ppw47GkHUgo6OEWI/jQ13VJJXGYGhIg/y9ChZR5wymfVCB0zWOhbqkM
FKha0EV/tCfAGVgPun8eZXy4hILuiDEZl06oSbqyj8Z8K2speJpwnPAXgym2yby6
bzaq679e1pMGWio8ZnpWVrgiONhGVT2JJGzNmDKUQ1+A2KLH+6WJI4rFm8jdac+3
dn/iSLNOh5SIWjMhwGBgWUN5cks18+NEzI1ilpfzh7NARoeshTyQrl80Tiyl/F4C
X74TSZnTfxLOV1qDbZp6SLTVGceVHUytcmHlCBE+s8ic5Lw3/fj8ka1M/NM67+1P
cGPqoQIjQ+/Ei9j9xko02KHjZwHrkiivFCeFqrq/7HUDVKRbevDihiI0HdBRodLi
MuvJMNptSK7EaoC9A+ckOSJUy89SyVgzl1ZH6tYWRbr8katija4BIDFTx487na5b
LeXC/rLMTPMXlpYib/6axVjlSMWmPwwjAb88yUG9dk/PDxOYvQNl/F+2EyFjokOZ
oI8VkaFKr+hbSz/UPEfTAiSG7eDIHIMyzFUSHrNIu1raaO/BQ4qVOwcvIh3lEF5o
GNWrv1ng/QI50eysVacZePaOyMOJey8TN1z9fP3jKx448po49kHOPftNPYyNbtfU
aXYtftURYzeL4XZZwypFbNYkwq22Y45Sl9Z0ggF+Pyr7dfLEbRcWKurR6hm4q1oB
gigr5z6qrzsgFb1acCIFS1M7IiXhFlhT3OfbgnUpR/XYjg1K7VnR1csF5mOYHzm7
mLcn3pumSjd/zTW/1w3b/c1QAOwNPXJ8EMB/PLV9ZV0Aegy7Szyho5x7Y44Psnkc
UprmuN4JlaSxDLMW2lzxm3PDkxltKS2ZcU2gRfTuYklxzB9zLc/+LiUqhB4Shxti
QEojPtW/5aZCz26FuObCvNuGxVcTgolIhqPFbKXA/3GBxDOgDP8ooPaLhZpqAz/6
kQMz2kiE5Un1sycVLLN2jkjO/MsOKf52Mp1VlPishbHsYrCXpPamW7GquSoPdkl3
Q0IyD0uBOPhrWIX/XAz50qahVtBg8XvrRm5qCTMNfpN7dpRLP6MeJoBWGEYgVbDh
tOLFK+2gyd1s1HLRUGvkH42xHx6sdrkdx0rFZLTDbZyKVZ0M4D1XnGOT54ANaY/v
uQRQUxFGeCKwHIeexQ3cxRlEG/fzb0aaBhJq9EiwdhN3fDUqJU83SS5vE8YQ6AGU
Ak9a/4BwUjgRF5DHrQyyoReBHcODrE2ypzaXw5w2bEhrRmZptlbREPT1hD/dfb9e
3ZJUOkHOOonrxkg8b3i/FPJWN9BzR0SduVJROK8a2+RJR61STBBo9I4/gFGXonuu
zjRPN0jPq4q3dqX9Bg/VAuQxA74Is49cvwTZeX3W3S3Errlbv7plSLsanY798SVk
fKlaAxVO1H1xHMrmPW4U7rpIKOYSWl2zQSVgq8qMloav01i5otMBeAxwFsRFZDji
JK07LMaqwUd9Tt5Qt2k2LRRGSvYd+PdBEP03DkJkyZcilBxt6vAA9o4xtqCjZfM9
4XlI6PSePygtOeYyZUhkpI4IcX3MKJUi9Ewfw+4QcfQW46upENrn2d41R2zkahj/
dW4hDi4xRQp+5nxW1vpMM7a0BINBIwrBOGw4WVfTqDp1MMPV/oB1Mzc+9dTQEUPT
FEtmc0vf/kRZOV9pnYcwBJKieI53FiVONKy2ZQZTa5jV1GOGnW4H1MrPNJ5f8Pw9
TRnU31L0jHYq2Da5s0SPs4lAUl4M0cKfeVqiedZJLeWOQpXVW9iX++eVNIgKNzm8
Oj96OGJkSkq0y7HjimuOSA18dFMNoA/L63ZQVGw8CtTCEdRE+7z5Wog0c9mJgCFq
R/V2RDp29zMArmJ/l15dVET3g7pJZR10jQaAat1jyLkvrHYNop31I867U/RtT1pR
VUMSRYjT1Ti3LNO5/nK9uFovCE7/oRObbLrmn/tDyTsF+u8MZDp9q7UwgVYt5pvB
8AxcMpmUlpbLjh7Wm61ZBPZ4AeHMLwSDtyDaD4M1yn2CP5fjl2Em739YH5KZ8f1O
4WzHpXVJxCcsHXVwE8IJPnt7+jPGK8lYQ8WAhpUzp9lmrq9P29IpDsp1VH/gszgT
jLZPpIEoTq2sBHfIhbibvb3HRf8fJP/Fa72CdzNTnv2aB9ptplLDy7ax97CSwKYV
FFO+Fzc8kCGMTXqH1U9gHNlysiUEyeMuTuGQfqRJVW69EHwCeFqkqIKrc4iz0Chc
RMTJWJXySF65h4Pc+ORghMMStNaV1IMjSOJLbXEr5U2l1AxIs0rwhZa+IueyxzTm
RwGV3wG3icO9D4JD6QOOALDLW/IoWV+hanUMSVPmkKmruGlxdtJwVCdy02RGQOJU
fPFEQEmti2bpLb21WoMboMO8nCN6egB4/RgNZZUnBddY+fKv7QvCz0hpFICd87Ji
KnMEDA86Pg6bCkDB+E18/FwD1FTfYJdAXINgRdaDWhdNr5pFoKcbbX/T8a6Ww1zk
rAH+ouu8+o2iCTUW9MwcBxNXEoXAInz2NKypLvArendb014Ms2Xfo+TH7sYgVSje
pHxC0UK6r/13Xok+BgynxUGagNn56Kz7SNqtHHpQK7R6K5zTjeNIkQep2yazebU6
fygIUwGXJlbZePBmUP0wlB83zq5pCAxsG2xFd0nwASxUNro/Xc5/AC/StFWGV72a
JSeDIIKKFC5qQ4/kK/NvifDApb4hi438zWNT9me8Xrdi+vKDRtfFCfrZYHD/MDq3
VS/FQ+kWVU+ZgDfnKfycmRK/TIEtsLHVT2wBKWD8YGl/2QOluKkSV1WIkGT0ldf2
VjvLipYpf3TeN2uNmQVb6/othU4klucP8E4P2O0JauA0EUSmMs9qBBmvDtKGh2o9
663dQEcEgeoHKFDSkYGh47P/WSUXReX9ZAzw7vPbRhyAwheSVte1HkA52iouqfUA
qDr2RkksQB5/yS2mCkVYbS80c/Ldb/TAa/4Au2EcP4bpn4ezuzYPkE2WkQ5yuVjA
QVEnAIt1Dt4B8QxkgnqvI6Vt/d/ncGicZu41Fs/zLX7sLrpoRpxltDZKi+Yb0NoB
UWIhzth9/p1nfbDvbffNKuv1mNC9Q30VVUWxxvwl7oXpxFqhVTZi/50qyfDxCxSw
mPI576Yl7jQb1JxegNjqwuftjuwzx+2iA80K9huTLty3tVtsjYDsZAEX7wl8q3Oz
93TZm1t98fKud33GY6W9zKa6v1rFdpt1GJVpTFNrHDy37GCC99Adf1igImyktFa5
STOzL3kpSvkl1b4cxv94jOfzsS1DnFtVZ73Isd51HBlkZLff/YwR+MCpdpIogms1
OgKLKmiG3PRe+IQmMlT0lqcHTRBssXFhSrscDm4nPPBikoM/SnlYOy/xUeZPui+o
6IISs1rVWWmTfrfOAH/3mqd7lC/0ccWWHTfAySW3WKcdNnxCmMo1aPYQcyiHgWjO
vKHaYqBKMoDAAyvbOgtMEW81clLQG6CTe4DuQXN8QFjAOboiXDKj1UUHvr6DOQgY
fPzN1Y7Rbrg02Qd1SYORD5hDi32mkLsl7I4jKffnbdG6IiWB/WB/mnVnhGvgI2cr
VQnpO7n0Tq+ZMK79JSqc+RD2BxqWTqN1B+4A1kuMs31YcqQZ/Kn0OVg85w20lsGB
mvsseWjy/Q6ta+nB3dAqo0cCkpoD/yz9w4ff4KON6N4AvchjoPTivzjyFzqwJw4G
9VN6ANLpVZnwtPO7rTSpX358jJ+MVvfgB5qvAuhp4jTyliwMkPiL4Ot6GQS68Rb0
NVKWLLFt3eghmjOzxWUmfnrSGiPzsiKd3Gdu57WPsm3GmJ1DTSKYY64gTzT260l8
9J9ZvF5y31JBhe32PTYPRPH+Rr5PriajYS6gEcJBjsU6oYpAIC64E9VISxYBl9rQ
vwVzyqQ3d8TjeD7jjzHqmj+9su8CGz79wM+pmcc22WB5saOd6aRYDcCM7wtIWQbP
1nSkvGwI+LlPpjK2K5SVJcw6ww8Cxb4U+3eq64NFaxx1JD3noFj7wIPgpYVwfJUy
iQ/GxIQ5H7+KrC9/aoRZ4qzymS2fuKCu+LMOUbMDJg6UFFnonagZvkOEJThgQZZm
CTA0SZLWk3YP/mnnQNwqp2QZKEzkYt8KHN2lWmyr8p1AECyMJuhL3s+gVc/bN0ra
L0tEMJ5TDVVy56aRjqesf26MxpeFdOM2pOGV1jpbuxJf703lTmsQey+Yx5W/2+0w
yzGbemb201EjKtsboP+TAYbfGwObRHEws3/i8aI2WzuHZIIPFNUOuLE261gNglSY
O9bhbyhagnQq2NlJh6tPYNGYHrpjePSx2EA/sFrJJmglMHW8G9HYp1b+3OXFsomC
0VEl+xXXAR8Wfpj7Rrc+wPJyiuQO2M8OzeEgZKYY6ealjLVVFh6p2PFZR+jhJPSx
Tbbo6ZKmMs5EiflgRB1Lb3+EaNsGZIBl1SAt8uZb6BI+rPgqP5Gtan6N4XBN3dO3
1NoaF18jeG7+SywEYw7OC0HuKFpa9kyFqSUZoMnKmMuWmoooFIV8BHDxbYU9uwR+
sEXjxdYF6U3w4Iv7qdvjNKhPQmGX844rPv2lDH7V9N8I+4ObWkfjWS2gJZ2OHPM2
B52br6lKLLaMBYehsQbioEEZLVg5NRg6R5G+FAKYEDOcMIBt6NdNWtdjcHCIANly
N+p+6zdX6TdbkZBlz6VPvfH+ledRIo7UVY/g2rrpQ9Jta5WfJ6givkxnkB8vtj02
kuH2bnxs8PjmC6lrNzovSsSO9eE6Mnpbngn1Qdj+KIRLVggekHZQ0mxd/5xkF/6Z
GZTqyAdCk9ElzvqXEDPwhl1X6ZJ4xxjLxlEpVGGo2KfhNAddEl/GukfEH6J9R2qc
YZJCUa6B2QmHqvdZ3eGOusQiS0RKgodcoyxNrezjdoTOyYDiBn9RHSPTV2GmDONO
ZiROy3h1XMo3SwMrcmPpxC7BOB3zIdj97hZlDnPHrVN22h6mWQwmt/vNM8cZe5DN
UtImZlWodX3hWmwGmCkPeliobaUaVw11WbHspOhfwuYZMuDjIJuffS5hVMLoIri3
+r+fc3ofkuwIY0tizT0/xpMJ+krmUUBqFzP0ephw2XrO7/+UZ3OfJLysGp/bvyFv
wzxZfD7EMRrqLksEU0f2VnP62fpyoh0GUj01Cn1cauFIYqKOCb0yWxrObb9yZUUx
FCb1YhhAQipNu+g0JH51mbGZD3z2n0s2nXpDWas98dYATNuPIBvKaMZPLtRg4esY
6SbDInq9HsEWJbNyBY6Uoe3WaCG58FVZg2ZUcrBiUx9M+1cjGM1ARUfZHMcNKi5G
G60Lg/pFij5jeJjwbg9ePLTvHUdLl4+jDmwACnb2JxdwFJv5IZ4ae+5kmqkxBdD0
Nkye0qIh9Y28ZAM4G4mdt9zlsiYV6bXKL3tO10GnXzMTZtpJ5Bv7zWWRyQMxYFbH
wLJT0gyckOI7alW12Fv/UKwFR+Ep7PahRLh2Y+En5SzeNrS02upzJZvj/tCMryFh
iWTv/jdnzbR3gH0ZG07BrN63oOXWbLGgR/nDi25iwGpUM8Eer3HZJ4Ahjuk77jL2
W5W0QvSPd+F3s4TEuBqYwa0mLuoYvcbmOuYHDikS4hQbpwRlpxs0BLGXzy4z0yNu
HMXgvDItLE2wY/wvUGdI5cuVom+r0ZEME/QUZ7M3hqevjpwPfj592tnk14Yqcn/R
zhngiiwHgJegQMYl3tXQYu2En6T9Lu2Col+pO3xPMv3TUetyYxT11DpzpJk7gbbg
FqCU78FYWqGh2NQ0JLzcbnWCEMiOwGsyrmj4N3Awov/C19ug6Hj2phNpBiAHSbg+
0isgVJ5ReMLjk1XxLLd80Lere6luyTy6OKJy6npvNcHaNr0pJRNybI+NG/zDRzwn
GMwQVpxh7JebjHLh7kOhQeVeD4panCjVajU6t/Y8ATX5Xd2vM/2fiO1jHjjs/7pe
xBJ8KXOc/Y7u5enjdK1yzCQq/h4y0rFpMWbgENBecFXTc7itr2Gj2IjQRij6bTFc
A75ESNe6aCHcAI+4A31pBZHmpaHDKCUVY2g1I0mnMWdHYriALKZZLN8iDv4mo+Uc
+YFv0o8eSn5PHf18m7FdRSmD4SaCxSaGoAYibLOxP6Bnemod+OZTnGhraukQXNUV
qojnyjpKksWukUOYsmTn689M76seLJds8ZEAP3Gy3XnkaW28O6bHtFXz+SD9a5QW
kLCOSC12qHYaQek2sT4pGrjikIfY1HMXQ6bJHUYl0hXWKSde2xqiL1flSPiXFZmD
scA84DiVvPi3yK2IM/oj7Lu77IXthNVX1V1KN51BcLjL/g0XNFlcYx3JSy7qYiOH
7sp6GM8QKbx9NM548IGg/vAAqna2MP+If4q9iobkDBRGRP/747c7+UWaml3EN/bv
ATtoo6A0DYwDYaaSIGMJC3TGgftz9muTkpb2FNUv3B9XtteM8afyzGT2SO+QraXl
fD2v68y+X18ZVbK0ybRmKgyUmoTieKMpWniyRszsallCD17iAYetp++B094lz3ag
6EVKf4tl+f1oXK+Xn7JMj5uIbHdSc6eEO+miCaGvdLrT824c8mydn28ea0HnWd9r
pkkb/oC5glXEMVzPLvOldFrSpulYg27YbGasTKpQcvGolcHfApxhE0DSK4+XGTrV
iwBpD3jViiiCT4VfSSV7pw==
`protect END_PROTECTED
