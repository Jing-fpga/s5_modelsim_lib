library verilog;
use verilog.vl_types.all;
entity stratixv_hssi_tx_pld_pcs_interface is
    generic(
        user_base_address: integer := 0;
        data_source     : string  := "pld";
        is_10g_0ppm     : string  := "false";
        avmm_group_channel_index: integer := 0;
        use_default_base_address: string  := "true";
        is_8g_0ppm      : string  := "false";
        silicon_rev     : string  := "reve"
    );
    port(
        asynchdatain    : out    vl_logic_vector(0 downto 0);
        avmmaddress     : in     vl_logic_vector(10 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        blockselect     : out    vl_logic_vector(0 downto 0);
        clockinfrom10gpcs: in     vl_logic_vector(0 downto 0);
        clockinfrom8gpcs: in     vl_logic_vector(0 downto 0);
        datainfrompld   : in     vl_logic_vector(63 downto 0);
        dataoutto10gpcs : out    vl_logic_vector(63 downto 0);
        dataoutto8gpcs  : out    vl_logic_vector(43 downto 0);
        emsipenablediocsrrdydly: in     vl_logic_vector(0 downto 0);
        emsippcstxclkin : in     vl_logic_vector(2 downto 0);
        emsippcstxclkout: out    vl_logic_vector(2 downto 0);
        emsiptxin       : in     vl_logic_vector(103 downto 0);
        emsiptxout      : out    vl_logic_vector(11 downto 0);
        emsiptxspecialin: in     vl_logic_vector(12 downto 0);
        emsiptxspecialout: out    vl_logic_vector(15 downto 0);
        pcs10gtxbitslip : out    vl_logic_vector(6 downto 0);
        pcs10gtxbursten : out    vl_logic_vector(0 downto 0);
        pcs10gtxburstenexe: in     vl_logic_vector(0 downto 0);
        pcs10gtxcontrol : out    vl_logic_vector(8 downto 0);
        pcs10gtxdatavalid: out    vl_logic_vector(0 downto 0);
        pcs10gtxdiagstatus: out    vl_logic_vector(1 downto 0);
        pcs10gtxempty   : in     vl_logic_vector(0 downto 0);
        pcs10gtxfifodel : in     vl_logic_vector(0 downto 0);
        pcs10gtxfifoinsert: in     vl_logic_vector(0 downto 0);
        pcs10gtxframe   : in     vl_logic_vector(0 downto 0);
        pcs10gtxfull    : in     vl_logic_vector(0 downto 0);
        pcs10gtxpempty  : in     vl_logic_vector(0 downto 0);
        pcs10gtxpfull   : in     vl_logic_vector(0 downto 0);
        pcs10gtxpldclk  : out    vl_logic_vector(0 downto 0);
        pcs10gtxpldrstn : out    vl_logic_vector(0 downto 0);
        pcs10gtxwordslip: out    vl_logic_vector(0 downto 0);
        pcs10gtxwordslipexe: in     vl_logic_vector(0 downto 0);
        pcs8gemptytx    : in     vl_logic_vector(0 downto 0);
        pcs8gfulltx     : in     vl_logic_vector(0 downto 0);
        pcs8gphfifoursttx: out    vl_logic_vector(0 downto 0);
        pcs8gpldtxclk   : out    vl_logic_vector(0 downto 0);
        pcs8gpolinvtx   : out    vl_logic_vector(0 downto 0);
        pcs8grddisabletx: out    vl_logic_vector(0 downto 0);
        pcs8grevloopbk  : out    vl_logic_vector(0 downto 0);
        pcs8gtxblkstart : out    vl_logic_vector(3 downto 0);
        pcs8gtxboundarysel: out    vl_logic_vector(4 downto 0);
        pcs8gtxdatavalid: out    vl_logic_vector(3 downto 0);
        pcs8gtxsynchdr  : out    vl_logic_vector(1 downto 0);
        pcs8gtxurstpcs  : out    vl_logic_vector(0 downto 0);
        pcs8gwrenabletx : out    vl_logic_vector(0 downto 0);
        pcsgen3txrst    : out    vl_logic_vector(0 downto 0);
        pcsgen3txrstn   : out    vl_logic_vector(0 downto 0);
        pld10gtxbitslip : in     vl_logic_vector(6 downto 0);
        pld10gtxbursten : in     vl_logic_vector(0 downto 0);
        pld10gtxburstenexe: out    vl_logic_vector(0 downto 0);
        pld10gtxclkout  : out    vl_logic_vector(0 downto 0);
        pld10gtxcontrol : in     vl_logic_vector(8 downto 0);
        pld10gtxdatavalid: in     vl_logic_vector(0 downto 0);
        pld10gtxdiagstatus: in     vl_logic_vector(1 downto 0);
        pld10gtxempty   : out    vl_logic_vector(0 downto 0);
        pld10gtxfifodel : out    vl_logic_vector(0 downto 0);
        pld10gtxfifoinsert: out    vl_logic_vector(0 downto 0);
        pld10gtxframe   : out    vl_logic_vector(0 downto 0);
        pld10gtxfull    : out    vl_logic_vector(0 downto 0);
        pld10gtxpempty  : out    vl_logic_vector(0 downto 0);
        pld10gtxpfull   : out    vl_logic_vector(0 downto 0);
        pld10gtxpldclk  : in     vl_logic_vector(0 downto 0);
        pld10gtxpldrstn : in     vl_logic_vector(0 downto 0);
        pld10gtxwordslip: in     vl_logic_vector(0 downto 0);
        pld10gtxwordslipexe: out    vl_logic_vector(0 downto 0);
        pld8gemptytx    : out    vl_logic_vector(0 downto 0);
        pld8gfulltx     : out    vl_logic_vector(0 downto 0);
        pld8gphfifoursttxn: in     vl_logic_vector(0 downto 0);
        pld8gpldtxclk   : in     vl_logic_vector(0 downto 0);
        pld8gpolinvtx   : in     vl_logic_vector(0 downto 0);
        pld8grddisabletx: in     vl_logic_vector(0 downto 0);
        pld8grevloopbk  : in     vl_logic_vector(0 downto 0);
        pld8gtxblkstart : in     vl_logic_vector(3 downto 0);
        pld8gtxboundarysel: in     vl_logic_vector(4 downto 0);
        pld8gtxclkout   : out    vl_logic_vector(0 downto 0);
        pld8gtxdatavalid: in     vl_logic_vector(3 downto 0);
        pld8gtxsynchdr  : in     vl_logic_vector(1 downto 0);
        pld8gtxurstpcsn : in     vl_logic_vector(0 downto 0);
        pld8gwrenabletx : in     vl_logic_vector(0 downto 0);
        pldclkdiv33lc   : out    vl_logic_vector(0 downto 0);
        pldgen3txrstn   : in     vl_logic_vector(0 downto 0);
        pldlccmurstbout : out    vl_logic_vector(0 downto 0);
        pldtxiqclkout   : out    vl_logic_vector(0 downto 0);
        pldtxpmasyncpfbkpout: out    vl_logic_vector(0 downto 0);
        pmaclkdiv33lc   : in     vl_logic_vector(0 downto 0);
        pmatxcmuplllock : in     vl_logic_vector(0 downto 0);
        pmatxlcplllock  : in     vl_logic_vector(0 downto 0);
        reset           : out    vl_logic_vector(0 downto 0);
        rstsel          : in     vl_logic_vector(0 downto 0);
        usrrstsel       : in     vl_logic_vector(0 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of user_base_address : constant is 1;
    attribute mti_svvh_generic_type of data_source : constant is 1;
    attribute mti_svvh_generic_type of is_10g_0ppm : constant is 1;
    attribute mti_svvh_generic_type of avmm_group_channel_index : constant is 1;
    attribute mti_svvh_generic_type of use_default_base_address : constant is 1;
    attribute mti_svvh_generic_type of is_8g_0ppm : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
end stratixv_hssi_tx_pld_pcs_interface;
