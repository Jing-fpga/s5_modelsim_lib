`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8IJAFUf10DYNYUh+/ThmBa/zoY2wkH/QuhMep8+DkFvXNhsiawSEo32VuDjxkK3O
t5mv9qZxj1VD3c/TGaUnOoG4Sv1qK/duap3vcgmEP17w17L+sErB3co7kNYoKEvO
dRq7xjXmw9wllVdTyFnUvvucE0nSFEUxG/KKN66oVxPLwHmSlxTPExxyyPf4eQUQ
EolMy8RJzBtb0pizitoMg4nvykbewtFuf1WGf2rg9xLq9IvKgn8e6GyFSchkN2nG
dg1740cVLry2WcOU1WBL2JSrNyuvA44hdGOk9IbCb1WNCAcwJniesxZBcQr1WUlu
9Lsvq37j03H15CnkuiXeJhao7LSDSQFZRRgWEJf4ZTTHY44btY3dTWr9h5KrZswo
aDHQ9UKRcqMlzUdhvOJQq+hQ865J/xPyWPKBV7HG+kSk5/jfnUmaa7EDHeUUBCch
jJotl1ta86iG7GdWF7bVIPbXwTheKXfMby96zfPqgDH06ynq7ymPElUTStE+1sCW
loap8G7w4K6QiCavACCMr4NP5QwrtSW8FA6LEidBhxsTT8CkFgm0aNewpoKNGm5W
F+lHxQ9zMVDKwc+UQavysHiB2xMHKMEsq18osQj9Z93OaxXxrNl2CwiNO3a2AU0d
/lSUcELGTJcMjqDfcH3Y4oQcIgoJ67hHs8YBmBh91w4=
`protect END_PROTECTED
