library verilog;
use verilog.vl_types.all;
entity stratixv_hssi_gen3_rx_pcs is
    generic(
        rmfifo_full_data: vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi1, Hi1, Hi1);
        rx_test_out_sel : string  := "rx_test_out0";
        reverse_lpbk    : string  := "rev_lpbk_en";
        mode            : string  := "gen3_func";
        rmfifo_pfull    : string  := "rmfifo_pfull";
        rx_ins_del_one_skip: string  := "ins_del_one_skip_en";
        rx_force_balign : string  := "en_force_balign";
        decoder         : string  := "enable_decoder";
        lpbk_force      : string  := "lpbk_frce_dis";
        rx_lane_num     : string  := "lane_0";
        rx_pol_compl    : string  := "rx_pol_compl_dis";
        rmfifo_full     : string  := "rmfifo_full";
        rate_match_fifo_latency: string  := "regular_latency";
        user_base_address: integer := 0;
        rmfifo_pempty   : string  := "rmfifo_pempty";
        descrambler     : string  := "enable_descrambler";
        block_sync_sm   : string  := "enable_blk_sync_sm";
        rx_num_fixed_pat: string  := "num_fixed_pat";
        rx_g3_dcbal     : string  := "g3_dcbal_en";
        rate_match_fifo : string  := "enable_rm_fifo";
        tx_clk_sel      : string  := "tx_pma_clk";
        parallel_lpbk   : string  := "par_lpbk_dis";
        rmfifo_pempty_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        rx_b4gb_par_lpbk: string  := "b4gb_par_lpbk_dis";
        sup_mode        : string  := "user_mode";
        avmm_group_channel_index: integer := 0;
        block_sync      : string  := "enable_block_sync";
        descrambler_lfsr_check: string  := "lfsr_chk_dis";
        rx_clk_sel      : string  := "rcvd_clk";
        rmfifo_empty    : string  := "rmfifo_empty";
        use_default_base_address: string  := "true";
        rmfifo_pfull_data: vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi1, Hi1);
        rx_num_fixed_pat_data: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        rmfifo_empty_data: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        silicon_rev     : string  := "reve"
    );
    port(
        avmmaddress     : in     vl_logic_vector(10 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        blkalgndint     : out    vl_logic_vector(0 downto 0);
        blklockdint     : out    vl_logic_vector(0 downto 0);
        blkstart        : out    vl_logic_vector(0 downto 0);
        blockselect     : out    vl_logic_vector(0 downto 0);
        clkcompdeleteint: out    vl_logic_vector(0 downto 0);
        clkcompinsertint: out    vl_logic_vector(0 downto 0);
        clkcompoverflint: out    vl_logic_vector(0 downto 0);
        clkcompundflint : out    vl_logic_vector(0 downto 0);
        datain          : in     vl_logic_vector(31 downto 0);
        dataout         : out    vl_logic_vector(31 downto 0);
        datavalid       : out    vl_logic_vector(0 downto 0);
        eidetint        : out    vl_logic_vector(0 downto 0);
        eipartialdetint : out    vl_logic_vector(0 downto 0);
        errdecodeint    : out    vl_logic_vector(0 downto 0);
        gen3clksel      : in     vl_logic_vector(0 downto 0);
        hardresetn      : in     vl_logic_vector(0 downto 0);
        idetint         : out    vl_logic_vector(0 downto 0);
        inferredrxvalid : in     vl_logic_vector(0 downto 0);
        lpbkblkstart    : out    vl_logic_vector(0 downto 0);
        lpbkdata        : out    vl_logic_vector(33 downto 0);
        lpbkdatavalid   : out    vl_logic_vector(0 downto 0);
        lpbken          : in     vl_logic_vector(0 downto 0);
        parlpbkb4gbin   : in     vl_logic_vector(35 downto 0);
        parlpbkin       : in     vl_logic_vector(31 downto 0);
        pcsrst          : in     vl_logic_vector(0 downto 0);
        pldclk28gpcs    : in     vl_logic_vector(0 downto 0);
        rcvdclk         : in     vl_logic_vector(0 downto 0);
        rcvlfsrchkint   : out    vl_logic_vector(0 downto 0);
        rxpolarity      : in     vl_logic_vector(0 downto 0);
        rxrstn          : in     vl_logic_vector(0 downto 0);
        rxtestout       : out    vl_logic_vector(19 downto 0);
        scanmoden       : in     vl_logic_vector(0 downto 0);
        shutdownclk     : in     vl_logic_vector(0 downto 0);
        skpdetint       : out    vl_logic_vector(0 downto 0);
        synchdr         : out    vl_logic_vector(1 downto 0);
        syncsmen        : in     vl_logic_vector(0 downto 0);
        txdatakin       : in     vl_logic_vector(3 downto 0);
        txelecidle      : in     vl_logic_vector(0 downto 0);
        txpmaclk        : in     vl_logic_vector(0 downto 0);
        txpth           : in     vl_logic_vector(0 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of rmfifo_full_data : constant is 1;
    attribute mti_svvh_generic_type of rx_test_out_sel : constant is 1;
    attribute mti_svvh_generic_type of reverse_lpbk : constant is 1;
    attribute mti_svvh_generic_type of mode : constant is 1;
    attribute mti_svvh_generic_type of rmfifo_pfull : constant is 1;
    attribute mti_svvh_generic_type of rx_ins_del_one_skip : constant is 1;
    attribute mti_svvh_generic_type of rx_force_balign : constant is 1;
    attribute mti_svvh_generic_type of decoder : constant is 1;
    attribute mti_svvh_generic_type of lpbk_force : constant is 1;
    attribute mti_svvh_generic_type of rx_lane_num : constant is 1;
    attribute mti_svvh_generic_type of rx_pol_compl : constant is 1;
    attribute mti_svvh_generic_type of rmfifo_full : constant is 1;
    attribute mti_svvh_generic_type of rate_match_fifo_latency : constant is 1;
    attribute mti_svvh_generic_type of user_base_address : constant is 1;
    attribute mti_svvh_generic_type of rmfifo_pempty : constant is 1;
    attribute mti_svvh_generic_type of descrambler : constant is 1;
    attribute mti_svvh_generic_type of block_sync_sm : constant is 1;
    attribute mti_svvh_generic_type of rx_num_fixed_pat : constant is 1;
    attribute mti_svvh_generic_type of rx_g3_dcbal : constant is 1;
    attribute mti_svvh_generic_type of rate_match_fifo : constant is 1;
    attribute mti_svvh_generic_type of tx_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of parallel_lpbk : constant is 1;
    attribute mti_svvh_generic_type of rmfifo_pempty_data : constant is 1;
    attribute mti_svvh_generic_type of rx_b4gb_par_lpbk : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of avmm_group_channel_index : constant is 1;
    attribute mti_svvh_generic_type of block_sync : constant is 1;
    attribute mti_svvh_generic_type of descrambler_lfsr_check : constant is 1;
    attribute mti_svvh_generic_type of rx_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of rmfifo_empty : constant is 1;
    attribute mti_svvh_generic_type of use_default_base_address : constant is 1;
    attribute mti_svvh_generic_type of rmfifo_pfull_data : constant is 1;
    attribute mti_svvh_generic_type of rx_num_fixed_pat_data : constant is 1;
    attribute mti_svvh_generic_type of rmfifo_empty_data : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
end stratixv_hssi_gen3_rx_pcs;
