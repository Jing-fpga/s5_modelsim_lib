`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fuun2GwgUA6dgbJxCXGRs18xvJRCpzyuW0OBy0fix47sy6RxOcj5ZaPAYGL+Cdqk
WlLnXop2nlq0c+U9CR0JJkd/lRwSWAwxW9Hx3LIRN6pP1fTc4OPv7ZBpC7gxl0w/
oZ+iAvIrhhK1g2A2K/oCBTH1rplK181l2P3Fc+LxB5pJCJriw/Lh4nY6RzPK0fbr
o+lJdWZ6z+/s+YVJ6ExGWBPn3iGbZ/eYG/9f+cVMDTv4wxOyrqsa4ks167hyr4xV
97GEPvFPe6IqPTHkAuO1d3/iUxoQWeideIB7P6RiTkB14KBPOEL+TpoqnndnAW1a
joVk//CTv1zyFiIR/3ydM1zX9vT6HhyyBEWHOoHHpqRUSMX8ZXzox0S9VtbtHrBY
rLXqqh90u0PxqcEHrOVj7zmlDaeF3wWIC1l0hZGpqrjx1SZE4VXO7AyZPcUmWAk2
OFl8lzznMz4jSxIFhLZfUZFW8F2rO+cawu7zdCaWAXo=
`protect END_PROTECTED
