`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fJ3zhw3EI/SHmEaN7EchlzL0OTRuQEfoVx9rQR/IhFbzSzxtQ3jQds4Zxhrh0QZE
ITejlX0BDX6ttAWcpdGqnxBMnrVdMRS1FCweXFkxIp8bDT4B51ttQIzUdVE7CppB
qSG/qFHStROhhOCZnB8Sz3XQzbMgfKZ37MT8l0nl/btuF8cnEUXT5f3UhBPlPypP
rj/sXaOktSjMhhb288itPz7l3FsOQUZAmw4bIiyP6s6DaJ6t/k6CXceUj/mKc20D
VVXZIodr2kK4rfYKnWj/IQ3h/Q9KAIQYWqUTRkXYU7oqkJV1MP8iXIfgp5sJno9m
Zjk6ZeAQpHddCmo9UzqCnEUVFTYmWfxJz7rwDb5v4ezOygLkDATFS3yI8JC23uEu
dX+3iGIcj7eOfFQHj8gDOmoQnKoVUTkVqkgJkRCR4NBS/P7G+2A58QXHl0XMh8Ir
lf8o6EpCJa3a02Lx7lBR+pgOltCRsOWrDhFTOoaBdc7gtDHu3Yy6Rkg58e4kG1U6
+VNOtlhOetJKFlUxQf5GV+PqZOS4GYHKZcny4nmXhOo1bUtPjDhmlx/LTrnFsk6X
mkW7fx/onpRzP37oHpCxTnmun1HeynUwE767n83JKPnRXE4D6y3RPpdoUfUI/5Sa
8kg9IWfhhd24doopOxhdjEnoFOzgPoSviT5F2ofngSH8pqgwIt1Zpbk7SxwAp6AP
saa5jyKAJ1t2hoVx01xAisXJWSSmOnrdbi4NsQXFf9UVYmIR7B/1x+nwbANyiiy5
j6hJV7R7s9qaxyF17cBYrNXjN4ODLVozibvqTKyqAQB2Up/nVDdBi/R47+5/tAXL
b+m5sABO1TUbjYbEQk5AEbbGj+UQvou6t/pDA6b1KuLsnhFn+9Di9wW8iIZuGQJI
nmTVCdHIeaAFJ0QmvYs4SJDTgk80zFWFhpMbvD8VjlCv5dBx79WEXQI072Icmdre
enfY6ZSoA6oUPD9mkxmEx2F0KXKIwejJoX7WXWqW5Uwg8LNKsewYvlfKw2SaXwJl
RviTA4GPOofcOauAy+pn92XZwnj8i39bvtlX9960OiLCk6m3izZCQ2tK5ll6ePF8
tSbmWd86+Re5qWj1OH48TSMyFV15aoiHiEEJz3TXRluuOuAf85Y1gBSZs8PXv80f
HjBrK0vbH5XiHM7AbAES94EoOzjGpw+2zJA4BKBgg7yX7caigsWwa2UI4yhLvySX
p7RrNIQF57hNSyknqlXLxb3r8TN90TRwQ9iw8TI/XaXgFomntGjOlEwar4BL88DQ
XdZt8s8Mtcb1KIT/DOTU0Hlx7q7lFftRRJ+NG03p6EJtiWE+N7WkSFyaE85TGLrM
zYJei89K9DgNV+ST1I+irUPNGgqqP5F+UlH6tLo5U9WO/eUY/pDIkCjx6ktoy4no
8EXXyW6iEaupELC1biq/HFFVHRls6ClrV2NfE6XnSWsUXA9A9o0tFIivM70jUn+N
XVEMb5fziKdr7pb+LbBkwLSiY7raX/9MDEf1JYyZT/2ekCPmCik1wdev/xSEHhxA
bpk7oYNqGsP6YATmvJP6IYPsmqzUUzyqd+S8eL1vsMCOkBMjETFtBiGHO6guMGO7
IOAyTnJwtufPq+b93DQ3djRJ7KTbaLGkJyddHUq/p727ia1ilf2I2RtrEahhf6xY
pscvoeNe3y1gvRzseSZZ31BzQ8jh16SISYbofq24EuHgCo1AXonaz/Yvvb3TL/bu
ZtwMFa9yealgHAxdTKfLg+L59Ggs4eq2WKOxGQEECBO+ujlMGJWM/nsXlX4LbE+N
tFx1ANboPVzUqHO71J5DUDS1EymBS4TZHjWLW7ANPjFd6NuTPkNvs+Puj4eSXpmL
jIOhZzslCVSQLM8qMX5XGrBnfRFGNFrEvX01tmq5usW86CB/Rzunu0rjS1mXZHbW
JIg/UpQkI8TlDp8E6oSOpkbaGTsTgxNs9KeUM3KY81FiPugnHbDBxHwJ6eRuhHDq
dvux7kZS5xGYQyrSkuhR/BGWR25HWeVGpTk6AC9+KuMCAEs13akJUGFnm0rvJYek
ShUJ0GU7rQEiiXvTwXn9MzIbnEDdIySA/1c+azWxHAy7KBb1ra2zmYrJuNdk3g0A
5FrV9uXZLlrT6uTNCfyJXUlj5LfQ2iflwR/W/swwfbmJQftkoGvY7VQ4v20atTK8
SiJAgVgupqSdke6I9X+/OxFN6iUx/UyCMdg6LXVaHN6FrXqrqiCpYoLbZObzvuSy
Np6AhP56CusMEpilGNMrFlySAZC/I/RtwdS3MoAKr5AdgLzQrUOLiL/N+pKR9YtS
8p4zIIScSGa0hClz+RkrLQ321pw0Yh32OTWffdkYo5ULXnqpaqr+JUa/KKiOoPov
K3NJku5K8WIb4tWkE3iCndQG0/7bLI1WYfepi55z2APEn0B174CFb/PRmViTAu2J
ZKmiYknO3Y5BSOWeLLrV6VvmIvxghETrIWB38GfC6OeGuMwQ+Q3/7gCGw1+1xYn9
2WY7eiVBAUqryMOnVUXiBC8RjLUuY97ClHPUiREf5xI8XJwfuMWpyhSGdjQcBOfv
+L7257As27o/A2GBcgtUtnt+UwDwkPVsEKL/Ezwy8xzKFR2aASOXf7syNTx91mr6
Fj9n6kZGtnYly/73paZnAQ2iOCR4+jYCb7+BkI0/z2Tt5nj+XDt4qaBCLS6utMir
yuIKJ2max3t3lrnzJ7TsFnXymJsEo+ZTJ8NrEgOeA69WsVdw0mknvFGnJIpwZK6i
Y7YRU1vh2F65i2kqQ/DyDnsT4fyqNPmq3PB6zuYt7po0fycduMOQ7TODP4wYLHEN
ggncKtdwihaiDr2oNe3DiO9W9ZxqNnmB+9BM5JcngA5BhflR3RO28A1iQN2OAZ+r
UqdGxA1wnGtmYkqXfOYmpIttWc/qhEOg2TN/fGauRtRkPVClA58FXJwbBbtLmiz+
Q18/wuNqoLo7ZjR4s+u3vIy1egpxzfSBruDgK9sMoWbU7npFTV7tBpUGQ1eSBsEu
bxUBohziyH5EggLraneal/ck9D0hCESmedNcwe9MsWcSelpnf89EsechFUmiyCUU
UfpC7OvNmbibTzwb9lEJ3SzhDcoH5iF0sXA+92MSloc/PkdSluV0OJISpZXQxCF9
HgB9y9HDdk8UsYwOAapGvULOS8qoovZQopELxyDwvR18AdxAQ6Vst12yWhnUjGXe
M3kLH7gvVp8N780KhhYVggPuxFD5KKcnD3gds9jbnpuYj6GWOQhDP1DthvURWKJM
nDdvE8Euk+HSoT9j5EyJnucnKzK4pDtBKenVk88YXeWVKO4yI2DQh+RY2nbtPQMh
e0rxZcwhzvWMY4mRZfJmdqmuXmdT6Uuu8NnXnvrCIifEjo59FqKOfK+/yUR3lZAb
O2JUxB/AFuregA1DmFqXjFfskFN2WSHXsUFT+U0LtK+wqFgL/5netMb0iBPFjDDb
JaB5Bq4Nb1FUbET3uaSUOiYFQhmbijulToyEMNxbQoyiZqtYMC+VCncv42phP77n
LiC9abthD1gNzfY1lO7gcS8kWy+hbVY1M6B1O1A6L66yRvXGUvckwdo4U/Ue92Ui
yMVGO9GbBMgDjVmf/SCdpMp7qS7UfCwYwyLOHJXYJy6uyp2YQcrfCGyA8GhGOFSY
5hTrfLmD/D9H+XQ4PmVwC/4n9zdbJ1vaG6e+4da+Mqkn5Sj9OLgXZ7bwHV8d5NtK
n8X0PgKNkV4IojbuhBhXBkNIz4hWHTsNYBLhvGpJRvn3lTmEJJ6EhsIkSuPNgxvz
VLwYN4NG3xXvr+VBKLLkiBTIY1J+BuPJteqwSNhCKlLoYkzJQ0qYlgZYA6FGHc/t
kMNm2FOEQhpTeWB0UJNqFBilzLSCynHxsImxHXt7DfGNkPCydAmcYd0k7ozEfTcT
MzW12u6Q+UF5mQIZv4j+jZnFvg+r98V1EJjDMSgHPDRgHJD9AKwxLKmEeO/EqAbq
VEHPhN4d/a7Zlt9kmxxl+MBbgcuUsUusBPMbvkEZb6to5kKTmNXwkdlMnxMWjWN6
uqlyMrYlQFjULVcZk4iOlTwOwz2xaQ2xD4mWkA2zCykwWJpL7phhATHq68wIixdh
dQoMd9PCNSAFL2lSh4/MOxOAn9LX6XPwwy8VpBB2RcgJPy2xdaIsSkJM+w1Vv6FJ
33c/l1DLHoI6G+Vf6uoNNBToGnozd7Uswb5VCCV9yhJ6utrxrPIwoszdyL76ZLZi
JxvZd+JijRqKg55eux2UODZ5UHVXYZljuF6A31LigiCMwmFEDsn0204jHNBSHp6x
n331Vjg2PmeqQx7u8L7a4MN5kZpDOVop86gJ9YrCdkuthW3yrSe3Ua1dovoIoV/W
o1pOclsukBkHSooXGcLsk/EAuwUW4hXWCX4o93qNZgB5iihZei4gtJeUVEk+ae8m
heg+ssyvDAxUCvTMsDtf0VA2LXVi70qKBemYDHS+MDcrUpgVcYKs//R1hzqtwS9d
/H5wex8Kg196P/W6K1jd+0U9gBVidw00SpzZRrbmUZwfv7gfOocselYbx3v+qbrF
oha9HFJtAiGyG96jS60YyxgUF09C/YlglT6zPcaAQ1M=
`protect END_PROTECTED
