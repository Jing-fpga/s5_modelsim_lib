`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PVcxFlxbQyXMmB5UDM0xJORIRNCPrt98hwOvmiXY2SCPF4bmGn6bIl7s332SF+rh
hHiU1H/C+32fRgy5wyHHRU/30ut4B/e0G4EgL/+k7U0kEO95b9EvvIVuAk4l6jQC
ycogUrehOboFJH2NVJl7uG3Lf5YelHTcjF8aWyU2m/UD8Kvt/8MZjRfDSlg5BCO6
4CTyam0V5zw7rke6LBaXdjqtpN5clnzL+Gi42QyTQ1Y8o+0I8tzd6OgDzzb9P1Tw
HqiY7eoo45t3C5q4wE9a7a0Ddk+KnTW2VFjZaBglpJyiFEFv/Y8UUQwGAbaEPBs/
IjCvRG896vSzKedObRzG5jJyxCIopLbhJHf1sq9q6ZrUcbDC0Tgx4FESTqaand2N
JKjMS3Ant+p6RCNUdL14jCGm+Tss+uTFfUiCOmdTn9tGO+H1jhTXddeNvF0iTfJD
WwW/6vE5L03tNhKDsvGudPtVFNQ8hPGEU5kRhMdgTVumcJ2s7u6Lyyv9sNF/LHih
JevAHpSKnDT9zOYazzATTH9ADfnrp33C6xOQXxl3q3GYZLw2K8Kj0ShXzOFNJpkm
jm5dji+Q1iEbsjgMoIWMdQXCFJBPYvLNXMpjQcQg2fisQDS3wR5megHi0Rjy0A69
lE3boS7r204i0oNf0cBaJnYXWK+q2yfOgMt3sMZNNykD9E0CQWbRB3BD3tfaZ+tx
x/BwFQ15iX6ZOa5+FPFGc8ZR0rNJY4FYoot7u0OWzwZNVuY8yOciXtzLQzl13BXQ
whlBp1f9dZq+3ou4lHJArxf+/Ffzey/izlnL93pBnROJ0dxxd4Aw38ibGpGx3eXT
O6/zjNPDropgs6JdXEdTP43o1PE1b6nKYfsAHkw2jiBpElcdMOc+Mp2Le1P6TE0s
GzD1FqK/z3LplkvYhySiUJ/4V+ks+kkxBqdW6p/3CFZdnaJhyngTmyl2XkUhOrLD
N1E7BZ+5jv0N/4xTMfUey1TlojDmRmM98hrHNBh2xBN3zCNwpevVcKe9fuNgFAvz
uW1wiFkMPb33xFVIxJJnPegm1oaKylB7J8pJiliwI/Ds9IsD6iRImNWE2lrvMWSO
B+i+ilh81ueKDrMH60y+Wzw6RGwRra39Lgf88bvC/9+4qLMM6GsIOSRQHk7Gye2j
ujg2uhxJVY4ibvuiBd9S4vqEz5XOmBzm26BbgobkOWQFUbezAr7IYsuB0UVVPSwq
Psjiw260af6Fm4P4M3rngOM3meDRvjYMv78vOreyFKXGESF5iKWmyebHGgA2NnrB
nF2QEmvSAK4BziPn/+cDjPNmUBBBkf0ODv0WgnkzYKkcFf//RF0aT/isB6miGg91
h9trBCG76JXPNgHXNKBRLFGuC5VKu2zR48UFKNY0Mt148nkXNXjv+lzFXOZyBcaJ
9JW4PiKaQQksgm+e6pl0rh7BC6QNcqVg5R6aHzQ9CKSsRu6dQgj4Yd95/Af1jpbI
lyemTfT6i3vYmevbmXH7xWGCBqIt8GO3DCopZkw2T1PYrqSfo/6gQ4dhWEnR1PCr
u0n3tFrs8q37G8r6qnq8BSNA/uQIHUjB9w0dJr7G8Pp1EnZjjmVgFnvPZP7TH2NH
RPETMIxen3ore+FkT5zTMyPrp/Zje0xPvlVOBdDkjKcEzWk/Wy4Z8sKbgr49nySI
LYplh9AKDH5Rt2Hu/lbo7nRxx8SadoSOT/YdZkAQxY4KPBuZnv6++MSK1uUrdmXE
0okwYdRXkic2sjxMGg7v7pHOksrOmWkac8If3EuUqjoltdSZVPzHAxvbW0moIuLi
m1Dzg/zHQ+ysAaH49d78iVjlzaO+KBismv+z5jb/in8vbJJcBUojLpJjVgy/KS21
pRVGPrbzU73DV5oarUDTODgynZCbUB6VgkchsG9K4xN2pcmg4JFIW0hi0vLyV9uB
sYtGzJrT5lGeDjCknoO/srQ86Nua3RMUygSfYs3EKu0Xu405olrMRNdG3kyYCwYl
a4akBX3AGbUgKO6HoOL1Jlb66dsgf/AXu82FABXcmJe6PcUCcgW062wpeoWdpcdK
Ij9fu5/VaRaqedzqTdNp82VhrI/4X4RiR06HA26cmdHHh7krlcgpD8qgzxK7EwQj
v0+V1cJipslWm3OD7vAFbAtsBbiSU0R9Kzty0SfCw03j2/MXW2PUykfajZK7VjKe
prnE78R8s/k7TnEeLtGIJw==
`protect END_PROTECTED
