`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WN351b5a33MmHTGaBSP8vbIRbriwonKzI3hLd8gZcvtGHCbI/8hXSFhdMCRFsQaU
RKWIf1oraLsGXJQEOy4v7gyx7d0lmXqhx/T6bCNOnKEw0OKxhxtjThqflQt1e3zw
vllLvCVZ0adZAqobkSz5cm3O33bWOCSI2SvMIw3VeV08QCOdTBkPpwO0FX8CBgTe
jl39dFTlXXGID6cCDytVMej5Xwa8wSGkkIa7wIsZh5NeHmW+KNxU1g7LOPI5gzAt
j3330gV5sNTMMGcgjdc6kceJuktJfLomaS/tSDctaQT3KT5U30fXzs7OHiGHGfbL
IvnfEPtcfJHXV12+vRTCJRH1G2shTtamyoZOLckCwaB3CRuwvVnamYA2NM8MUN5P
eOkuzvAuMsp2I/vYZYApEf+xdOipDGrWYnFLhUGSmQf+01sgD0dwAY2Phk5sUm0E
sKk0ATKxYjlkKPSqr/OQkCai5e0ahWMsajNogA1eMtAyBwPokurMKqG2q/cLSp4q
FXUaA/NH7pzqgqS2c+BXqYLX4fW5BZIxDhrNHtboVr7EpjnzB0I8oae5kpWD/eyp
k97iSgjW+gtZJG1pqkyT/ifMljA2+QsQJ/B0YJWYYo3DYSH5OIPrY65hJtvNwsfj
w2hQtbBsHJhhxWLS5YCCq/fw1mTUbqQ4ND+VqaYYN+ysARtp9sj9h+WQnpepG2GC
O5KIqjlhEJOVMaCa/5wQwYqdiI71kVJOmCUPVOxMJlSdz0o/f9Gr88hWZh2FBVJa
sAVnY052bRc/QCUdYaWDPT12ziPNd+rkTG868CjkDgywNJmFPjpEbX6KiOC4NPPo
6kTSW6b4iUbHtW5vsDqJAFp76K9HpZPA4QdPQYjhOGxqpOUsBIgJDeEdLhaOeMC6
ihEJuof0ix0/VrgfDACMjf3Bc5pXEqr05Z8/9FCDnUn0+5wC7CF01VbvZVX50/Fb
Ux2U98Uh1n3vC+p7Q2ZVk4dYmad6rUwzEulvsDAfIyXibskHWSgvO4dC3GOvBu80
fUtY1UYqZ8icQu/dNcRFPpcfgzEcLZMAG4GDIpRLzCGkbcfNp8HIRvd7KSrxE1Fz
z781Pi9IwiY1t8ORJqoYvg0xgI8iemjfsDxukWj9iHs=
`protect END_PROTECTED
