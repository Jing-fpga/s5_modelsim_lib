`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w1ikahRQf4WOvi4bTLuY8l0loytTWWijtG8JvzWykmBnDgd+S+fg7swRfxDVvGcY
gLrcgz5T1Yt9RiyVsS+5NunxwuKvQG0KCY5FGyJ3q1FZC5A0ndj9t6iloLDUrFqH
3oOjCUSrxoA0esNeDJ4y2BRfmf0j2we9ZRA+OsMosJbJA9wvhpTJVeU9jUddEzUx
DfBtQldTzSbSsfmcIsFh2cLTHmh2wKSxUTpzdvSmHAs5CrUgJjm0I9lKBIRHV6ZH
VOlsrGF+YLhYtWByCJg3wzgIMZX2J6q2mW5wNova+zvyb2KxbS8ACVuXZUHbc0hW
fjQS4N9I+KLO6d1/6rwgcw4BdSQ+1HaSOuHto3NIguP2IRRmiQrYuA1YDsCoZ7oK
vvtAt+8B+or8FzfFeLNL1G7g1KGIzC3uakR92FDGyYmXIpiUohxUeEZSXOx3iOx+
7a15oKfF/w75VKD7d/LGq8hL4Vyfd4kDdbF9ou2vNKtCtNM6x/Dt1NdMjMG8xGWy
P7X9aYLTK4SwnVMWZl0IHX6lz7133UUWjR+WACjZ7PGa2Q96GoiSWAnpE6fWAll0
IXFU5ZUjZjv8oKvkKpbrnF+osj/lxD525Ia4q3J8eNQBcby/8kxFs8JeII5I6Giy
euVvyVdSXtrdXGnu9Ov22ESi6t3a8nTYXQ6FG2L2mujHipLcXdSvB4xrFWiO25m8
dXyEou/gEubyGwffyPXWMQCnsEp4dfR12HS3Z1e+f6w5QxmSv6ma2dnb5tPsRv6S
NfB+/rHdRepZqR0SOvDDPv/VEuxeFZ+UmnGOkunZ8XG9Ju1vVhWGu6/c0U3Z0M+3
2vA2jz0G/z0r1j9MVjnKjPSLsh0iFVvUHMrvl1369JkJdgLv9huB9x1PhFVsIh5i
HephB15dS2Qxt5T4ClYZEw4k99pNfPMEOOML+kS0YBMeyav9v3SoLHETkLhXrd7d
Re9+KsZNfhrhhaa7u/V3VD9DvT+AFk8Da2vckutIv9i+q8isyNx3pSYe6oUZr6dx
Q06+ZPGfgRWjBOkMk1LKiIL4j7IWYHW5NlVzKwzWPafOnt6So5xmAJ9HIL8zxC7m
QR6mBtglLu2rjNISdrcrdt1RQ3RKNdQCYEZBiFvIkfF1R0qUC+K/uMLYXig4oenl
UfKA4SpHs6fP8izlHd5VYbigJ+UN5f/9XtpLWAv0mp2OAidm3ALziPaOu5hm4rQe
rKKlpTp9hek5+ynusVjL63oTKJie7jKJRBfri+kd/jq/u7f03lzeoS70CdkVDPSh
E59QpJzCIKTsenqogjI2jl6caXhSCEaY/TuBmO2sbQhk3Omrhlc/9vZXhPOMYHGK
97s5jrJxobx5VXmVOwB1vIaO48aqvk+6Doz9UuNS/i+DhQD/TpkVfdfsymBPs2OE
uYEvSCqtX/TthjTk1OitV9+bPZ5d01A1amqZfzLADcfGbu/dfWoBIVvk4r/3JQw5
9za95o9Wb60J/RQHXkhxWLmaZSJo1n3ZnwYucAMMIjrYUCIHPWHyzWwhtyo0j23m
NiryiBC/yOSJtMcckZZl9uGKqDn9IKq7Gz6ln/zyK8QXScOIGHIbm5zh4htH0co+
lOUNI5nxYhGN6QDLIcsPdKZx1Lkdz8cuqWNtnci5vTuklhXPd7ma79jNmDGJe1sh
iP85O5pOb4HU6kKJn+c3Z4YyJzuI9TWZKI4m1BX1iuyUhWbGx1L2YJIrmK7tqVSu
G+gKcRZMROXuAf17SZgxkPGugTzSqfG+3wiC8xRnQ7Pns5pFHuKuu14IRzvQcn9K
+RpnrGIagVLy+s2G7J+CKmkFhvQcKh6O7/YvgtiF4INx2/nZFFCvNc07LEZh9Fg1
AVoRVZleuRH4C1gZqOqLwGnUURSYAt1AQkcoYE3YfxZnx4Slkj/o87gL3WM00X6N
urtULjopRqxBLhJeazBUyyoCzFnJ6fbqKFYJJLnKdJ/F3cRRWLChTSGtA+ysFDKg
Z5mxybYIniPKJkAd5AR1/k5cDWgio39H48agZdL7juq1LO+vRRYS633IHXiYwl6z
dW58tPp84cbsAGm55IVUVK4GfRRGL/AL8yK47H381qTEu7M3JEUj9Ouj1/7gMzZu
bSuUQpxM1auowW4+LXvHCcQMyPAl/s7hTJ+78TPkH6FLJwqqmRh4G/bZTgIJuSLa
SOfiEtw3wN3Lb/Qepi7QK9tn+v1q8CSJPdlZsSoR9JMKywlpkSjyS4oY5CYtoIkl
2Li+ShtpwlK8eJneMMDb9y0m8lMu96ec08eNZcxmQiLKfZZM62mHW+m2cIZCFFY5
8hGp5djkusmjTcGgv3tQNeVzHz3luSuQJcRsHZYm2/fL5R0wB6qO2HlkkokhOmql
kPmsM5Nn5JyjKW/bg4cflBQc2jtgGk/R4fFOXiUbHMtqy5EBrEFtFj82g7uYO7LT
MPlymLRaGUF1S7//w+A3aNOcJwqsJC/1kV0yFeUBoGNt6nlp9f9R+Vz7aluJxNYY
Y5GiLPYIc1LgELVnqpLa+U2wq/sV6KW7cMGMzCaNeSIL/fIb7evVkriCTU6ouqmT
FULK3RkjqFaQHKQ68pYv4XjM3ocRNlFI//rhlS7YBiJKikFz8mdvbkMzNAQ/tQkc
ndZwED3ds/wx5OftTWUA9WoqHL2sKGQRSlmrYd2ociIXRsJJH/G++trJiq53TN/u
1GtcsqgV0mxw+B4czXt1n+brRNTNb+IfOJBdCU61hhSCD27YhX4kmNmR21nh8ihe
rgGDN7ipIG0aKX7T2gs3vvUqiQ4uMlgPnEcwz8eYUEbIvIImmdxS4fZBFf1g5kYU
wQ+uPk0vBuo4nofyrMqRIaBPAYjj49ZPcCNHquGXtUUPUF/U63sh52CconH83PgD
II305DacAMjPu/9UlwSnjCbZw2wh6YInMheQKl6JukdW1rsldm72HYhd+rb9Q/AQ
mKslHynOnrvMq9LNOQevjoJlYObwmDIQyDzuhlL016WWj5x8wNx+cf4YB3EEWdzk
+xT25xRSm7R6KVhmF4SSgt54rypmRNA91AzcftBTihIEI4M1MGtXBtNu8dkknVrV
dnQJ/amg8hPedXYcGb6bAJe7uGEXUb4Qmp/FWdAFYsOGTB42I1TprIKkiYIRKzfJ
Go0eH3R+ux673xXBrVOmsmV1+SOoWylVFKdOg5AwiXmkAIYZmTh/r007qL9CgALu
/ym8/OKqPqMRmhXoQVTrTXV97UJLr7ne/3LK9rZraTcUbN2QDMUO40ZC7pf75JRM
E9qWhfwmBNJ5OxTmha/vt5xZewSdNfXGsfPSQSdbAcB70SLCgJJ7/kqKyl/hOSAL
5TgV02UUMVfF8iIUHLHBSR6R5yroz4vJtPWDd9lEDoF8w6jr56Nyxrrsz+fZzyOG
mdUTWTWd+Y3blF2zCHhOQ0HLu1LugYapdukFam7PXi/gpAnWeIHodFWvKHZ97u8/
J1H+8Ef29vqI0wxI0ISeTB6bgXcWs0e3o3YiieSDiVS8Q6V9t3fxcdodCaBq6Gjj
r1ljALyue52wyPv9EMGlEflOP/n20KTxKJkpnYE5Jqeeu03jIG7uEYMGAMdEoa2P
oBd/YKKo4fToA6itPh99EQjESt0o6rrzgKrZgu859lzTmmOn/TFqhk45Thvn3pCI
UmpoPy+tjLuslA+SDGlRg891743LRdM29MaLQ9b9458ycP2D03gFBR3cyiOnpzUf
r7BkqLGkBxt3A319Fb0JziMw6qdBj2IfEUzXggDvXDmIXDqC7yAK/Uhpdam+C8qJ
EZtnvcltmvtjxZT7sYs96Or/+1Fju89QMZBU2D+gwvwU9Tsic412Wru2uIG55dsb
/wBIAdS+fcpvvSyaCIInnJTUzcd4fP7Tz7ETVzyHwBzIXjzF5tdxLVjIYNXWkRlj
20wpTq2cd1T6FfvYY5DxfafJ4MS4wOphx3FmqktrJQajgBgkgUyi8tuP45Y61Viv
o2Keml8UvnTaqODyoQpPKaJN4AMfHbIvQVsSh8imVV7y+lpzB0q+QIeYGvM+UDzx
AGIDttuyuwF6mBFqzRxyTKtiNcCktN34HALxBgT3kKHAgzklFzx2ktkafZgEwsxl
fk2NbIotw4u24aIF3rRrav+ndJLMizF+z7UZO59j80Lzll9NMxaHr4cI42G9a6q1
s9fS3Z13poJ0GRV3Vedeyw==
`protect END_PROTECTED
