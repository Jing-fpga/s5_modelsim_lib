`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XHpzxnLuHEo+noM5dIqFOaj2z0hOVi8T+stxJGbCgZ2i0QpoGZiDqp8VZUq1Wf1P
UiJYPkaG2M+6GHE4YuAfuiXr/O7/ItQPBgmrsHGsCp8g/VZXPgFBxqJl/vjSBrGM
B0Wvrz4O1R0cSYbID4hnuhkidHqntdC45J87lEKXpLmhEKK50ZCb235e7XxKX/s4
Iev0ckZd107s+MVPUUpFFgdvovdh6ErG8gNQFFR3VJltV/LlKMFBCpaT+q53oWx/
kjKPm/52U7AeI1IvLqvgG0l1asYjN13jwrOS1ZbfuRl8MpXqZefox8+haLtojY8x
ywyRbDbqywy+sLYZD0sa8PxyAOP5LXdnZchHv1zHTrhhcp6BychhPw11vZ76G9iS
`protect END_PROTECTED
