`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zQbGJjjpW8ZquOXTBZsw75ukAzWNwGPXQzxJx5vde3xTJAZVh3kT9f/5BEhsElti
mK5Rt09MIsBjSGzGFwtKYECNB1usmgTfhL9AZR5yVYQIFnsTSc4bBis1SOY5s9M9
0169IyG9MBuNKdmhSI/p771kN2Y2SGlSXIW1fzbOwbyRc4WlDK+M48y0H2xqaFtI
4v2K8JkzHboeF6lzaMNUACpSnur3EKGOWRBR9R0N3sDHp8b107PsmmrjfYncDP3x
8fkUnpgUIWuBAlSNplPZpyZNoZ1ya4H0jJ0exTE+lw9E6UDMP+/O7Nx5QreMbr1L
Tj3seW8U2Kxg8xBHRnH3KrWIoDV40F3/uluOKQ4xf9OYYQAn3awCNHaZzlGXGEz2
sEYsq41AGFWUI/bKSTJGlttEPj7V1l4yFAtxkvHsCycpxl4Fk4gf3GWlD07Max1F
XSlCiDyEzBqM9Xly+OXHs6p41pwDGJWdl/wM1uTGREjgVaCwEK1b0J9JNmuJrssF
CpKLcac/YCkO/mrsDAVEEQ==
`protect END_PROTECTED
