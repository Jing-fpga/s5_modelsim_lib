`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7EWtpd+AlO3Usa7OQs5neIIM2pyBcRVI29tmphiMjmb/59WEhMHBIeiuPa7gOnX0
YtxYQPxLCxao85+gfxYg5oKMqN72QRil5uImjnalWpLFXWS8cDkyE10mULonXC4r
vTrZkNTzMD41vyi+2p6uXpxCAm7m+R88GsNcd2GLsYdr4AXVxt5M5UXrf2AFSMEE
QU/oekT8xj5Rl0YDHmKqeWXEVdkMZmYFdS0jnfjk+2Ymf83/Br08ktVoBaZUBGGi
jcrQW+xebNybXXBkg1Xj1tWwGhk0D6NgsmzZ9b1XirBW5xpnO7dZsGkitFuU9ET6
ZorcoC2VVggGC97uEBA6zHIyAv4YAVVejy54816+KXsi4cRV83cUM5K/DAE+xPHD
Xv9d3aguvgZ42CvVJNg+KjZx0yYad2nzUMRwm6vMPItj6lC56QYn5CHiqneJELpc
zDTiNpYQ6Rm+9McMm/hU/t+ewXxIfBoMSyK1xlRGZpOoLIt7L8JhERtDnlalyFQx
qNpAgdUu9Q9oKjAPZzJwSqggVYFakhAK8iW75tzx9Cjl8mPFMCEA7BSBNYOP0tvP
oYvput0FLExCQMW36Xympek1/LPrqBKYGEl1Foiw5p6Dm9eDpWKU42uA6Ojg4Bx2
ZaqYU+ggQ2quvfGTWOy2TfpVrGrZZ7ZAhuFQrc5Jx6PKb4s/xLDkJ8lSgDtGKWJo
e3hpLhWEaSHjlyn8F5Fgr/MgfboVnCC7zhkrJJUhqVra/nNllnY4tbFT3sTSoGSL
obWcW9awP02uYOzDy3CB7A==
`protect END_PROTECTED
