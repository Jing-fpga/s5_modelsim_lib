`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y5On3dlnNdfKNw5+AB797+S3EsOIj/x8SvnZkmc5M9m4syv5fI4M2MjfWRBTeMra
zieRNERE2D+6S1m9RoP1IRDjAm4CXOk0KeUZygFE640mMMbJfl80TiyyPT3+fx7W
YDcu6vI3Hh4NodyzKpkJ5LE7Gtztzh+88Rjqlt0/Uv0dkcR1unMtqWHxjTmYuKFF
4krW1Et3CcocVZNrOKQG2LB6PaDS1m2r0Kf8aDYq8nOiG3w9etXjd8oVmwWxBfU0
XKjz/mupHJ8hA/VGjiZdMPAAlnNu9bofnpWnZDHuZ/0D3Cetj7jnY1fcttX24nnW
N70RZ9foq5PVRW7dcDq1JPQEUKSthlzJ4xS5Pefj76ZDbtEOk2yfgSJk/OnShy+W
Enj6zYVbyEfq02UdyhtSiyPt4fgWAFq/UQuVZ7LCFBdirn7SExQxD1XP5z5IL0xy
Y0nA0V84JYh94ldpKYPrhYtLH9iPHQg4uM8M2pDy/2lrJqw1F3A46WmY7dbczprr
XyWDsyBBESHkUeTtFpXwMId18X4mc10rYt9qcx1vVgb5T8jBNGkdN3tjk5p3lK87
z4Aluy8vKqfLsqGa2uqdeBO+bWRVm346NWV/ylRM2Ch3rIa2QjeRD1J5hP3A5YWD
Ju23iMnq0VyuPftmpzpXNppcek1iWwtLCigTEkTiPUS8obQxmtRyqrfMGBj07A7B
bvNdnHsRNtS+FJTlHMSSR1uq6EE4oXxMfzuMm6BFz7OvscTaH8+82ttTfGloMGpR
jPHN/6wEsD9sccRAcbPqd8MiG27QQzCwX8LV9oZV3dOI36+HwldQOLwvF69HeSKX
iCRV0ydstOIhxbs1Lqqtxuovqe300lnnkJJd9HCEZ3KdMAmQALLvAAWgnxPfaack
VVbt8gnCf8a7Cd4EO55AndPoAfv2b9Lh40Riddi3nLfRLhShXR226ORD/mOVUpBt
0KUCTLbFZKPYVQDa/jjSD9jAg0YxU1CjkxOjGo4W4Tv+nQJCB8d8FzkQsK8wby3G
3BH/ZSEf8RintCulgL9v0gQYBnlYThbI8b31uuX/LVR4Q2XYwc9+shXo2qHtc16O
1v5nki1y6gbwKoBYQNCS4Z9Xk8d049vbvaSj0eD4AxiPLZFJviXIZuaVaulkBCl8
+9eJLO40WHCq9uIcwtjwUKgmFbntXe8KFeOa36YBZFOvs6VrtEX/l2lLSDXAliiz
UB4pq+xCg/pJbkzaatzt5Bw2/N5ajhhPLkEoSSDBHw4B3cvZwvTScSuIEH/Kk2cf
pasl+z4YiXd8fUdqafN3JT2xOtEOJl6v41a7ZZEabx/KR4KNs55qynYRQchQwru+
cF7r/ybfGdEhik01hA/TiQvZ6RpNhmS7Od2Pcka/WpE8w/HQaQGGqIJqA9YzqeTN
CqqSUDu7Lf5pgLOclM0eMkCfbqgMP+5fC1kngvjnk6o4trBQSyvMffg0J2kzAT6y
djKZgP6vz3aS5aa0C4NJfoJ4Or/OUW04XDWHJCUAyQje+OcTng31G6CNKqt9azVz
1ElD9asrTjRTVd5zxRfSkt15/DD7q/cdXkx6qYHUE2WsmPQbIbfPZawpe8Vz0Iaz
bSRt8BiO7JzveOLKH10FKu+CRhFKIwWFKO4ccRmMFTA5CQE+KIh02Y2YhHDw9uRJ
YJf5OKzUP97Zm2bP0Gf5rDsPybmzE1QXIK4eWjQb7KZG+nSBBCq2/LFsXNwI54WA
lHvBwLRYHbKXK8AjXbAy6sb302G5oPZKksc42UStX+bEJtoKUx6TIRezyrDjkhx4
6kKGz5hNFBixWj6qpX0YLxKgwiXOYipmO0ebWuZVWVjjJqTpYZv+iKvgZAldjfzb
+ASLnuL3ECCp+SBBBLFmRKXUaX9bv5qY0mzj9G4pyen2It3vRy4GQzhtL/t5Jdf9
3Qo86Dk8VkZ1EnlD0jXoeWwckk2YSyXslm8FXgGrky3zdVkWU9mBWeKS193/YdYd
91d7jQDzBiAq16pX1XwZjqEpIqPtN0JbCAcIv+oeiwDe3ZJ15xNS2yYah/uofa4z
vvgbKA0yQfS9LlRNNsZQKx6Ml69Xo+PyQfCe5Sln+blrYsyh+yql8w/fYAgt3baC
I6HiTfSDa532nO2IzrQmf3A8N8i0p41YmWTFt5uDEApYE0eYvHnHEDCN2Gk6dqMs
wVepzezGSTEfDQXla7YYsiGP/edr8q9eg2qdQE3UG1hCeRIPLgplyVKyS9T6Yk2C
vjS8YwPgxeO4W7+grsvp4rqfCbcwABF9fdyIO3lF1tTKmfdtyxY8H/tsk7aN2vSm
ZemTAfV/RWDYmMMNxS2m2TS9msnG3kzODOVWxzVppXHWgv0W+v4wFmWYqkf1YcCu
EhWHCo1FhbJvLaN42+J0UWshd/cUI+GklzgtgnquWbPriFYBLMHTnuLmVKJRdRTv
xIKHYF5RQli0V4p+mXDr5ne4srTNpiBTI9kRYhew8jtg8HIytY3LJiG/jHsws9L0
zrrI3x7VzQMcVDs+o3wohgPsLBSA/SYH0dDNW490AjtXE398Rvu4AUE/dApc7DEs
4oqfzMrmSww24bL0rDesRX1B3ECOSRa1Ebera1eHuYi3qTl7o4rOPWt8+xaZSlJb
fN9d088rF34zhjh0/ZShykEnL9zNOG7VFGDobPCPzkUzJWRFQ5LU/QyMhLEJ18A7
xFCuhGiwKzjG4rTpj9aAaaLI+9WHDtUvXyJ+/egyTbBTm02oro/xRaKlZGGdoJZ1
zGOwnU+c5UqI+6vWAMJ8tUjQoikbdHFsje9PcbSaIrArDKyAWbqAib7kSMsjCaju
exaBlgVpSKGpD1N9D2f2Jw+obstExb2OLr2sVymdlcuczWTm3BCtI0Wa8iWQ+ypQ
bs+rUHVPp6pzGIY8GrY+M784lsg1JD7oNGdo7xpGanJm+9wx/vYtg7PofdAQNvqx
DOctkz89i5KyxpdCeHNPxRqUa253i1nAZEN+aTt8ZwBxbtiZWTUqtWCzTsVxPphF
BH1zxiqBvbgvActWkkV+Wc21t2TLeBb80E4XEEwwCTpWn60kVw6zn/9CC2/oKhwm
GSN2URNqolebvz3L7Ifj2orzFeZ8POlp9vIAhxvPU8BZwUju219tSo+rzirlIGmX
jNRnfhIAarnF1lwY4azk3ttK1P/MbeQDXOLZ83MjUJyU2WXllzLojUliSVb6I3ro
5DVX7f5LaLoPeEPabKfE0+T4SbosanZv8OilNv9AdWiUAjO57oiX7nFfOFMVx9Nl
XcgZbbU9vjRljd7ntZGxqDqgmA2Rmex973r99RnrvrgUakxcs4TIw0bsHL10Aks2
cdHFerbJNCW7fTuqLrwlgm2ifqPlNgwHUELqs5S1g9hjf68+uX6t0K3hv0C/MNWQ
BAjYGxUAdLfWL+TkSyQEjQZqge2vgB5tRgxbuqQ6OQwAOdLFcyST1o3wk0YTsevv
sq5i6xkrkhURw6xj414u3zzhCHflonVXl9o7OChKeuiRm5bhqdU6XqsJlMUBUpCG
vEZXDIbQZV+/RLlkpRu3jRdi+bHPm2VOyrvemtXmkYb8lZ0z7j8VrLLf0mrQgtAK
o3lZ+CyPHFY2XUQ+UKyCmqbcr9vSwBcSQCj8eFSUjnSCcQUkFA6kEMifQJ3BqT5v
UcTPHwWHvuGZtLrT9K1E5FqNSqy4g69W2BXKY2qhcRQ993LTVmKc0Zz+tqblGjBE
Wl6QRSyevyV1nXgF8Jy0tkXDVQiWqolYQCZjoWTWH0m46Bb6yIHCb/+pVfEm3FVw
UfS9R/5t2KxgA/T9lnA1zmFPfgAsQWCr9lSmkJIQ6pLecK+9Z4bfSbC7T1wu0ftJ
hAj83+dVPGVcYuaJftemP5tyrmCwohse3f6//iqMaySj7YN7Q2RlPXDtOfgRAC2y
Z/zunPnwWimDO2vW4WBaJDUIqDptPQ2xrybdnswtb96IsRV5zynetc7k3oF2jU6L
qa4zz7qJ/xLSyI26GtGPM0oymHSJRlZg6izl0tUwfAncUqneCALUOP7VOebgDVDU
gfGWowR+9tamBEGwunv5T9dlj0P50Z95r2NQGM1ydCg2Ui1DMk21oZdtxd9+zVuf
R71u8pcyV2PJWAHcC5XWz8PyozkPG2UN7lH9f2RN7i1oet0/Uz/DZNVn5U8hpU4H
u3qIOpvZB++0VB5mf9mDXlGDxJy9m+Lu2KJ7mn5HnMBzNQ9unFsnBv268sbPg8w1
2euT35EdGcQObV+UTdBiuI2LcBKkLllNrAH6Pl2BAdke62x4YcKI3kljbsL6FDwD
2UI4GeEq8P2SShlEUbSJsjG2tnebM6godVedK7wVTnFpyxIRtNjN48/fzCHYJdus
UQTOHFydmsy6ew2DP4eB97UeJ6qU/9TrAPT31z+lalhJQ3qHKD3L8AJLpCD7pFx3
TdKYAT8Sjm26aGVQLIre6aH2MieO1yRAfzO4JGzmXT/7UeqFxd7IEK2kF+7Uudqh
v7/BPN8hdKADrcC7FwsyLZtOoo9nvfw+mWWDxorV23PF2/LGEhk1abAMG3E6fnuq
Nge9X5mGnHo+JCFw/obGPF9a/Jm+P1xXl2InF9hPCAEFHcau7uZ3dKENGVAGqrGq
p3Oyvo/XTtwXKWf4yymRA7GjGOGtIhlxa52STWxNQJWjh9DFyKgTTJRb7F5C3i7T
KHL5FjNDvrZmgfRnELxM6DEBg98avggxPFxWyzhAEfuDzOfpnegbIDDf3CiP8Uim
iGYjoZdCYbLOfhb5Yhm7ehlBz3bAhz9L9I8CfnhpAyWtFfY1gVR6HhlQO2RCVLrM
d8ccUQjw1CAK/jWv6ICf/5qUfjosjU44vO2GCskGpSqtxI8Lkg4jXoLeocvhsVl/
48FBIRzg5bPiRiUxbTdwvuE9vOcEgk3MIySJIojo8GQkbj/7DimrgaSnv7eWZ5t/
1F8QoYIqYKLmCHGE0pOdX62K1Gd2b6B9xUjjCETiScnSEtXkU784JJbXMS3396Mx
C3dcC8qOkviNo48Qn9GAbM3BeMR84fbnE72SlMP7k2MsQmRuQRaPE0mDzrt0LasQ
SgTJW5I30qKTYCrCUT628v4wg4FgTdyEKvHHYjjIsR8xRUG2MUBKsDBdbuPOaj+M
34sv6p1WGL2rL/DVGMCNZ7vHJUfSJ4IRtmgSTDBTXggCWCFNbjPzOHqfI0ZB0Rla
LhMnQAkNqRY9Mn/XCQS1PSoRhIt4V3XrP4blmkVJObjZ32I9thA5SLNXYxQqtPhC
/vK/AIWON0OClq2LX+w5u86rjzK2Wvtks04BaFcvwDA/8ZOeHpAmdqQUZDe0W7HW
0AVA+8Nh/cR9J54PjRo65VcQMHPHUKXHgHkmZmlRqMe4WGvZJAgFuVNHpBmRk1m+
kEGxJD5xduYg5UK2KHJq1HvtXuzfWmyGnrSfnF7goDDAn+6I32laKJM5FtTAEK3l
grE4ixMEMXa8JWmXeIOVjS4smShe/mySefWzymTkRzyLEJN84jp5ovjfg3/9AKQb
FBMPXFlkTFPLLcRgKIAAA4bnxxIfWSYA/kqFuNnp/ge5h51SWJGgdR7xTAsJW7DO
Fdoj0IZCK2OEjXCdobittMWdbnygjLjJ6RrBnHivYiykd6CEbtoRnOIAAf35ZVF/
VQGegl/wjPUoxdo1xvQyiqyN/UcodQu+6zaZUFLSiBuMhxXN2y4nSi34nEIYMgTr
M+1Y8ASI79qQmcx+rynYMQcQLl6PShpyIk/Li20OPMnRM0A5wyCUXjHe3z8og7gY
f0Xb7tNgv3gJwoFzibZj8XREo66hYCPjeom1+UiCxq9a1k63Kt1PDGmwEsZyJi6s
xL7A56KpQugtn49vxBKRfUEUmuAgNmbc4X7S88J80wEe9i+Ot2rucDitihKVCBmu
ug9lvfKnlnU0wYofD4JvnIEnlwTCX4jPOKhs8TmMHz8ehNXTeZGb+EqiEfZNqIpN
7dlqwXFRK4QKAaA6Ta7C2WO/PBoGTAV/lT1j+T/nCZwTE6qypUMqXVURt+PaHQCe
ki3N2v2RAPrOYWx0jTAeDm1Kl5NSfx1DqO5DhJ5RTe9hAeRvbhYd7XBj9Yg8N0MB
xUJp/zHpmy4K5hDD+2Eyg8hXDoG8/iAleaRDAMklLvdhzqbvpp5ObQISTyDdsz9o
vuUB4BN+8kQ9ap55IcVWREZ+eai/w1V0XOpkpnvLz22VFAtyGYR0MX+BIrS1ZDOO
O/B2XuCPDSoEt4sn9BkzRzc+3GX5sEKXlSPJ4Mqc6AJnDSO6g7MQfbUwHO296s7U
3K6lvpQxTmzk8QVvye5et5tlGBb3j/giutbLCz95nuCTt3df8/kDIzgK6mAb1Q0d
UPbIa9qfZxmjEPqmUe3+8/42Km2fqa5rw/GqHT2jDruWxDOfhrbb4KtJRfLm3CV6
N4zQixBJCmmlEOm/n+2eDyOXhdMfwABWmH0ItAW2EBCogb2Opsh7LeWl97di06+N
VZWENx/WsuTFPe59uMUY5awvp2D8LNgR+f3ZEP3ZiuFWPUuCaJfG6lxhiEyTaYBj
ZZTKU5lO93au/D3y5cC9lPXihD8VnubQkoOQqXfnS086gcJMTwI/ebLrTIoLXqlT
PSCQP1DYwLsK5g54sU9713Qb0T83kYACctHd6/Hb+g2y+0NybtknmtrVxQEKW449
1ae7Butb1ylM4X7NbAGwXCWWVARwdvt8urZpLOmNJRpku6eLTOPzmDQIDctNwkJZ
ebYY/V5Te0xBZ++9bAi0qtl90Ql5v+Vp5mmncUoZtOnripB4NxTsFmDzKBokLw2S
0Mx+UOEd+lONSzRB4tY58QmxdbuSboauwASYWzrxeoh9XeOavRrhhhIHEcnHHJzB
MZtPZoMQZ4aT4GkpPaKvAku5dfZnzxXyKR6xvKs4UI0yNnIhRzLzxb5XLalhyUZZ
5n9cAcgcbwuDlnl2/0VXTx1UiEHvpj34ajfzT5J9/o7PF0x5GiG75SK3BI8QbRne
QQslXEpybA+t5Q3TmcuqcfuaJNjgE0cKfJLqa9jQrKSgmgoozxuC4A5C3TvuSnck
QTLfzJr7loixQC23TqsEnVIwYYITG6PM3izIFJNr1HN945o6yOVGy3XpjOfAr3rv
W1lSemzdLGqdL9H6DvmcTEAWdPItqexB0AZfcuFmPoSFTYnpMuiXL4GrllaFeQ5t
sRQ4YQtmwCLwWXnlzu7gva5CWpb/BSZxA6+ShhtNztbi/bst78YIhhG99zVPuEVi
4x8EklYCqvJEop1/O8PgoaFT8/IeMTQnnYcV7VWYweJP7vma729ZS8cQLT4xwROI
FqJP9dJDii8xDVunfVg7M9sV3i8IWWrpgQyeONA50racicAxfOfyP+Zx7h3dyC15
aI+1p+Xzf4oGNpmq7MHwrrHc/B27XCD8svVcTHQA6zWE1bIbFQF7uS4GimwTaMT8
KZKy4vugArXppb2yqaYthyE+LJa0lsHY23L3Dl9MBj/1AOZ68SxX5RdR8tw5Ygdf
Vz8KZ0BxKnKsg0AQGqxOciZamss+t9h9hhcNkeKZ3htEMAXvdc1J8uDh/ZsTEZFV
lDk7cb2zR2WMbvx32LhpOgDtcVOpgvaeL5OXw7yEYrtFwwXMB5cnCXPpZtvA8cwR
hiAbpHW6xRBqtEIENKOA42lFdS6e9BvKydnYYcPciCzjyNNJEXHmI8GqR/4HfRPl
Ie2XGVVRu02qpuMe1CInQGnfJWJdLc2hwCcjmB1CZAH3IgHatcC4o9vgHHlaBMFC
9NEsBZbi4QFFE0jPBMVOcoHC95FjeHBdJeImnb2KBqYoEMUZkEPGNdL8Ia22ce3E
a5xSowZcKxylXz2QgV1fa5eF0DGkv4jQewoHRKyrxqImYUQ9S/Gz2RNFLfr3Gcv7
pQNSte8p9t8DOb34ZlF5CCFJcKNcqwDL9oMY6tmx2Q+fvmwUc6hUzeb7FO3YCXc1
OOkR3cn4F40AvsQdJLMIIHsr0W3xjUiGDvikzgBx81lY597u6rrhp4ETwXdnD3/H
w81mS23nEXpmgE+vbi7D20MKCWytaZd9ZfJEZ8GlYo18N+rmQ+QimbM8Skwh+iem
zDODOkJVD1p9GN9YZM9sXrldOvcZpvkQeJwKr+RZHUdP3Jw+tBIdA6s6hS58VDPW
knJgIZPIHyHMLUQWybOzJtiMycdbZGY2Grl1amSww+6bw7bON1AuCOsR6a6FHADO
TaJwQdACHgaM3+2NhADNtEKi0xC7VOcfxTRt2V1hvGUcdLCekDVqezkVIjBe0J7o
OwBcR1dluBp7Cc4RPf4Pl8GUgG4ZEEbvspKnqEX4QTcx4C3xOXds+EPE7mBLiqmC
qC4pNjQLTa4rnRrPe1Za1yCr4cqEWg57Ghtr4WlneCeXvrNsCo0BG86ktbE+s9OK
mEdH8rsj7NMngRQPUrvBB3i731ubbMgBdQbG8gQVMErqCiLMfN4TDB6H94BHWixO
Mjg9EsMaHkRHcJCaPpJgXX3/xBeZKAdTsVDFCx5560NXg7xkiUFirYmoH/r59p9Z
qGEbMAzc65xDecwOJhZvvZ3iNd1BKrYxCfDWMg6WEzMakiqGLyP22QSyTFedyZcG
QhsPNMS5z2Mm+Xgn1lw1ijHw3qacuO20k8PKG3xhmKjqI7UEI29K/h7BL/pUZmn0
kEjwMmiT8f35tjvwaxoU9nOmV16bzdEHs2LPAtHYH7YWxd2tyDvX+7j71I/1d84m
leJf84dCkc2PtyaEjzRkRTuxrtL1Pm9MufhammOBkxvtZ5ukGMmuE31PUSfA4241
fcp5EgQdZm8bIZ7Q7g2H5VVfGKaFGfxKuuuojOh5blK/Z+Cd5gBEdLwVffG8TqDT
gTgxftgEM8DzzNyaytYBgyWcpG/ZyNV8fngUeLjvBV8w2icECd96dTBGIsbRC+5j
jXo3tOqyLso/Vv6jUU6K5Mijul83r28OCWxxhVAe9bPnb9OxEL8yGd862W2E22V+
CsOcQbO7J+fCKKVhxI/PnDdS0unAZlAsjMJsNznffJ1y1kHjdlPmjZCCfJbDR55t
6KKqroNO4NsQUlBHT4GBcwhD+QnqgdFC/XlKyBHVo8/b7NGHxq/Y2XPPai+Bm35X
7OsVgVC9YgJJnO3TXZosPXfrXqi9E+CakNeuCCGsiW1kuW2YmvWcOtBz4orDzd2F
Z7CasQpW1bufpk8Nxfk896AHLks9rF02J5XMN5l7FQz7XNRTb1/WrsWlhrgc/C5m
qPhYfsAoB4klP+ZLiFEwt5CC9bc9tuFp+T72vDPu4tSPzy0ylTz7T4QWcaULI1Tt
pnPdbfdtk4M8LC1lwcS2B7mim0O8tIE+7/sVI32WQx4brOBROKnHwd4p5Psvvkhh
hQq1lwxmGG3DtGG9ykANefTb52H/36RuG8RKwH6xhLdXvtad2FVyfo6Aq4pArT36
83IOAaL75XK0XSOs+oIyO29jKrC765zE4nECg36LR6K2gjr2GUT26Gj1RMzycqGO
JW2uRqIWRwi+A5WplaCysrp+LTEQAzeDUayHyw71MEBd9zgv5YlLYd76FUrcA1hL
dOIgsi3xXJb1gziDWo20Pr9nJdg6bzCiTCxDunmJs1vMRXeymNp6hLyva6P19pR9
lWzEG2lVKT6NysmiHqJcySMZszSMR8UgPw7M2XdRIyHax3KhzX03vNqfFwn2hUM7
L9hix88nEVLOHf6iX+/ghnPqTfshlyajcxF09PsT/ebXJU00r3lsjcmnNHYyp+hT
pURIGO4Qh0fMOvf91REhpIIImrngrTnpPF9XmdW6VB1NLpwvRJEBgGG89ofUq6RH
186ubz5MwxYUUXQqJYEktoTu272ZwfgcfYJZ3Nk6I2o/XglF3GcbwZbBh8tcNx3a
Wr6huK5F6+ZkLFVwo2brQhmxpzSw3IjeR7ZjFrqfHPV5bBnsLSMTxOMIuKyxeegv
pFrTsgK0QvDAgexCAQ96vFRt3/UPzBcdFpSW1n99vO3eMfQLGjkjNvOttMJCmamF
6MbU3j/agpvEILrose8mUo3dwHMHUQcBFzh9k9OJoL8vYKW5OTzoo4QezrL5fsxx
hJ+bmWr5XdXlaBcEbEJAh4EXvPLfT+2q5v6uajPQIjAJtzLv4jR+84I2X6lenJPj
CHsopyC1gJxu7bUwiUXwKEyQjRPG8SHc3FmiseYv1lenug8xHxsKEZP5xUjUmVim
vBLEJx2zqEB/MPg8XYxyecq3zGKmY9TuNUHtDTkMZmiR/lj7cIJtOARdVlbqnLBs
ZvbQNaYcy9cqzAlBGheZwMmQGpMthBlBU9pmn74KA2+9kC+TMgBiVXz31H1GU8Nq
6h01AalXrr1AGF505tgBJjcA1PSTFByfHoPVo1pXlUFzzGCDcBxxnekOrT+vHQiB
RKUueD5xwGbR4dOZV/7G35WHorjfm1whwC5EcSqZqmJZm+A18K+IiEVH7mpZl7g1
rz+00i5OKB8gCn2oA5x2wANKyCO0NjcTHgq59rzYQtJUTDup/xs32KDjF8cxJgFT
UEo2Itnwkk6ow5Ei0qps5CYsLHzinvXWWCAAOmvBdLsinuwCVdxWWeZzduBumEfp
7v+qEcXvoRcIzcOeqsxq7oYl7gIduppUHdBcqMzK3I9R+ERC9lK4o97Ob2Y0F33E
GTLwg3y0gj8CcUA4YG57zpgGJtyMCulOamKev9N57yuuj9tdId9kn+sginAbDoZ5
jSsxnYeu/26aok6FQSn+/jHabKF2NjsvjeTpn+n47zHKqfnlic0oAkwr/ATKZESw
/mgbRf2L9usHx40YOmgk26CxKJMqmEWchtcki4WZrmUOo0wxkzL5/yL3X38o08H4
5oP44CwDkdl6MTVyHHeIHuCsFbwo6fp5kcozsqu9ddYPFAvSmd0/dhac9ZBPghRa
TWMUZGz087G8XffGlwbjdJcH8kL0kVaDZVYtP1sEEF+ic3GnXkdhlmibBef5xPbl
O1LzJx4j1vEIDFwh9+dSEVAn5khP32wYKyt+t5T+wooq4MRab0a6+hkkyEEP8FEW
cRzmlSSGPVL6i0l0C1MHBRQIbUnOQfZLY3xIErrf30FSwnCQFIctmYHPfnSUhKSe
9dHfAwL1yd3SAlX27dhipEdi09zRo6Fj+UC60lh2ANrYtrTB7Ge6I7M0jPL021aI
VfT5weeR8x835aswD4uSmtBNH+GY1DicpmW31a6u+rq0tVgC29KBm7A1kYdydX8h
vTM9Mk7wZKPsJhK+jFPvxPGonjGLM1bdUCFWaaIqtOPT3aJdrAzR4wzHlcwJk8y7
RbtWnSbjLFrwEgIFJkQpeofRJEH4JxFS9VERVJi9zrkKUVTiNYMxiZ9rNKIyxSqX
9tFGhUCTGzx+bobO9mmiFcYL4ftFRM/yJ8KM4fMjC09VHl2wxsBugk2MxWtEGU9R
g+Wp7V7u+LkWbeSaozdH4MCj8i9pVBaCtcU7mpA+hSQ9Nuukr/8AM7TZMwamPhao
IrR/oWLbYcmac9kjSObkGnoLfaEMnG4yWfSmOQTqs9r8/xAF8ysiPoSDGv6YSKfp
5AYKIrGuK5zDLJHmWtpK4gqd72qDIpd4xVpraHFM7fX6YC4XGpcNUw8iklBp0z5m
ag9rKH8KIdx0iliGOhqmkqrSqkvlrLTApO7qaRLL8WR8R2c014rwdI8F2tIzUaIk
icp7kSPBXHgdd6dsrd0W6Xa4k5zcW6RoO3GJ6LMCtsJa3kUaJJh231qRTi98kZ9O
xS07t413bdMKzlEo6JvegqaK6eUmG9s/aUXhS8zG1Dj1KX1u+Lvsh/l5Oa3wquAP
yhR+6BXHcRzwMqYQgUoKPmUXTzuQqWLNbN6FoFp9zwg1XNXQUTSMpfAJwDOvG8Je
oC2TyrAI+zvmTVMZuJ+mW3pcve+RA/vvp43mUoLaM8pHZQ4Gsysw2jsDPPmWODYn
Rmt4+w4eQUHgtiWBR3ZEzcQ7npNP2SBxuMOlXAjw+CIL1UNAfUwmSb0Yizk6xzR6
AijW07sMB2a5iR0HwneeORoJPursOZkjztErBKhK3+DMwDQaOQqvkx9V+BKENuiF
c2Y+t/WEczn9aBeWw0zZ2vHU3AkSMMRfZVYcv21jr6oyj16efH20pJYLd81BJzc6
PQ9ov7JYWUCPBDPTtOF+BOCq6ATJOiOM7xSNOFNt8Jou8QXI9rV38ejDuFJUWVOa
5wcLt4I1CSwX/gngEZxkT0zzxitEqwhvAmvqABVh4gD3XS+q2l/1qBQd89IG0m5B
S8ODl3CSeD/+dAyQ89IPTgXUTlGb3HgAF88ka6JXDsYpn2qGzhx0qqKDcotocZfU
a0JSbXwTkW78f32sEL+HSbbFIjh/cXLjfxAEL0jk598TortY/9r+5SYtGbsn5WPX
D8UrBlWkuk1rZ7p4nWamEVZRqC+4/mNLdeuBfv8p6NWE9YHlTSMt4fJTmFm7S2ZX
60oO4+H3np6sG0BeOQZ3xMRgcTXcWM6VT1zq4gyeOBneis2YH2m7PC9k99gRiFhu
rTvsPBNgaYGnrjZmRY55a9zcUrEWzVshrkHNkcW/0YZ3mMiVLBZnUOpuNASyd6g5
Z5SypQReeGXzHFiDpH2skDJg1XzkXj7fVoNoxFv9jMFbkGz/TtgdTm4d3robxyfx
Liu2v/p24tXH/LIUOGshbipYnrdEBqDalrVKr4XGtGVUmo1Npia0cYVO9pmNxGfl
5zhUeI1cfz816J+B8ZOtPZlKbHVa6mehA4tEUHC5MkveBHh4AKckwddI7KTKUYj5
c0d+hsOmEf/JOGafiy/lkVHb6yXJgfVStypr9U98VBfmmtknjeiaCkLFvEFnS1do
oYAZ8sX4i1ZiQkp2ohlS3L7APa6zjUJtWzRGj7MgcKhY49BfakZMWCGMFnaEmZcX
WLV4IBSMgowK3vzmQPBhODeXS+/OWWw2KBJh0a97n0NHrk0rMItQxEQiu+V25sEn
T/YRrGCZgEbNOScTcQjySGZ2JuYdUw84kclgqWPV5kbilmJ/z0JR1JPB2r9f8b4u
fN5X3vZjICOjqRLUTiRb5EzqRagbjrDDN/ahe02mdw4B295qee8cTM2CesMM4MRS
2uYUFO/Jb8MbroZ/4JwczNNCP0FcI4rukBkz7DCGo81hFttn3ZoAKE84JErxSaNm
MPmrQxSQ1ggUMnE3nkvYVbeSskxP1aYzwFwTMaR2fKzPI+lgc7ZNvjZHIaRfPacZ
jvKRcWDfl+q7U/MzQdUKHdF2BeRiIz7qiWGSiYjq8E5SqU1xRkyrP6D8hMPWHEwP
Tl4BZqjOa9HQFLKKAmvXwwzWBW62oSyNfTgFxnpoGHX18FD4wDcol3dqzSZZplZ8
ArOutEzQS6fv5tYiuKsOC+uMplNqamfslTDnZ8MbjYYksm7kRXHn31SmRSpnpRFE
dQeOJXL58vyE1u/sOC1Yg6coZOCQOCRxGwXSyZVMgAHGzSAZsybMBFkIvldMwpKO
bIiqhug5NJiYKy+snZBrzP+aZnlRkWJ50vkIJ8tjPCLZKZfrFk/Tg6AJiqANyzf7
YNv+o9sTKO81ZUSoxrWi7HdoXjp2b74Y794ouMMjihXwljt+9At932cioYvE/52O
t1ns7GgAeRENl/cT/H71nnZbUvKSxeMQvyLg8aNS8RUaS4X+dxTuvQF+XFp1qkwt
GZvUnWt56dugHfkHR5OQlEo9OMurzBYqBkKDlT0AggKDugzkTHMmzZyvxeTcnRHz
xSz7QmxQZCKH7lTh67/4PPGf73L/xgLy6d2RQ2Zid/DKA0sFIUmDWGyT8K12RfqO
8FS6GJ1h65Ijn/TGlshwSYqomwP7ujLTEC55080Xl+RkUECK/tVVzQCVydFUbNs2
7Zy16veo901FwlYIVpOMjpew9Y+1ABvYfjfHEehVchhGUq9rbGyTJAbHfzYI2hCJ
T+NJjSBcP0A0uugXdhJ6UJzuwh42b6npgCe1NnIQZxYbPF+Kd/MPZkWC9Yp5NGOk
IYsMBRKYxoaJ+61098LQRV22yeTEGxtGMPful/mi3z1qDDB8Cb/mkgiKk6sLtzs8
860ichHqPUHHfZ1dNHgFQ6oMGDGoULHhT++k7vv9YZ1gEXngi3LEuaRIxLze3n4a
4JR7RAitzJIQVSynOe381o9CnHG6TxfbQQgAujixYmcKAQZDYp1zr+1C74WB/ZmU
+HComn0Ke1yfE0ZYk6RgSQwDK0xvDHPkfIPp3nKL4YYu2+ZpHIG8UdIh/npoPgRX
3QjDuMRd7LR0hSEBFnxMFQ7FsfYhdeJkmFGaZtFIFBcG2S+bV7NV+yysTm0itKSE
f1gIuZQdJr1ZO3YmvgFqFv3ArVXlUILGGBREKurM+P8Ov78ut9AVVpJmyPtihfol
z2iSkVJaL1MhSZy4N+NwOKdwuWFDQbW73FbtNeLACUXHDDwstjM7L/WUNNevoGTs
f4aSzvXRj6jR49Q6DWOgqAGxMxQB+taMcbaTt+076E1dRO7kGM/spNO4Zwb1Ga8/
djSjm8G7ol8wqfTxtkQpO1bFbM2hGqgQ7BrJxplSRF+A/4KUrpkb56gvn4DvO/tH
hfxK4R8UuvVpo8vn4Xnay8uTw5HYgyJQbqoRy4JuDhKc4RcrSay5xm36xZQFhQbe
wy8fIouBkHW4ldBcB4TuGDi1f7kOtDtvj6x/VudPkxTAHZ4O1m3Wdgoi3IiXfafy
xLLpeWUaw5KK84PvblG6KOgVSPZ5jnQjI86qtxW8+4hse7/YzQ75eJzU2gyL1m4l
xIivbzXXbBgghi7qd8Jl5hkeO0+5tf2+O9+l3y7zYVsxIpQCdF8Xx9klVAs77CGp
nAtzDJEZnUlIf6A1L5RpyF6kz/y34fJTqE9yXM2KfVY/S1r6BL9T1ugFrTH+RKwY
UsOcNwK39gMwgl1qr+Rg/qaz2cH2p0cqUlLJtZfslSdZcV3EMInTHHOmd1OiGH1q
y2GhRflGFFGt4AtUZZGCMTZZH1W+VWXfss1nXDoB1wu73ztMcXTcOJ+5FkAKYLQh
mSR2NVOculZIggOVN4WM274m6qQjlH7EUB6ucctVHf4+sGjVIFGaYyDpcfvhkm1Z
1QQx+NrXygrWPvKvlydLgdZP6pBzP9sUWjt5zOCbYc34GFP0EcZ/RRGoV1BR5rwP
wWJJAEqoRYDCC4ORCt227UZohqFWi59YPcBgGyquQKkH1DfFulUPZkjRzUNaT7nF
U0/4V3DjhMpvA44Thxo/5S/kSFVBpq3YJpHXszeqNmiZybN4XKGafruQEF4ZozLk
lEKIzsKD37hM1Qk57ZywK5jNTfDmdgoio7LPYKjrD03KM1iyvZzzmOAOry6BVYit
SikQ4P+/d70nBHFj0eQGoDOU4JMfrlYnzXLXANf+9F7iSRbjMZUWwzVbT2ALcS/y
SrMw47z9oZGk+lVq8rWY1dxEJItbjVF5rRmZJIGAalFHius49yiR9QFIXU5ra+ZT
5oq3V2Ql38eaJEQDdGj55nEU/dOHfDb/u5r7+ajBAHJiEhs4BOrNAa5+H7l0PDOs
eabLfit13a6r7mVCppbDC+zRzJvpqdKZE7BHQAYRway3nb23q7sDl554rBkIm42j
/d9HkTS4RuyJl0RxqXbNslafY3SkJBp7d+Z8r7TdR2JAPxvXstTghU7F9GCzALpG
qdCFH+mqk3hSKnnsrn/DIu6MacpXHBX7nzaThr5zNs9JnVszCI3/hCn7veMaaQ70
Y//6uVl9cQoUPQJVdj79HYIhkY1r7RrofmZAwDCYlFVxKVyY4k71Gd8JHhhyJRiG
U85osUlNB+Tf8k3iE0Ma9mN/XWvJugZ49kIvC7rrW6xdOFa3NLOBH55uxRdLwzSL
v5CAzdEw7Gn9pYih92B0uMroHpmcxjFmdwJro01mKvuyVhUV9+U6KmkLmmyXDOsx
Emfh2Vao0lreqyKgBar7WqcajkUI43nimJu0Kba6SXOHcqL3rK7ou06EGe8dPMHw
nAMVCWCaWK2+A0dDp7TgTFzvk8eu8qG4QZFUOoD8NIiBBG8yBVuuZaE+RNg7GBsc
d7wQdmUyBMgGvUv3YW+cUdRWg6+INQVn/tIWIB7Y8D40nY7Mitad6VivsbhQugfs
QM1Z/srly0u9gSxnPOhVb5Sqc2a/HfGB6Rlcl99fSCKDin3Bsc/J8/1jBnt7qSBL
QZ/Kc7sZdx4eoBMRozoiptlQNXUaQB0SrBk+oX2ShF9z8r+zziJq/RlujWjfHKpz
kggES0ldiemqwugReeTho1J7gu5ky38T/a96AoAEYMixXeaw9cglH/l6aeyQSO8K
A9PAqUU36atB9j99wD/UUtZW7gMoHLfLnctIvxevzLE9WGil6G/0840XpB+5BLev
qB+mcSx6urFTx1s7XuS72Jqbv+a/lr+Kr4B3giJXKuDdpH1D18wHS4jmPwRFMW/4
Wh/7lpyqeTsikhEWPeQT3nM8yzZIKmrY99gA8aOWtvUmk6B8cTqsm7SawBEyfCPH
g75PTsRUmgUW8v9pxGrnPduB3kMPt8YsdMagiIahK7iSeAInbqySqLIQUSXWbG0E
butfghT2oq0dzg/BSueJS4RKIHdL8vuSoTawVi7KK6uhW69JGF6nrVgKKAzbxcKR
0XsSl1wbUQP32tvCgGzWI9flp0o2RM8cOURBTc7v309xtR7TPbTiJz8nV8D60DH9
BIGJXmI0xm4kLvwkXp1opzfCOznqENI9P1hkNZSPDdI+AyWWqlPOT5DY/dJQW3EX
xlXAlxw0FLJh+TvPhXV5roL8HpxS4HSfpoV3CHkrVGJBvK264B7W8x5H552y5Y7q
SneeRkQWqdgjsSFrEcZi7YV2y4VeG2rgUVzqhhSsvDJ+8It8jrle791nOEKRXoMH
Ro071py2YG7p95vbS1L8e9U9QsO2uvBgnts/X+ZuuRvk9c0qW1dved9u/uIcRY8l
p1hZfu9zViCT93yvRfztKy1Jlc1GdCpbyqpPmej92RetJ5JwenIqf4AZon/mCqdS
BD2SsBor3DEVYqYHWPvPbA4ZS9nCzgms8pn0kRG/mA3cs/1zdI5xabUCwCW+vWsC
jwYgzg186lq1j1/a+eV1JCn5l+kpbk7AunUiF7Iioi4+W9J/DXNs8QFiiWy4re1e
`protect END_PROTECTED
