`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Gk4WYtQY6A9g1MJxgbiBj4BVzn1+b/RrIQBMNHyoOXQeRH8bBbvg3C31Pm78uLu
rLErfOtK8gTf3Nhx8+1qtlDX4bz711AJtmlxy6LEEvccDMhclPjizxpJfYgEFTbN
+7zjqIcdysz0bi+wsU7cxeQ7bOOMJ8mjVb0pJBRHa3lgA+k4D/nD8EH5i4ouoqS5
0zhgdA3jr/ZEF6pC1aGHHq/IOhUGgTtlyvSYzE0iVDxW1N5dGxN71XW/foPILcf4
DE9u/sgwce2yDYJbTfhY2OUbSLIdnp+lCbhZzj+sIkIrx8QCn0Y+Ggy2QIfXb8W9
Dv/K4eY/Uv7fwgxpInNqi/MSpCkbTqUr2J4wxllTiQ739L8NiJXlwMUJtG0c+2M8
V3hrQLolMOSuD3lZCOapTR+wohW+tn6iUhjUmeNoaDpEUnfIHi9z9tHk5jdf0SEt
ga3h1H5nrkpJK28mfFLMWXaZ9TU8hORRAutoiQK6anaNCUF+6rYTJhEJY0//EW3G
73CX5Cw5VKCwAxledtrW4QtjJNuLGTDTyKsm7v4IkCKRVbZaLz1+TNdhdzM1m3DL
Bk6BskSTq7HLgoWj2KlSSyB/H1LUUoPiSsmTSTT15Sdho8xRaWmMuoIWlkfRknLw
9Q2yhSOZuV+UQpRQOvbLYAy56FqJyO7dVtjKjGK6o9iNB4f2tmX38gO6NT0MGoPQ
K7lpA7bJvyO+Qeo03BLk0lcCWsPPDm0AfjvKywMOCJ1XjRwweyfyrJdPZUPIUnhQ
jh1j1f3g0o2M9Yjsxg/4yz+7FXKQqc1H+qG2LCl3Xg7RHVGt0E3W/XA8E/t8WcKn
jqMe0sgl7MZA6YX3X/SADPrxrNIvC9XuB9kB2H5YjMN19kZO6LROmaX/s88l9CLc
ldmntyoDf4SrYFaeNgEXFqDWfgb3l+ixtTHQxlftXXwS0IrAFoEpthkWaqipZYxo
JSPMVWTTQ7UFLUEyLa8PRk2vSGX0gpONWqeHB6n5XVaIWuPRryeLQMaGEvZumsRx
GX5ngMgqk/Hv/XxsoQVHy+26sQqeGgmEKKkJc+KpImJVraU7oTvVT0uEHidUuhI/
yCQjY9sZil6MwKSYN2SfZYvIclj7F4GM7xPMxlLjOC9U76thJcOS73/C+45Z9LQO
UaLyuw18oxXYZ8P0LJJhww/qt+2c9e1nd3oDWA+cxBOWOhlY6c05Squwi4aCo1BW
tmsQ8PDq2e668dNeUMbsxUdiRteF/qGFth66KkNJKCPQWu/9uossEn5jGCqsRnnz
04JJyx5oAAkG8GOVRpsah9HnSG9Z0ueXLS8+GPqltoEWw4yHesMsFkfGJKzXKm+F
85y9dse27+QCBVdsI6SvoQhJZSklKf40bELVpW6swPd91Kqc0KQZXqj1eupcAf9R
OWEF6gUZ0XfzzvUfKj+zVQ/aeHXFbUrA9wrnHc767pc/cIqHBBt2i9I5x2Lqa5oi
`protect END_PROTECTED
