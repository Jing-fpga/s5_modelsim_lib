`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bJ2Am6v1rMlQeiOt9lRCfOs1lykZ+5e7WgE4pGArDcWrN+VkV9Qo9C/pvFofDpFt
c3Gf2X1J8JeeVMYG95q/iUIGI3e5x52qEc5Wt89z8ARdQYv1O4VpU6X1XNkMEadz
rw5BJHva27M4AQDd0HYJBVujkoghEL68PyyXmizgt3lPG8WDM/G+LXBNhZ5L2bqA
e5CS9bzouMRRoxSldzBY7J1ldOtAtxzEcJ6zHrgrjERGJl7rbgkXXLyvelivgbTF
e/V4RBliKNgSbUUhkgxpsgz2gowQmtkKnqJ8V9LBzxsZ+++ABJoxCnK/eNAIkGzi
2l9TUSbBCvnggGlQd7yVkGikOj3AywbW6xteiORhv2ZWUrONB/RA730owZRbSvKw
bXVsos3bwAIgzvPYwESOrDWTdUc2PMmCouAhRwCUN4FsI4CgXh7+H9UM/2TZ+10T
GpNn2x+dmAHhrNX1EH2NbDbFXcX670gwNa6c0z2bWGXGSsOQ9N9ssMRusvCGT66a
td+nXzU66G8KPQmhKXIlhvgatjX9KWHMwI17/cQFRXLrdDwf8vhIUR85ecqRs+eW
+f5tqozTzuT1TIS2zzyVFiO0ouS1/KiwB/8N+Zz3fz05BTadwMKN5V1jhR910qmN
p+ozmnF/9DLIMudtvstrRTqK/y5Fc8mgoXYFpdYAAKZDMPOzBM4hs5xdB+9FOS+f
nsa1AxHgv6PisCLW9yZDlOOGbMhu4ijkeXaKUhDgiIF6s0d9MUS75jknc1Hat2oT
F6GM3ROchpQbU1hlM9LNH+AIF6jT9nfwntdKICJTlv+Fz/dP6TVCbk48QPz7VjvI
rqUQ9hpa+HJp24b59JOrkStXI1IrADHcwiXwnVba7SzzzI0N9P+h21ysQJYwv6QW
nJffEGiQcRFQDvf7Qoy+r9nhsXp1Z7XnzZBfU7IjHk6tam0e7DH/jHwfnzGALVUw
fXxusq/fuKESv/yHwUfYLAZcY4VPY/CH7gzPlawRCnNQtPhyHxZy0mY5SALaog22
bDkHKYxGlrAXlWeEOieWUrlUV2NTM+z7fYOJyvPS4qcf566pzIky0erQ+0Oi1Kpc
496hW3lpDv7McLv2zdKnczXIg9f8VUaqqe2FWCs66kzSy+t6KuNbMuYNxfKwembD
+6q2nnHvsWlOk50Zm9Cemk5dgojz1kXTny5jif+jxtX0IgLsnO2SUQCykfz/WEEd
3E1KN9UV/lAvodZ31SCvEJC1hbk6Q1wCHaBcMowITkb5JsgkcBmge8rv2xbozGkp
xqxtmXM8pdv0ElVYkaYtmOPsrEBHOFK8kaNL0wxWevB+dE4Xck6I2vgeUH4fLZgI
R2JrEsAsYKLTOqZ9sElNFJamo31n+VXoZ/3VDrU8pMHy84Y8Rqwq+zTESBkBJ9m2
dsGRzmm8SMjagbTILUrRs/GwQC9KQDTVZkSpIwO9IHyZEXDuboBeLlDGEkiimEu7
LliuGcpaQDt/Ds/lLHP86k395wDOG6u1l9f+f7Cgynu5Kk9T6mLetl1wQuFI6iWu
8w7KwJ7+E0pMpy5YTWxTRG6n0HS3e4kG4FpKwPEJsPS62fpqxaSZ6vfs/DCwBF26
8APWWuLuKD55Yw8EmKHpsIQ++ZUtAdSpj2hs5fERHUU2vm5kB65H2p3yWd2y+Uex
g7qQ20NRozyp6MkYcneLtF3QFMP7lwzLfduujH5QF4uGC+2f0pgvxcI/sCR9TPik
4tBSNzFzPC9rwK+lEFyhLCllLad0878RT3xKNYMqbghyCGkUaJAure63QyEs6vAF
MEydf5gWIr+ZVd7eM6n182Nf0ZCxbyRz80VCTR7XLnlR9oYbJg/WjcwpGJg8Xdrk
4n6umgLCy/tkU3LfbbpJ5nvcdd+Us2mHAX65aJaAjANpwvRiDoT9hx7AJW8y9a96
4LpT069bdXpASSfDY0VgEqe10KfeGjsc9eGjjVl39RqcmrTlIU88d+mpeztCXLcB
nZnXTh5tgsXIjD8m8Dliwr0FmVYQMcIt9IDOSHO2MPCCzjEikJgpo+0hQB1yLU/r
+Wya845WgNbjDfyfQt+83vhtRHAbWokcVFmi98xrOYbJ+SFn7xvBuhwF23NU5CUz
SZ33Rewa2aabpGmF0KHvhrewXS2hcGhaMM+T5PIHFzaRMrfaSorTbWP+CL/KFPMg
O8axIzHZS1ud5YDxuDrPipJ8PTiDhYgifKUwa9vqX5jqLsplrLSwJPqPz/wY+z8C
Nt9iRJEB87mKqhqr08Db9EuhEvYf5uOsE+phZXerXUOgh/ftGXvAI2G9H5upb2w2
qPUAy2tBDav1bcwHA71DhTZQhUrTyhsWH3HMWqy+8ZibaKW3Lqp09qKM6kZfTPTU
Vwkm+dGwY3M+MLQI7CdAdQ==
`protect END_PROTECTED
