`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4oL+bj7tmiwpLo9SWPpoUA1Woi7nVnB6eZzFHRGH2A9y0+PcP2KDw7jCvOuf2g1s
wzPLh07Z2gWaa2WCfUs9AiXPQ9KqKA7FxQheZ0Czej4yrQFUf15f2kqqoyi9bYrh
05zjo6YLJBjOIX9N/Rx9EuEJSW8YO3xJ3zveD9XzCK5bY/vSCKwj9O1P7aUkePLe
bIdieQ/2cp77er4znWrRpytcCpQnW7hhLPq6eFNCLlXpJFyFwWJDUi5pHMJSAMvK
CYEhpK9Fg6zgIFaD7XuuI691DU2hV5PPXXwSUbSsmvXM2wFIyzbCPwsVN8AnARL1
2o3ybi641z1fufo2N4BAfA8t/m1rpZOiqL18Eh2MDd2ZIOuuMqtJXqP+U9IR+kKs
N+kIa4QcLZ3St894JHnxS/5jKgRzm+2eYCgSVyFlsnng4foSiHQrDzAJNnqbOJZk
K4asy3yHnNfxqmpFA3rIthbLgfqqY0l3HgpPavXR1FmeEhahgzhHcmxj38YRqNrl
h1s+p7aVSd52w4OzmXIBZh9LiyF/zGbzA5a6zAE5p6s+Y8el9amuke2pzu9+njhQ
rlPIC52+Qkhhk6UMh9vjvSElwyt+Hea8knvBD/eyL+525VASd38L3B6VdEAOs8zh
3fTkiZHoytD3dwYyS+UYmYpBwVl/79N5CFD/TUFwEqidUTCzST8GjsIysEuboCnj
BDdxrb1eu2/xeiJxSk+yn9hRzPlG0aFKjdITYOAT2J4zh2QHf4XzWgmznij3iBNW
Iq5GXJz2Onh8CZye1O0r5JEuZCrnFVixt3zRLa/fAH1peiqycPAO6c0TdkDWP4Ek
2cdKYSPEKy5XsR7Ib2cZo47wpqdfJdNKuFTxmr0NtWlV3XWfwb5N6orab3HqoYwQ
bAtwd0EYehX3C8+1J0v1kGBJouPD5PXjxfINfO7TpLUzDAdb3tO+O4aSu5y/7Bqu
ASMujUd05uOMsPIHI9ZspY35qfWflmZwxpzaZ08HHD1qYV554gBoBAC4TPIYjnQW
xx1SHQCE6eTnSg/N4Qc5jYIIy1ZueQLTSD2Zojm6+QuMxv9I8veTeO8OR+V460C5
nNumIz0U7YI38wUbuGdiEIFQhxhiDpEpTqzpgDpcSz8BclQooaheDpwi7HhOvWfB
/r74GUUgJQVWp65J/vcgjh1wRM39gdysDQn84wDPXMR0JZia0aIaoSnDnA77K4/q
fKZpxa0vnfdVTh/MrjVpszMNtZ9cLSK9kcGggaZebipDn7S0hiqyPZoli4EKtUkZ
Y322dokDPsIg5x6c9CypFhVLiWEB46NaMuCY1kPzeLrmkE7IIOMNwFpNMQOiOQ4l
RITVlUa5VHTZW2Ig8YLBwcVRHrJR5aauu59m99PNCHxvKnZxsas5BVZfkpWstci9
KnAscfmqNM8V5VeiGUhtFRyshslqjyY/av00JbHFK6XPOWlSxzz3n5HoCvk9s0UB
aGUMtAZFqRErPxix8B3Cv3810S6C2eX3lGPFbqhepiTGmXEf+fu1JZLrLPBVokNo
yt9oXsN8uswZGQNAOEmiTX6WjTuJZumP50pjJRdEgTND0+jz8/Q6eGQgyH0+d8mT
1nhnnVLH0PGGPbx/PV/kjKfhoDFRjQGDwaeukJSESwvhOKdSwpAXCJpDXapMW+OD
TBVI7ZtjGZwz76b4XC6EfVBsuKQ7m4eZ4KGb0AM2saJMqDPcaH9JyWdQbNEKohZh
fVc/BhmzEU0bDrBm5kERnzD+Tv6wmcWewq9ruI89hrvA1yGUhCgyOekMroLFAPXv
mhfhM2ZGxBKnNRboUkeTe73lsCWI7Dn+kOB47hW2AcZVT3fKKZNX8DjCZFUApd8L
5uJvNpOSuGfLJm9Ljx5KvKBn0OP8yGyphj8FB3VbQOs=
`protect END_PROTECTED
