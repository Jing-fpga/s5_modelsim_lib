`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+eZ6SXAEfYOS8rrBCjZn37aJk82pU7MpgJHnfvomsWnwBiDaDb89ziZAdzf8HdHe
03npmg+GgoDxVbfro4ywaeElIQYPfpSo7e7lnCuYAdeAaQMKkDM/dHCgCoqsWsih
df9uovB0z2etJyyNCRg2jtR+aYRe6zO92E/KocVGRsUPzzPtRW1yN8bFARaEbMO/
CDIGsSjeBMWgnssG40Xhz1R5G9+rNNXjtwP+NOyEXZdiaHnC1trXpHuYzTZFxrp3
tVEhlJ24RSvN2wKA8aPMfA2zMAfD7IYjd6KpeEPjMJ+tfe5NOblW19Hzz21skcAp
16oR7J15lxqqDbhZQ7KbkP+6iCvx3Cd/rYDw+eDP2lfLsBzC78/qpeWgmdzSyKhQ
XeHuwzfOZISDN+xoQH7nxPrOl5/zRPzRBwdMBTghxsEhnI6vjNHG4UzgoMXWTGLI
D4Y9QsEbcZ5Xpvawlq0KX+afAK7U2XiSR03G5BZJw4z+UwHWNqyuQW4rcQba3sE0
p53RX2tB6wSw0EBcvysplaJRAarhpHaNt0trF3MZnZ71j9grIcz3GQsur9dhNcyV
JhMzHxIVt7Pg8szcsVaZQk45k4IOFDuxfSKUMNLeWls71+H9shVQk1dmZKqdKFbO
Pb49r5dEYOzxp4cxPf5IohsmATnYztDaxb5QbqmgzFlLu9Kq6hU3chL+ur0dIVyL
DG2pxw/9nxcGH+94QLowoq8QcFH8tRQ1V/ccJamo0wf2r3ALY5s7c3jjeQIgCw/d
JMXRIglJDFCDuYWnG821ggorOHs2GdsM0MlXWHFpH/oKZ2PC9nXHRmHTo7Qj6SoJ
Y3yQQ29Kw0itpp8IJEr8LpenxWQE9dxjXg9x26b1B/Y+VQixBA9AJw2s+uMuL6UH
co1wRNuCZyQxEZ8hjzXamrwZ6uvUxX1G9GzfJtjFIfN4x6ff9bxqmPWAoq9oln/c
g3hAmZDMHeuO05ieJztBp4uAEb5qQSIQDkYfyG3qkl8MB+ncFJbquyjl2v/qKTSR
fvi6kuJmJKGOJQ+elwWfDWgOafyXzN7fA4RyolC9/y7jb5Rk1Nu6qsyzO+z2OI5s
Z5gfJCNz1of+BNTJKEdBGCux7gYzanI4u9Z/rzK8Db2keyVnfPRRTQjYK4lY1DGT
amq1L3qU5ZTy3GVdIKn6AypzevWOQbkJOctsE27y/nfefFzylIo4Fjg08YmQIW92
auz/u17OmAl7IWR3wc9dB6K/0Yqef2mTu50kXORfM+ulEIEFzAfJN8esvm6lRA6J
vy423V31TvjfMrrnfeLe9AUdlj7Ik/fJwtV+oF/89pvjBBDik1tgmpGXPwUuZh64
cwBuiebvabE48qGtZHMfXGw0bC4I0MEmBDsngC0HF2YyvI2Nqi6k+ji3t38qDYdS
LptEHND+0OtI+YldfbPvnM22VX8SYEa7sVHIvcOgsW1FTIvlyh6hlzWUOA2hMGjX
jkZbs4InKVVP+w45kQ7SXsOAkzT4MJK1kCrSAmVdzb84s+RUQaBlOg903JUp+IE3
yaPMM+TIFpYBuCfDKwrLfQjjvuE5dLvX0txf7J/2KJHOHvkYLTLYSGq/sPTwlOOX
C9JIBVmHzylmugInF7n5JaEl5DeLUWWGDGFa9T7AkAaiU6pm3+tsmyZVJNi+IQDv
d3QB0+uZtrYWNr31AXfgOzuN9byQwPXnZje8C6PU2Bx0RlaAvD69h+RLsOh1hd+z
ZgmXoHHPSY8ich9WgTjQV9nqZqDEnBImy3pnWvEfNpxoc1Db2YCBvRMJ2J0FdiXw
ArCJWIHSfIupiF6chTPP69V89kt/FpwnktLWNuQYPJWHjt2y33DyslXd0cJp/77O
8zrAgGarKZnGmdteStFSpZ7zgPbvdQkRBrhZ0SYkw+0LA64p89hDzoyunX6gDI9D
LelfSeNEkLdlTHofo+rqzqB9CLAda5Y8jFhK+M2C067SnXyz+PhZGyhsiaImX/E7
FAB4oAHf7+36XWA7jqV114eZUrQNbfMaDnV7P0DpdiqzVjV5CDBYRTb9tHC70TpZ
1uEByiwFfiH/n7j+ODGrNX/qwtp9c8Eav23mZMhBwaa0rSMwkJZdCp8rVfKk4kMq
HRCWazXCY/bKd+jPFVWNhZqIXc9dL7kMrLIwGuVJPMwrPClRmtX3E+a8yD8oXbQa
BbxcLE0Wi8L06/wAMnTv5tOJGsfDJTZZpX8G0sGzxnEsKtBsre1ADr411cEjcVAL
3SmgzdeHFj7iMi9lqkwylS3zglgstxMkqn6QeVfVfwH2n9Ug5JG7ov6lgMU5cqP1
zaUX2T3iRx3Q7V+89xZKpWVYwcCJYg+40qdujeVuRbCFK17Ph1F3RE3f7vZGz/6x
cuITvBVm9gxLezHs7M5mYLEfeYOK6hyNqVTT/QIugS3G9LNgAZYjFoaZNQJn7cyJ
3oP06pg0mfBAwnlzsdCnTEVFfn1g0ruSyQkcND3ODTs3F3k5lYjgYcnM+2imDpO3
iFoLqJsdhpwI4btVUQOpDiNnoU5UTLoxVA6m1GzKNQCmZDpeltVrID1w+1ZgLroF
YQ+3Acy0JC3FTQg4GAp1UBioeOwCj6f7YHXiDeeGBU7P4i7/5uFHjpwPxnIbc0G9
5yHj9H8+iA8unp5JQcf+vLJ3mDPpLiOgZTgkLux5fTM4LD7Gf8VFLMX3SJxvPS9z
/7y+GwoiEtFcKEDXipNxbRodcgR5+nd5c1NOZRHUetYI6kdATUhpTXCP8sg/R4EW
g0aeMj73xzxOhL2RQQU9tMVqOJpOktlhLEavQ/XYA23JOSrasczWWI+oTyfQbovD
6g0jESXN6CJYkwQi2dvK2co/OY0n0zq9g8Je0uTE0qesPnDK9n+sL0BpWx6q4aga
0MV5WlKf23xzyIqcttTL4rg9D/CqQMEq1LBN/Z7y1rXzewEp2KVr3h0mXSyQLpgP
0YVuGaxcWSHO1qEoMyJ7yw==
`protect END_PROTECTED
