`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tzimful2uEdBE3e5MbMlC51loaUzLD7WduAyZuuonraKMmn4W43hjyNzEhSlQE5J
YT1xcc9gO0A129QyENzYaRm8AakNA8Q9rnBPFEsNxIGPfogPUB0S/hfL3bnPTgnF
3lPJExH7KM3aFBTusk0J863BpXcGtjbxG5X947mThCKlfPfw+bD6TUaqpLMae2yi
mHFVcXjBQ7il5aR3KvyZTJBh7Cliknw4wA7cWmVynLgbLnqNRtJHFSKxP5sKzIAs
GmpGE5ygrJ1BWoQpayeDIGvILBgojoffYm84Oo80PsUiKAB1kmAULM6DwS+xIxya
oSWfn6iNcgMz9YDJHSMzpynYUUp7VBIgV/bJfWqHyGPKLR3kDivTbqCWr3wZ57Ye
CLf+Ui7ra8roSZ8oC9nbm1P/1t9RJ2YMcjwGr88c58e+Ba6Kanjw0TItP5gM1M1K
jY+wB8dNoiFO3cVRtSW0Insum0AL18RFUyTxLvWdItZMA2imSXn8KeBX+K7JPjGD
mxE9HUEPHv+XnsTsLDA/ByJmEYSFj3Bm1kb+E93sjG1VmL6LgutvGvZecbrGvbjp
fHcKQL5FwmEfzs5Ao7+3BzR3Gam3Wv0Tgve6spgzmZpIfoIG7R2SUo9sdSIDHZEc
3XUiQAtt6s5oDMOfkHDPVGsEV/xDw0TEO+F8LCaEnftqlRYj8xW5Wuyh95hXofLM
/BHULoifBwkjoWTeNuH2lKsb3VcfTHtwXCVxfV9IKhFGkJlda97qy67sMMC/J9pf
5QrxLcnv85QCDVp4NVpLmerB11zZ3cHrTKHE1x9JhUPQ4O/njkrGXk9Ejb9go9rP
4Jw3twMGW9jjQKQ7XLidVKvuzL83C50wo9zLhxxlme5W0pn9FcHH9VsmsWQmsbmr
1ZZ85hqwOjWrqaIQkUSU+0nKF787fs3HlVB8vQmYLrDPTiy70lfowarj1lq3SfpZ
TSnyLwYOirktU8qWezvBjUVSU4/4FUYCSK+t+OvxPS3P4puFvEOxjUYjG3kMz5ml
Ei0a3Ws1yzKCYAa8L6bjZENX5/KmPOcJmPWEdUdMGer+urzhDmwrp7UQCTXd34kL
`protect END_PROTECTED
