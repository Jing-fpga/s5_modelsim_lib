`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VzymhryyZCyBNXMvKAWEcO/llV4D/TPhy6i94E+RMctrDtSEE1s4dKKpCUilXGII
t64Nj4bEnTiJooe6Jy0ONWEMg1NSFDRPAP4C9XenShzcga6cIfWwzmFCjdgxJMe/
lYzJSgiNIE7X3AZmpUtXCaNRDb+Es4M0XIiY1t/7O2VTMg4FA5TMSsLK0HTKm7K2
RbZiuWA/wzqav7t3IhiOva/AMmzIzHMyHsNE7KyWftgx94IfLGvsoF5j+RGXcQ2p
bHhNF5ZX1UNkn5lSrRBhBw6kCSzwFcvOgv9X60HR7ldfSAfm/AQlGDzd/PNtCdpN
9xkz7SgB3ZUE/WoONthpY0dQ8m05tfuu44iXqp6PZd6gizAMupgpvz+36Emq/hRO
GGa8MwwNsBtD+/Qz+N4wPk6scRV8kryGzBgEajex1lkWjq2PUkXMaCk4WDqC1I+o
ocSNKrx7tMKfT13zeCd3Jiw3H8PoTRLB60bUPS4sHABd07v1E+m11U6WqOR+7aIa
619dWmYsTLYHD2UPWg5a+jc3izTS+KoFwMA+knh4GSJCUmFcjm1naP2ydEJhiDz2
Ce44Ms655q9Cgy/2tgG0K1u3E4bNZVgwYH8w/rezFQkNi1fKzjMPrYfB6U3cYD0a
swJEdWD0xzTOI9r+ru2oEhUvDNtm6n0sVh5q9YaNFl/2jkD5+VjXGnppftbFVtsR
hRl7a+Ke6kNX7iy7EmwfaL+ifOW8VsbOJaELHK4pkNwCHpYO3xIeBtpDbISg4Nag
4wrM8s9r67/AsnRRQm/g26AmC6hB1YmzYYTtFiD0LUhSLCc2wukZvQ8Cvalrwvr0
W3OhuIa/UOqRaaxM3o3FbrcOpQ0X4NnU81wjGR73InFrXO3R3KkBSDhnIdBgY1kE
PQsqDg2XWnA1aHWcMLnUSi3NPtKM0Pth8U1YKGK6EiQ=
`protect END_PROTECTED
