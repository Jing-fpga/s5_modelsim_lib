`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZoRSAfNglba2XBrA8EEQBQHPaoHMtHp2+zoGUcVurueT828juv+8TGlceDwYP1mE
uYivLjEgBc2aLtkZC1aEUWkdGzFTepvsTKgKLmG3ltH/cZkh3kRGq8ECOK7RJCMB
8zGtXWapCfi2UIbke8XBRRy0hTP5X2t9s6arWyLwqEnAgL+RvP7/Vi1EMBFIzrsv
+pDwlw+e4ouVj7GnYjwu9KzOotmrhZ5u7vCnk+SxkdsydYNB2zuVH/qSNEPojxTb
8z12NHBa+BNwruZq1GTYO2TICVV4seeu/92OEeMmM46TkUXGy4QlNePfXBlU8vSG
VrhZZgk4Un/FyqCbg/FFag7GUknw7LCE4swkAPgY5VUycO3sGNqxo0lY5AWrJcVH
sn5CT6vmE8MNoOk5/IiN9TXnJHhlA+JHd61ySQSO0c0nozp8UCVDTKcIpMogTYF6
yxDq9wy7KBvXJPm8GwykHfP8a+Kpkj69DB7EzKfM/Z0pwgdNdF3UpB7AlYDePSg2
vs7Qgcp2Uim+gep1I4a2h469KLla/iyAi86prQ4yT7zVypj+ChcC2ltJmuPXK0BS
9/5I0v3v7WCMPLPpjweOL8OpR1qy2tlbHxxy/ZJqctAz9qC9ojuGRQZbtM9U/IX1
itu6gQg5EI3G3G7N/Ly29LB4o1QnMusQ3oMB0ZBGHNwYx1imGOpAi1WfRbTfI433
VpsVi2DBn5J5I2ooDkEK8+HfTJ98V9XOrHj3og5zgHMkzhJfAEkGmz1RdELm5ZmY
PyeQcZhZZDHruW6PR66lM9jSUSXqThTgTKbytTl54qLMCa+qtP/AHLjbJlh0lDjw
NUe5RrZc9ndJQGJ9G5fbP4MtddA28NtKIAkDXKPIfJfduelRVaZ+CgocPEDKdPoI
i7k+BgNjhmaQWyJ9tr/j1+IIoczC8U43GXjJBw3zmcNYenJRS5CnwS8cKO//AJm7
WT1cZbPLNmF97uEt/ijWCJXZwVw9MVShykPpLDZSQJuPn7OroDultaWT0lYFYJ5A
/ID7FPjbTLvK6+luJRtj4yle7+lq/9wbUs0QAijXPb/9fg+b/72lfvaI3UfyjlHi
qsGnKgImQwpCQhj8l02Gdnpl2sTsku7/A/XIM6dSj/miXX9A0EWsroD+5xqhg+5/
P6WWua/hI7Gk8aJK8ozaHGpN33L+IY/wjkl63ojM0C6r57GER3fWYHWDYdEBIEIJ
1cQ9tm3MOj5NFykuWLZtsiCScUtUNxI2BOUGT6YLhhxifWUXP+iiiRiBc4fc9WEp
Hf5Z4LpGG1JzHuRO9ikzvyhk0gWaGDrzX684YwPan/nSZaW0Sspr6WhF5fqI2yVQ
vzyF2WmEXJUQj3k6ZeJORxaI7aaN/YMSDgoUdWU5YUxqHQurudkhj98mtq0ioDLv
nF8cdLCSpYs5RDGQ5kzjRelDesTdKGfNql7pEeIK3ygFL+m3D4viKZaGSGGo9iKD
OcAffnoM65L1AVyu2uS3ehcjgnP14KjuzAXsH4nelsknmGpqnF/+dxgR9pzI0nXb
RcjJUXt+b2iiPZduyzfNuB+u60Tg69iabqwZ+09w1vBkzX2NS7s9Dxn7rtyIwZhH
GNhkGPbWu6cWa+BiGXRZDkyoPY5u6wkBiNz6r/RFPCud8cnxGYYapxcldOcTEryX
5RHLo+IeQutEe6EagRzNQQnY82XpeC7o98EmV9Kn17R08gs6ZsZGYvzV2DRWbbBK
sqbHvwTen5iA1H2nT2EafKE0B6Y1vW1FXRyBy1q+CQ7qPA9RQet/kyJ4JQENq8F4
hHdjuArSZmj5NV86GRqAD8GHrGLO/hQbFs+ip+qQ2NwyPdScg4l40GoeoZkylk9y
WsFgg4wnHzmomm3g2xw1vyPY+y8DYwVI+r5RVgxNt3cDy9dWXmLmL1kPccKnxdGF
bwO66lUHYBYURseW02ngSYlKjqUDWnCXyI04n385Y6zQzq5LarMNLLUS8x/kTW30
27ymmTrtsqhPsldnmCeb/lA7U+BaWEnam4NYiTXceepao3J0aibhdo2y4v5z+JgF
rJx35J1+YQZmYrP79zlX3BMRVWv6nlb3e7a+HsQOn3LnqT1UwPKbCejy4bHSU9tv
ufF8x3skTeMIFNV+OIiW+np2I4fWEaxEuhCPYqTGjWEQp1vdShIbKrcam/kmIK/7
84e5MyVIEWNDfp/uXy3UffrsB64OaE6iBh8vooSu8NJGuON0GRZDvJeaQXqF9Y5m
uQFhrKI3/wl2Y73Q55xG13yGtfM+x6ymCa015XGAohXjD7pqDobKCYM1CXmsgVgx
4zfptUVtuNYns9dReSaW+xKREHYty+kKIdR8/zVogyqCHqpN9TprqsswlyXoHr9D
dhld28qoTxbwOJpOMAhZgO0WTsVrPIeRKNJG/GDtOfYfhSN6STFnz2OXMNtOPXUU
0MeIQq/KcuPWE2lDNOZeRWQcnic2k5cgJ/UKxM+tqlg4LjdOeTmxH7sGDbu9x1Y9
aQ0/XsMUK7fn2veIHHMiwM9J4SJMeF8WpTnG1nsUOOij6KNgPEuCoeP10JtjxMLF
7t3RPC1cifnMwl+YH60a0eYHoTWP+RJVejysPqF5NRN6hG/JZs0bZHmFavIyB/vc
lcUzDDcP+O8AUDgiPgzP4rUWnaA1Hv7Ha8ktiOOufuA=
`protect END_PROTECTED
