`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wPFvPpwUcdL+1Iiwv6CPEw7XyWRieDXnCKyy+C+x0WKz1Djh7pOnNnK4wYRhMNff
VQD410nbCIOL8krckPsNi4fsUjWUpcW75cgGE0cLkMNL6QO91ZjnGx1iZskPRjDw
P6gSdhN3zLTENGZQ0ZvqkoS8jHuz6D1wN6dalGmuHbIdnSUY/3Z2Gh6sXLuRT8MS
/mIAlfk3A3Id0y84F4NbOAbJqcJZiIi30aE2w7fjkZ7JDnz0BzsODYLhyZLanxBG
lpHRelUCNz5XNYCcABhYx4Dn21Iukr8+brDZsuc3zsl1i4OhG006wv5m6jxymSyG
LUtpjTwiq6iqZ+h/+9g+V5yGOKBkez3XzbcjUCiZ30+EfvqZaPFkUbEZhch+eEgL
XA5h3EbMVSONLwCbTtNdQNzLHwwGo/bDGqe0KAyGdJfWxcoDmqfYsMQKy8dyLUv5
e8AYbI5/lVnm++tFmUhMg4LyYku3CtJY2rrXux4Z6gqgaP6xwAMpRu8k3yoHvG0E
NheduL6eRljRGnytE8rWtqWnx9fV/LmnHnqkWmI5EnNSYw57O9oSpHQVWpOKsPsP
13nu6abjVhyNFQDS/Ghoquo/TmjGxpiThGCQVF4R5wdjdpaVwq28GqgbpOwQ8tWm
e2tdsbv4pCpz95rnHMxVYXrfQjiyKY5MpzwU/Df3Ulrpp7qA6D8TUfSGzBGWagSM
01mM0TugVgjKSuPwG6t0QP9SN/Bgbvgj1U4p2dBabAHTUGsfT54g7/OiiVxGqeUh
lavexEL1a5z0MezQeQVd+cAbX6/rOimYenE6T0r05IoN7b8CJdyTjDuQBQHx7Jy8
HYh+gUcYeLw4sb7U4MaVPhRIh2GuA0N1I+eGEVDKuVK23sSBPYu7oEtYVDXSJkv2
N0/ATdion2b5VHY6NCwWgeC+0eCikJopyAa6yZu5u+hymgpHHtRfDHgC/7ronpz9
K+9yFzavlvqYm2Ek9pGGDVStIUj6jEleugSJClG71M4ua9CMyAIWIR6wVxaI7Nsx
cgUAJ+uXgxzDq9HACD7EmPFNEIOgNCMrQ9yqiaAxan79tNPfYa12swUucfLRmwGX
zAH0eNzUw7G7mHHntMKxCbKNdS3ICNY+VOnl4aKZwVDeBdvdxiSbhxg6SB1i/LbR
BiBS0vCAbBYIDxifVmzjCwqo7SCTuT1HveS2sB20l3Z+Rl2CiJIJII8LvJ+Kb7bl
ui1lFHAAJ6tlycn+JkvQfwLT9Fhxzuj4bP1D/jsRHroP7rdwPrqcIveyljNxYPTY
H+XYI8ZxlDSH83kivdOILXMbvdaptK1951o71S7UhOV7exa0raBopaqlpYL+wA/R
94zfOlSNpjtQVjATdxU0t1lmBSsBXoBsaaGvU+5pIq2KeVCZiyV2myGgXrzgImva
IIdXxn2A90kSkqkBkVjJvog5zPsYijAQOQ5A2U8AI1HH2/3is/3CXPoNpjgq6Rwx
PXi1NPGAZmYsY+6RlVcLdiVFPfC6XstBv2Om9oN+XPFhDnCQyyPI+GvAIzGvF66+
+jACYUci/Pw4i5alyl5N4AKJU7T7jwE1Eq+/UNTYez6xrG1k+OneJAvjGUtP6y5J
/CGzKU2QksTvb0SKLVD65CLo9dwe7N4iXEeu6xWvbal6z/FKtJXjt6s/JnB30Sl/
h6FnpcDVB5p1qh0l0ypJN5XjAVjdUhAx3nSgQMjKDeUWoqY8eRTQmoozp5P/9kAi
Bb6WYTV7bcKLycBjJZ+9o15oL4EWHqLsuEutUyfIMAPT1gzGJjjbuhRsywgxN711
8MKJApxiFQeIehfysZvfYeaLFN/oCLFh7Fgdw5ha1Sk8KGmEfVgr9GW2Toy+rkch
bwbaxuQlAH9qnlxsYN7IOvoYDAQI+t7xZBvpFKKDeDBl85taZUS0EOZ8etuh2SDw
P6AN/Q+ebwYBtoAFBsYI4Mhrc/s75TZlIPzfxzQYxBlXmgsBRFGrq3wK1Shpj+fg
/QU9/Qz0GtgsMoTMjQ5Yhsi8Trna/7vVkuCjaDO0mHg+ThQ6osK1emQBG9RvdAR5
cJaZlHuO0p+OUkjedbbHCaP0UWdyqKcHTBFtj2y67Rt3TTpfPvYfVnM0DgI4wU6H
++3RKzNkCBymKGTu1dji2+EDCa3Xc2Krn44/GoCWgLsB1nWRKnWuboBeHRPJm5QZ
wHPb59093BrU8RTPVtSr7q7kNCT6LsmzNEX262wXwTqbqUETLMU2LEf1wpo8+Kjl
g++76gqkTodpafGTyH07GEGuCDGqAsKyQ+zIV1U8spTXfA42DFl/y3mlohtZMWj4
6koYqKKs/w1mzgVewGPYnLUT140Gk2gec3lLQCX0rsGeaDS+KI2Xf+yunAJh7Q8X
o0yizw1A2hUXpo67TbFD6p7HgpIy6eia98ENQayXuOiCacVpL2xoj56LQCTzqh7U
2XWlE+phog0YFIHZleqUWuN0TGrVglQ7HqE/PR8EqYrasYUpLE+vcKHncFyU8CFI
vhrP/CwwmvQbEUufGC/a+lluvqvyXqFHRweJYYjPDyq5O+CWZOCZeSbVOyTzFf4g
7sxICoVO8Bn5NprXRmxT56EWA9Z2Le2vlY7AGf8EaggJgYOX/hQTUZ+lAWmYCjlp
3Goa1+MiZ+rW9hBbsPGzgEle87KqJw9nm+kFkTNL0RnMHeXq594gDEpsg3SSkUoM
wR3QqpHnt6mHu7nZ+bgVYJ3VW4G0+jowW8iBEf9HGI5+UE98arv/T0PspjsmdAyh
PeZrjGJEK5ZK6uV6uRxiGWNlY36Rvb5ibGJfAc2IwRgyskO0mLxI1HA3K8ecZFPq
zTdo3uXhRRh4eltfwoqckcrJzAOHkXJVh3/o4l/8v8IydjyyJ/T1M3hn8kKyrC8n
m/Nm7XdiEDMyVzgZR5L/rRdh+jLkk2VZrDZYihouK5nffh9vbq+lesALwVKin3xq
Q8pgMvQhU+nwRMEDdZOojQXzBKum4L3R9IVMAQ9vzZTHD/HFfKvNt7wPeQC7siBH
5kaCRmosIl1dn6hBA2nrdlH5jUCxX+OJYZ05cBoXqrI=
`protect END_PROTECTED
