`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xBG/dxGmFt0C1+yaKza90bgUsYOn0Dir/kUZMMkV4QlpQKroHNWXj7NR7IbkYIEV
ONgjNI2M8/fBHVnk4V9QeB5Szv/I/hRjkE0YWmXHYFVfx9NuAitYrsmOIrSEAmT2
6Kkh0SMiF4jy5CwJfbp9btoLpao73ZD1sxCQ/IDafBYN1lfPUdITwDLJq7HnX1fm
mv4O+/GLWmDMM5I7BsFR+dVCaHv+0VoZvodlLXmTap1DE/bJiXAewud9h2kynaxz
2Bkuev2l6ifFBxZPyAgwyNaTxowXinAcgM6MuqyXZu4HiEqMeyPC+FrtPjgi8U+q
N9wZvSOJdGcDqnCTCj4hYiwdh7pHQYHjKJTY6fFce2qt/E+CfgDH/C/yAiBzHcBJ
JFy7Am2rH3N17rDV7dEkI9HrawarlVt9IxHI8BB7hQULmwO6tGN/tIovJxjNXg+2
/7lf1/BgsxLGlhQTNon0G4SZtkwCiEHyC7irXJ3dydsxspYLdc9waSDlIQ/jA5YE
oFWejcVVo6r65SdJjZ3X2ySTARv/rlKKOpXwl7tfqClE1LWFPqy3uQ8ZG1IHS1R4
zMWloLJFG2MOC3pf8lZWnvgX2V3D3/GuQd+fnTbG+wwM0L2sZdZl+ebDmSMYFsrU
unVbxfCdzhdZI4FFTEXTL7DbjF5sxlu6HRSz7zFGeaU58Q6pyxlouB0FEPWKN8H9
`protect END_PROTECTED
