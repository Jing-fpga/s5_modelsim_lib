`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eXXZqm190LhvpqNy5hu67k79PaGbZVaLb9dwak0iRo+O+LW1K3j7cnocLdnTj947
VcJgv0GQ8rkY/803Vz3yt7vMXiSg/OnWTK8XYbR6TaGOfr/Ygu49hfQ6KAHzsrg3
u9uFOF6aTNUqQfwqIyNrghB45vtsJMEV6Hk1huRPxiyGSsBpjpBfCM6z8gIPI5Jp
/kzm3AEH9xSeck0xnIjp90//ZH/hr/BDetwnnfNEvLS1RXbz9A912stzPFeC0Ij8
bDu5lofS7WHPCFg5QuAGCRFonFmTi/SXlgVd9y0u2hCvFkjfAZ28iuoWHAUmuieG
s8PJDUCZP9rLkFlVceiQLrxi6VOjh9L4byKL83biWorwzZXb2fPTeCMAsqaAM59o
D+VE6pThHhrhIavD8v9Eg/xXP4279NQgpXQPw1qbW4CJo5dh0HxPHhkl5PE3Xgtm
JGyjUNrPq6z5ZCzR70byWkOMReLOpJ4m56oSfWpD1aRpFxS/oDJrHtZ0Ear80+Bp
QcWopPrqX5o8Q5oQfFYOeNC1yfwJEbUQgCb0BGuHO5oU005UVFcosjZumcAsJG6U
HQ9mupjLKR89GLEkcslNLtLhb/UB6XxmE+JmAfJ/+QIrcYBPvpb0+bqxgjI0T7O8
k/AAr0K1pAKCDGkfM4mwChcCo1PIiH5ECv3otCPQUnS6uyIi1CyREAQliFwoFHi7
iMxY9XAml3PBv5JdLz3ZpCJWSjJvBzS4YwijrTdFtEhgOwBwMwXNshs8OaJs1cGL
H11AtAVXEbcJ5z3vliELK8WtY4WiKmUQW3APfcbStyJTTzy/NAkw8dzBRwdBlDaV
2D3nOqS46ujR/IpD0E1uaULGoAL5iV/UXJeHSlsFEBpcbZBeGDAWZqaagpBJNSz8
xDYIaifeEXxyEcFBNGDrUHen4TsZpDkomNygHOfwuY6v67fO8E11oFlwKEckORzU
/fYmfoWwkjPqDYwdabqPPEF6QEVmWBvPeiyr8/Qoa4eMY7lOlu8mjrDoy2PiY512
niehj0JnR2gaxLkamxbteFoZQXmG3nnV8fu158parucWSnhXc5wQ23dwB63QwEc0
j7aCglCLcnWRStZnLUK3FtrfydSmv5iEWUi3cHy59ymRLl/MWTSxi8R/VXuZrjN2
n7aP5n7/TF95SgWB+gpxWMHdGvw52xlawGP02Cb/O9LDsieoxw9ecAojfGnoI/7D
wZ5xuv5bCkSDY2IcGZNn1943N8S0xSgNnpSySQl63obXWFJsjVSaOwMfWMtRRHi3
P5UyS6abQEtR8t+xOmrsOndahj7nO8sx7/Vhm3nup2lSnyjuasV7rItDjFpumg+4
5+W0Y3Inx/e6Rr3cntj7wA5uvuuLOhFu8ZQMwSwOx7B/ok3j8tbzHDaVcMnz2a5l
XU2Od4r9RvnmELYLzpaDjrENJvZMkJVm1OX2uO+hXKqYeFca+P//DRRdHcyQBkFN
OypmJoS4O/yWEdGLo+mGKVZQQwYf04/EjyW0z3sBiEbHaCvOeAK8YF9/ZqeHRpHd
DsRLXLVPrINxsY4nJcVYIXInuQD3mqxLBWIR/3rnaL3d1C0Pf89LejOAxz4RxRu5
oNqhlkqjUp1bOA384sky8JPLOxHSHaeYXTmOSH9lO3WIeJ1v9Y/wxoXyPcEd/3W7
sr5KksQUk6laBYV56Jfrxgd48Vk8yuh8Fx2OM9B+lOv11TNSqi7nf6rZMvY2orZD
gILSvB61zT0yp4ynJo703d6nAdb+Pz/53L0H27QLScun8DH/zPLnF/3PAPyiX21a
mDdP6D+I6HTTvCsBO9WT5Frpp/X2tL9A145qd4VfHbkeEXlZkNfJNFlsck+p9Y9k
ntehRcZlEARiuaX11WLQw3WwWVruhw//RYWBl84vzjdbC8g0ZEqThNU+NngqmIYU
3gNpAFQx2PtvPATuQ2jFNNNslnRsH7H0ZRIc2aAtvY0CR0Lpmli7SkrTHxdfAowK
LCzhOzLE5p3R8xwm9+NsbQC7NjP8rLKVI4uiKrU97N++doaNdxFk4tck1AocpEpP
cyIFWvFC/3C7A9Nxn41zWhJVhrcLo2UrU9HDDPYLAjeKT8HrJJg4q/0tpOPbgDBB
UG4HNMgy04HO0+JQeyuube+x9mWnwEKb+ozhwZyEz3s9plIQySl3apOTg6PcmAeb
tQHb1buIn8kVllvb1PmPJ4ZjkcMan6s0KzNnGbkvGBARzpKvKybhZkA1TNVRO++Z
LtZtCLlZKODg13WN41B1Yj0c49UVZFzVJLi9wfk1JkLja4Exp7TDMyLmAZUc7pav
8aQMhG2jqZQbn5X77mk3ua18dqgDbPU5Zc0u0FiJR/BjeJJs0itCRBkD+xInYG+0
VH7E+MLI2E6d4H79RTPsR1yCLAgCfNEwZpugAiTfAZxVbN7qQrmq41o5qJ8onmyH
Jp4QCORefrI65i6skNq1rjcRC+NlejrAuwyil8EcFX+h1SkxwpbyaXph4bMwRnIy
HBoHl6eAJahgGYWuOqJUInk4EozrYZFM85I8tnd0rDGEWg+SjieFkxFlQ6co071G
rgCGBvpY+vRIbL0J4KXJRDCTfyQjpQaVV5lwccdvx61ipZyFJBsan4s4HEVfSLWV
+4Xh0/MJKYcGbDeRCALfgD/AIMXCZ40CJVtUngLAYQX2DMmfHpSyGC/Y2mb2TFJl
bcwyPeCvaD8xuWPsZBMCt7baFu5hRRDR9ZranpDAqXU3YsASzaILe69WEDspyjeq
RNhHPmhgwI2GcM54cLFW18T2cn9OqnmM3nbnHFLhPX2Y7nty5DK0KbHJFvAlf40v
xh+nJFBh5XnowVEBDsGuk9GZFkOsP/0Uad7ggAGXKzicF7JdbwVmzGiwPD8FSc5N
OQWsCSmCWph6VVaAUCAr2lmDR/Z2/ASKWbbX5nnWP3BgjHmBkL1uTScciPaHOFJB
pjI0xTPyyMv2M046hdy9Pn2MCD5vQzZRsGp9Q/aoH2GfL+ej7TGAaepe4H0cjqki
aJBmt/Z0xL8JYa1Vxmj2aL5UHHl84bNgZYP3mwe4tJOnPT+5Z7XAbEoqIhorkx5M
kWZ7SGA4F9lmIZZbZgPtzsnI2C0hsN3Z/zaa+2QzYbmrrDOYBzxP6zAMKV4NUb0h
rjpazpxSw6iSe8WYV4jQ49bYjefsxEec6feg4+Y8/Cz8FZylW0PSC1JSPQQS0/RX
imBgru9Ktghz8eVb0A0fLP/d39Un7QvHXv8vT7pjFXdo8z2YPWmbGRqFZqT4tI60
W4Zxi6j1AB0gipvfHiL/co9Zrbxx/JoBxhisqVtSwJPIF0T5tGl75FZtsE2XROkb
bH/a85QdNGzJcFILLhPvUBf1Ju+K2aLfFX33Nt90cXk2Ms7F2U/W3S/qEX87PcO1
pW3za9mfZAT8367Jho6cB4MADfZ5+jURfHdi8OEno2rKEPO6ecac/RP8pEo5zQSw
9hmKLu2cUKUGdeHln2Yp8uJpx3DPWtTvt0znxQ7P1R5oSNN5oZRqCwbL4kwHd1IE
xu87fAhWM5JsC1Ac8JAi2zZzXT076ZIipbo+5nGKX0VkAGjz6dckqbzMFiZykuJI
fbOIsqf5wLq9DkPEkPAXMMF2e81j106pUu3z+IpgSOcPQU0fOl0tQf24rrSixOk9
seE9NtgG0+4OS9J94msII7wY509wi9HrzVfHcWY+ZEg=
`protect END_PROTECTED
