`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FMwH30GtxQxE6MaVssEM5g/o0AtzlUgm+2SY6Zvf1urpl0wnNYV4H6Sq1W8IJdss
34zDfgAQBBiVgiDRSq0hKpyQ53SH2mxjqxPl5PzVSBVgQ2dweLuwb0PLLUgbnEUi
JM/lYZTi2XUegDP/jl+1cFy0GjaZKrA1/gQJQXUk7OyVma5RV34EklffEMXZE+LY
BjIX+F+NNVpf11zqnyLgX21R9rT9EYtRAuobL82oqY9QSxYD+xrUXxA4GA0b7ON2
oUprmKaWYNifmDhhAtf99CFF9DX6EISoHNGIA+ZHblXzqMkjrM4pEji9crB/FbH+
84oyfv2pbVbonPgX9jvao116rJ8En165Z6NkAAtYJJMPyPNRZYIi1DAuKRwFy0k7
+ypwmyZlNS7Lsqgy35R2sdydtvvwBcsONHOKKr6p9Y544n5ESm1t5zJhcdh2ofBr
dv4INKFtj+boJRrXtyfhkosbl6uQoQHRaUdcZJ0fUC2scMLU8wlcaXebmO9LXu2Z
hQnpOxuquMFz7eK411cdRXy52rpNvy9UsdBlnPbFLAgWVKh3pl3RtCsdEFujMyPF
AKrAIjl0UpGECMy0d9/81WH1DnS+C6p+NTosULI/LZwkqxvHxqI8y+6PPkTqcnQI
ioFiHOXt2wZ9IT5jUVxMHKP6RkU86+luUsdUIZsTcp0l26Gh9M57yzScFnalhxFy
RnRYUiPb3YF7HBxLiry9KkpVc/E3Qs8+AZQDeCQNOTw=
`protect END_PROTECTED
