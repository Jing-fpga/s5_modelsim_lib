`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e6a8wrlADH5ldA/iWjS/5iTnBukCtZL8i+8Xsu4N3Dj4eJw5YwH4Zvx8mLYQiOUp
q9+/dlHuMMsmTD4kdkYJEQcku7hCIPiiCWS3r6BmUJEKF3I1KuayRvE0qqQu4Bi7
GJwlGYhYUvwuPwKUdsVrmwyCZnSfyzRZ1UNwoNw9QHxp6DOVSQT3UE5Mh/kG5fBl
EptDC2ALGcIfy8lUETnfdOyn8aEnXwZgQKVnJo7ISARLcQgOccok11rtz9Li9Fnh
FN+H3mm9z03fhxz0JrR/7csR9Z8W+IqrOM9Y53nGnlgmf3HIBIJIdbZ5dO9rlXuL
L/XbC9xQWu+Y2bqshkOBefXgWjrU7opEWQW/xpoNCX6rnh7UVnB2Pcowt1HpyVzT
9+aGuPwklY4FHWG4w/yg/OnZ7G+eMKtYRmqFEZJ5Iq4rK4SkBUxa6qzqY2jhHPc0
C/KMbd0eEvwlBE1u1TOWzUFQ9VN/gOvA6x7qpfm0DHwhO/mJNqLDbruPzA4B5NEa
cEu9Pa7LEqY2vupsbgil9e6F43BkdqhDL/q4wsGw6rm2ps8WMJsGG1r2ah7F4vLr
ZrTDcehAF9Xb6ZRntSf9RxAmmK6ugopMCZL05IJQq6hHjDCxSSHyu1YTWOTUUt5m
C3fD/9mwph2oGuUtcvYDCJZSiLYNX8VVfudtO5PhUrf29PeIMXT/FLz/VXfm/SmC
Aq1JxT8bV60Y/DgAiplL07y7vkWUF6E68JtLgGQ5XkNMclsxeacd6cOo4ifvR5fa
/G17stHkBBoL1d5RTBI9rLroN7yT040cxW90/K37l9eBoFBXn1g4NxXzkiakYR1f
weL1gQKj1o81EQ6ZAzWE8tc7p+YEDIgX9hzRqL9jcWBL0eOsLNNSDroWuk3pejXY
t0XZs8GhBEyO8nQZbcMgklDz29tVmzgADigTI3HKG3c9oWtEoCb8Qxlw/8ciwYAx
WKTSUhdwdiGez4A8HP43/Q2PGvfQIzXlY+apccfh2HwO6MCUchrcJKFD1HMVX0n3
/T6R3jdDtvTIyM1+gPzpJhdGXSMka6SbitaJusiO1q9PgsCUV/9gUZlEIC9HXb0/
3v6oJ69Y5leAvmDpx1MkZhPSm2VOINxqcQfXJN0Hk8skpbqMPP2zJCGqJqNGqwl+
37cgsQIp6KEgaqs2BJyX/aq0Hnk6Qb9ao9QzcN4mRF5ir62svJAaVY8IDIWAndJQ
qOKipQQgDy3r/nGPGbn/miJ8IyWlrMgUnSj7P8CMcnO2FtDe2dGUzRkcOe+yBtF9
ms4XqI0G0Rr/Ii7wxhqxOYjP/sHK+XmpseFEKshAT+ghLwW3f21QCkVz5zwt6iWl
UOKUCrhOWlaTqg4yiEV3vUhKysqiYJd4HoPAWbzvjVNHSZSENMe4HQmCUv9npQhf
kfnkI4BsUk2O0uzt7SPO3t/UbKf5H3+6X/3kDArqV5Zf4/h/MWUFRa/G6mDlpEVV
1JYft9slWteMN0N9Cip0WbBeTswYP1iDC58m23Dk1HrXpgAixAo/uY4OB1ftFKs/
xD/n3Qg2LDzb1tbZDk6Xy2b51nB0H06OXEQRsI11l0nGljbiWuXgQEOIEqAWUmFB
/BtR6OxKbU4qMxu+gproWp6LgkHQy9HlT/+6v+him5VLtpYd6yXC2x+ALLOjqb1K
VaEgyiSaZo3uiwjvy4U0Gq5Ea5jkgL1cCSKXBqK0FfR8qxoCGlz1pr3iFL7+rElC
rfjWE5nxIUf6rmUX2Br74NPaOcMVNCICH8vBmMq4emwFhbLr6hS+ucP+InIoJnT1
YVjY6m5UV/zgIGT4RvqfqOwXDbGvG3H6f2lzTwmQu34oiwUoWziEtHUbShjezZXh
madCoF1THuYbHqu2psTOzfPn2JstZ42LOjQ3sK6udOPhAFLX0vI4zBnnkGwWLwdj
ZAdglMmHUcfpZ/WPFzoFftvrFhRhMJnfdTubJdvaXxLdpdKqKjTeLIjV8520vEHD
aIWGXQweHc7gzY9BmESMdt2sJwIeUtJXjNT85jrNogQkR1hb35cWpQQcU48pKW3X
PRAxGgL0+z6MuO3b02Thwv71Ej4Pxm4S+fL3cN/zSkApscEDbXH13bWs8yscCJtp
IcXhWP8CIPze9B2Wpt5ZbEQZWgU4z6Z7cR++Lx4jIlkvNOhPNj9rE3cM35yLNsca
klwuCaNyTOuvSlTJ6O0J2MCo6bnAGzh0MsjS1R797/aM2hNazI/CVSJaCoHWtAQq
8iJclwDL/Ps9cjQpSeFumvuohFU2TrcrspXherZoxilmHtXIiWbtxGcpiUYnRw0z
LozSFqGCpV63td1eLCDuzWwKqw36QM//3yS0i5yj5xOtaDsbpxX4BwGTTBrzshU5
sG2KAUJHCiDpoD5bAo82zRS9ClHHps5/R+rOTmvduurMDjF7+ars34SdU+y2ny+5
gSU3x12001Lkpul7d/CYgz+p/KCSKJSVOr74O6rRYa1cULnnuujfHNkcCI26XD/U
+/Xi7sjTY9zWI6jYk4GNGMqLgvhBGnSZkyC2n/cbEvNc+aMxyZo0OWxvtTZSob7y
tQjdg+TZ0SCIAVr3Vz/wv+8JpM1PARHxuUXUgVEz4f7f5/G0Yb6yo3hB4fMOYAAA
MdK6s0MDUjworibuhmsKZXLTPSHXK6updM3rlfW8JJTEzfpzBQXeRAlmZgBy8Lpr
01JMZ64kU7+Xtc55WpzB+kK4UnOqRdFy5PA+KZ03y8jydubOM4jMRUQAvlYPk2wr
3IfOBhVL94aAhdbvANnIwBFdbm8KBoj1GPqeF893g8bQU8TUer3wpaoVT5U9VYfM
h1gYCJuKM6SdSV4OE5DbbP7mSF64U9lajkq6spL2CjxmKByRWmnEGwzsUatI/Ybi
YUK19iOgDU8rBCytbplfS9HpHa0O3Y3ZWx6LomkfanmYTiiY3UfCnjAqFKIkWYMc
XISxuNv/0n41JE4V5rgxnukltlZNdrp90DrXNhL04w3kh4nwSwPhpAD6A/nu/zx+
cSibjSFU+W0EFbjSxldZXwCQ8hu3XqKPGvp3TGXelsEsN/nxGvPkx9maKXTtIyt4
P+lunnEl4/GwaSaPSfZxMqTeDIdmo5cOU9ChFyvceO0GsDm6eWSdukWW9JQ7bLCR
I9lQUZlvMPPSuGw1fiK+jeBok0483SRYhVYtVzW9LDmFml1NFceKFMa3yzHYp2dH
lCcI4Vq6N/L3u+yJLAC7UXtM5pmZFTH28cuCCEjj9GrI+SK22bO2bdLZb2A2gwMN
oMZbuMGzCF8Oo8wYJP6O7Ep4obImtTHRQ9PP5cUnrghxdoErDl1L4pFcu141mEWq
2rf8Rz+E5AVDlCPWTvlvceTACUhXstJ0hKBFOsYJxMd2+8Ny1f6MOcgCNNe/AW87
zguUNVdXMPGVRzc8iHJjyikL7IhSP1Rve3nofRU1CAylCmsL2DSf/RZId/0ez0Z6
L7Aoc6YTVf1AmHKjk+EfWFuQOsZ50nkgMJ6mKl6CT9QlTVtgxP5LVIsAqBnXmp5Q
YTDkrgywZBLF1PzCz647q/Aq1IWU8Q1h+c4fKcN0icXvs9beOI/ksYb0YZzVUT2U
1BBQqsxBqIwyZhnzGAedeYAh59RDZX0IIj6Yt1K5shAKmEjA7qB6GnUDuMcSQZ4L
lSbEGYVcIZ0Sy46M+F116BSmcOkL99/yblqzR8t3GfHGifFSjG4loxv01aEVsCcS
cpelZhfwggMd3FIQIoqqxQFOuM6KkwK3dvdpfRvgLx8+ofXVRbHbOKFNuBEm68Xo
BDAw0xsBPYrNCcyCnU435cvNZXTDHZcY+27nFnbw60dR48QxwI0Mf6V0zlcjM7OE
QKEnZWBFph3AFJLDr9M9x9WBb8Gyh3LwsFtInZiKhXVmqnHEHybxoJH+QaYCBKJ9
qrgYIcnwnsi8zNgGuVXcEnLSukQ7otgkyPB9cTww3k+1pVq+d/uo3fij5RvFDXTH
3WNyuOxhzIOJaziFYY93RwIoISARHiZhlI9gLqkN8wzshx02YpZm3Nbm9DOqsUWV
OoHTb52ppnqBDCZvFU4qcu43buPJNCFNiKrct8aLm4qgTHDD6wqG7AeKf2KcIHud
MPUuqi+cJOg8yBCdDJPT/n5ygBRX62lWjuO8lE22MaXK4Uy4Bpe4Z0tKsFJR4reb
p72Fab9AsBIZV/p+vAYLYVkt4A1gquyTLgRWoVIGgkUzjW3o3J1pGp27Ei//0aBp
sZbKuyQOWEWp9ZVw1Mah5MMzUQpQK1a0rWwLHglACFyCDEiN1f7FRiRSUJt8X8BZ
q1Y0hjeCZKut1wtmeIsa6NyAx061UkmYWTwmsPF4f6ipB1F7vnQ04bZfNASbccmN
JgOCG6VLM8ah3mm7+vWYWPyy3gonJBR2AfAe3CU07r359pAZ5DE75K2+lk1l2C4u
Vx0B/rfFoG71UZSFtbzmIk05YazPULGR06b2Wl7IgkPDlFWOQ50Pz/zZCi7GM3Iz
sCQTJEbEz1CQ3BgEcUHLOKBySic32dcDYfwT/BS3ITFkV2s3EiZ9bTbEZGlCOcoy
VVl3CRUrPbwfSzNpGq5gRZLcEmjyjmPBMW15o6bs//N3qVZ8rCXI8gC/450jhM/i
END4Stf08uNyiaGu+e5PlxG7o/PMgV3ejVWW2jmtrsLY0oKgVrnheUzr32Jh3yLW
9yGuqZSrhzImztNQVcWZqOoLK8FPJEpgiG7Mqvlrrr84DnHwYu5BsO9kyfAHA9kJ
YQhdxVz1U4YtJ20Ju+I1i9xRoumcW4sKQQlNOIbQcJx2k+7SbH9IIku5rxBdzDu9
jTKggccqDmJoTHzBPmv5oXOEf4la/O159YUkhGYaT4Ref4cLzJuteFc7A0WVNisz
S1jjNauQj+HPfRDBSJM0FpWYAhjeQd9i4Bf59BBWGktIHv4uz+N6OMPEmsP27u6v
01xYW3umLmD55tq8I7VTvaesbDUO1ipQFBAwInRDTdbwV4DjElzCJYET7QuMRZRQ
Ep8A0mWib2t+mTE5SLF9akkym2WUKCaGadEYwUNKRbqqc1GoxbhnTFgyvrGRKDT7
/Jcdgy89VUZVR9PzNqIriXJt1LmE5lu3PSmTE56jnicK2enbFrkr2ahDpOdE+9Dg
1geeoV+dP7+E9hAg4Vj8JifuzrJMkaUuyztDs3RrBXx67qHzssKt/5NdngJAKhzZ
cYQKEXYFB8UfnmUn32PUBIIRLaNitFxeI3sojILFDAuiZyucupOqwnLmKWema/hq
LmqEv1xosHH2bVVGtO93VT7c1pTkT8tFqU13S9EOMHBcB0IcbCzx2ecG6ZlfJ2Xt
ryDnKAflvKbSXEHd6pdDbpRfRG5n3PQl76Vm/YZwyUemKMFDwG7PKZqijqZ78psa
vqLYsxbE6/MkiEtCmsaobHIXp4bV64gv5eZ80M21PxVMNKZdqI1fJ9ENUB5VMCvF
+x26cB0H7+cwyCSm3n/zbUUnhBPCFfa5DZU+qHs2/rtpaMK4YpwJPGAxUCTLN1gQ
gahutkCS6pzVeLcpVqcok7u4sUiITJOih6gLKHkgKsjEVbxLZXsbHTSLn8aUEauO
J0UxGp4VsTtBS9QcUBfQ6zy/UZKFyhJ5IheKnDln5bY4vTD10dzR1r0F/z1n/idL
4PjELpXCgmrzB9aaAmXS2Yfl5MahrXOe7wdQ3dqPKKBMpYZL/eKdTeonRXZkmsuy
FQT93DpjGxH18fsN1q6XFDmWPZUpt+HHQHeBd4m9W4VW0nqg0+Wqhyx6NrFZq/aV
l5JpxI9THPHuw9o8GQ/HbAYiXFOYGTi3lH49vImwDje9ma3No6CektdmfoWndIt1
oB/exLzKibkDsObSkWW5+EQ5G5z6/f2PfwYFAMPC6djn3t4dfCzcSWFUIq2R96FK
F/AVo1t+EQSAEkF3IUXd0PIz6vgbHFCrD+/CBxHryZ4CULWtiuskp/KGORuQu3fc
JTwp5H2RMn0lLOiy6pppW//zcWVK4aaaRbQKc4SOYLxP1A7KoWcxBOtpDoKshqj1
SEnzq0K3XZfaRn34mHQR9Ur+3ePGgPTMcarXqXsX/UqmqunWJRpC79eLGxG7f3AL
l81+Cr6Klwu4kI2f63ecWrqECS+dV0FstBvil59JGxKy9urqir6jckMNj2x6PDCQ
KqEvYWH4838nrukHO/hmDld0+24SXiWK83GMvPU/bAwEHdKGBuDVq6ldkQCo77xd
Xhuqjf1umY1Dl8T0UfgRG7q78M5NuXYA6DXw+2u2QTVjY2oSn+yPkpnrKmzNe6fa
UqkaL/equmG9WEoYYBsATm72+y0y4vgxAqG+IHKO8BKxauZWuRBCBDKuvtyoyQd1
tba625TQUDkB/H07IMYPpeIRVIQfzjeMCLNddO7B7JNjEn9YKj5IvbhHO/c8pWK8
pT6qSmQm5h8i+mXZwxqWYOoBfJlz0qyMAzw90QlhI7yRX/RmSxwq78+Xf+uoJ1Rd
H2m+WjlRFsssW2qm260dRkaYBEYt+3uImr9Dzb2oKsalUQJQ1nfVfsgZkPYZ8OFA
EoA51aq4f5Z2UCb+KytEfzd+X4uq7Wu/uqsgMrMz+fIvg9BYX320mjdZDT30iMMc
0tpLPoyso7KRSV2giodtYaI0804sfU8d4gkeF6cHNG/6OACJAqskieaOXx+WXC5x
Ja0qF50hJKuvMG6IS1a0ooVuJDGVLSiNHZo8y8xf4a5wT04Rw4CT5U/yFmBSG3n+
cFqga+kyeZBM3BlBEjtLs5qK7HK9w8t3WrRpNvir92Z4dTm2hMWwWS8ufGFONJw7
7KpqYVisPYDKAOt7hqZjtm1cJi6Ep31O2JJGp3XdJ+1xmpBs5EdqnfuJuYiuZbSP
w5yz51pRmUc0kVFmkHLULQaLiU6ES1CnjpVsqBcLXjHiw5BG7LUmM94mEGRkDEPy
CVF/hNL7oOsfPdaghOe5NGrss9r29q/JrzVBTNMfrQ3g0FQRhbjXREuMdlyPsWAS
Caw7XpDkjrZnbZjWf/gl9IhidXIH+SefilG4XM7V7vHWPDcbqwENGL7eL14auw8h
W+cxo9W1BmMRpomeykSMK5xxpEVaffRcUB+or0dHxICxf5Q8JcKW6Vu3GAezWPr+
WdVqYZntEv/MqoQ7K+YXHef6a7kUy+tBktM8pE2yTZmcDR4lINJKMTAG0sBVOM4k
KAltqJQrMYz7MP2LMoJQMBS3Gd+UlDXfrgZx0z3F1jlqA14sLER2rSQSvPfjAV0e
snzyYRa42DgsxQEbWImGG8tJrAsgQve6sJMa0pAy6+/2D+L9GbIuxybTbcwMeAdU
z8c/Yrl8popZFU2tEkfc8j3Boa4rjQEwhKkEf8fiQ9zAXp/0gF5YAQcK2OJAGni+
Ohp1ez8xKT6snESGynVUPvLVo6iihaD4Mzuzyq0eMKOmuUAjl6SmMQxtUkkaKSFi
+0224JhCNmZ2SOI2ex+oE7oUeuo3ToMRsAXyXxPSL8yzx1QRjmWa0H5TPmiKQJX0
SNByxgCnKVo65kBwOnwPlXKBG4YM+MHIWEJlaGdmFTeP/L+aosVmUyU+ND5/w54Q
dRjT4O7jAbG35ZpJKvVFGW4veL5cvdpMUl/zsdb/dYt8M+/CLjS7+rvofyp5P/Op
eSa3wS/NTnzh5rBpl7hkg0XlzIEaQuXOi12+QK2lWgle/JWFxWhgYR7DaTDSjLWZ
HIJqx3ub45ZauM4kdo9kaKf9g5LPpDnopxqZhCJYWVhI2Phi7XuXXkFd90jijCH1
iB1a/+SOIeMXIsSQ74HuGlQXAXQWf/tELQvs8xAsL/GA04Idyux+KqA/zOxDhUrL
1Fyqse2PfTZaM+kDm3NOOZhy71s/HSaXIu9gGb/CuE7WDmwYqBrVayI60Wg9qw31
aUVX7JdP/0WlcNbcpAICgpY5LissSrFQq7zF/i8OWinEvBvzs2t7MNhLlvbR7ogf
KMsTl8+Ip/yilkls+hIUioVunGcEIuVIYtSllFr4B8swg2C5ShabHF734J8t32Z9
HCpAM7ldDgD5EQF5dY8KI4NCmXuBEc3quyh7rBZtCy2O6E56kEaX1Y8Yw5E/OlSG
cBkFwf+CbgoSFMlK5kdE1Nio0Q4VNixligWSRw8wk0unRrGQ4gTZ2x6FB5XmtHzX
dCE9hO9xfcb1PPzsYhFIaDwZ65o5QvvS/USt28ZoXIl63fr/lj7rswLFPvcUN4lg
FshmOmpsF3kH5DBDZ+8aKo3EtqcnsOxRyJRNjUTqgTyzrHoW2+4Za0Hh1T70hZbK
MYiUaBSARSdIkraLS2Hs4b4/Jjf5Rk0AHdKszJOKMyw48cxdsNo+rcMFcLdd2aj+
hPEwuaJxofT4coMQNvKZiYg45PQ0MiHVcFWJyW4TqMDQdKdsLj+iUpNA4fRfP29G
ZVDKxdsMa9fud3/sx7WqV+3Mkxqk5JTszKsqgpK23GRbYcWYWphrVFusNj+JhrXs
tx1Km2/EKdCciV9rrpg+WgG/pphGOZisqzT+Eg1X2avX2r99Mu33ZO1Yds12hZ5X
sAPyYjOOxt1pTAjhfdPc4tICFfAp3gyre/RFJebbdAURRscorZypuQs+Y5uHqa8y
yqwtwvCqCESBpJIvgeMmRHUjzIt/HlW1+9kwpQZlwB3aozh73taUwTSicBOs50UN
ZHa8nHDWmQPjP2gI78mc7AKSEPdrfF+9n5W8XmFRrZN9emrcmXIC5Sb08HaZm/eI
1tzhOgJuzgi2Mcr4/npX549xC9pM51rEYxbltUEf0MXiDjbER1MZHCT5kdAjnU3T
uI/F2wFpNZ83f5axQI0a8IVmiLtR0KPF7u9e+JhxQFmDrgzgLr05pMPsvy5FXF8O
eHWAntfcmTEcN0urI3m/wQHw+OwdnEO7t/oQiaA7Jewq63hogp7NtbdOZgPdLzFz
pzNsKvAZsO2gvMGwhVn2HdyJjXPLPXxqqTxlkLOb0DYt7s1ZKPL/ivA06SYOVw95
LARVo+fQnjtKgzCq1gHD5RX//eS6K/FvrUn6Jz7xrHoRpM5n+ggkJo8SDiQ/6uCi
//dJeE1c7IO9iky9mCsDmSiLW1c0ulSMX5mUbrlzqH5pQM5vQ0uev/BT4Tn0RF5G
6v/rv/y9hSMGZSy/YmynuNnKgavop/ELYKROQkcaMFsDgdA6exHIlCUqk1wtlNfF
hqy4j8lRnxPp0r8sqYHhzYdHN6a++BclZR7AWAoeoQ623NYtvcA1vxBkTws+hNKo
+9htPpXHMOiioMVv6okqNdJJ426uO5tn/gTaplor7+fayxRzEad/lqvhGeu4e9EY
I58yEYcUXxYWGdW8dRC7FqiJoS+MZ6hOEZIg3RdWziM=
`protect END_PROTECTED
