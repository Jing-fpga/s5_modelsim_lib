`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y8+rGb2B2kG8eqaMSc0nAKqBe//7NQL1nL/2JIDRBl20FCo87C94oLRvAaITC7zE
ddw6fKr8OJGNl+denEu+m0oh7iZ4e5JDeLS4rOY0iiUmE97l9a/u+hYMxn3r1OeD
Nw6acdrKWv2VR4/Uapz7eE2WiPo07UVfX/Sqwd8oFn/cJy7bd4ua5k5TCkxe12b4
uakGkiiYKAvQ1yS+L1Cudv2T9PxeUdOF+75f47X/3eCUlHx3IfHCOuM3MK9S/G5P
GW0AumWghSuAHyoqeYZWcpWyBZ3O4uSf/phYMNqg2uugGcvFZMOOXMKki/Un57dC
cavS81l5flC1r4wXw2PW5vnoPbbDDIoN8pHWBepoyziWCVxSsobDWT+DlBjzFxjm
QT6ae05SlYqHNeS2dA/dIowVlpi1lVW08HLfA86o5iaoAii8WjCppRE/Dz/B4Bjc
Jk3xVmJDCbKPc2mN5+ONjas/Ek89nM8/gMlT0O9n1bdAOZIMo4DTx5j8xSejSzZM
9Ba0L6at/8Nf1TL+Ixq7J7oZxhaDpaC5WTGf3ncO4831jblJy/Ggk334HRDyCR8+
aqpVQww7HsxkaZBFeGtX+zsy2jfjrtjMe/EtaZkjc2Augj8QP445tzrebYJ88QVP
K4Nc0WGwGqfqp2yLf3Fp+ILkh8kPYK1rVoWBaBiDYCXfxnuIaJAJV6sESBfdWrvH
mMPbCjkBR/jIkRVSWZ6OjhEAxCs6u0cxpVT9SCBpyNRJcnxiAPxZ++dsi16y1Hu4
2LwJK4M16jtXeRqWJA2ltt3k/JzROOgcjQ+on/znXgOoy1Sw6grUUcmLRGamSbN6
r/6dk0iUgrzrbQMOmU9fMoJdVYf8CtT2Br6v6z5xc5UaopTMZmHwvjSPQqbpZjSQ
m70YlQxdQeVK++6K6VSdfBs5QJorblnQwyIOUrr1/IiieW9Ey0pBV6zPCkbZ3cKV
q0LLkrCt+Qc+sMSvt7yD+EyDOIx+zfPN84v5dgew/xf1Q57N0JBXI93Y9WCW+WD+
LnltaO+mZw05Jhr4W4koFh3ZXifumjIvsDzk7CQ7ChZz/3i6VKiON+WE0bhX22VU
X2GsHof3lXv4fHXker12fjH5dCDcvdkVSYGyQIjvb9QYRmCrpnjXEoFefhkr6Wj8
uC6iQMse2kZQMDjUtRGHiw==
`protect END_PROTECTED
