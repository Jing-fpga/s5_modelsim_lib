`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8/zGb2SsFUaRwXclV1LGunb0oFc/+Kl4J736zbAywH8AZYWnDtV6aC8I+91dGWjG
xA+rsvNVQbdjQavxcvwtCZEoVWe9qstNppQBnKYSzUJv7mUyTCYgqO7LQ0nd1F+r
bzz/1E1WjeO52IrFMuK2C/Sdvx3U4hTd9oIzfi7dg2G5DLmyUVnb+BV10WTFlytO
08YEiC0ozKIDN/3FZfca/rdi9Vak9ySgH4cO2rKfp9V/+ZliSlCxjVcimYb+ROed
MoMYZZadBTFqvKajYMuBi0CsAOeW2zR1ZyOYALsRuPh4X+RQ+tnG+BvzvH3y/0s9
vBKfcZpD9fyMFmHEkEmRjCWiNwnJpWLnrFceOfbgBk1OPAThtquMQFUclL5S8Wt0
rCRHYKsUZndn3xwrVWdEOcEPmXkJ598iEIwyqa7BJFZaKQq5u4KDsFB9q8ENuMdf
sCFgCgV8QhE2p0VnwCoXNTXEKCk+KkAyWkna/fn1oqx0OqIMI3N+caciXz1bPsqb
zZ+/VNYkHcdQ/NBrx4Ejx95k7Dipm51zu+1jGQcX4um689jD2lwjgC5+HPCpmyoV
7YmmzTpBCl6tBnyWbkBCfM7twZsAh1fpE9nV7i9eYltI+2lfOfUOwJfGal7TuQ9t
Q3gTQuzmyy/K2/7zY7SJGpFyzdP7iAuf3om7jaaCtE3s2tvI8juvqGxP9XvHuaBw
z0a9XJNsXU9E9QPNzqPHGkzNwyDc36032Q9HCDqE9m6cvfeNzF9MN5SgFNOfhs4O
n7bqADiP/pnFW9L1F0UgaNtzeOYsTQm5nd9os48DqWHNvPbM2+0Epf4UgTveDoDs
yLVKrhYEjLykuFCw33cF2g/h260/N1tlaoubuTTALeL2wBoPe7rWXpbDKibwlNF/
KqW9kVbs4EwOKG5sugE4IZHhTK09XXLHwTWmLzVko9qDyDeo9tzsSgmmWHH5HMs/
JFQuypIMn2OH7AXmW2c2Z6sj3pBo2ECBd9wIuJLneF1nyM+/FsPQrBCLH+IsO42F
voLUMjjxVAL5SW5/ZD2EBLdjZPgcadM9964hYKy5JasQVZ3SuN9mInowWj58baRD
Zi6k/7yRDrUQ+ea+q8xi0Z1Ds8/xk4NdHMQ1V9ZJp/4GfYkmvTj3ObvON7m90+Ba
EKaIbO/ILeUVOoKkAPIjlefz0TtS/4q3Fy6H5f8L//J0LAoP3TS8gW/zK0L4/Ng9
i8+y1MvlDRBUzc3xD5vGpNMYmHKERwPOzv/WFct4d0EMccncnoFSh80Im5pOucKR
12Z/bAptxJAXeLeVcbLXTAKmxx+JIOkUUBZN4gh8p0jSOg3eolGB6WIn9BWaL7Fa
aZvXzGI7uJLvZOK0YY4gxuEogp+7fQmMkWQCl/tqE4xfxEr4CzmMF8El8LyQBU98
te9eY5itboOQGlrh8I3RIrYSHI3Y9MMO2BjkTDTBkckrGZt+Jqbzl/8p/g1W4/N+
hSU4WMiem4/yRsCJ4OzsIJCnDAIw7mUl0KnlCQcnI0ZdzbIq+ZmnEPEWSYHcurdo
NHNkeexOSm0AGYvEu59gSn7C+nc4HNUTr2z/NzJYZKZSA+aQhHc05wUv0Juco3s+
6y+R1wMabyuX7O7WmjYV+C5njUi59qzVGmcQRykRtfKy5AS2hGgkUSCtPXtMInHU
qf6xqh/cfmhIo2HvRnmbQ2gAs3YyUzSPilAjER3UZYo8uy0AUjuWEUKM9LlB3nzn
OXSrheVpM4Ks6i9N6xSmpR4fsscR+pk1oSf0Q46LEM52Z0FJy10R7PckCNmpWJBr
tm+JOjzV2MZh+4YQCCrK4LsA1/1CeaFiI9VRJMBKGijZVARWf2xv7TgcpouhR3ZB
SoPgOoemu2s2QnrTjXPpj4sKTL/84k5AgCaFxqTD404szQbwRDDR4A85nPOLyXHm
z2EECLfDYSxMNwZfZCnjFtauqDXBU3uRsJu76BfesbCcCTKrjvl63l7e5XDo+h3R
ce+tzOPFz21uq7WEYVA/F0IKfkXq5CQ/JOIQnSBF9OPvmDK1eaS2nFifNW+GeiRk
gKyZoVIuXqwDLArkMUKo9wirhMhN9D3n6VYEHJbrYPBjRrixMlkj1DdPbLJvQNJc
p87y+ZjXiHum0mSFkn4HYuiD6XyksYLbrbIp+2Wef5iQIxnpvgLKbfjoY0m2b8vn
da8inteAaxFzOtbhxPA2S3jzcZgiWSjCdDOfF0PNxnxBjgSPg1iO80yP8d8dX07V
J7HzAL2eRZjfQ0wiKCR+pR7aGvzFQN4CS6il5iyiECc=
`protect END_PROTECTED
