`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PaXHyXWFOwNhjOw+zlNBNQeCpeq4omHOrhziVXk/806ZEbD+Fzb7R1RxliYTCnDt
fW6etjYZgq+3yNS3/BGdPbHsXsSAuoM6kypa/SoDb/ENTyYttvZmMp2Muh5iEDmM
SLbCvSABPpWx2htsi1DsAxB1O6NKn+QGn+X4+zf7JZzcEKX8+RSWHDw+KP532H1+
B1ZJGMAr74NxKQvpTXYNvAjmg1Fbdl60z/PIUmVCqclSUR6r9IIuMsjrsK00WQU5
YE0TtYz3/7y9lu3qFSREzeKyW2B9Z0RqhF4MfPTrV9idRKYajcrbufMns1gsiB5+
Z+TDXdXNNSpVXdaeXmPS2ZKJhUCPfMvCUcWP2PNRVE1lmOE62X8f7GAvUOOfWHSp
pmCPphkbEzKdKHl4x7/5AsBLyG0iiyGZT0E6BoV5fcJDvFJHT88C7en1NtS3hK2u
Ugezcp+ofpk5afccCIatuM+fqLuqYImvYi0bzGYJ8NsSBMuhlmbJmAUdzODmAUrY
4bFah5+PbTkXmj9kFIYovYA2Ia1EqjVbhGayW/MJeOY6zNhl2DhiIVP/0JlDec/u
+PFzFDRvFBfcPYdn6DLhUnM2CcRUToHZeDIjs6Mq353w9wyhu0ydU9CQ93fp2kVx
JkLbHQ49ZH9bsIzk4CWe9Et2Gej7SZZC1S78U2Lg0f/YwndSAb7xJJ1hzD0N4q/Z
MMmDFwKfvQ0/+nWX1IkMc6zMIClwrsMdbfPnFee/EzfY65k1SSGJyitPpC2U75NN
z4vU3KWH/qouGOdIoGl4MTzEdwLTjXyIp9J559NO9my/+jEfXBL+LN7IgKJbVVuc
hPjQC1Q9AlgVJXJdO722vXXAraWwu6GeKHYJpcP/VnksdCvCyHd+V3YOzkQbEeIx
2F6tVUyAIvUigBS6OqNjfx9R1C3FZ8Dy3IDCi3Kk3MlS1Qvad5ykQWBqljWAMFUV
ZcsKCoUPIYzI6HZwrN5nuqCY+8ukPzzoYI2xu3AwENTeAVwYQtrJPXlRB1mwWvAm
4x/FDgL0z47gRoLw94//sWZyxUFbrKNl00hPYo4BM83j1hzUbIaCHcBF9oL149br
yAoegbI8WVuUaSkefL2kH1aCy51pJYkXlxH9bLSF/DMcALZcaL9QWBPtj/RZGP7q
PZADAujX8L/ZJMrtsd4Q+BsyO200qfME82Vs2vWtGSEF4WRG/ajM0+Ny/1wGbMH2
PLrCZITXjZKK+90qJHI7mOo9GD34D7qDDRLwuHHWw7YYh2HFeft59x0Kj1n9iPnh
SnQDdihgorSLNxL+EofPhIpVhxEKVHlyBeuw01Qe5zsPEnI7nQZhKEYvDb7Ki0ID
CLAFSCbKf4VocwS9QinSneAvfSF7Vadoov1Ej61tuv4vP5QSn3SE266oha0WoL9u
OctwJg+inr5j9DEB7T8aCY0KDMukkvUdPQrRGQMSIhLvILy/QWLzlMwSfXd+erEh
/keTYP5rNehtWDlhoWJ9NZKTOIkIBUTIGwwVsmiXx/anmnHe2RFh5pU2B2ZnEIZy
k9UwPjWHF+fAsNG7EtaR3tTQOwX932hdQPFi1VE54/1ktUaeQdRNVZEywNINH5m3
VKV9mNpnowAlGARmY4iZmBMVaAu/rG815EsrCi9zRxo01QV+V5xnXuhmsyrpLUeq
QJ5+BtEYsAR60Svjf33xzIrtxyLTN0mIIn141mibQCVLkOmJXakBgCzZA8jLNO5l
WSJkxY9YzlNgkGKMuC886GJlfJU4mA+FoafKc97nKgb0UuTMAo5qGQr0KZgt7Qg8
/KsAB2ZlHyfznaYRiBaIR+EjrE3v5gwl938mxSOYuYAJAurVgEC5q5Rn1B3pm4yd
9fDY8XJd9QI61n3QVv1ODgMNXkqvpYIXUb3rdYELckxbj4tNPLKICR4XxZ+wlQgw
4x2XPx3LBrNykr4vX6uH+ch6LpbEbGzHWI6IIFW+0dPNQ2nVBMXLebNvLFiG3uf5
vQO4AoLx4v32TArEtSpxvNCml8UWUrrCbgrSc5nMxFpxaWdiYufPIiZJ1Pd4GPbW
R6qAn/O2pCPLnsGtb9LwoilKvKn1ojRZZt+b8RMwajZtFPRtm2tFTsG7vc33NMnf
W1YTpjESWPFIjVwlUzwgeOaW34WMXdaIBK+BqS3dIvEjLibf6KUlXpj43TaVjPzz
8aMRHOQRJHDPmE+DmGbgHTElvRMMva81MIhkKqeHPI98Ju1BuUYxpy/jBIq45oq6
SQ1phwQddmqQEFPqux+kEzNZtGhZVrqyPF3nX/emaGY=
`protect END_PROTECTED
