`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xdYqq3ojXpozbnL1JCBx27gxNYxdIpxSezK77TkuIeTHV3kTMCA3IRmsvk6raEEc
HAioPacqpQ+J8aCi17O0o6t7VJI2iWcsjDYHFK84zZqx9QI2YIkVN5GCdJhtCmop
bCHvXdpr81u2+JJmnhTiACB1AGgBIAQtTDBmhZeSNp6rLRGwl1r/3P1SzcoETNsT
yq3zHtg6rkcMDX/35wFWuyPHHBs2CyiKHz3i946CZzUd/9GT7DMXrhrmNmaMjRwk
WYECW3e4QArge8bQMp2Cglupko2T1vI70i/kMh25aRkXVyq5jfoyDnVxzF+Lf7fL
8DQqkSCSH9SNKl1IWxyGgsmN1O7p0so7moLq8amy2z53lQw9RmUU5stCROCqn8yP
ks4Xxt9XQzw3KHWZqUe5qXoUbO8oFxMx+SYYCg/FdMetumP/xbVaubaYttSoqQJh
CVoteISzN0RWI/nPSaze3Sg5d0Jdsm4/cgSTbyOiyV8+sIo1+3qBW4aG2vX7eIRZ
PpDSjHtk18ZGIJYaI+P4nEj6iPfJjPclhWbxlAYbpYfAwpcH+QCvbu4LizFZJ55f
8I/FUhbiataJg7xSj34sL8lmSy+YBrE4B6ZX/tZrIv7P7sqQfn05kTZhBUKAfUPn
aJ6JtsK9Ypr1XG+PVAPsV6bnvvnwOZZ6Ll0uf95yi6oS9KgcoGgpb3+W6BcCcPxT
GFbYw+DCNGPuQKQ8BL5yoNlqidTPJCRUxQI4K5thSWCdqzd+4bfKlKPlmHLK+Bwr
VPGYzEf8ZJ1RwWh0iUwAUw4sqkYQ/xG36kYUsuRvagWez6946yRKsq53X71jV6dW
c0HNjhbjSTVkAJnlEAUU6Y1Hn5vFjWS6jvd1M04wv+TpY4a+BN8fYPM+37Y7WsR0
A48qX+7kLa6AB51FRHySBMbbPCn5UI5UmGABnv65CN5RAxXGdDjb8/XiHX5SeB+7
anla43OEYI0EKKkJewlWNO4+l7fOxB0MAgSr786LL+iMBtQR9d6A4+QqMuUt2FMD
JkriMxZRxTOVUVByQEAYYYvdaMEzTTp+D41XJbVF1FpO1a/WocSl2NOpuB+kH6cd
U1/dj0io110oMsNvxJoLFJR1Ti2SpNwRLbCPblRiITgFXpFycAhhB3E5lxBujnpW
0umtv37OB7NCLUu3D/STltrD9qH4vgI9haNNYEilW4iGkdVvJevXJ2XRmcjMWR5u
0QLHomvGuHmrIwgsj/nGr8VF1lHbLGE9vOqHEoZbunlAESV8drexKwZee5+xk01Z
ELkQOs/0midSwbk3q4+zEvl8dKmLzvH/ClMNiqAJxT4j5RMbB+QA0hX4d8C9qdVW
njBdfjL1vgSRcQPOe+6VoG9z3OR8LUVidYlvBTYawCNH+vzoFnFTnqZpa5aA3ZQc
jthYYM0ZQrbfpSnhRehvEf9jZt/TcTPCRN2QWQX0+p5yr/S2hxoGsYc/JCbdywrB
azSdIO6zaFo+HPq64O++w+5vFgzFcD/Oe0/f9gvoxzHw0MLhUJrZ2z0ojxDBFUJ+
Ud/TwlPv+MrD7DzLfShmvn8IaWUqrqxRtoUFefvnM9r33e3pXcw/0Ox2U+W5M77V
OwjkGIYXRU32b3vtmlLKbSoncIufCDFbujIBs/20kjKM9pssts5MGyWBFhETM0yF
NzqZ30c3g3/VMSbwEHidQL76vfgmaj30xdZlYXsFfOr5v6ng+vGWp6NNNlUgUjpe
L1T8tK4i/ExbSFcprT0CFjbwm53pXXkFRqe4KxL1ew1w6qOB1fgHQzDxUS2Q1MB/
d98+XnEN8lEIWDWfmE0Dzth0cv66oqPdoHJ+vOz8XNs1L+PuC2Jc601ytZrngyRP
SC80lMyYqX7i+8jOKy0G6dLKExoisZspo6IqDDnnufM7Tec2hviL7XPtWU+z5Rbk
0nBU6e+xtVhoAu9G/T++F4LgAAQjnoZ9hCVtvc+S4eCibLyCKlWQD70oHC7jyEzC
RSSPuLPWt/mWUhD+gfCeKHO/PMbSGL01kJpiznne6O/dB/Hd9Y1pzW+f3GslJ5aV
D322kyiWY/IIYP8Fo+ezIx5mQv1oroaAKmdbAejFIv1gG5VvB6P9IZsppfvUS1QK
T2rD64i9UiybqmUHIMzYXhynjXov9TIjHi/dMitfY5iPKlkHMPVjs5fqL6gpSGqU
R7XJOv1rXSreH4d1laE4nAoGUEryPQYptmmc4dL/21w7Lee9PS/eVe6KVKXaEG2U
znuGjh5PxF3cUjfWrA9g8DIL9E+FWQzedGTszCdnoeaZ7rfWchZtqnt1fKakkl9e
XyNA/zacA0ZngqGKY72GXQ8qHvzubh47khi1ihgtlF0=
`protect END_PROTECTED
