`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tWaRpplXzlAg2dOxU45bc47oBilM0fMrwWEGPiStukcOIHm86nn2/gpPxklnS0+W
CqRPRx4lZcCThQspihZAR/IfIonQajqlq74NatjzSzv+FgZLpHm/pVgkJUOPjnyc
vsYwFSD8OOeg5TgrN8Qx4dGJROAXrfMf9GDfY0SLOps0fMWW1fkYNLndsQbjxPb2
tcOIdo9Uo/XnOcQcicyyhwthpPEPMLsxJ8ueZDV2M5Sknv5GI8fIoAZGa7P9S1Uo
HaqN2G73VPOF3z+gMOqIrbYS1KopiDwOVUzP968+gdXCFEVBINf6R74PpVKibcCz
DNPHpUHj0LL+98N41l6jtm9oBnmAQNObnQ9YSWhlysNv0ke2tvE/9fRRuwOK9ZF+
mQJEC6ty3DIlEqXiCSyg9RgdiuFOFgJq8nPLbJSqkAFGfa9ck5yv9rDWGAN2xa4v
tIVNcotnjkfWh/k7A+kOe7Wml7WPXi5EibYusUE0Uk+/Je79eFWLA8dqxPo34G6J
ihGV+mHprGj8T79DpKXGElMnvD/3ljpJWxKpFbHBHqTbAEya3wUBf9s26sfH/LVi
UC+MHbKlptdMNJZKsvWR01Za2YfFHHPkRCBNu/FlxeSMIYxHGxp6JubYWPkQ1nVL
KwTX53LUzIZpXB0wz01IOVujxjyYC43WM3fh/7J5fhubEek/nK4XkE3D2/NzEhjv
+uZTux5G9+eRBsiH/4dAG2xJIqQyj4/vnvlAs/DOb7T0IPijVhBWfD/r5od59jue
bFIHjJclbR1jAhEnHl39n6AwhYm9db0fY2LW7CsZux/3tjEBM082sjm54g/0y6NG
rHDph+XSiYs60VSqpg1oyCfgjpciN3YSrxs5BX3/7v/5hF6Lm+xRZxCf1XqnW7GX
CMA8fcb5GTNsXsVvvx0rJ/3D1foAAUfuFSgE7XoasRRzXTop5XimUcS4XXiIQ1KP
3lghF3zveKxk+f7xApIKiZuSsq2m3PzTy5uaUyOKeJwv+DALmZqTUyF9Nxa4JR1e
MlBgBA9ojsNpuk4+Fiiu62dDiZQv4YyHLqUUfe+2d9v7JQAae2y9LP2A+5GODRpZ
pEM1GpJKCZcrkkWn/ZS4DuNXB2wr2qChWQ7y3usgOe6tU4P8vAEixIxz0oz8sqWk
yMbrs7dNdH+kJWrWeGAGZP74dhCOrV9ucgzmrDKvPCtgI9MA1CESsoU8Wl1BNagx
wDBfnTIdPwWjQyXQYGBNwYJ3wNw66fQxjsJqA2Rt9WxSwgQEIiIBGB7PJxVxjFWs
gYN9VknI30ljkjcDivbpSJideTgFDVEGjDLYama1EfIoZhDzc90qEj3IWptNMp7v
XRIBGsesD8+jtKlkimY3kCPuaC9yRlzuAi/c5NdIE0veTtWqWgU0oOcaddJQ88lZ
u8MnurzsvVLAYeFtGyW4WVXYx9cY4iQSsvU0DD2nHxwhQO+VPD/d572+qPTMdqSK
gXLbg5PO147gseaw6rH3fFjMAV3w+9oB1NeEcxX/PfgJazIgBvYMizADlBZdc6/v
bqwjcc9re8kEtNgRag08/CCC7mUSYbSbPRMKcq83Rg6dVrGgPpnHWK/P2pJThVpV
dMxU07nmztXUh6rM7sCn5rOznSZfsfAT38OhBdwfPg06+TLxfiHvWbtrdjabTxkd
/GFkLOLO3I5XGiM0OqtTUSp66NXEnvdP374sRt0QVLjRD5CPD4djd7Fr7h5asgkd
zxmQfkOANglzk4UpkXRBBT8q7CElYwmBygEPYLhin4kXvU3+D320YAg6emi4R9mq
ekiOXEmZmo7nyCoCWtgFkRCRwKfr0m761+qfvlW9+9EObXtUt3W9smGHopM4ZunS
ar3HlWmmZgalxXSXA3D7/fon8Z1CpkC4Caoz3w8HtuRd1w4zSui1lfgjnsqSZltL
TELNMYkpo/O2g0xTymEA0IySXrvzd5eKfdPOIcG/0XBqSUKZ21zxcU7sOdMBUYLb
4qsGioFRHNQz9ovdQo2CySTGUSCwGsYWHvvI+6fFQfy9ztvC9RjZfuk7KZhWWKKM
3pZ0eHHu4atbg7e2iOtS37DBLi1ovZ3YwKGCjRjN9ZbuMErmcOasK8upyeLMH2Rc
bjYJcZAFGyP9KP2R/0MB/h7iYX9cPWHcvUTGw0wuxWEgsIxOGea1vUSrTYbJ2w1B
vqCOYuNPEXs5+NIankzCLx2KPkPtjwjwO+TsEAIBnITlqaD3hP7gXK0FsqvewYNB
x3BNhxKJDb0R6zxUqD3fsSrD6YIqvBQ507DV4gixWzGoSOD9us9SdbfQwRel/OsY
NphtW8XF98zJfkKc/pp+KzJaeemoi0BndcoIqqfAa7zdH1LBu5x9oF07yUHY8HRV
mSnNbLpAROIl9EcopJpTYlOXyeKT/6kvCZuhFeFJyqf1s1anQ5qwGryfBajrxxQd
njn8mgIaokATzPeweRlPZRhHMAX3pk9PmVam7l5xsXWB3ORV2Ixy63bcQd04WYVn
EvYkcYou+43yanhE0gQH2WcHYMCbomfnwxXrt/7BdmkioKhmiTpBkknwjVSsPp6E
8rF59f3f1+tvsR9ryUUczSXwjCCHDljwDHiozVVbkdXpBUFidNJ9HimGG6ae1k7l
kJARqumxeD0CDamFcJMBnvWUrEBUJEghxPcnYYW1f9ZVAxYU5kdXXEGShX3eLS2L
zoVbe0yPEd6Q4Fjt9aBgu9oWeCiCUMmTooI75XTrqYxC30q5+Y7moWlxENkGZj5w
FFMdcMENCsDHyCXf1aBcwXFr6GtwvlzeHVNy5wt2AER/FxY4eos0IeyshuSimeoX
iwQifq3QFhMmjxXbC4YRLmh0qfBtm4ZnuJMsA8IF29FzfRCvDhgnEDdshUWt6rlY
XNDD1pfRc9GMFlzUDebzvaSLcjfbmSG73+3hpDyfIS8yr5sa9sVG9P+Zhfh0uXdA
xS9U0zIWoymv6JP/01wcZRzVJzni7saxAKG4DXF2d40HkjAi4H8AaNNMUWaKVDbe
UbjOl+HMXiPotTMkGc8iEmI6lEJox1VXFlLcR2RTurnxIAMEYJzfVbq1VpS07LBK
gvV7xFLfwqyd+ixPcY01AMOky8DrCcG/Sf1Mf/VD4+ZYiwkJg7yjNXy4T0WzD8hp
WsGWdjVZ59wo9h3ttEIYPPbQTvW5VUS1pU7+n92gNGYE3yXmpnDe3gTrfyWBv6SJ
ljRnqR3iIM6cwXguYSmFGBTH5ku4mpP+Ee+G4FerpMiO6b0PI9T/zO4WC6BinQRW
Lv3ZPMhWj+F4B40xl5R1SzU2LSHyX+BqzF4IBkjrdlGp7n2pSpC3FqvVnJjOSYVw
QnaaHjpprhK/N0mP/nDzJ1FkYdZgmKKZLG7+HSI5MhyhylWW5kCOWop6M3EKt2R0
3pyBjJyfRFn855Jdl8aZpcoMngbP4FAWozWUoUiFuosoivQimHA58TPDmve/fl7q
rPAeC8ys3QlKHGmx1RekQUMoHorlrAQ996y8+DJcWJ0FLtEY/CDDy1DkBO4CcANN
TixLfGVamIeuMj4ytNR+mR+ZiSytTIuPpGOq4n4+59PhA3SEPZ8csuTLdmLTmwgS
yyfFxR+HSOVPRHw2PWx7Q0QB3CAiMAJMny92s56GWoNjV4t6ASyEboD1NXauu1OE
/HSUhCUYaly/RDarbEKfMigG+uMbs58haReZQ9JoZYRp411zsFjo4t517efDlOFO
KSHNr2umgiv3+Nv4/o+Ci8yikKU4w5XxXznIo7It2Aqh33Qy014+TOxuaTPC47Sj
QieXbf7tsW3Y9C3ay9KwQivTgbj2Btc+G4pZ7Q+UE/0FEc7qxzCrR1ITOIDr+Rc0
dEdUphaKSnSEeMoq5ZvZinfWsMGI0o7hh4594PVM5ONSwvYo9l+X4goWM4lztpJY
61qWtZFKAEpVbcpkcyRuC9NPjB92AdqtYuYRIdK55I8yWJfV6CkkzFB6ptyDuG5B
2rgHlq07GciyXTQ1ABvOochqlAqw86BiK1CjAPQH5sVVGXmVFffCeX5cO2JhUFCv
6MuRQEu298q9SVboZGz5dHvjh4J9GKnfxvjoPOtxcFQoGs6cFZ5jER0sAnQXSgDy
M7WY1J2aGqGxAP7QIHAEhMWqnE1QttAJ3LLLYzNPSco9QPBIvWLhl9bGaBGwxodr
iz3/7I7AiozGi1JJESfjmGFrt0z78m4Kn9YzxIyDEZBRuEr1pekSRnfMmljgSUr2
e7MrowR/6eWCRxSUM66zmhPTmNxd/msXGXXnl3ehbJI6zd7pIw5YPCl6ehay2D1A
hNFu6FK0Lma4Kvb44y4Cr00hmZ2h6Xd9T8Gtd374MC6jOVuVr/udLAql9yxsNnhD
whI5VSF7A9A/YpIRYfnfdaLr7VLs5m+zQS5T/oA2hNdw8nC0VAOrYiYYuo/ko1NN
vcbzlt/WqwYoDKgnz9sP2z/4/YNhDcXKAufDZTmPoVLEvk0i6wA34yU0flEbiV4k
cKdbq1WQk12naIkN5DnyIGaY2BMxRIdu4qqpxjgLD0gpyonJAkEU1u6qJf0vY5xS
D+CVLgnDO5RSKr4jVvEMUJfFv7YPeSw9+wK8QJ7p76ZCrZEuB+RU2g55p5EMTkOl
yLA9OpPBrpelBZ0vKfxXR1SXuHz9vQWQyrWqu/bvyQqQJnHjg+3gGECE+qskIxiX
Ch/Iq4J1oUxVz8CgJzyNROLvjBhGsD3yaL3TKySHrysdzGhNg9Jipc21CmaQbtJr
F2ehVkY1an2JHAAR9v3ldULGCtBzazprzLJo5rWQ/uSWv+shWnWlyu3fS7doRsNo
T48KDakPmdbdeHAUL/vcKHtRVDN7bDy5pGMFSUFbkLRq1ms9S5WTyqNnkLtYnPSf
3YzgohIoy+VxEFXg8RjRmr+XNu6tIl8Acap4jt+CMTCsgmHVxZoDFnjtRCddX4KQ
3l7YEFKveM0ji5EuXWI2T8hxwj1ZSj2cJsY6MLhvrDK6xuMZKOGN0ZWgorLWSFaX
juiE8SBxru/n/cB57y/2qH+0RIRMGkFKvCu4FoS3hIUOuzPkI+A4zW3usVsbv5Pj
Gr1Rj6UkH/E+zv9GhU15XXoHJCdGKgmJTvx1HzqbQrGWfCoHPr+XxglcgygNs8NT
VAR8MpoBRx+AGkUuF8v6tKZUTKp7DbGhgQjb1vWWEkzs8PyfLBRpC4hTc5uQbc9M
aBvBL05BYXXgXgnmuWLfLXvBRzHnZQVElkKRZeP21cZk0zOhA0gtHRyxJn+p+fbB
pBeWDBlWFNuuXB0haznL8VTGQ3m9R2it4ZtUkd1iZ3yjzT1Cl5m1HmWx9t8vCBlD
mOiMgVFvyy+q6MJscIv9QuJVlrRpWqM1ZDLfBNE3n3AqytjN3WHMJNyNV4rTz7Bj
XNhKXaqvs5DbAtPe9iUjfciheoufy5Tbu399DZKfjywyCptA9REYMRRx7TmYKCdd
uivZhZwBHS0UkC8nrz9MtVNnSRzFgQrxS6UA0xMsZ5a2FIwoLglc7JJxuY906yxp
mXDnXRBoKhtCLpy1bkxHOO6sEJR16XXxTeW7U9Xlwp6QNlIIZjNjx0MacJ9t2O18
O84eQ1dBUJhM78gfEV+H9A62CEelLgxlVf/ns7PsgqLuA/94n+VSZ36spilpJrvK
R+0U8eBofxc7G3mxf3uVFzP8w63oh7gkd3bEG7dHn8QuIombYgCm3gXfEkuOr0t2
YPJ2yM4yx7thr6iO0hCunhhhrONe91VFaNGy+5GWG/EnPgFaJdZMWs7jCcA6l/mA
juc/oSWXcwmiaMZ8n+K4aBYvdsf8kFNKbJO8UwqsSuVKMItROcKeXB0uCuWMGdxa
8b0k6havcNY6f5x/MAn/u9t5eYA9ajJO5I4ELqoCubJbfSWuqf5bhdJq6YM8tc4L
4FBWXWSh1+Q88IXu8bvK1F6leEz/ypyQzsaFkGYtsPdSewvSGPhk4RJvQX+mvwyQ
jjP6Ye/E1GlL/82Tynt3YKhiL94e9fSQqwCO/HrBgU19VmegZ5aR30WrLCKgdeCZ
Km1PYSNTRV6p79QT3EH7ZawieQGudT8zV+vbnwPIEDbOtU0MnXw63tQb3g/Dppmg
YBKQgU/k+GC78fODNwQFeKFom2WPNRbjJITTp+GmPcupk9s2MgBW5TqBjgxfjg7k
XOWbzN0WQJ7MFxHG8LByw6RHpLs4GKf8pdNjtBvPkW0gBQaKEMlGHqdpDmd8W0Ju
vFrDoJA1fNyQEW5lFjrbimM5fIuKmhZTwImOGFcd9QvzCMfZva8moN92rWwF/pkN
INaxOhBEiinpG7jLhFvey5M3A73xw0nL4BAO7+BvpRg54O36CIczActihN2YSusa
VxzOn7SbWdHCb4xlObi24OV3EZIDS2yoM/qHODy7ulX6ccQ2YB6S2YVpaXn24Vw6
0K6tbbxDAI89tqrN0j9YrQcUEUi+pmHhFwNui5g3CO0w70KtxxWTiMSsVg+C9Nli
lJhKCHlGKXbyCniyDCN0V8mZtSqTKMDomPUvvRzcQiYA8jZqRpDLZQgU1PNCvGtx
Q9+bJ+96VKov504/+M1oJpzUvc9MsgZytm4wdYyudkzWKk2jTwFMWbsXjjXulIDn
d/2ON2ASrcJsVOXuGKthJw/Mb7UZZLoTolqu4+1cNDbVR7Nuz1d8G8BGrVxaq5Sl
XlmaS6z9c/yTGK0Cg4R9O7kNLUNciYDLRUgYlQuq5IiLpdkmRKeCx+BTONY/wpAa
6E8ZABoP4+NvE+9vtI8qT6TAty8B+Lu0wdLG8W55GvN16/JAiMuyLpr+ADMp/ShV
4azw8F8eaiv0CdDrcqI8EFqZWQLkKULC+Q7hhLkt422veLovb4KiuDBKv4K017zK
9/ulDgIa76QSxNXCtJb1vVw1DRLLQEBN85heT5VBB6zHAx8lugE+ZmROh+K/Oe/Y
ERW6E50Bb2DBpM5EscRsYrJwR3l7bqyw/lE/BgdsUj3bIbfNRzSCJnBAiVBGOLfo
0ZqOk0zn4BesLPbl8TC3NJuVGPJuf3p45dJiqTFJH/LZpE9owyeeTGjt4Z1JF/6V
Fe4knk60l2DFgzaXoCj732dtJFOPcC83X3aBEh5aMpFpOLsmHVFwtkTrCx6ohXNZ
mvVNfnbRbwcbM6Lc6OH0iaAbUWjGDGll7vB4/KPtv8n1c2VwQ/Pez11LKQ3N2zTg
EO8yT0YiUrnbhhvLbjOAN5/mKq5MHsDQKiD1T2lDwG62RPXU2WKkfb0pD8F1k+lg
m8T9dJCQX1PKBjtCsSqIdeTfh8esynSU/NnNsNsVKzCNOx4o0VbWr4KQO3udJQVB
oJdOQtsPHbJWqWT5wWQPnFabsiiewN/6ikj/VhPQhfvroKNXwoIk0NVseFzsZ+py
j6YuJDJdjinhwSxWm+LRPKVzgH+sX1ieEyurzrQRGOa9DYyZwJqyGKJYSb6K0jFN
lbhlFMp/wD0cqO161bsgLbHwok3ldyslr7OGf36kG6Nv2G+vQBAibuVKGWJjKNUx
4olNHNmS2ojNDT3an8f4avwlujQrQE88kWcQjtkQWukdXbEW9unDBB88uV7Hz0dZ
RCUaBAdgLyvrJAeT4KRhL310xeiODigcBOAhEO5XEjfBeLmhQ6M23Kfcjrfg4+CF
8VqINoPrn0/EFzKlxadZl/ligcNj44Xm+pSpg60mSbuWLFxia1GllN1YgLx9BJKN
lypfXpmG935lHS1JKpm7i3EHaM3u+ooTEyyJJPu353c7JUZOqJHpKUXW/7WqX1qj
eBv2YN0Wt1lUFL66/dvKAISkCgxkLX95mBIQhH++FWQWsGvhIr0eAVr2DOD2Rrsz
2D126lIzg+8L8zsjrbkwelS/meSyP6d8Otl/6AvmqsCjjRJSvvfdoultZh9Pg8ho
wfXKXjfH7epXo5OtuR1jFZOX5+36c3Ilwu4M0Z5hCVSXOj2p/pbR3uHd0VmMbVtC
hmBpAwT8PTxeZyhbrSGPqJ1ukX2RrJz1pFznJfDiXZ8zE1zXFDItNFlpEQw39/jP
FTgGm2DHBoJHCL2CeUMqEGzbGSophl5GaHdmpKoxhpTMp8IWH/2m0Z3T0nA3AprJ
USWeAEn8DO0e1g+O3Z3QP5kvF4fLH8kZYiS+kusJRbcw+VuzSwpLTgcNPEMg7t/6
XYfD1AUgQz3nrXATJbL9Ai+0H4raLSKHKjkCwn9lxQZRhpNPLBYVTcXtNmV0tMr3
Du5FsHMIj+eLTzN3S5+eG6g8E7hLCcsQ8VHZKOPkQ7+HGXtA0iwsPIbcIUgTUXYX
Gb0gni74moe0Wui1C/Rc/Qzt7WcRNWSdHfvVjXaIcw829B8zO1i4Y7pImEeQYtN1
cM2TmuV9fKe9wUhns+Qyft7tPAT91k8lb0av40AppJjhHDYG+a6zpnhwj5BBImsr
1QPaDQNZQWQu+j1d6u7mR/MO0+EDUp2iNDzVntfQwJP4UcWUtj4a7gyGR/WGOPeQ
ary3TRsBgNJ1aU+/yCZ88b1bLQJDhl9kcCTCB6nG2OVBXH8IhLyIu+EWRqgnT2J9
1XwVAsLhnYov+JUQTW+eGAnDNazaGUqLfxFpU1fYTjkvcotkMIU36c6L07AUk+xR
dlXteOhXrPDHKL+7fOSVKN+HMggP+VCQ9dJbLrEsn9edG7oCL7W+imEGIvkp6Y3E
7x2miYihhPtI1jxSzJrsglNPfnkAOuxCSxCBg3tGdr6Ctt5xuRSS0uhIgOUjX/tK
IM2yWsq1uw0q4PVy27QfLw6WP8mYfQse2iuZpBTgMCaeinH+CTZMMFsCol0i/fc2
P/QsRWPe9inzhWvm+ARM0brVo8dUaAUFk6CMJUoGb45LrnSE3KhSH7Wqyc1RoeYE
lONYroo75le6ovgdI0ewg+ShX2MBDnlLaVSdBDyDvZLzAADF2H3j4++o23parw4E
AvHwtVPq27s4QLH7VNwUUU3uAJXWRjtHzNKe0vQ4/LqldGjymSONd9y65oorySo0
15Gfp9wmUDoBgWf8qvro8eaP/y/DvJR72aivCnu/xm327wsX22P/evmpGAXJQhVX
acw/dgm67ms+8VlWkIeqWwotxQXvhPzDuvATe4dsmEp/Of6Vwddm9dMprlPpNGNp
o1qwhC3Oot4EebyjMaLoK8SecQ6m/4XlNn3NUJ4YCleaA2BG/ynXuj5iRYyRLW3b
usTKYog+JA9TWDOl89Z6LkzKJSsGGkRoZ5a76CZb/amDmRk9TFpxtpYXVZLXAyGZ
9Mh1dMCL1iAfZuRGaHP9pjlk2axvE0rf3QNlLVFKf62Yr3D1cLYJi2HsO3/RSZx8
5Tir2BwRfpT6E+Em4zydIEt91O7oM512WfcvUgIv29IRnpZh+h6GelgJINdPfnzA
hKmuf0ReKGcVtDo8HJ8V5K6dGQSL+TmlzoVE/19Zfb2H+02AGftyu77AMZoG68dx
B5FHKBY6YvgtNJksW6O49mohps7QPcOE1d5uF1iaO2f4FeTQM69LfYOKyHuhJ4ru
3haoL+0NBBaooQtoCygsEBYUUgfYGzG7pgs4HN4oEh3+1uokGsObpedF/zVWchFn
8YGrgbGkhl5K3lqwB9Y0eD//d38P1JCuT6NMg3dFhwzIxwTM7I93wP4H1WHlYgt1
1iKY4RGg3gaNakt2E4dyrgBR0U1OMdpgxqNdmumHDYkFUH7VMACidKRoWLqujM7G
V1BrDxuqDG2ycM2yHK2B2WaFQdDVm+/Pm2hizyp2iI6elGGRlCaQBdhg08WLm78F
RO4hDEWn/XHjSvQtlNWj85ignwWHmJ1d47jH2mLmL1U+7pPoXr+Fa3/5M+rP/G+D
KjQpfcVYxg2ol8o9pQl4kFkXXI2TKfBVbxFH9cmgtziWT+Bz3DTDeQpvlEIPL+vF
3XX7QDMs3dO1clI0r3EI1GdbDP3UnizlTa3k1dJ201HDde3PuDCspxTep/e90N3E
ODMdtHOGXk5AhysgtAwGflUQmoehxeXqneLHrR803gXvaQknb7rsSGWrm2D4WS/V
Ss3of/e6lfaGMOZZJj0bXxw5n8FwtVVkYTgdiDyAeZ5y3hP0x2oL/uiBXygVJWC4
D2CA9VTrK6u7rFsOw953WFyzBHWVStKg9ezcBnCBKEYDLOoYfVqLgZu0v+rIcxLn
gDbcWesmPHoFFSa0X+s84cqrlHPbVYnNw/dcGjT3erFWZvijrMR+v9s9gEmaFLCP
7b5YJoxEQ2XNhlgYndIFoNToQMsvX2BvYEfFBLUXAbJWG1zK2NdF3Gz4GAiYMjzr
oDCq8w43BsxTYiCdW++pfk8ocTO5K11RHV6m5ZGNIh1XjzPkkuSED4isRpZ/Bpwx
bfNCXxIUPEqDRoi8gex0bNQC6SihhATHIDaCbx5JKmZCFLsWnD+JAIdb2n5NwlEE
RYlwJBqDuFDv3MHlV7akmphaBY1zTCJzmycXo/CIX7Tzh0Z6CqLvynMzZuSKTEYX
zc3RKDWB7VVMOoudrRehMm2EGPru0zAPGKg0MCxiB6K0WJ4SnMU8+RSt+uiZRLZH
cNYCxj/d/5bFud3CGspiS6YG+TNBMXCd31R0JP12dqIvAIhuxHLQnedKjXPE+kPi
iN05udVtuSy9lRoWcARZttG8A4VEj2nKmZY1uOd+eHvLsXV5UbbNpBxB1CzQJwJP
/JKzVnRGI6GxILt5pnBzfeUu9AAmlCdwjR2qlcB1qwbO+x4WDH/vWteFTNxQJful
0t/5ZHWSynDKKz2CeuUOKWceIIsbGu3WDoVD0nsZDcWtg7bQZZLCOGjT9tmH8qU3
qRSKfus7KVWBNZhAV7r+sE5/l4mCDsD9cArnschXw4SVtWhJmcsbo7eNcl7CDnW9
mKdANmucyruIkg1ph/I1lhdJY4g2W5rQbD0AymmpifW+pfngXSACkxucO6GZs7MS
kzw3o0Bodp6TY6vSTmMC9LAbR/tFRuGQ8NK8ktKH5juMujQIcYBczp/kJU7m5B/E
jM9eCbQmm8ELIWcEuxQH+EoizCi912wiva5cHusPP959yKSu7EHJeoFjY8z5LduM
Q9rmezuGV3FXLxEycTMB0IUK9mQc86DfPLVyoAVOmZt9NZk0WJX3b16O4g4SIInz
GTtte+mBImqqMW94vfM1h9EiA1XPozyuMBftI/Rc1MZ6dbMv4B6JU7ZVklY3owkm
dpxpBww6XnVn0qQvv2a73rlV8phkca+Gi+hLsSPtSCuyX1221VisZAc4P3Gc0mMy
HvzRsbdwNKW1GUmWKBS0Zwl/r73kFtek+h83aB/RPX2tNyH46UILM+cGqM1MhuDV
rTRLv78bitghnKwgvztI7w2MXAUlGLTSgg8ON08gbZGfLYG268VjHguc5oQli/EC
B8Mca9UHc9xxlZpgvVhjIg99hyHogP0QqpNJBzHt3GjEDxtWW1qYg5Z/bBkVjTUb
vGTkhk735jUuK8mttKKqyeq/1h9qWkSXJxU4rRCgZ+JHPWSRLjwgHEVG4+W9L0WZ
mhAlkTmPvnwd2I4W81/A/CyK9R9nwoZC4SiCHqiFtU20IYX3+0PYdfDuRWGV33o0
i7Ou1tpT++tW6nM7ybRd641CiQzOZFxgmkYWpU4W/rpk98tTDsAPcoYIVURIX8nI
fzt0lVmBubl1E5O7QrUamdzNLd4GLwj0ejgntzT0ikYyeYNx2WsLhj7eaLJUDaz8
rOPVwGG/allufCjb7Ubk898fNj9SxFctDfHa36Wfa2Mi0y2ViAv0tXBFeFNukBUU
0ifQfEHiEI0cB4nJ+Bi3L7EPksGo0Ip25fhSjhwk2/j7LTMwlTAPyplhkC8TyXQi
Oujvw2IVUkHEPzJrUwBVLEkQrLMiAOyeLZRF61Uj1mEfWqzTogkchF5B61AbX6GM
53yzhYMhE+C41WHvYYTxdLO/sjSvtNUTA/aRVAHUeqP3lF+RXiYPKl0GKjPLwvFF
MtkE8Rizo0q4dujx8rNNtaGX+W7YdBN26GcxZRvnPU1tUoxCZd9J/w5txCZ3keT1
4zaE8WLpLOs5NLZ+lnCKunbSwGtFjIRL1ulYdUOZxv9GhRx3rH3fyGSV7jdEkdLj
eEKko/8/FUtl7ugvOQ9QRl6Jvv+cu6HwKyTBCJ6/NQTEevV4vaoW6EijxG3IeRVu
CemhgeiRo6MPjHY/m+HOX7AJrFThx6rJz+PaEBXXUAD5mfsDqVFJFa8YhPhM/PUs
G2HHhP+3z+MYWDsqggdoQQHTHCBMy2uCsylqdnUYA5ISBuQEpPF2jCt4EYC6/JFQ
l/YiFpzIjvR6KpBHbtnAhOGRbRmWUdB2Xi3EhOSNi2C1kVc0cIPpw32EIRDCEmx7
QjoBOFQwG2Km/NKGmsTp5I0EMzPjpYzoGRlYCinRILhfWjNRuUFXqMT4q/XP3qrH
ZzIA0oXiuD11nzKuB+SWSgfdfRxdwW2FLHSsQeVctB8Hu2zI/gioL+IcHThTYja/
pfydDrNB+2xFaqNa207FPENyS137Jsz9nZmf9rXhmjBkuSBoDjTjvWL6Drz49+fu
UuY+tiaC8dL1LB7m0OOjOpD4G+Ks93sfi84ltZeVCkJZAxbuGt8rwrDpPBUcTIoK
QettoDYMluP5w4jRzxyHvk0Ue7QiysCJLKoex5Qr9glrAY0bdesdJp+MGHihuFHr
5X0MYOiCBadq54rjpNria68u0htIGbSqX9eoC7hooe3STsjZsUEBwnIV+1OnxhAj
T7RvD22dUe4moym2VuzlZRK/FucQ8W7Q7wmH1uKlj1AT91UBvWFb2bggjariPKMl
hf+tQl0qOxFN5VJOQqHA43lnqG16nA6VNzLM6Id+omEchdHh03eAXcpnCyJmafr7
euwQtetBoCZ8BiQ4SLq5kHBQUzH8UDzBroz+V2u7p0S46UhzAg2IcxoeRlyC7BVh
zC+pl2JjXQVtLSh2oDTQK/xzFZADbb2A4DVj4qTnnq24w/Z2+DN8GVq0tLamgyff
NCozHG+70Ahco/BFL5kSv/Da8U3FmjZQW9PY66qd2dZoKlpp5o81P0V/J3RV2T61
1WKD99viQURld1auP1KLeavS8GkqRkr4yyG8MTCVpFaeUscskebRZcRqRq1r+D28
7uDEAAh6uChj+cD35dOTRWTwCfhdlpykN2B0BoWxFkQTUzaauTfghVrNFS67cpJO
kRqWyM6q+Lz6T6KLW7/asbFl6MszKRNge+hk9xctZ1JjP30LezyUqs8QQwodtWt+
v2WgDT1Kp+V9Av6gTIAyI359YnhwK64YdXJvnfI8edc=
`protect END_PROTECTED
