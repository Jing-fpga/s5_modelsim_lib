`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UYYHFRswJNbuTlzhTntpxTYRaVjWy5WfaG31WPREWtWPwPS7qQp9nhxG05x5Mjyt
9ivBLoOLGY5AUtAtrgYAvcTfAtpMAMSQRDU7H0OsY5xiCz22lRWaF+j19/5NroFh
6L635AOFvvC+nl++qv0EDC6e+wIPYDdoT/w4V+To/GDj/p/RMEtj3aSJPb2liI8U
PBtc8NaQNXFzsBt5BlViZOhtR3xJ7wlQIu42UwAK3bcSbNNq/dPVlVFDw12f+82b
Ci6YS+q8/zRbJ8ZKqCx119thx90Z++/jhJgAyypPevW0HaWIyE/zD75DvPrpjunq
SV8APqCohUlc75ct6EZw61wGYRfMPuflK00w9tYANi27KbKlsl0y5crh3bn1YZop
bTWEK3yipMHZNzJVnupZnsJEJU0jHtaHtQ7ryQQ5w1bqGz+24KM2HxkULlBZqxK0
9/ufppV5WyEqQ2cToqsgWV0HsthFaxvDVBj5YVqizakjwuLTgaqcSoZcLVywURxq
ohx79SxXD+t/YGPH6qsd1xRZAuM0LcXAMmSOmJosgO3d8KRVSjtZ0ttHS8l+HyeS
QeMVIV7z9tjTCyzPRx/ITUiKduOKJTcYwTfCQe0Pm9I66HGlna2N3CX4454H38Y8
2LH6+p05cLdCBL1DV9f/3gW+Tr7oPlCIPEkyD99KvDqfFcyjHrzwT76ZHe4E/VXu
3N+uBqwvpPbGaEOPm/Hk36gct2XGh6on2At9hV3TSGuLeCUTJzkDTH/fWD7Ho0ge
WF1/qHOHtujvSvBcr9CmBtOhKE//DjpSCUENUrvmkN8=
`protect END_PROTECTED
