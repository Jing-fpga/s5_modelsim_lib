`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RXJPw6fP94R3gCckGe8HkgVp6dYrqBae5/q3zXyiGL58AMX+Cy//JeU08DTCuIyy
ogX2AxeWN9Ue6FJE05EHeE8Jh7cNfKjKajGjuLMeF5OeciONSGgOgo+bnLv/eZFw
DUYnEk76k7iL2pJHYx6EB8R6dLUOrdEUw3A6SGTwJKLS3mIykD7qN2Wdna4GY53I
JdN/5JapLu4B4fNWvDT8Hf2HYM+EEjIVJhcWwWiuWsEC0dofbPUQ5vTDqIVvs9SY
jylggcBYz72ootWi9VuTUkADso5yoc+YMjUzlCQLug+HxO0vYLaBS0JlNVAbpboU
Zad43aBb6LrynUyLp9qFGFkcLIb9Yx8Mu1AF5Rw+7Egc3IVnYw370/lsNe+6iY7S
64K7i5hcC/F1JNFgL1O/4o1JJoyZ4rHmE4siPFNvTyB/RgfN+QN7Iju/1evOhWRd
bNmc6G0AB+A7pvXNBiUBbiUf7lKeLsGe7yPXWE1Wcuq5ltnqWJDt8gisTh6q9UIj
Q8XC/pTcMRI2fPo47Abd5uNreI3cBNs/2ofv1ZSzHrxMkyQiMKFIzeF3rsDwZMZZ
b4yjQoANcAcAWlzGYXQFVxtkXSIOgNHHhXu0gsJDH5cFHmH0HjX9WaKpoDz0ExGo
d1al/ZOe5Of9AvHw7kaxiNc/9BLM2umwAua9l2hQ9WBr4keFERnsradG4EvBS3eK
hqBtUnAP/xyYu+W68vDpz5adhRmDiGWRe4LA4y9rTJM/0aVPeNHGFNb5XtEqpcZa
bv8v+nFucxpKiw/B9aIE7zSZaPf84F335uUkAd2efNvHeeFR2dm3EraNMnSHTlcg
VKNcJzQP0eoE21d3PHAb2FGKtu0R8pWtYMraXORcf505KtYxX6ZKJqnpJJwkxbpy
P4deqP1m5dTAxPnbDfyoicwedENbeNa95Du3gltMEgHzpeQNnumBmYoxblUlCffj
Mam3ZJK17B8vXAKZZg+wn31J55+uAxFrP1OG/gOjzcUdHx0QCTPGyISkhrfJkCHU
p4Ok3Sv22i9R0YYXM6B8f4++z3tUJE9BjMpkianm5IoX5L+te7IzDp7KQ7pmGU/r
FIMKwW7gWIj+32pDeAy09SH8pMFkqiTaFsp+e1lEy1l1Zg3hLM+dC3PrrRkPom9D
DDNcOw9bHdHU4ek5NcEewtr8fVI+LJ9EmcwttAOVDUK5zPuDWr5LIGCPKr35MM7w
yqIzkMQkslTXXNEh2q4nk/1T6B8pnnvM280+ZjVwtGOTb89C+jmVxIEK2MhCGT6a
lewoam86oSvYiEXH1mSGB7zpKwSRaTBLp9eQRjCVLEap6A5ZjVl8s7povzoctYHx
WVJieIlOYsG4GhC2I/ftROX/l4aAjVbjHCMnigdKEvMum65SYER7eORefn9bPVEI
eQgILwX5BQULRMQFTRUlnAyhKRx6gZ/iUiPtX5GzLAKptD0UhT0lLKJQWSsNdEBt
BLlBNKaZbIHLJCPiei5oS4bPCNiOQi5Mg1utzUDUBj1qj7t/8A4mKxvMa3fDOt/9
eQeAnaZT3pOYPTomaOoY+Url9zP7wkwOtfRJLOqEA/qJfGqCMrRckCwRyoA00o1S
Grtr4wHnfBgZN2hhK6xYNvYIYrZcD6Tm3sSJgSwYcjvky1PMp+2HPm01fHeIdvDd
HANS+Fvuv6hLOEPyXJ2j6glm0XaNDhfs0NCazdc03JQW21OTHZ973GYhkoEr+oqz
3eplrg3ASDPrX0tldWQj9TFFjq7nWOQEOM2jDL1MNglBj7QYY1l9VxnxBm0S/IPC
J44flHldEErJmFDYtftmiqs7RxlF/4mo7axTVgaUO9+UPErBK8ljYWArcx26icxi
1b2M39fZc/ClL4mKs36JXddHWOoR5tgBqwcLnCytAuTyB05drQEfEJHsKZVUfkR8
3pMo59Eqpqkw9pJXKJqB54mDprunRmvm5uUeGEI0Oyf2du4uvDZsXQdis8f5wOhR
cW+ksnDnGFB/Y5VpHMVg8B+a4Z8llTmv7QUXvt59uIW/zUhjNsO+/wzxQjmOjza/
k0jtHPm4ELlAaPp8x2OBtfC2k2ZQCHLXNyTV+wGutwVrKkQPMBYoKZr8lVjbVho/
`protect END_PROTECTED
