`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X93OIx+LsJzf6vKHvz7czeEAyjx26Uk7LewBrxWmFDcq8yNaVxsW0feK57NRAQ0G
7Kv5y+McHWReSY/SOKuL8TW48AoUMbkHcuxgzspZTsrGgdGVRqRFLvO7dNerVchD
HSJ3filSqVf9EMYhfr6Lty4U2AXZAAx2qE3855wRoTVkEGzoLWwqrphBx4b6UyfW
fgJnEBK+ONw43VlU9NuE2nFz4wTlWTT6Xy+Lb1Ro2QISGsyQpfMJa0LUxvZB867z
P/los3i7HAGK/LMq2EdYhBclK4z6a1zXPnj/IoE/Md3X+aFrbprzk/VgRX546s0U
qdSeUJ+i+eKYm9A6izfX0qWrEZtA2LJn2UW/SzivtKLpGDzILo3pvrmRs2E6WPxI
54gk9lU6o3ROik1lLUT0yqDvrgdo6fzno+KkVoai1dNQ07IsWOTj3UG+QmdffA5x
lMR1r8sw1V3186/YWAVIiSjej3FkE5t7HMA608pFLESJhqWACcvsaP0KoPNaiQJj
u7o/gp1xDZVnIB5LanYxsrU7qavCu069ESyjTp4jeLKruw78PjH6O8xyGknLPwu0
99f0M19w6pe9KOkWlCLB1g==
`protect END_PROTECTED
