`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1C68JQrE7UvokUF9a/kDbcIhPNhyXt3/GRdD/q6E6gkjfLzly1ol27ZJIic5xqLi
jxqzsg+iw2UzZ2iJ21mX36OPfpG/WpcFu0xeeLdYgVuSPsvnhkVlGQtV3dppN2n1
U2IrYKl5EKFWxLE4QjdyuyHjovpys4rny4nDZ9BTqybaB5oQDidQotAGQ7r5e17W
Y9i5RGvHb/V6jKYkJYmwGtSbXiAjZGCupx1VgIgx5S+MLr3vjOake3qnrX/RDqBY
/jWFC4fzoPcJ96QbRhfdaPuu6R6NqqZ+VHYdE+9pzVSj8feX2QsGA96NI+3B1w+d
JrznjiXcrz5nCbs0wvwOFAFFDQ0SRjFciUoWKiKa61jsgEWCPfAauN4jPsdbOoqa
mIdiv9ibRi59l19XtBYwDch5oFqy51OsXQzxHQmpFKk4Qyrga+dKjB/1DTFiScg1
lbP7ai0oh0fK6+hwPTxH1Q==
`protect END_PROTECTED
