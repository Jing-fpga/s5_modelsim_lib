`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQG0QUDFBdVS43TX80gRTXgMAA5Px8qOsAAhJ3fKY5m4Cq7F9VyC3u44H1QFpmVX
dMfsb1JL+zbPs39ANuXyQzvgoFENmY9VGc/jEqi2/KMJzbPF8/49s0XFnJswMKOc
WJb8Mo7QsyDq20/1XdwhFPr6LPRA6KcALFO9xCfcDkThjWSLnTBl24tkuc7booaV
25wuXMoJP2O7nEvNkN2oQkPPPiyFRE/uj9MKuiAZd9onymgeu7ZKiY+uf9kudDQr
c9Lru2okxWoSJP2ZEjDO8FeUWjgs7x71/RL21ery4OHWHQd2T/Vpt83oa3+CSQqi
nzORZaRXh901tsPcZbKIwbgsfBK7fdM3aPYr7tJEzcn18OoQy2jSafRDkx4MP5NG
niJLHDGmJP/3Fn9o+JRL9L5XCb7eLYrn0xJ5lNJHNslgRmmEHn+LeJEjwcCvgdLB
D4sWwt+xTbmFtTOoCD+lx9N8UIyD3CdkBoxwnrLTwjdAe/EeZCdMEMYbwrKg9Jq4
XHAntQ9Gf+ELFpde7QFjBcojDjyRwqzHAiTCDSxAIM2nbhQrE5TAvMCTnm8B0UZC
xgzE11TIRR1H6Tl/4mg+FQEeOLZDlVcHj+UpLs/idGOHMjLH5KqoniemIhHJ9KZe
Vz0vdLyUNCOeZOAoPuSijsEY9p5kfGT2AmpVusIiEesvefmPljckw7EfU17Obeqi
6ya5QfZ7JYHdqYjpuRyhrS+riksBqnwqAOp+XA5Z1tV0jNyyxXlsdid9OjMHasuC
`protect END_PROTECTED
