`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZlhY0OiTinfQhbYBiyCos7qnpqCjVmpmf9B6eIy4FQz8bnyJj/QrpNa8Ovbd3mL/
2mVqk6e+lN5qkyyyxWeBZrYGYgvCy3rh0e9C9BHlLogmrBwqhpXaGA0EPSoFcg37
intF/5AvxgqEJ0lnO/1+wmCCXim8/rEvK6bKGK80mvuyV4owZ6y5u6dBXpPl2HpW
NxfC8pl2W9xA9n6Ijvu0BywEN0bBH2r0p4EHAR2CnZ5tKd60SxzLtmuzKdYtIJTu
fNonJ7xYChcqlTl21rrnsjE3Obp7/egusPQvhYaqpWIpw9c0wn1C/kbpkvgGHm6k
9rWS/vkNCmr4w8L/SVwkmXH8GdCGyN2vN6VdBrn9VHZQGRCMa7Mm9Bsak+J1PHLt
Z5E7zoTtD6Bgdkn582AcAGX4YDWcHqFACCuCS3AoNQGkS/SAmKWn1fr/oOY3f2Sq
YDgbpe1VtmOT5cUWWM3/QCBt+1/mhiqCQ0F3TXriEMU=
`protect END_PROTECTED
