`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TvmIZeeqDp/9DvFt75eiUH7jhzbfSfvdpvrqVb/Y1KHUlZGCX7Yczv0lMlK/5JB4
wkxBXH90lYUQpLqeXw8O1b6VnLIHMf189DZc5ErfCUpYhr0fWJ+ed30TxEGcyWDh
OT2V59xFiMzN42/FQdizsgcRQOhdj0W/KCIStubL/8V2M1RpYfdVO5Q6FLbDsDYe
ivvVWBGcOZW9OzvFhQTwXyUd4HdfGXgS0LIo6IET30MLKbPsK/g6RJ87R1te6twi
kUFtNMFWxzh4+odKixhCts4mpm8kQ7rY3ptTZxiLD69BYq1eL94ZjLLQSU/uCOBt
f3MxPRJyGlw57JMCDI5SJRsj/H3cJw4GulbKSjDkFJGaWjmBJMuEWhmjr3Wma2n4
TdnJRf6XwGrYsWv10FNmJ5fcugsP8q7B9S3jyygs+ANHeN2pvXEvWiS74s6J0fue
Qe9MnVvVfdvSWkX26dbfIdSkCk0xqEZICmfbmsw+Q0wVMyJHt/7CgPQNx/20lTuL
EPYO7X9N7J4Ccm0XBogl35IGtqIUkNf3kGGP9XxzQEhVTaXQ75ovKwqzdcHJzDtE
ThLYcVT+Dck8mfRlDXYBhU8T3dUPvWuoflCuyhKEz91acQCSpPSiDsV0II+Bl9H/
MTrAxFtL4o1GVdRnUWnui0m1JCj9qQcn7EYZc5S2lL2vkIBZZtVlRGU1lk8XJ/Lo
17OO0jF8LPVlskYlx/22xkrGBjnGG/FyXEagK6EYNivOuEgAl5vwNS/XyaYmFApb
R9QQ9tSlrVSzWCRUik1KwLTX2G1xnTN3HDD5yU6gKOiifNxL7W2yjgWUtWvXtASP
npud7T/aaY8XLtApLbY/XD1RddVpm6yi4Iyk5Nn/B7pMHKk6wclFDnxZLhxWDff0
G6MrPx8IRHXloBRpS+BbJeO2uLALXqP/BedLFMVSosUgb5dWLu4vhu2v0rnhybNt
IpRntRHai5zMxP8WqVm+HLqE936M9V+DCH/pXcWWkEK5fA0wv7fFmPht7DynAV3G
u1hH2aaQdg6bsamxHrWIrRLRUczncAKGCL6D3vZTSeNgYhQAyY5zbAZm3gkYYoDr
seQOCREz2KcI38+leWCXP3OSJWZtH+kP9QgxUCxUSOPBaqkcXzWNibwyZZqDJAG2
JtbqC3rCdeYtgJtNk9myWvsxziLOKMO8/NuSlJFjSRHc6aTWguIyb6TaTzOnLJfs
gLOoGdjMmnPHdT+WVdkCWSnAXPnl11fK9krusUNx+OYnskqtjB8/L0zKZYSXjZJ8
XWdQT+LB2+01yDT8y19vxd6gCTkSL8lc0zHwR4HuPMs=
`protect END_PROTECTED
