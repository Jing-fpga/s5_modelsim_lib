`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E5yFkcsen4WAPRm6AoIsWsFfbr+OfCTd0fe2h24CoQMXu7QN2E4kypifpHi2HoRf
K+OFWlLy7xndPYVsxMd4UgVFcWOZIz3dhgRALu2T0FMw6iwhQzfYzc+TBBXtktRG
rI1eedztmoOukhPlUvOS8KNOUrM6PdJYH90uegbGbvSMozY+G5shgxh0kCDpeHcY
5c/dmT9q3qM9tdpd2QkGBgD06vyyeK/ZoC5aFJlymI+QXdXKSoZFz3kzzrlIJmT7
R/vSXHk2yrYPyilqW6Vx81h9dXm84cp4FjtR65zUPto5H8ldxLmiP0y+ZKjBBGaY
cfRKUJHUVR7OR84bLEiOScHYNA0if5AKyblUgawDXCKiAicyPo+9hdazaJTEFro4
C/gaFDtpV7ArfO2SLUbJbVc0spC9HFgExKAbU0jE8qe9qf8hYwIrVMKTpGmAsrZu
tcHlYXaIP5HXkcd3vPvu/mJJSxbJFRQub5XPpvDewdtq9ys/OWXwJG5qB5i+tMKO
Dngm9Df4Bi1jTbsTfinGZBbCUlShS/r4+zxAEsPTjLyIbAWEHdFQ2yDLs8DLyk8E
/TbFYAgKH7kUqy+OQK3hflFco1Ej9nF9HH7nwcttk+kkmz9dxdvTu9KD1w89NQYG
ZpFySkkHeeNygvw18dC8kx6kgCXK9vbA9S0Fdv+0N08yzmTHsddyyPmVPohMInL0
P9fPAv00RafFt96FsSwj5vBvpVrczN+Imfq6DF5clNm/oKDTcWM8KrOk0eazsH3s
XdhcIen+RSJ2pg6F1ONALIxR2oZvoFW/8mpnpWrcnvJLO9NFU5eF9tM+3dX0B0So
kT5ZJOZk+4lXZwaCSSmAXw==
`protect END_PROTECTED
