`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L6GShUvzGU+00l2orbmFEQ2TX+VBV1zZnl5YXzJ2G90xOm3g3trtTo2+SH586TBe
vMsbqsI1qyGVXqoP1JG8y+vwIdCf0MBEDAVLShtt2ugDhZ27I2ZljF6/0+WN1+RC
FZJtJw/dtl4hUUUzkrlP/RM36W8/6wMKYUHrZ27+S3K44LV7K1kQCmjS0eoy9U9T
BTuBO0HvYDpsfIRIrI5miGN+ixFpIVI7wlAFT2L7gHO6Loe0b4nnDQD94oEhDrS1
NCZUtCB+uk0BNPrfSJC/WRT6aiaC09Se5R2nO4GULwBiidpP+LMPLMeB6hUNnEKX
8qXUySD42KgCd/1lY7WOssPj23plpDL6ynjja8ynGxnafjjGCCSuT4HSQO280HEc
+UYsQD3wRTtZTdzTVu34IYClH6OGBhu61LoquzAQSCzvJiCC2QRNUKQKRHMQJqS9
E/GQZvVQJeItWVvia7HeflSbvtsAqn8tHHwTL4gqg5TZz7cvz1d5xALvxrDXltCQ
82GZfnrLiwOfjwC05rLBQcN3RRRuG0my/W7fbS8nA9GEpjaIpKf1i/vPoFUbkOfv
tAmOLfBc6gDt6IOdo5DeNuk7yPXwTHBhL0E2iVsgwqsMUp8H2G5LLXLVJ8iVUmLs
7BB7ivgZwL/cMDQrpbIHdaoudr3y6+XdShvIEPskPW4xAIuoAISV7QqnQT5tlZZI
uMkwegFjd1IX9R/cFLs2iCmqrpbjfos7a3CL3G5apKwqLL+TEAErS/TzsEOwPUVs
53f8BRpGqkvW0qG4NIBJWonOm0xZ+IErgSscz8H5Azgk9Bi8e4RgZxDy8U5uXBei
I/JZYTep4s3Cr2D8HxUpWwzKD3Lxrylx8TM8VzqyCMdD3gOiDqIcPURWP9HjpE/e
/XJnIN0UnlGc8JTdu6hsFk742XjkZJKQcsUGnd+zsJ8yhZXeFXU2ASsbi7Mk0i8m
`protect END_PROTECTED
