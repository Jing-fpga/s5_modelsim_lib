library verilog;
use verilog.vl_types.all;
entity stratixv_hssi_pma_tx_cgb is
    generic(
        x1_clock4_logical_to_physical_mapping: string  := "x1_clk_unused";
        x1_div_m_sel    : integer := 1;
        mode            : integer := 8;
        x1_clock2_logical_to_physical_mapping: string  := "x1_clk_unused";
        reset_scheme    : string  := "non_reset_bonding_scheme";
        clk_mute        : string  := "disable_clockmute";
        data_rate       : string  := "";
        cgb_iqclk_sel   : string  := "tristate";
        x1_clock7_logical_to_physical_mapping: string  := "x1_clk_unused";
        avmm_group_channel_index: integer := 0;
        xn_clock_source_sel: string  := "cgb_xn_unused";
        pll_feedback    : string  := "non_pll_feedback";
        x1_clock5_logical_to_physical_mapping: string  := "x1_clk_unused";
        user_base_address: integer := 0;
        x1_clock_source_sel: string  := "x1_clk_unused";
        channel_number  : integer := 0;
        tx_mux_power_down: string  := "normal";
        use_default_base_address: string  := "true";
        x1_clock0_logical_to_physical_mapping: string  := "x1_clk_unused";
        x1_clock1_logical_to_physical_mapping: string  := "x1_clk_unused";
        auto_negotiation: string  := "false";
        pcie_g3_x8      : string  := "non_pcie_g3_x8";
        cgb_sync        : string  := "normal";
        x1_clock3_logical_to_physical_mapping: string  := "x1_clk_unused";
        x1_clock6_logical_to_physical_mapping: string  := "x1_clk_unused";
        pcie_rst        : string  := "normal_reset";
        silicon_rev     : string  := "reve";
        fref_vco_bypass : string  := "normal_operation"
    );
    port(
        avmmaddress     : in     vl_logic_vector(10 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        blockselect     : out    vl_logic_vector(0 downto 0);
        clkbcdr1b       : in     vl_logic_vector(0 downto 0);
        clkbcdr1t       : in     vl_logic_vector(0 downto 0);
        clkbcdrloc      : in     vl_logic_vector(0 downto 0);
        clkbdnseg       : in     vl_logic_vector(0 downto 0);
        clkbffpll       : in     vl_logic_vector(0 downto 0);
        clkblcb         : in     vl_logic_vector(0 downto 0);
        clkblct         : in     vl_logic_vector(0 downto 0);
        clkbupseg       : in     vl_logic_vector(0 downto 0);
        clkcdr1b        : in     vl_logic_vector(0 downto 0);
        clkcdr1t        : in     vl_logic_vector(0 downto 0);
        clkcdrloc       : in     vl_logic_vector(0 downto 0);
        clkdnseg        : in     vl_logic_vector(0 downto 0);
        clkffpll        : in     vl_logic_vector(0 downto 0);
        clklcb          : in     vl_logic_vector(0 downto 0);
        clklct          : in     vl_logic_vector(0 downto 0);
        clkupseg        : in     vl_logic_vector(0 downto 0);
        cpulse          : out    vl_logic_vector(0 downto 0);
        cpulseout       : out    vl_logic_vector(0 downto 0);
        cpulsex6dn      : in     vl_logic_vector(0 downto 0);
        cpulsex6up      : in     vl_logic_vector(0 downto 0);
        cpulsexndn      : in     vl_logic_vector(0 downto 0);
        cpulsexnup      : in     vl_logic_vector(0 downto 0);
        hfclkn          : out    vl_logic_vector(0 downto 0);
        hfclknout       : out    vl_logic_vector(0 downto 0);
        hfclknx6dn      : in     vl_logic_vector(0 downto 0);
        hfclknx6up      : in     vl_logic_vector(0 downto 0);
        hfclknxndn      : in     vl_logic_vector(0 downto 0);
        hfclknxnup      : in     vl_logic_vector(0 downto 0);
        hfclkp          : out    vl_logic_vector(0 downto 0);
        hfclkpout       : out    vl_logic_vector(0 downto 0);
        hfclkpx6dn      : in     vl_logic_vector(0 downto 0);
        hfclkpx6up      : in     vl_logic_vector(0 downto 0);
        hfclkpxndn      : in     vl_logic_vector(0 downto 0);
        hfclkpxnup      : in     vl_logic_vector(0 downto 0);
        lfclkn          : out    vl_logic_vector(0 downto 0);
        lfclknout       : out    vl_logic_vector(0 downto 0);
        lfclknx6dn      : in     vl_logic_vector(0 downto 0);
        lfclknx6up      : in     vl_logic_vector(0 downto 0);
        lfclknxndn      : in     vl_logic_vector(0 downto 0);
        lfclknxnup      : in     vl_logic_vector(0 downto 0);
        lfclkp          : out    vl_logic_vector(0 downto 0);
        lfclkpout       : out    vl_logic_vector(0 downto 0);
        lfclkpx6dn      : in     vl_logic_vector(0 downto 0);
        lfclkpx6up      : in     vl_logic_vector(0 downto 0);
        lfclkpxndn      : in     vl_logic_vector(0 downto 0);
        lfclkpxnup      : in     vl_logic_vector(0 downto 0);
        pciefbclk       : out    vl_logic_vector(0 downto 0);
        pciesw          : in     vl_logic_vector(1 downto 0);
        pcieswdone      : out    vl_logic_vector(1 downto 0);
        pciesyncp       : out    vl_logic_vector(0 downto 0);
        pclk            : out    vl_logic_vector(2 downto 0);
        pclkout         : out    vl_logic_vector(2 downto 0);
        pclkx6dn        : in     vl_logic_vector(2 downto 0);
        pclkx6up        : in     vl_logic_vector(2 downto 0);
        pclkxndn        : in     vl_logic_vector(2 downto 0);
        pclkxnup        : in     vl_logic_vector(2 downto 0);
        pllfbsw         : out    vl_logic_vector(0 downto 0);
        rstn            : in     vl_logic_vector(0 downto 0);
        rxclk           : in     vl_logic_vector(0 downto 0);
        rxiqclk         : out    vl_logic_vector(0 downto 0);
        txpmasyncp      : in     vl_logic_vector(0 downto 0);
        fref            : in     vl_logic_vector(0 downto 0);
        pcs_rst_n       : in     vl_logic_vector(0 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of x1_clock4_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of x1_div_m_sel : constant is 1;
    attribute mti_svvh_generic_type of mode : constant is 1;
    attribute mti_svvh_generic_type of x1_clock2_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of reset_scheme : constant is 1;
    attribute mti_svvh_generic_type of clk_mute : constant is 1;
    attribute mti_svvh_generic_type of data_rate : constant is 1;
    attribute mti_svvh_generic_type of cgb_iqclk_sel : constant is 1;
    attribute mti_svvh_generic_type of x1_clock7_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of avmm_group_channel_index : constant is 1;
    attribute mti_svvh_generic_type of xn_clock_source_sel : constant is 1;
    attribute mti_svvh_generic_type of pll_feedback : constant is 1;
    attribute mti_svvh_generic_type of x1_clock5_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of user_base_address : constant is 1;
    attribute mti_svvh_generic_type of x1_clock_source_sel : constant is 1;
    attribute mti_svvh_generic_type of channel_number : constant is 1;
    attribute mti_svvh_generic_type of tx_mux_power_down : constant is 1;
    attribute mti_svvh_generic_type of use_default_base_address : constant is 1;
    attribute mti_svvh_generic_type of x1_clock0_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of x1_clock1_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of auto_negotiation : constant is 1;
    attribute mti_svvh_generic_type of pcie_g3_x8 : constant is 1;
    attribute mti_svvh_generic_type of cgb_sync : constant is 1;
    attribute mti_svvh_generic_type of x1_clock3_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of x1_clock6_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of pcie_rst : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of fref_vco_bypass : constant is 1;
end stratixv_hssi_pma_tx_cgb;
