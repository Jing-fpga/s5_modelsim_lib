`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SONmp6ASG+P0FpsZLmDUAaL03RCaK7XY2clNpD9Ehh6ctZ0liL3JPs6RqUFCU5vg
4EpdqmfjC7fFtHeynjqv2+pIpb5O6WDyzyrf1D0Xz4D40H1lWtet4+yjyaYQHza3
LEJIP4SsrEaY4MX/9RfiLpYj/xhhGT8VnFQZwV1P9c9eYisFhwLTBuswXa/GAOPV
cGsAsH+2HAtfCcOp7OBLnPvlqj1VKBScpsPPYcVWXpwJhQM1aef6N9ItkluYxzhG
qYH14x5myKquiPHLv3cptywLUiUyxC4jU5J1p2gK6BRHlbyvT960GYeTH/pfl2mP
yggoyQZa+6x3aO2XAuAxOz+4Aoz0tBR/9ZeY1RFxTV/43rj6NL41z2yLp7TeYm/K
hvpvHw1yWzQLlBEQcTK4NRsB7nm664AtRhw1pbbibTc5hvTe8ePgFKXEyZwBj+E2
Wu4ugKNIhLHE+g9vnZzz7PLnVeVZAdyvtb3/HCC7LHQv147uUkqAdO37B2UUWTDX
rumfJudMMR7FubNz8cvBZplGi3u0m2Vbkx/olhUXVj9oi5MDrFxKPdvwv4IvF4lQ
ObwnvVqtJOinVVJRwlrKQDayE0+gpRZjOb7HxVhghmyflKnq/VFE8wvuMPyhVyzL
3tL9AcEKp+adW56HEV2NU/UB5l2kKDMGx+Dp0i2Fh35qPj7SR5rLLiDbpI5KuTlo
2dgitTF893xhNQhxaPulCTfdwezui7Kes+2mP8+G3O8kjvYh40g/W/8TiIBIAwWz
ashoQaUY6jTb0Fg3fctjyV1W7Zwf+taNljAcUxqr5WLscmE49mRSPskgAfJHPXbN
`protect END_PROTECTED
