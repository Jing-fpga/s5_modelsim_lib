`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t+5N2WQH0IsWyexiQ/QpcXXgHm09vJp7DxoDMW2NS82qrFT6IEssw1bcI63ycZOM
vG6be2vTPGppd7DrexlUmlGo2T/gHiCuJ9bYFjbpDx3D/ut4CLOp43CJPJ9XQxjn
MBVy8tJmjub+ISzv2oUa0JAlC3sz43fYvunt/uBKoDWSBP54GqFtkcWX5CKnkp0B
xNAWaXU6/KBUWyg/GUV6TY+jLk3uVy05Of1cOj6uuPN5ttmUVoE3YiMDK/y9jwZ7
MEKMEcRIpOXNKj1CCpCN/5yfgM6a6it3f02ngIvMNFVHUJWMqKLhXN1PEl5Cfc+b
WP3W5cRy7IjN5hcmAz0dFSdZ/2bH7DVQdG1sQD2Fe3AhtxbbAL7FCTmkVL+CTvyM
ffGPHSArB9urHlOi2xP2aC9/Got/LS70TU5IV/93sU8mFtCXVNw0UcjGTspxQNjS
A6Gf8On4njXSqj2R1aDNUrXNc3tDsSPmuPBAMkW8PQG/bAMmlvCkDwreBbL95i0g
VbPWCXvGse3PEC4rVxvVHRgqDh2s4yg6H4QBcDtJMr+158W1ri1dmPDnemaRhpJ2
MFb69NHcx5AWo0EGiRGYqHBbu2B+XTgSEWTRJ0nUrrP3LqLZCmqVJtkvbQDAh3w5
bLxCgHIEYSNceJTm3KClp9cV7keqB3bvyNOu9BTI/CDBx7CQp1H5qeYS49mczLX0
oCOH36V5iFt5H23x+C+my0DWvSyCO5J9Xx7O6THqIOT/TZYJj84rWX0GYBeZb6ul
SUyaaBawaxv2C/bOyzZHAMWEmTVHDB8mYJG2tXoz6zJBbeA3mR0OgqapC0Xl/cmr
aLHjiA62xo8+dx51xOEHWvJ9M+KF1I/10kVG3UFCYh5W9nGwxXZzU8tpouCWz7Tl
jaosGWboYWSUOIEncKkyEoeP39Wovd3NQzfZjaVL8P+Wvbqunb6QA/HcdqHqWuvh
ZmvSUjwuFKF6uVh3rdZF8chvM0Qaq78A/W121EpXkJexoMv7xz68wybSlHm6Bn8z
fX70wc4yQk6vHchilwnHSgbKuSRXGIQ9K6DKnJKlOm+9aQjm9olAiDtuIH4tnm7a
T0u+xKfxBYeXL7I3c6oArwUydoEdi/5BraRTNxFyo6XDeynim+DNa8zb1fJAk4QT
vL+b4U4YeYIY28KJDNpBpLvwYCtP1ll8qzQlQjlYPqou7gltvV4OAwcgpCPGCcZ+
2cHUASOZosSvZ7OoldtxRIELGZmrOqCYH3ZBbz8zSslL/+MH/ryc10FU2hCSbvxk
cf9q+wyL/x9OwYbcixBjX7VVIECP6Nhaki31X8/DxAmjHeN1YQtyCRVr5rZiW/m2
93+zvKo3MTBLfRSoLfvvO0LXeMe+rVTLfMDQVZj5Mr4oaLlq0gsplDix8SnVDpsR
GnH+nJlfEpr8jxW2aeZhPdL7eYx8HkTFs6/dCHf6HbRIy11wFrPJkvr32XimCRH4
aEb00+afQ6LjTMMVgyPNBZre90m+TiCKLhYWLk7bnN+KVow47fxhgRGBfWfmfRYz
BYWNnO7OKBFL55DSs54uvgzmX/dUZMfIPNQvzVXfkeR76UAIITTYS3g0WIjDByJq
jpWCFAMoXqK+85ZUfvmeFHTlI+a8cD94fqZWulZZ5WofqEZNMrZ6OQRuarNNjV6j
9xWuwd91xxAqpdgL7LIPdT/z080agrB7Vx6y4etmKSy3LYw2hTFFz/k4j4WzkrqA
VzVi+TxkSlXutgoqGiGEi8PamM6F0CM8OG0WmOOfTx+PFTuiwb+xkDCjddTn7wnC
pD3S27o0ocPMdHV37MCoIB5YdPuSVRuLbmUkngoscNWzC5kj0yWUwaVfqOp2CowO
dOQlJaPfK1aY5nnKsyHOnHu+s27v5iEEcpXMEhg3J5RG3k9IE7kxx0zURGCS2l5T
Zs/QaLILCvh0eV6y16ysqhBviqAC3Lp8fdi3GZBlVsey1bMMV1oSnihbsJuGABNY
5xbzXpCkysluIYK1584cxonhWvGr9JGLK2rSTJL72/X0HmoMQ9JR5snLWDMb5Zd7
r1ANLqUjNwvtjrzH092rlHkfk9OcbDFancnmwh0bnkUGhbXGBwrZeqY6N3FQCmax
FlISgKMbZ8xoGXqwZo7MqMC+WCJSvko0A/DbcITBQqrq0grtaKmvFYaJX+2+Q+6e
uTS8Br3MAZdEDUudLcwJ+ZhQ2C7TbYjmNhF9V6oTOwQo2X5LG0tNa2bjnjDrIayr
YDNLzQ9TcmXIZvCYTmxPj0T5RsCyGS51aOs1r2WCwmL2NSmkVeJqxfkGo3lyyLFR
h3uopSd6mifl18fq2MOqEUdZ5TSDCD72wAN4fftKv4ynn7jcm4hizFO9I7WwBBmD
PwoQOUb+EjwXY4bPeZV7Um8j/A8uEuroZ5m/uNTomFQvZvj0f0Jj6kiSmrMkBuyv
sWA1wOTd4GW7ECWjja7jigdzo+PUPjCyDZqmmUIusVq4TL6uolYl4AxDiNuEyr9O
Lsj7DqDS9Uow0ZkSzFtAgveVUTeQifG5ukK9nsun8USV49A2onjnV6RxfhED3KHZ
pcsncT4SIuxB9Yetn5DAuhiH8ae3ofEk0E19T5o7myzgBYPWo7MQBNk7cKcbdpqN
5lc1E6+1wuolHdNrBIszMAINl3gj3M+syyfa518uqWbUqzQrSdcyh7c7mFbXIXDV
bZypYvKAlMVymGKRwm726Utkj/5itx+rz51VF5PguHpszp+ddlXswOu8qecnI9fQ
nppg+ex0MG/RNkgN7mjtfJ9wCctIvGBZvRoIPOSzpmNbSVZgMh2GlR+4+Zj2UQbR
I2sh+a1oaQrUENSV/58suvj6Z0j2cQKKswQ519AKlwyJcbS+uqSUUeJ9OFJ63Ta+
K2wXPAP5ZGyhAVf3wdFNlEmPOHkQEv2t1k7BO5g0sJdzHafHPCxBdXoQwkbvJ9OJ
4NfLveNADqswSqHvIsjSHFrjUlymMbpJ5M3R0ksN7VaHz/s861isnObevbG3rNMk
UHhpsozLgFIG03PZMez+JY8rBT/mXSToPhZLnwtpf32g+petPJ899hv3H0Ej8Gum
XS944nss+GKID+WQwm0n8zhQYaIZUh2zVt+Qf7mBlghHXWTTu8djlVzq+cjUdxS/
WYMrf0GRfPPoL8xKhj+kMMwPbsYqgzGMsrakM4jKNIaxp+6mR+z5/QPe9QE8KdYS
I2FS0xHrjDfqEjTuAGJdd29akpG3v3sZzAO6nMHc4aMJdH/absUQrXWu3OFCZrR2
A2iSlSeIs3ROVRl2CibUiA4RX4jkw8lKZ8rFcbE2nPtmj/TbnUdtq2a9xijuzjjo
Ecz9nFlnvddj5EP+DDqO2iZpG8Lel8e0/qZjUKlK6b8Oa6MN/MdIsqRUMqEWbZGD
WcdQOUSDZSj9+uY25V635JGKCa9cbu1RYiFzSlzmMdjg/8ut7zgy7Gdc6gNni4s2
HB+ulcP+DcKqDhb/kaS6MrlvH9NT/yhGU041XQlZdG0Iyb88Kt1XbCtqRUC98d/Z
T6/bwnzLxD0ep9KvqGc8FL+p+80N8l1xQlIwdG00cMO3y0U6XWfQHfqXqttE3lYG
o05kx9Koc6Tf8AZvhU8ZNNaHZSI43qFLq/NbeG0G+WAx7dmq5HyPHXNXHg2jvHlN
BP+j7x7dtU5vaDD1c0IHqcmXKkDnw4XaeexM/+17tKBswko02fXxRTeotDi/WqAM
mz4dRIjlbQxnM90gjnKD0BxXQhxaGdjowc6EC6M3N8r6LJSXp0LjB/snDAz9wB2k
fHO7wVSUP8z+IDdRO7TZzUyKkD0Xi3VzR9Yhn+kw9pzA5S8vsAc+cqTTDGVTmDix
72Q+uFcwUevLYRpGTFV1V2HjiRbAZdLRrzCnow8d92TST6mmoRHHC7Lr+YCm0MJR
Y+40+op47rw3PtS3WAu5daEtp2GogkQ8ZUi8r7K4UnM3ONwZSvNPxdlNtgEQaHt4
+/4rHE9/PzyFJbQlCZ2JOByfN1zQN401p3WzN2PT8Sf1GRZcUfixMtjuWxGpneM+
XPsiGmibdMF1eTbsFfcFCeKqARgdaEVjnjR1LiY/1USI76xUbqgisvIVGDIx3AMU
7jMkFxY0X9kmqfRZmJfQgUiRQofGNxS8gUNKrKx+4bz6mRCONQ5GUbOoLq3Sj3Qq
Af2HWHfkZ8fJNXw3WLF9dHDUqlQ2Gtg0a7MA4/MYecDMlZlSXfGtKF5ltoIdcSb4
8bOYbTtSFm9BesrkHs8uzYcSzG4b8ywvLPZbaw26CCjnr2rBJc5J+hVRrVZy55Rf
09K3cK3iuYdsRB6tWUjg/2Y6ta5/oCJFHV9SckmONJlrXgHtSTJbg0K0T1nxabM5
+SllifFpgFlsYQoijBCOxa+LbjRf/yoEcdnzMheTnVq/CeWZSuGSi8YcB42J0peo
VcHuEoVbnTjmGOzXXPb8lS9GQXsu2Zi+tnLuvF3l52uY4uMH3J97fsDDoLQ6kJTh
ZcFFW6+4rgCVm9ajkWJw8EBIZCM9TIr2cwGeBmO/rd1alsS1HhiqoxQ5FlYf5TTf
in377Z8jLiTaIQm+NWUVyJzICv4FqKeWKijjJChFeOLPEwQdEuTachezT4JxLUBR
psghp42r0pXLMQgwY6OgBt6j35X90aH3w6qo0k97O63FdrX+upNQx6fIozVZnGll
S1eTMGIs83ZJgzssu0wD0qCpkcnmm+0CmlldYKCN2YVovGwx+HnbU6AMg6HkQBXo
oj4/LqTxUF7AApWK5U9rg6DUUmlb1z5ncfFd01Q/A2VKYffO1X54qjXb+IGYcmdE
w3AqZVSFa+Rm/p+Wp2moh3ElGi0tZ5pQGZQC5MNl4gTSxcVkv0xCJlAwoan0psBq
xrIW9iU5UDnSLAJnufgC6CLxfOzL9t2zWZeVFjVTD0QWadq462jPk4rMdu7Ona27
OzriacUCZZSIZ+70meo2updwKUnzqilj3lBSr8ScIbI3wjwJebtqWwstPTP8Okgl
WRXMSwC+2njNoN5NOVVdhkSayCl/9USIcxb3KLpQ04xIJWSNx8HHosL2kSnkAw4X
A7HVrzwmpnJkxMpxzMVobLuJOSLxXHRE2yTATvQYhDPMPDYJC0q9Cy7lMgj/teL7
pGjqODviaGrxfPpZfkvpgMFvaxkyuq5KzoRow7BrlOJkFav3kOSXce8mEMomQK//
+fIwjyY68MAiRXadaZBQ+8OcDgBJGKhcllK+yI37xN2lTGsP8BvcK3usYopBoR0o
Rkg3ICgv3Sk002wHpWhAK/4GowOjxCUU6wPvVQ00iu/9CQVJtEUC7O02yY7U8fln
h/O7VhLVWSdGJSnUECulbds58df0KSWb0BzYgV96oniDnSTjOJOg5pQzLETg/OPE
HwuW03sQhmU8PYxQQoWgMaVxE5U0epjF6t1sl1iReI8yGM9GUTB4ewYWMVNLgy0v
NMHCIW/7vT9+QiT0E6m6ofxo68/qhi1RGIQozklQ5Pf8i0t/P0c90GV+GPmka+1Q
1yY0LTX4Cj7+7a9FbRTTwlpS5GawIYgK381e860ZPLJe0HLHAU/Omm4t/m10gBkO
YAtR6uYwCCv5VQ+Ba+fkZO7cOetaiVTaDTVp6QBbDeNv7A5/okogHh3/C4eMFn48
WBXGeSzlsMkeiFkW2cW2clblmYyirCnrG802ooGAR/Q2Vcfo2yTsHETNCxrhZDvm
RJFfd+nDOMrbc599x+JadWn/Qqr7VTcYjzuoAz1Id/qf4PmvcS1MU5cUaU6EVPra
JowtK8s/gpfPlqf+lvgdjWCJdVHf2CYuv8sxC0b/kgRfBbuJhc16XvmQoD41qGUa
zy7ZG0PHndTxZ1ZVR+L+7sJG0i736LphfjothgjgHJYbqtGGpaIBqATcJ0eC0aGe
5WTFx6SbgfebeMGXAHuYnZInxy19Xo+bzwILI+Pu8qZo8HwnFCR3HapUZUuZlVuk
A8Z6Umrsa0GIjFgn8pt+8cw4i53s3JZ4bR3/vejom1MIrd/T5rskY40B7zziye45
gJKlSZ/AiiQGRRJFzKy96F+Nc59ZgTtMd6fdogCzsrKXLhA6qTj/Vr21DhCxpZ0u
/s+MFiPpbKBpxHw7o0f58zzb+AYfrZc21Ppy+IAG3RD67WYhxotMLkyyo5p0tCFX
ycdCqFrQVT1pwPztrNqUZgFdeCTCKx2qssJ048SoHz8fkwrgxc1i7EKrOykXUUe9
SMp0kM2rV8WP2zouBwWMr4QpLDMgSWJ2AYMThnP2SzfTaxc8xLh3WSsw8V59+S8r
ECR3S3UG1abIroXKdlMj6bU/hx76vmxvywj3QZJv+BnQ1IrtkHSogP6uWTv2sgw+
ySuLxvjBFVBoo0GNOgxx5FAeTIyd/lhFjH1F7XHhOhQrfc34Xan30pGOQJLh9CWK
VqvdCoUSERKUK1ovJmbFbwP3Z/fHdqsCW6b0Fh5uh4jaXK6yjfKIVk45qYPHx+0U
XI6pPz6BnEe146HWuPGw6RynpugyHFykO7lu1fhqrkZnDLvIsNAnYgLitBe3EtLL
gfqfIaqQEcDVJtluac8v6hLiTFi8t3RpnmOOcMMhKTPwb4fV1ffCftDzUEVEGbW1
9093GtTpKcz0iZHrVTDseO8W92fotiHRCnJLPRMMpIWReARjWdHJNhn1m2u+Ecpx
PSlZasOFFMyIIiyBAVTZTov7sYIwtkM9mtQOedHnEdYmBTR2pnOtnRXPIAAyWp01
Ou12r2Vffj4v0FNvtDu7xQBxuwkvfvlv1veGfZ0AiI1q5QEnWDTndLxbss+nk/2Q
pyfEKQNDKw+dbl8AdrDmtFdD77CWM5vRQWalevCQAm2UMcWTyJQtCx81hHFkpfDi
LH5fitEwWuXqe87TW64rZ414jGUEXK7uXwTWFk3DWIn5ya8Cbf95LM6qsJSEOWzx
XwKJ+lf0a9tJEdGzTd8OHrxIIVYGevRbBsVG+h5bES+DarzvOQ3rW/HRcDQ5nqNA
WnJzcuh+tH8f8UPim2ic4zVQOD4OTpOrfu/JVVio7rP/FOXxDROW7zR7GOBh89+Y
S+6F+XcT259wZCN4ppLfib/l8jd8dJUrohWSsTw4Fd+Va4mKPSR/6aAR18fkB4rh
z4P4wIGC6n7eEeTmYeHj5O3Gz9lzT5xdzMih4tJ7ws5+rpM8CtgeMbVgZc1xoLPz
oJuScfaKiTp1pwlJzJJTRazSUbZGVakJGmS3wsKKqJ+RJf9KYyixVFmdXTb6+IVD
8K4oD1uat+vmDBt+DDnFH/lork6cRskAo80HfX7G9aW2u7djFIXpl200zzt2Berd
mcuMXzIniEET0CQb04EoVv1RIea002+3Lv2gQsFeQcsNQ9RriDPEIPQnmps63WL4
YhrIWnMp8kybNWrMQOozlA9iiEwnuewrLAKeoTFwvgHiIqMQ4ZBK02jT1ULGuzre
MeSD4spguq3xri8JwDY6A0YwI/lSfItc+2EnlJDaN5owe5pocCfNPQdD5dGEad4v
/84knCKdikeN9rkZtvVBas64MDTHKolEN4PT7/TuCrRmv3ic/BnHZNrsGuhmhMv9
J0c+bid1cxRUV+svsZbh7rCNMjtaxF63yDHqycBJ/iJewzcgB7p6KhBZenE2HljU
8CvuxWPx8Uccem940eBRQwUyCHv72OZiZIM1Vi5XxAyqqBtpiFcYSTGm26IYTcHz
DX3igYFmTBoPRv35LM7hZ9llLoYrB3LNBEqzLugP7B2I4o4F17/J21i4hnnrytGH
k2pfT/ix1j/C3x1iO2VPJiTn7YYI21WXExL3gH/DbJ5Yqllx7hBr5GIe36+Erq6e
rgixI8rqfpovM9ZuG4aDdG2rXCjcRGb3t03bKoNMQn3uWkGEZOnoranvOnBGwHbQ
Xkbzo1vV7mkiiHhoKPVFnD3boQtwMEmc6bWiT4lArBgR7xqRz3VwmBbXynDtvQXl
2nOpuuYUnHiS3CMsYJdDTlTsnD6BueaV9qUW0JH8vzA1gbP6E9IHjqaGogzb16G6
f9BPUnfW9dkHop6LrWo4OdXXzZbh+9Tm/NqzJ76IFJPJ+vkrDQ5BtioUDVFKrXuv
BAu+11YgIfqE6vEOr00VFa4WXFrrFsuVzlXSQeTNLvLx2N7ygYuzzBZ/5nI76w+z
ZAE6+NC8ISCDqekqjblf4fedEXCzl3MI76gEMri6ZfRZjSvRCIHxFx93yeHxzNmq
5gck7L82PFtWNLfhYMsYOLim2bdYi/75W5VlJEC38zkV1C0HaVaFBmFVhCu3hV0Y
uc/0bF/+FFflq3YZsioXoFgORICz0NI+MnRThvUjxQ7fgEb253vmjmWhT63K5dij
DReF0ZOr/Sr3oRhhP0IMlPNKcx1hxCo/POqDIYP4NnlGb/+phM5maYSkxjSoeBKn
XH8nwR5XbpCNUtX+T1INatA1YpJ08+2hCdbWeAj/v60FYxAI5PcGxQ9stw4obTvU
Q2wIHY7dhBoaQTKkJjVGr8KF5cb3JoZuMTZcamNTxY9w4S9+ZlvHxRsNVUJ2B5K7
RlDfqHVQh+owgHWF4HqjHDtEjsnI5kLYXU+A+tl6fAPGYpcms+e8a6VyOJI2LzLL
3bCPfOAxEB+pD9hmzLA/q7c9C99OXAZcGCjMXcA3zCAU5UC8WCPH+0ErbYr9JnTX
m0G0skZ2UWPrnyLbKQcWlkaOAnmvLDhAyx8mIhZaDfxg01a8e87D6/hTlnXoJqcj
Ry32RkHLgURaf/T0GXGiolQs08VFz18SX4PNNbj8F5WjbYm4pqjUyy995a6AqDU4
oxF/w+TEx+1ffkjUBBZ/25jT5RK+q09cpPyCCxtS2hyWN2aXJjSZwTedqicA256o
HjxixoxWrimfEL89tSMj4iMrfPUy/g/znVVmTvhWJUJXOJcINJfSheqs6JikRYZn
ZxYpt6ANzqZ4pqN6jgpAEhZgEyMg0eRVukgJ3roDpTWvsBhXEAoMCB/ww+iOdbRv
7XTYGIohcYh211SUvLlVk1lFCVEEXJzB3wu+y3+LO3YtI95Tj/+dpHVo08Z8bq/y
ag/O7OgMqafsTJ2Vo5JVFzJ/Xc1wv2ZZMvtuEg3f1pipBtn3tXMMsmiSzVLldP/2
tBrqR9K0AD/QF5d/Tb4s050dtb51+N13kGi0Ym8MyIfo7iI6hLRJ6Bx52BugZXD+
j10yM3ZH3dksI6Lm/WGNpH74vP1j3WRg4WGc9s6nfFAKziPDaloY5FPkj0EwlkJJ
vbF2ET2IExwFdxznV9/BG0K8iYiyj/uJA8ktD1eHAcTr6YFTq8j7H8CAVuNhp/1T
BVwgbwU3MnhAtCxInX3Zdf0pCqTFCFmOQ/FRfHlEU9djEwNJwDxDfwwOz6Ovh7PM
GZ1q6KhIFR53ctDO2+//+g8yRo9wx4DgddgiapTdCDimLmnrLQjbRpZ8oAG3nZbD
tnrTUl591N/rbUwVT7IjqLLYWEE8fiNlHghSdrljyXhvWAyo7MpU5z3n97XWqTIO
1/GkkoSdwl/GjdpFI7oilrBWCw7+KCIbxQu9m2dhNRgBa809QRctS9vERoFqq/Jd
a4A/b6BxdFzwJuPcw0tiuE0JOo8MCTSACiVOUFtq5O9yjqp6j4hqgwRdG3YA4rpc
1vKiHKQsF/6SdgqAOvxEEKg3pYgz41SeLMAX4hGwAgv+VY6h5SWqIwU5ZNSzh2wL
XZCrJaBoqHFqRnLCQWVP4LZ3BtaaD2ImoJm5bJkb+H15wFHgFXmR2UHWGccxx/qs
1LdS+FoOU3WN3bgSOiHQFSLuTGap2BZbNqSQ/k/qDmD8huH4dQQ+ws8AkCcQiK27
sb33nG6xdkaDUUN8gOk78Hz5PJxRBs0SgML5ShIZQxXNQ+sbPXvjJXJN+VyKphtk
J7w10CkswXCE62ATlMX3TsCsBcAFoKOtXRQBvcGWagP3TU4ceiiMuQf4TQ/a5DcR
Na0Nv1ywkmfGGQMTOCHV9t0kpiTZn0plagQq5VfBJyW9aQnQb2+wIyBCacLH9+j7
VBlt1KaDdxQKRz4czqXf2DeYBJsQXTU8QEkLHw51AhiMphXNcuOukQeMnsT4OKvP
zzqd+SYpj9Qms381HtSprN3o0WMyWcWoUZ+5zC0Lf0M7Ghv6oI+1vJT8tJTkwX43
zLk3n6x8J9S7bBqb/aBb0Q==
`protect END_PROTECTED
