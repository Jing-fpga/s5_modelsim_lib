`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hdzJSKhHc03s/tvJZRJlzXOUwn3CfhZC6m0ECmQAUwYIBVEBZPROAip0T/beQ5/s
c11YNvuz/XLQ/gED0EtirN6weULA0m/1AW/5kClVSnbIpGJPpO1pUtwKmSTBbObS
r+cQ/4r3+dfQfyJu5Ir+bZPVLp+ChdZ5oMQ10yDa5skUsBFs4uF04E52kQ6kMlxG
mp7titenFMTbOlmIUk8kyyvrRWrHG6mBJ1v3mSqQhcLsSEgItgzglwK9F3BLP18f
4O5Twa0I+s+m2bQSszlaF4jbj1thffdw5hFeBAEz+QF/okD1ki7tZMkgAq/GbDwd
tin1fs/Ypi8B+nJXyJcsOUMgjqHuvvbACcznoUeQAvTqSuT8y9hzf8PYRUgNtemt
3KjR05EBHw/hTKhMTBoUdoUgCaxuFPmJRrpDF9M/uLOcJv2GqllcB6KL4M6tDQJo
yH0inBGIYYTszxdLHTsW4xF3H5kanimRlGCBcTudhgfSR0nXwMCtsVOL9iN3HUQO
/vy2l76Xm9/jII9RwQcJQzqQ45siuS4E4PgQ2aAvlgE2IBuEcF3uK094aiy4cS3r
gAlvLFTKKq77xlZVOZh5Wl38A6h9ZbCC9M2XQohF7/I=
`protect END_PROTECTED
