`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l/Cr1+h2aoZxErKDO+MqtwpTPssNX296eZE/AgWIYGbgsBw0ZyymdPxpJI1A1ZtV
y0GcAQjw6gvO/hLL9IMX1euDvQSR5yWh7ZAHg0jVgzDYOXZr8aZnhtgjcV+TmxtS
KYtepFJeeyriz8QQU9kQnSpuDa20eUKkJZhRm8ieTEJ/I+1C+H3hYMUr2IjWHyLW
BVkb3CgGTSnHwSkFlIND7mCAm7+qeIKHyZuB4QbNL4D1szBt60xmRcu2IwG0m14C
GQw+srAtAbQYHh+HAp2jPNqkJzOaTWdsHYp//OrRcsKFGkTDAOyVRnP0qfXafWUp
1Xuji1ajuF6VyVNYTTckiy6TxPHiSOBB5DJY1A72z+GX0c0DjChmC/pvXjRmkV/e
8kJoSHamZXxFvNGQux6g7UFdVgnc6g5zfLdYm4sRKCQvt8tevPQ8hkrP4pZuTcBi
fsIoYSZHB9mxtgvvwFleeSGHYC2O6SGKQTXdUJCB+FSCrmS9sPm2cgGtPg5pBra6
6QFSMl+buT66oMwvFSsLlly5M/l2pVRMor22LGPs/t9wuxI0mIm+FwVCBldVwv8Z
eTqx6Y09sSlsq36A8lgtoQj08WVULUoU6Uhwk9geUMQIZS38W1rYD8uiusH7wIy+
dFXwORoZ0ot3c9fO7wltRJuUWO0GYIxQG2W9MLX3FpdchGohZ39LRVr6t0vRmy9L
VNTHEsSX5Ja/LtX0IwSazNJu1OJUsob7oafGNmn2h//H30pPd2MYWkN5Hpi1cKoj
lZhCySHlHqhTO8g0ObAJMG4Omhl1sI/7rUYvIcWVjJLXdBC3+1K3uqTuu9OAsoUG
DfVMNo+Uf/iq/3N4OWcMh/QHEd6XmYOaFjD2Vio/qCYok6d0IDJWeqmUHJlfV78U
nKL9EW6ygE45ud5OouycqsPSYCNcNoNkjZYLI7q63i+JUovrMPKjhLL814yk7JZ3
OXNVvDDCpnHvlIa+fy8a3EGTPKLqPZQgrtW6NTL/9tNfb+J5sGlgMEhLFTXmrHsw
PAkXUmZYlBkfpNtONcozDXW4Gh3bWusuuh+jdu+XiXbL77WN1dyPLncnIrtdTdco
LyTuCRt8nU4YSfibw7lF2ZT+Dxsa7wvdNqnRNpOr8pj7AWcq71geYvcBjsaurWnh
YFE+kaH2k9mnpjziczUyPz8GO1AnJ1Bsk0TvfDwAItn8+5IHJdGwpgOXVrd8Cpjw
R8t+D6p4yVW76aCwzgxcqswzIZqON0Z1vK8kBuIoovqMVc+QZxH10+5IBuwe+kyQ
feLSOp/RoMrXikoPhG/jgjT+E8peFA1Wk6nvlTGsChjuuuh64m/OPlTkNmHlp3dM
ayyT5QTsePrVq+n7cH2DKOPRc5U0VT0U/+PVYaveaL6pWLLTAq8CR57aDQ+Qxzz/
m8cIp2C4PFF4bqNP5ONL/wCUb+l1ic9jI9OY4kKSPfs9Tqtyvx6SQ8E4DBRbP+Tu
/jH5HMw/FRD77viIx9orRSMlf7x7UzpTsY2mVOlYkCNEgfYpWJoD4KssdbDK2zLN
YmTKe/s0m9fAKXZGOGs2lsAu/NY2Y9UUTIuRUwtPn1zuLBBsFRMANRPGfrMEEkcd
qhHZqZlwB5Y421bQ7mbNpE+DWxVgaRBYhc0l0B0OUmQL7JHALz0+wrQeUu7f+GrR
KuELNsJ4BbReQUpsBZKugy53a4/2XD7RJoUrZ5kCu7CVzwb70YPZIOWMmoZEXF7w
Kr0qjkL+fSFlWZjaEQpoFd1Wvwe+jdqXCMeh0Qw5toGwlhLxxMp1VbwiZfEnLJt3
uN4fKKXHJzXvLiKk7Adf6XwrFjIFCE/qjnVLVoQFlVqsT4sdZOl6jkfUJhr7eKZb
brUM7IOuaZwusTcSETmz2tbFZ9rApEK+jwmwTp78cQlXjGjL/h5UvhLL7pY44h8a
4MVn37xo6puIHwU+q6RKDoGViEq2HPaaeYGDfRDI/CBwkmMsAF7Mjy59Jh94fiqe
AkfhpeoTGMYh7N4Kozi+u8kzeh67CkuQV6REPAc9koSjXkhP/ur/fQtGgtD7eidD
dJeD5nCdSM5cOfb4w3XD9AVyWKjHbIPM7fAklGuYfgHbQ2lD2CyAgKgHN6G/PJnI
mp2GshnUH7cIj4hyErt6mpHR6klaFt6JuJgSQxgFp52XhubxagcwzkbhAuWjKu39
zQeR58RrbAtTRQczcliHSQvKoxL1aDdrmbWoD9KIb+wbKpEjVKiumBGgCsayzqn/
6FzSE0lrxoO1EWZq40igrbpdbKUP7xyTkjjF6KYsRlLgfjMixqOL9GnZeeZ5FlMD
WmuCc9mFPli1nn26ZifMqMK5MoaFS8oXvnQYsbd3GyRknrtefmIadap0FOiCwN+3
vz8V8A6TdXuD3mROCGtOpsh4W/7i3vul60wL2j1VpvVxcz6+2Sg08UXR2vUg2my7
CjwN3N3sVdanoM/rtM25hcG3P76/+kuXmhkFPjBq5Vh3/wy0mb8gGb6XSK7QPe6D
Lz7A8Hy5XrX3X2PQXHMHVvp4UW3d1qPZ+Fj+BN+ScA79yJNGuEKIZTSoTjYZFFhw
Q0dLSPxTu20EFe2tLEy77Fk+lzVCDdJ/Grkoi6eGGdntMpckstgGcElL0G8gq/0y
bEqcj+zF9/Dm9lSmzcyY7BO246nMQpvaN6596c0qzMD8Tl04T78I5sWYoLEZlTnC
fdMFcBr63wOV6Y1/z1Twx3T/VqL5Yd9benK3JYdX1OvWBzNE5Olc3egJespLFOJN
NGePShIaPAW/IOsX80V+9pgG5DiH9I2Yi1lgoOMboXA4yuq/qbEUyTPu/xos9M/P
M7OaDb5rYqgBplyYYeewCjtJfeN2Dy6N1VdGv3w6trBALXRdtsc4RMFVJFXNKTYT
r/LNFPy8tRzPzGP4ySQxqHJd18qZ4JBqLNz+pdM0hqYUi0S3vb/JWMTpLZavZpD6
/LlE5YZyOIQi591PiryJ3WEsVN/Gus+5TGOWOp3cm3qXJRXnQ/iqC1KEG83u+vSR
kWAslrAMj0SGd5t48W/8jJgRKN+hZMxOvkRWn5KrxIgs6A+/aG2Kbj4T5QdLTgrA
rObp/EcNpi9iMfjGnl+R6haM53mUxkk1suk/Qb0E6PbR5ywrkeer2urxSNkq1DPE
Me/CxOjSTMJKsdAwj+JcCkt5M31AHI3sFkbm4iIIglno4zjSJ2V5EsUGcK0d078O
I9DpdMghcP6UluJub0YUr6PU++KCuTsE+zANStx7CQceknA2UjzmYLRpc+IgqiDD
HBhRMxRiI47lZVsQ/CGkHCOEZrrtkXh2ct2rCrSEtX8rg0D9E8jmQLXJUgw4/lhJ
`protect END_PROTECTED
