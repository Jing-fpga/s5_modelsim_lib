`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zwk1C4kzGdXqc759YQ2F0isR+bbeqE+kUkPvZSzwoyIogJSsrsTPZ/Qe8kAnkTv7
VsiAGgiXPxMhtwwdVrOOC2vlHt4A+xgrKEZE8LGKSJf4QEHj34Bn1d62hpCY53aq
y2CwvE//8/DzOrf1lVTYxnk453PAW6vTX8/18PalyBj2BvUBtdcNzBsVlDgYxaYx
196KQ86D16hP4bjOpU+NWzMHKBh/c4Chw1FxryAkOG99Zs9il3pDfkWasxdbnN3Q
y3kGikzTGp4XfRsx0J+PqFGTbs4ThGRKee3iMHaZegRRLOnNn6SrXbRtxUuelUGB
HL32Z8IjzfG8n1YUl67T/kcwxWfVVR5rOgFfOYJntcvHu6QeW+ToJ0jTnvU4Fs4P
3uDozGkWG6ykUpMHKHuCXojjsVz+BVoZYEfU/3kO/NWyhHcRTZQi/a60/hOR8M3l
Jx8Ocx49YFgzwPgT+6XyiCmIZCtrzQUpm4mG3ZNJ2HrRoK3lOZyLoz5JoOUM0hLI
a88ClbD1hSdjS1l7GyVgvULcgozz30AcoDkoJEZhRDzPPhO1E3U3pcdTa759GOYL
h5WLl1fsZgcvwBcJamoyDvJkNlRgDaHy+THnkJ78hrG51FPO63Ndw38zFfc+kodv
`protect END_PROTECTED
