`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4+5LTJwYACBoU64btQQmMpXoHDRrDltmTfFbA+SPI6TtMMViBOPrs7+Y+pbuwX9/
a7YIoJ11laGc9ZlnUKDw6pzSCeYKFIYFjd54Oqe184RNyts5Zg4JdICjl5DwmRQm
JwzhHQ6KvZMrPW4GYZN/dsF7NvjyrNrRHdsOIQQ7YPp5hCnMoFUXEYhiLpNvfUh0
3AAyan86Y7I6gkmTVRqOO9K0YmU0f/87WCJPRXoQyjC64++UaqzzqcJagA/1Mjkt
ChOLf8jpmi/CYFZPy7tN2QF4swKt2Z1me+1xpCUkpQ22P5LFzt02JR/Xt2iIdBqi
4HEQCetBmsNz/0QXGZND3SxH2Wj6NFWw+VW4scH1uDovZkPoKcOHHfRIhsZHNbta
3uoLEPeRdddN7DGJVewEAiNRpSQs7sEoDZ42GJirnkO3IQplEDtonCWiInc6EQlw
cNvciKyYt+XRV6ruMzVpZAPKvNgJgPWLX/sJ3Xjts0to7NFwhdKLotEMNLSOdnXO
gQSbJqWI76tFkfefOLAEZ2nplRjNU1ItCdfiIk+VySeyLNK5Xt/+Q4E/4FMM3cJe
gLp9KG3AyzBxUlnRJm3ZLA==
`protect END_PROTECTED
