`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AqLGyjtXqOqJwtHa03hXv/b4ghIn8MIb4lDIVXwCo8lb7hyJFI77LSvRtpoGY0F/
zhNoxcMTyJ5Rbbg+icSULirZ67OQqH3hkoYmxS81/yY5KdXQWT5WZiWGkRMPpHKr
qS3m+uUd+ssTlHZ/BpIf3mBIFDGfw1HIoZO7SMSYbkESQyK8BuUSZpFncsuLo3w3
yC7SImwJspjhNqbJXVftsDV6zGh80J/gvG6rphQldXKVxEBhJ5NAJh1L0LKBvbOj
TOT4Er3IIvO6OXQBybLHtDBk81GRq9prGTdPtxaVjFwMNTk4iNwD/eeoz42ACeBj
Im1KTBzqLkHToN/zuGuX4TS83IPtsz/L9oCqFlr1KGCF3Dw8DSFl65nFQnhM9Nul
cG6hZbon25VQQJoXLhWzGpEFMtUNFRxQc0sf0f6DwYf4NjEB6Vb02nCS7ShQgZw5
SRfTJBXDzIacaUHYmVjc4MuV3CatkVESQUrxmbveq1Cwx6mhxN21AmdVbUINB78U
5EfhLIUkneLTRqQzSKv5MFYy5EIEPJBJn2DY0SuZYoj7X1B0SUuFJYpOfvNzCPXl
Uz4nbEhf3siD3V+Auo7oqQuYA+mugAYnT5Advl3s3gnDgnf/29XIFLq1qgQ4C9gi
qPG66bpfkyCMgiZURV1BO/6uNMWc6ju9dGnAK7cRsRrE3cJp3tlU1rtak77o9gf3
LTme4Aw1ch1/cddN4U8Ard8yiiQHYsbLYVuBHvI+Nz89hPCMKl/V5PabyZM+NZVx
+o4THLnVBIDqWJnnDAxRLNcrFQFFlF4sntuoKb2Vi3TCilVYMZbiq/f2VdkeWygd
KMS39nc7TIYEmrGo5b8QG6ry60wMX99IJE3ULFhHLS06GbZDCBSse1Y08LJDIH6s
PhqE+KCrQZEjOXU3No9lImG1+iWIwxuGzOs8VVsYnllGoGuoWi9O4XrmX8XT2uYM
nCccduwYoKUVe0rtujiSzFGO0PqBK3YQhQ4lJ93J7w/RHLtpi/2rCK491Dp/IH0Z
7HZFfpv8LW7FbeQE/0MuQ9MrEgSNVd8AulE6JG+YU7tVEnl2lWFwUlMxuYUnQda3
P3MXxmvAJ7zmAzIkHh9k3Lhr9AqT6p2GdrxoVH5agebJW0aehHh6+SnuO7MZefGk
oBZwBFbyKgfouvhtw1b7PTQVwuxTzkjjfLZi087oscxJMj2LUTtvsAWUKNf8lmPY
Vl8R39qBE5zJCSPLC/pWDj/5pFsUMWpi7Xu3wqIjNQJTn6P9juelViVRFsLqzBD7
4M5thpCY/TDTP/1AJDwtj3LAs08qY/+pyJJY1Jk49IE4htPoGt8jQk9o47AjpHLl
F7lC3o3Ao/jcid8tnBnC/3C+dx/8ER4DvDkDKw0UBHP32vZtOV2VfsfuMOmg7oZ9
LDNq43uVVC3MVGEtIBYwbbpmbv3AsQv++kyiNrSczcsb8j80opk3mbLTUmz4YpWi
/CJrdFfO6PNbepZxRZt6Ncuz5lov6F4My//1eBew2w/ZQ9xHZ/d4I8M8M6t6hVeE
RyL2Zhb+fcCYXD10xyX5ywiielIqFwfQr90D8mcglzvzaq7muqfzwa+0585TFz8q
lDM7OHgcsTdAdNpiX5xALPurGjU1lqr82EVqU8D/IYEdRR+gYTcE42wYztx7FoYL
Cz6h1PTRjy55I59yyfUuyR+M3e+jI4cNZPK3MvxjvXP+MsGfCbDVBhM6JLoqTssv
BbG2W9NIhIlqFToPzX9LHXUWkYjekBo5ZXZWz9XWe4VZaZp4xuFir31DjYkorDkj
N+XyS5bQRvXkKvj4w06s+KxecvRx3WxI7kQvuzAxfeEjT6ly5oRmrSr89ITMH0LH
Rqk9jiEvkw1f0bDez0wnl2UpCyZ2wUMzl6Bb8U0Qp7pH8pboZfanmsEIRn+v8vPj
E/7lrXc0MD9VgaDeRc7pnNLj/9LrgruupHohG/ZDH3QkmZj5vcH3hVlxMmA1mDiO
UT0KFz066jOMa1HqKWRc2pzU4QfurwjrzhgXIahPQWkbuAGGXVGqI0hvKKqRFuga
7eMN2eQFuWJXsW1sECJQmAcr1FW3Ypdj9UezpDiO9lFJgGSQ2pq3Ik4qV/bqiwAb
7pwWne/K91dJS2B+NGHD7muZhn7p5pixTpKB9/e83Ec8OUToX204TNApRRaUB5pb
o9qRq3RJ5/OHHgl4Biifp+AcoGUQ67/IvEcDfobmoukDLZEUERZtS7C3yJ3PSqKQ
BuBwh791MxwUwR8UGyCMvxT90A6qrL/LQ1Ll3qgn1BpAyUM0vRoXyZZN6YE2u08r
crbYaztIweY/a6bWNJST3hXi1p5q1gt4Dm50ODhMyeGjqyQWtKdWDexX2PrulUSJ
p1YuSNlGwgo1BmN37ocbNr5Lza7X/A5QkYQgRs21Yrnlg62mEsvd/RIOOwGsKbJE
FicbyXDk6Hu1KWmGVjhcNtkwH1wSNbJV9UUVbTucOp9JaYoT7WQ6ReNMOfr/OLJB
PeJMpgQoZG9i4RQjyBEdsgoVtk0VV5nwU5QPZIy+bQ1OCvH9VzM6ifTP41vWvvzL
3wvWHUQOYNY6AzjUpHNrL59OEWJYT5n5Lvfs7Fqt6GhxCMUaecvBCeVoX6lX3Uwb
MJH93PY/k4hDLYqXe/ehAM6O1/KszudBEzHA//iUDXNsKerUTzhEocDRsxBTGMQM
lbbbA5yYMzk+hZB0Z0RKxYS4D2AAubFKM/G9GV9GOpIzCeUN2eaGXF3/fl13NPsd
vDnXbf2NQ+K8v5RNhB2xLTRa9NY7Az6CD8VB/fEXao3MG1D1tgY9itNBdFPqHISm
o4hiHy3xRiuHZhH5urkylDz3MBMQBbFhiX8/DQswrg+KcoJIlIh42enWaEV2vMp6
Yh8+s6AF2zbd2wzH6jYurxpF2N+6OH+uNsd18n7Wvn2VJO90YfttbJCMy4vRWy0u
78h6FJWRlUP7mMOAPQ8Aro60QA2EIyyrdMxACwfUwUZYTmEXfiq3V1gGiWvXXgwC
Wm/6FwG3fAX5K3KvyGR7t3DybABFZvGL9OiuHmreWlP5hIGLHzRIcAu8MbNJV9Yb
wFEBPkfhFD+8D/rTBulouLFLKdgpDr1GUsr8x+xGeWFE64vJ98LPYaskt5wTw3dX
hzPQBDv9IEDPie+FcsVgjvdQ+2ACi7QW0j9qLqJqdQJKGiXxEL853p5vpBbPLBWr
jYdoPOgPbMP4l102Vdq95I/pGCYLUMiyMaLCQ16W0sPDnOl6FmTLhb9T5KqONn1e
lk0YolUDYrM1V2H/ZTO8BSzSICRKr9Njwr12qgA/eceP36cNnJuVcTBCKEOookqF
60WbXs0eZWhu9mZfLKI2bRe3FrMDbIXHeMlrofyKUU/IYRgQrgJXj6G+6fMI6p4D
Frl3e+UzbED1jbFVW5cNvAYBz4VZbhPLWbS9P2PFQ6tXcDKnRRtKcz3i0H8dmAna
lmux095dMGx/XUqJ8v/rsBxNHYXA50mV0Y+jbZyUD9HtbUMke1UkObRiuxCG6f2e
BB7muCllrBF0NuCzI6KkrWTWCuu/ZIGRWC4e9xjB5txHqH0MO8WBm+OS71bWF2TP
yTApXUypVz4TP2xq5D9Mj+2tL31eQmhO0B5IWplv2CO4ogGP3PLJs8U4SZpWklto
/vzISdbZLlBlxvWIgwrS3jdvrhdcewRuRKIT9D/KC1fq6spXOUfOjx11ynEtZna1
oXskqHN552eLYQdtYs8tPUMwh3j3o5eNVP1JYlRiZY/KiDsTbrTt3wD/cKF94z28
SRFOxFeZTDUEbZSVRus+vm/KtMBkxd578/XT/h2nOihOPqwxMuiAYJ+4jSxdu/TS
aRtT/8iMf89DbGEmCYQThLM+uF/MUeKWj9PpgyqKrFLf9TvKb9nyQdUvGx8VqzQg
mJ7upPSDZqwzpRVHNS/76eIztCRSGtSXosdvziO/MCitvfMd1mANDNDZrlGLn8Gh
z7D3IcEJ6EiFQ9BUD5hVDfWlYH8RKQj6zPGN1EEjLfd/9K7TgRrwzi86h+ez5b99
D5/N0t9N8RNCHPycKzoCmBakKxcO3oFYb2Ktvf7ICH2kAUEmbwZXMDxRu0QPT1T6
vXdms0PEI4/1VFkQDYWv4W2Gn10jvYPGqeVVZ7mMREr0hJhMrK3O2YEkSwSt6vlP
kH4ljyiXOEMYvL7LfsL3ktcoJ5pPOUj4H38V/COZze/1YmoXcBPwinP6B5CqFvvl
58LEm3sTY1hUorhJmDlomiFnL3XrcmIGiRLk/7SFKh8JAgUBIJhT++GEdXWu11/P
e6y7k3w6MYnYPa9nCVqlJcFCvynw4aBV/5MhRnVdHJLhqIeyurW/4R8xgrbgFAHR
jkEb4/ufQXGX/VFYQCIY2osYN2YlLHRdiNeVXcndnG1q2/qiVDOI6vMY1hyzT/Ru
TWys7ecNqekJYL6FBZCk8AF5/Jw9ZJ40VYoiB9iGGwGvTVWw/rcxhbaFracEcUB8
gPAF+KUNUyHFHmvnQWSOzTr2yDHJEU2Ll5llx5QanfSyGtUaOVmmv6J5+/rUE64J
wTNXABmvDfRYdKIasVnYle/5K+7nSm+TwQ1Vsv1ghcy0SrnLhX6hOKQXiC9EVQLg
78u1mzexa676e2kXS0vd5inUGIKjd4E7UnJ4scTGskmizGTYMARK58arG3qiSN10
av2c+XR1G2x3m0VQpyXXjg0F0uSvCIScsV2udmcpH2GE86JHWuxl3X1XsGwqwAWw
cilFC5eoAJuJHH3PtpZfomvDcEqHkw27YdO8Zq6HcCh3G1gm8LFwl8mZ6zNOLOML
CTVYDiiJrXhbOyPrgN4j2RD43avYhH/dHI0qPf1dy/KxVMSChJTNhtuNOgNGGL8I
JWqqSLs911QQGsT7e6FCWduP1NaMH25wCpyOYOuvW92DTsUnn1C+fZjj40z8bNNk
p4V51mmEWq4ZZH02HXcyBZddbjjmgYd3v9XNMG+tcPhSDdGxl02ybnkPIoJkiq0E
mSxGMWdRBO33+vFX7ADqi7yttVFs16Bm3W7Olpkg737dAt8YKg/Gsh3PXCFVrjNP
Y6qG6VZpk5xHoKnqRG9tZ3Y4psRNMSAq9rHZScA1kDWqEOoyLNql4d/fAKAV8Nuk
u0P6Cdzobugg4DmJ8zwXIbgAnUj1p3rviMkNKBPVm2f6O5jLbSJtTH4J+Uog4N0Q
oKpZtvbQYbg5SlH71WRK7qV56OEAF2s+xQEIMuHyIIhFa4R9FUnG+Jp13i7KbqIi
UZ+lts+wnFwu1GfcQ2nteUcTqa3ad8DtOMF7EX2wCiFwNRvGD+VGzdGKDPs31It/
MJYVAzMdf/BdqLn0+KNKwcbGBuJGEqx0+69r+TVm5JoYYJgybJUsPwL3XPW3V1kB
O4U7v/JI8XIxhtixLtOyfqH4yxTs6KP9kIPCLKjoce+hVkkGRV/1ktYVNn3XkMMo
0ul/Ytz2H/474bkuLrPm1w4AHKxhbJSRzD/8LzEaCqVmPNjnoA8rB+VEnFE1fCj7
TGH4d8alvI1RGuzaK1Eb1GIReu8TuXU312aSertm8Sb0JlrtUwKL0gdmyTfCJZzj
Qag17jza209WKYv3zWwwsDvm7DN/czuMyjkfNb2k2qf4z4432uc1aDVw2m3CHUsp
j2/3x2D0hvvf4d9C2oh43h3nwearmL/uUZv+zkO4t1FnkhZtNbNt6Z2kw62ofMZZ
ZFAFzff++eQYJq69ItGaQuhWPM5TuJF9WZFap1ANYPYbA1BP7rPLm5BNq0VF9I0x
f7QHoXPWu2dISB8zPS7Za9fXO7GutJoopgXZxkpVR72Cr/i5sKOG+W18V8XLV30c
IdpHv4y/1WoOuu6EAyuv2F6EK68Db+fqzWL3NpmgxcOm4qBb3U+nXSDah4lIEG3A
mdcqSIHXvTgytSU6Y+WszQydRUHy6vUaJB1bNfthg6N6T64BDBwxwbTnCe3w+/R3
50CPahAg+4D1AgyGakALZ6mVuTjITp7GjUsmT5E9xW1fdMfmKq5dyGKbSmUFad/X
Z3VYBn81XI0CmEAvOYQL492T4iTGP3FvFBql0xy6Z2PHiNNhtPxpi57KR7+mYSqv
upu/+4jwOG832ATbWV1SKajYDFmf+2JXNxK40fs8Cq+BJJHSNyQdhKAunleTTyCs
7VEH9cffGRXAUOD+kQGvhkn0UpOrUhcnJztGZvsfkl45qjWhWFDkzb8MLHna8cK2
zOWrmp3GDs/0jj2zFzsz6JPjqKUPYFjhCnkmKGZ0KBSAeltbtxvSekXW4t1ZY2h1
K+Bxa7QD0pY+EG++phxYqB0zspbZJkTJ9Rbu5N4+1J3oMT4q6c3voWw1lmEgd1WG
845CBk2+IbXAanfjBDey3T32bTXjAcIj2s2jwOrthMoKg1ETrAf0htXAB6Qv70tl
B5d8ku/1ScAN8Nzn1FkgH5XQIqIkLm8zVEN6ge8DNArik2InqgYznuQeFJ8Xkufj
lGjl7fnlbB0xxwXqz5VdwoYkh+A6JnSpakvVeT/7bQ4hN30l7lzpdv28iRF+gaF/
Uu2C6oI+UNWFoO1nKSB+iRNDZz7HyGX1m/kqjAxopgjYqd5f6ch0fybpxkAsbfor
t3+JRR90tMYGx6Ki8ZahB+clU/MAvlUqvwn5G8TtFIYsSKve/J4ZxpyCjV9wOq8+
G7zFJwyT3bnvCwujdv9A98Qyy7pqRKdvsdJTwf8X+9uBiU6XEfPwxydnVRau05Fo
daOCKdDzvxyNKjPbpnRBe2XOKYHo5lYxQ+KxZ9cKm5H1h6i7Vc/5zLrf8zpw4u81
I/zQuv9gpddliLo0zaO3NqGMVXNLefeodZKwYjUplLiw8V6Vj98cd7iyYCg6qW7R
MMZcsfhq+/6eEJEEBxbaO6ZjpGbWrbDrxRLasbhR2mUy0BQqvkYzOiqidvvEoIQ1
MBUq8g4X4Z6kmv5z3LwngFoe5o63LBSibFoDcK91p7rGCfLewv1jjxB1Q8NHUUvC
DxdlbYvO27/MlPn7sPKHw1iA8FLbPRDnDA7pyqoTUO5TdzLaJSklDt2R8gF0NZuw
iSFN5Kj9Zrq+iSCvjhpvQ4NqRsqCgwK1VYoS9EO0dieufWgD31lwsMZmU1r5Ppwd
Vso5lLrJMNtF1WJL0UYcRfJqNYFaSOuGZfHJRNbrULldRv312mWJBTFRbl/65N4y
fs+CoaDG5uMetc7JZmBWXItjfTJDBswD10gogappviyzzEDqzhdCiwTaFHuCh45b
4GC0GaB5J4YwqFhofhqew4ZPFd/hj44KHvqVRDK1U5k3PmoLcnUnUt4XRO6dI8B8
bgC5YScCsT14wIhCQuwHGAMI1pG9f9qcbFbp3l0BFDNcd3XdxA/UlHlEOgl25fin
w/CiSaEVm+aHSfyoqZ25Mcw1jhSXLAdVSukRZloQ4jpo+D7146DR+52vUdj7wKUn
jPHdIZK65r20l8RyTZMAtm3yZacEmB4euv62vqhBItkFpkFcu/YxMQbu0XpMdHHE
5aSo30gfnX/Nq3PJm7rcFz7xJWSwpdvFfOlFNt8gV52om4YGOlLza0HNj1OO6Fmu
kgId+2h874tsUeMa8EsmoLPUJG4Pr7n65fTNehJQXRGQYVJNqayk/Pnb92QI3uVx
FBKfaSlymvIaZrvkQVeFecn84HW0KVxafDBWZeHQLDEV1KqVnJQ8JTMaXsnWDYIG
gslT/Yke4w8WNy6/Vww4N01JqqQ+qp2S1QznVmPCuf6WuZcUTPeqjdYd1dGjAiny
/zk4s1vjqkwoOX2taLsvKUxpCoeLZmEYantqFaMyhlsoM2dyXiIRPkjw4c8B477v
B5uNGpnLBBpQoa3NhWYRTYyg65Yi6DrIxnaE4xfQG0rXRtE2nsrpK05W+Tdbz3r4
j4kqqZkH7lXBmDqu5rePukSxdnBevqY8TSU8dGq76NoH4KF478y9z1WfCLH5XDx+
AcILLWaZwlPUrwFeLQukVc4V4Qv7OFLKjME2l3DvASrbAdeZ+HBWFC6DLTq7a9yI
Kz1BYvmKxZUIxO1Nl5jfydnp+CrLSn/zlycUkHQkFPZQulnKka/8UwqmLAoc0qz2
sRSezhXByxy5DByRlFuTf8KIx9H/wb+459KrlbUlN09sixepsDk1RUtnIYErni4D
vUyJ+zMQUpz8FAQ4OhlSWMbgYzqymiUySFIxReflD+MEzc65Du37kDXQZrGkSFEV
PpkEOFmwlX/B5/sjwWd4NLX5VCDS+BnZydhQSlQyBX0=
`protect END_PROTECTED
