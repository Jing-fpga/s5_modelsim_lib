`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S8Oqs8hJynCtilf3bVJTsNj/A7qYD+lEcqRFLdOMJ4JpWyQA4qGjdTy/IbhbLVmA
s4iH5xwxdmgNvr7kfT9biQVDhmhr6eI0G0Xs9OrgJkSGyL0kuP5bJYmr/jPXbWYq
FKBMB2wWxTG1krNBoWH3J+btYPD8Fjd3pYbdhTbyI39giP4ew5wVOkbWiGM8XxiN
5LIYhznfviZC9Kd67GtZl+EewvYV2UZUnPaGL6gtNAWhV4wABNQmiNwow1enwT/C
m0eumx4AQApO3zWtwHaAC7opHAR6T/Np00mPRphUIOlflzTQup/zro4eWx/HqRWc
VyVYlVAa/s+VdKGHQbczOxrrrH+ATVM6cvO26F0e5lv4YqXlzbNsjDXys36vnmoY
a2gV21GU2cR/cQkItsVcSnVecSnqM2495CR07lf1/h5rqHpaIpW0F0dzj/GyCasY
GV0RMIB0MGR/YoKnRVH6ztZy6geD28mD1cEC+RtYalCT7m1q8LDKTn6veJT05BHk
FmwMvtFVwrMJUrX/OflTiR9FvnxgsCK0vPTJ2Aix0GfF1muY3nArPLwYqD9r/jac
OkAuVyXMu6quzMvHT6LuhA+1zJvT/sCh0gF7igeGL9sT6J5FBkQy6xqaDj+i7a98
+n9S+fRFOIOnlzpQLYX4mAicpG817ZV7H8PZp4GmMPBxDiv7GsvTEd1LnYZ6/Lba
5DHIm5KO0cXsgoqYNiE1G4cCUdKDZcG2hYsRTdrEZGHf3n5ORPCs1nK/xF/s1NKI
JG0gh17GiY5iN/brSgPYuFK0bxqj4AcPJgjdZqlJJS0v4ye+7vriLG9Z0Lp291Oe
NF7ASPhlUHFXRySjSi7frAVjpWVuxv7DLdjYe2zFywARg3qE4jySM5rp4XE9NfDs
Y7w8TPMbYLDdkRSAddrD2zC0oRjRbGq/y0AOyErFbqxHcbieeWE19e08PTCQ1ePZ
qAfO9Hdeu3jrIQhPYc6u5aOtnx7QPi/289pCL1+pUjDc+XClonaobEu1m4b9VGGg
vWnIKhIbsTUP/tRcXvadmROsP/pcv7Mdoe1SKfVic+o=
`protect END_PROTECTED
