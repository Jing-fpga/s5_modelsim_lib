`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GbqhA47SesY5obvj8zI+59XmGzlED8VruMS9aNhwwM237Qx8t51ybuXlot11JqJN
imd2cF35riqcAx/1PRlADzFhP/vRLWhLdgdVCpKwxoxNKSxiTzFwp+1/KXbfU8pU
dIH+FtZ6hKtr+hN64rvbYSM91f04WOEGi6KkwzpZ9oDpPw74QS0sqgjDHRsrUXMU
gWf7QRSQA6oDJA8/yh3FPz85yl0wfBTogzQwMMGjnqQ6Md+x31Gm/EgiH9JytVtk
1WV02OqsHZ0zjT7URRGNiTtq5jx776CaluD0mXeMNF5H4naQxOQNMmhJPvU+X5VD
2RRKkr7y5HoKli9MOTNvMHoaZ/pw0czkGO3G6yHj7rB1Jc7hhMRgjJGAbTJ3qBwW
s2HtGcv+LmrsDdGIMj2pHKX0jV1Qbzm3pR4O1VVnR/3C9gae2/z8ztV0tuWw28sd
HqYzqMf7qBgM5RC69BTxbRCis6xjxvWMQzz8bepoXv8hhaitmLta4pWfzE1ysyXI
pj/C7N2cp+we0G8uLpHFoqOZhBlpR6IY2tts9TT7D/nNF7HSngD4kEHI8gSKwDg7
X5Efwdy4tktOS6bFJ53zYlSmGMDvKaYBzCraJm9kDNCTbH0El3561CnMj+TyjvSd
MP6CuFDEKDPLs8ZW3zzHxQxXw+vw4AoN4XY4XuLrI5nhryI8X7v9NvZvYx3rg/rM
xVZRFGV1YaYfWbmnJZc+lPwGuBcfOfWklcej2KL6zTHH/mMrUJdhVHV7drPVqxxU
UKg1Mbr0iu01eYOcVRPPQBwR0r7+GLwarjAbwhpcoxlIk7MO7fS7nZOvMHr6WQ10
1rjt06l/CPQahgQJWdK/cwKVJUykEM7b1QXIJQPrclzZDgNIiniN8Q09emqkqnDm
M4w0+B7tEbabd/98IEwLEzVXbp3S7nnu+u8gSoHLfV564vUAocz6lFE0Q/sMsUKW
oi7ZiRnlPNrMenuxqo2LTtsXApGXvgxuOra70PIE7/J6TSNYBJonpr5dzCJVxlIM
N9LyuRuNWjvNMGSfCgK3HdDFh30YKHs4tT8PgJQlhfeMCt2fCYZA0qnFzhAjLFnP
X4C1rb28sOTtIx7x4of3m5Bo6JzTy2iZeEWwaGh/SaQI71nEGi99Xiv2UTCsIpKN
sDpQyBpDC++cEONdK5hi6269YSsCEl+2UsVoKCDnNf/6+q9wEdq3mj8CZQ4STYCO
SSaarXQOylBG3xt0Bv+5li/o/rI8h41F/kS74fcdzbQDfQWN3OrDf3wuscS1WFSV
H4txCU5O6UnQm2UnQaYiqyHKze4/u9Ti1BqopqYop6REUrkxyHjT1f6xPjdL8d7J
OQ5jvNTzfjw9lLT2f0kydvqbeWDgypGfnviLOyGJWaOQK3UkIzU/ryN7vyMxPLs0
o+gKeeV+wCpVe95aNNeGrYVuLNFNj0undpZ1wbFycmVmjuZpEoGfwD7CffC1FGFH
l01J8GYOxWZtyU6jsWZ+mzfNlkuS/ewpcaANhgtVm0BQ464Hyq2l27okBL0Eyz+6
bcVv0RJfMi9kGwkHIlKKj+efjSbeyBdgDDfa57zqUdZ40d1lRbgWF4KLl1UhKTg9
Up4AjiyBhbE+5sNmg+VKM2sA1a6loGQMLDpf92IygPVDhvykEA+HwF+ERkS8RTyO
lGbfAlCitq6l7rnIGlr2UlkjsFqaGPe2BZhxV9n4csOSwXEQT8W8EBhpZu7ZngoG
LTOZZQljgaMTO0IUqvqBoZozE3EQ4ZgtkECee4aP/SfEXJ//lCq8JDAYd2G3kWpb
5YgX14OIE3hy9AwIHqumWiceKi9L6DCXokjRDJhV+g1oY6m56wgPuQjdcxBEyb34
dpCxpR09v4kDj5/dYjv8v13iBg809WeFiYcSsTeCA9/A+ouqxDZED1cac+NTspo6
5+XnbOTf4kvr+Psos9gTVeiIndPc0N2dkxZFr7umuP68lmWjC4xYeGLzNu1rV79x
rZiT/MB+Flkq5sTyUZTPf8rRWySkI3oMHO3bL+jM7aYRTnI4BwwxxPpRfzPOw/U/
qFS2+ouHysbgDHfXIk4nPV+D5IamLZv5dOmgMEYY+mOwbnzzY1HHzFcqWActLuUc
rPADfjTgSxmuryEi6WLRSaLwwvekMOzv5mz16qCFlKkMq62ZMoZh1EzBK1ArNYTO
f/2HdnrWS0jLmi49PLecrHoi6142xVE5AeOfhsrjMB7lZ0PTqTUl+q3u6FxPnErH
enuLLHcfetluRjR4e3xdCicaqWEEx4J/745B0Xm0GoYu0cVerGrLY75MrIRhDNez
GRY2J8EmX/rbKnIbBkwxL9uEmjGftYhVo744wu7mX/g8cBWYig5OA1KAyNlAqno7
EhIYRdP28yEOcpWN8F5mirxjuwHZEmbGqpKtnGiEZjWDaYAhufKuzxOU3HZHOrNy
Jwi2cKHgpjDxaEvsezWOW8fht9ttgqPm1G0FzecVERqnsYgHjpt29/Mnj+nXorAC
ZxgXYVGJJsAOsr3Io14mgulWc8k451aYAT4g+0MbOz87I2xwCkoAuPR1j3OESALh
/eOFYzYMS5XlKUbf93zkTht9OCTTqIDJPuz+Sojo+FrLBGsbipFntRSGfNfEFwq7
c5A8PAxKWPtvwf8QAQlxjBT5aFekYqVo3Q9Q70Fgb7AT0m52fsui7n6zpyfdW4S7
CDxOIK7rpnuYT4Y8NA0tme1u+I2u/qHqJXXs5VyYy3374aWYllFSRyw51ZYuBmLF
bx52zrGqO+A9jfbpsJDIhnVYIvWYCJtL8ewq+oyH/hB9uiuvQr7pDqFV6P2FYwdu
lvzeexDatJNoiQ9zYc5XsLOPR6BxLe/g1KlG1cZAuvBVzrbQzlOtQJLTSZUyIz8u
Jnp4O8Ijc1oWO39Yq8bk8v7f+UpEmzRm8gGVdV2eozHCKdqWHXlC87MBiDB0fTmk
RGnprzmRsooJXpe1Tr5+qcci8Kkj5UkRG3AmkZwuNX5Sw+UMgoRcKouhpihzEMzo
wvrhBK48jjTfvFP+54xuh6TVRxRH1OxkD9i/u3yUx4A=
`protect END_PROTECTED
