`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1emtOXU1AKP46cEwjDjiOZHbSffXVKd7iELgLdiwrO7ikQquAPK3jyuaFrCFwoGc
dDCyVsRdQPzglCviZC1jNAKY/gjym8TBesRVAoqmlb/IFNZSuS0pK2+cdAPMfHVE
W65oVbAZ7jametqPbWkYxLdNq/yhQiO580exUd0kO3cEK5BEhJRHprfI4Y3w9NUI
7Tj7CzeoGcBuyD0G1u6Z6vx2WjdJI4nDtOyOqrQOt676C26Zi+TETiuNCKES4n9G
lje/afrBnNpHwJY/t+2j4hIpg6dnx4PF5vRNOFgRhNeCdVn34gkZOy18gqwmfpBj
4/sMX2akJUtKUd1owCm5nSjj9B+b6VXwTGkpe7uYMy7GQI6nSToLuS9XDdTsc3Kw
cYzZG9iK3KsFHyGT9rlwYPpV7jcBgb3sZzsWjZImocBLiPXocBAOMTaXgrRV+K1s
KYaWr8kRMt9cCBIuGYpv4AAjNE7Kuwb+VnOWOLuz6FFt9Dpk9SViUNv4qB3g5LPX
g8jtjyCJfCi7z5nT11HUYDanBsQ0nIBn+t7BgYURwdfXnJgMR48oF7uxCJd+Hb3X
lOgaRYpi9sm2WadZQ/CyRc1lqH3LyIDh0ICQg0/YaaPVlqmBPtzPTCuCSe+U/+Jk
KSKMQng5lD3fii8n9nShh0/ocDgBdt7+5ZOtynjW+ptiFSQswmilpRXFI1owiuYz
4zJxZDjqk2UzvZlUwWWUK6dtY0vOMRLcGboEVDlEWcrDgGU85mnezoGFKShJZA2Z
`protect END_PROTECTED
