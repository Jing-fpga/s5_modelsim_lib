`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kcMKpWrzx+kLGAISnzK2uwLLwo7WryrCuqOkuh4Tf6cy96TOSyZmXd8DcoLb7/6J
R9IX4ltcTisvNSLXjWizbQsMAlSzfmNXGnmA8+qW4Khx2O/VY277vxIfAWOD7rgN
W5x9BSXobQxpworGoPUm/EFyrBSetVigb7qdbS+tewk74RX+zhkvzabUuB6GSbxi
nP1dcQpOuwZzlOXCqSeEwhX70JF5EUyP1r0/LSumlZHX1JQDFk3nkoWm4i3Y7oZB
FhF6uyjQJVmercfP/fOpQumN643XTTZu6GhWvDq6J88/9hGxcqUNbes+n2iIQXXS
UlzzqgrMorAfSmIwT1yroEJxkQCXUJJQucdXAyH+aHY3tLZrO7a+ooYcmMOo0ywM
HsC3ao6Brt/oTSrQ6+W1xX27n5g/jILSWOb19Wuwm1B/OhMjNap8UJeoaAh5EsGf
scpGYE3sJ19xpYhK2+ZcH6nwVIWxrkvH0CPcsJjOMi9FUe1f96czJaLOAmpeh8+1
B5viNU6SLCAsLsL6Z/deZDViy0Ixaq7JVilKVwQXPJF3mD9IAga9duYc7Yk9ltJX
nO+S0KKmuYWB+tJyeVS4sw==
`protect END_PROTECTED
