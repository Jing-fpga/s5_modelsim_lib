`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nfgmfp0BKRjJ2iFhkej4Xiy2EKvgGgFhTOy2lWyRHfhLWPwGBYN7jFXEFE8r+IVY
iRz57RiIV7PsdSSMCPFKZTHadoN3987K9wNQIc+cjCUDIkUk8WjX2eVsc9ysbHs3
iKj3g93tDrU8HxCSOMhA6tufKnMkocS9sZUkAKd6xdiQQaiUf1CFrRTsBdz1g3EZ
GeZLxNB55VbBoYoLLpfw3g69sa6Qd10PspaTsxLhKBwvLTA9LeiUb1gYqeQMgqCe
Ep8VnONV3V8NtBv+eJ0MVhI2pFp7jfryWYwpCtG3mL9ISOilPFLDhD2WnnIYUvdC
5UlHvQT8rrA1qOy11W3r968u9ninB+fKGMBo7jNo1neX2YRxAmYXajD0eash0lI+
mnTtvRg/xlVt5mbg3IPpk8zgse20nd4yfbRUKUTaPfl1IMcwA9lF1LxWn8EDTqng
t1wUXsfZgo3DFf0CjHq8eMnERSABdSV+gvjutoW+Nn1Dc4BPAEFB26WbdhtwOUHw
TIhnBl7B6zyjnLPGbcs3epHyTarE6Xjp9bAaMdYHq3wbL2PFH6Abq4mvuBZywSL9
xvYPzyBiWbqhQQZEMauEN+QhyftgWDSfjSrGYuqLreNgu2+xjBrryykD/C5e0Smu
4gXlaanDP6ibiY45FuyzAS02C3d56B0x4Htk6eq6gMQThcxXw0jBCa4T9hqWxIP3
oY5diktRDx3CZMoiBa8W8XDWFDBaSkxONnzsrMKSHAPa3SarMPVf1tGwR1Gl0b0t
I+h3Ca0dPUk/ySKFgaAr7FOp+ARkJfA6hIdGzVub1c6g2omAGOnG2k9lpPSVoE/7
Qs/NRXNf+TFE2pY667o/iNCXN1A1ILIuIByfYqfcSXLOfWXww0mMAy6J37+sXo7i
cTNwJpNNjPFbjH1K7U76LiDxpXT0I8FfKuB7YGqu2BOWxShVS9roHu45bHZf0kBe
fUWJfHDXFvbhk5H8Hr2WEEY5SS6eQtYtuWF0lmsB7k7Bx2SGmWv5x9qSdZEZrJIh
dmWonRppfMCE7udVIAWSuzFMRBOb3F7R4/56RPwf8i1GyXBnDFxjnQnYZraQEN44
HXW5eoKjEN8NJCeA+seRGjSff3dDW/2N/L1KB55k1T4otPtGlmpcwfp2Ibfu1+ri
/t/rMugo/tFHWVrcsdHPp41uQj/sn9q7KTsfs13fDtSAAwuBV5dIVhIH/gRZ7sIH
KuakLlqg/SV7rkP3IDNQhD/7/2ELaGNfYSpIE9FocwGY2yXcMrUsU6YXJDnKtyJ8
JHEn9xhicQH0HrJrU5onPEVjr9+qtnk8aWEcMr+jdKXWvNJbFrXNh8t8tKAW7qjk
/mwSRj5exFyUAOiOc7I6fDj3n98HQM/i31xGK/jjMJWG8sEeENTDUnll2h2UfhCn
LBfDM0pG1cRL6MW6gcB7QxED1EtUrsDeVz4Q3OInTrkwAhyEzuy8Y8U4906wFWYf
6lL+EhI8brw0PgjoP9IFW8qG/IpyU/02nK2Q7E7WVjd6W5Lf9CxPiCJ6z3MZbifQ
sr+P3ydZ5mdHQWWF7nfXxxk70vrqouT7ytjWUN4yINPEDOOuJQSaKhJeKf7q8ZiC
Fct9ZyD9gM5maFN8UfWqsYbauLVJST5/ToXPeaT13MhvmuxHLK1bVPXdqoKj1qIc
/MEKBdBt/ORY6ki+DiNIQ4aAlutyjKQ1ARnNuFp2uG5Uc6VpgxW5sQuLBQS0dSTI
beC/k1u/9dh69n+WtLV2VlWWtallz6/CDEC8pJUdK33foIMVpnsSdXwauYEXxWLj
xTW2kDiBdXUtVSXFEX8Vvd/lYOlxtCPv8bZi7v6wCHjAQq4P+vzZuccZqoaAYw3J
V68IYfCEq4/RFu0ljW9yDmPOZPKrQvrJbDz1Ih3Jm1yEKQlqgwyVjwJ0Jb3qgwtB
/XsJaP1jWMKBA1Fm7Lm2SvTnHAK1vw6tQaokICF2omZI3mEpRrdETRnKRZ/zTOCq
nAbDAY29ysHnbLzenZ1sniqHHjkITB4t796i3XmClTRJG2KxciH6jdi47mzH1PBH
S79R6VdGTo19OTD/au+8uEc9WT/vMBmYaVdj9Kmej2lm4tlJbYbHo8EjnCrzESoG
8JsWNJ4d6iCseO704S5U1YLk/0EFbsZ3mZBI5JkvyNGQgS1GXHq0PCibw1RMF2l2
UmZbgnqW3U7M48hK2AIqFumY52E/yM+nPvow2yeUhO0umiOOe5TKbqwKGCE1HHCV
UnV+JBiEuRDDwUQkzITDK5gkojkjws31CLnlDP4rRnG01giJimEADX79mpRzgr+e
I21qpDUHtmpJw4GU7yITR4eowwBoucMbWEYxmN6cZwr6O/QJYRobALJpGAV9ux58
ZqHhX2arC3csjz1gZ9WDnyBDpbDtPwCmVj8SvPa4SVli0F2zb28jK8j4p853s+0Q
tyTigo1fJe8WJYDSs9uFUm8RHUmXOKriBGYtJWglOlj1q6ajrMG6GgTpPRIKRku1
r7dCsyld2B83SPtMlHnF+5DnO4VsWNqsZCq3LhI/OKDMiBRStH4PSSzE+m8DYQUT
AqsQsqjdSemJYCHnLGj3JycLi33UVf+Lv/QqLiR7pJa30ke6CFr25iLIydrf07/S
7n4gGqkt/171JQUXcWHlmScVPr2ls19mzxQtFtsDfDHNHOoe6tqIqGDgxTmy/H/t
THC9ay+d5bRdxPNV5trwXQBHRRQbruxsclKB71HQaB7xQqaP95lvF29ccYfY2gMs
wZVCDRY3eoKa3lImNZiu0pQVxC9eH6Atm7OiPCdlg4FJH45nwl4hi8b4oxAOTTq6
WMQ0v8l6o262IexDJyv2+IT+PaA668HDrQSo6jq1CbqmyG+FdyF1znklE41/laeJ
a9ocbh5/LnlbVRgBc6+5px7NwRWnG4faejPBfOgIenFerpSaRM8x/5l7sl8Sjgrl
D9TtQMT0sNwlVLcDLhXS2jYhzfR3LikPjjh3a4ouj/lkR6YyLOwEUfA/JLIUFe9n
YdvmaDWcy3wbhJMDMARY2+jcgBrkU4xR9Dl6MBSTgXt3/xVF/Vjh+khNXYXKPLfJ
qFxsFiXL7nuvpxMPGX+iH9FTRJwD1R0IK83CJByTHbtrdaiPFtPk77/lSwW/EjAi
HmjcBuE7H5DIMYlx8lThacheKCBUotE0gtFzKI1plA741xLbLWZuPAtykopw8xFx
piUsR0tmEiwV0JTI4A93j756hK6Df0SGi+0mrJFl4tDl5duV96VVBLoJIIJthopD
8NBW+az5Dh/5X8RXzDfWAC7uUmIG/TdV3m5fkRMkZ9Y5V72InqYylg6fFzXJA/e+
/vQ7yNgMGw+W7cinjEqDRnBC3MLreL2un7/TuN63aB4EuTZsHs8u8hugSOE6ATrF
T1gq51kuKA+ckWWpczd0B9zRAgVOcCOaI4RPdLptK2LU6l9UaljSqnyv0H2tlC8w
KKow3fIqu1GJpPFEzb97zmK+wDurjb6WAltG16JVtrMODfp6o/ZKm7LHwVxIarLm
IAnHEI9V/jpa1mb8H3RxrblFOfWnA0DnVM47VMIkjprki0HZFVq+cryRYujz2nEP
7e4APa/e3LWCsa4+UcclBzCCmdmd1w2/RpzUBbjhC+5K6DcGc2RJtV0a6NHJPcv0
wEbsZe/ZTF3nGgJ5mP/lgy/GRI+zdhrGmx7A2ZC3XeK+jEQUpxJpDMm4bbLewE/B
p1mGIHARXfEXMOHb2hUWJLLMG5h6Wy8o+pW81HsyQuW59Shm1a461Cx1tqEIzMyp
6XiKZmHuBepHW0gM3cepq0NMbv9xQ5kLWeuwGb29fjLn25O/wShc9btsvIXhX3jL
/n1ojA7vj9Nryfh+v1nA8equUsrGmSAqDBRbRdG7wcyq+TfPgGDl3/3hVRC0llvf
PEbexD+F8dqxgRRrvIezdjjI61Qk/EdL3btDd6lgzrKI7FgQ1oM6z2OXHUW9ceUw
1nd++dYfv4+1UOfTCWNPWUzaKEbkgL3K/ek+V1swH3rCrBnKtQZRJ/c50X32cmkM
57ysYUdaqYa5j3phWn9Z6xu6DqdeaWaf6iRJKhtMYB6dYe81w4cZSotiapHzGbYM
uEYUxUAw0R0Ixf7bp0ApKAH2eKjDV5gsrol3POcU36IADQmkzH33TzCqOb15W9c7
h9fXj1QdaJiW4xVnasK5DOcFiPellJREg6pt4EYbXMLozmFYrlwque+CLE+yVmLE
eGFV+5HHsajAXSNuEtn9i3wsoiIYquQeYxBfsraTCJIJYEkvN+0fzT6dvLW9HEPR
QYGTA9uSDOS9X6qCJ5NMhMypZ5bq2IKkIAuE4eKF8r8C0OBB1AEhp3pbYnSG537E
kZCWdlkmuIQ3hNnFX/VGhVdWB6NxAv/Ld3msL2ibI9YRg3vrMbdKqtMXZ7mP4IpB
n4Of5gw83Tua0KlXinbxYfnkBjq2PgHKHXmVG17DGB7jfhP4ug+v7PBDSsKxzPGG
nTeJ+NVFROs63CS8d+5IFXjQIzk+qiBtYbxpxarFPzSGrZJnQcmAaFI3tjjG/WuZ
9TNaKhuq4cL5bugJYgH6LhMstCESAzCWwwRHqt3V16h332rFF8/EBxD/O0u/CcMI
YS3hgTtZx6T9rwOrtdL5UzAR3qg/EJQ2S7u8mjFkS0Htr1oomCOwV6uzLRuybl0W
6aYuRDM89lrtu30M4Iq1l24p+Czgs6VhbsFcYJxlQdN8aQaRldK95FkqkoLgG75u
k1uJLU8zP8759Yz2Czjo2guT0t+5/veyEPFP3+YDSNxz4QW5nPLc2cghOacnXZX3
L/QxPiQBt+CssnNMph8Kxr40YKqfLN8QCbPzdf28UlQn4onyubUltJZ7LoAsEuX0
pAvJ5Ye9aC2885JJAN+4dYwK6ZTTrGox6QMMWEV2AZBmRSfj+dtPu2nUUeBqjUW2
FVFygCrpqLMhq2Sf8N7Ctm+Y3nRd9Mrzfpgi9wvKwnLiIINAkLmzm8UaZ5BQ+fbJ
gnYYMcb4wVBdHYAmoKt2pq8kV6sW67iQb6gIsPVptZtdg1I/68yN1YXVoe2O6OI1
y5BsIRAFy6WnvJWAQwfkECqAskGZlZ6159cMQFbctrXXQB9cZPUzitwZBxMZtkcp
o+SMOH5eujtQ4sn9h7eJgRuSWCTp9oixVi4aEhLpbX0RhYnGK1flFCmAXF8GQYJH
gN72zAkXJq3WDhe0S5QtMU6/7lA/3aQWK6BPeVse7YtulnAG1K3ADFB3WKdMCNNJ
t8PiMzNmZEq+J5313j/F8DKSBvJh4qpgzZBEe8PovyHH/yTL+oTld5tNVwoANw75
LhQmdEBhZkY5wphr0cQEPVOVMIOSefCibrHZ6IlN72VJouEWB9Om1e8xcLNjnIDL
/l43TH3/Qa9nuh1vLRrONQixGQvr6Fzafx24fNZrnYYjqrPiLVrJBbdAGnYGmgAW
rleC/RBh9uTgaa+8p+G1rarGl07033NMM+BlgDB9MdjAzWr9ymRUTy+m/dEgpIM0
dApaM8qSUPxr915FURPUr/BrrYFoWr0kTDryRtNdXXnmk1IsU/TOZgDE5AjvCEtV
zEcAjshvLQfpX+I5H7GfKyj0+tHq3RXHWNg9hJpgU6Z/8kpyPwNmLOKpOGTpcyGo
ITZhS/dgsZtzOM1jZvHRkXDm+MtbxovsPtT68zaiXAVcMk7T1qHVWkzwvn1IDubi
DS07PNxIWy+T4E/5e1K/fNzm1YXzEPBVHJt9a/3Op2BVWQYZcdtmRIJWwKivhjR0
ogQ8W0AlrITiCQNLIgfrTXSVFiAUuaaJ18i+3GVDg6FLkfpa9w8MZkhmBieXgRqb
sDrDap3uw/MFIb7wOujdwSEudH72MNTU2SwaEnnwxZfc8mxlaBzbPSzS0aHhme+E
1ippNXcaAkLM0HV7fsl5bJIXVnqYdXuWbnnZytKhv988A5WQbF1iKnafnNKiJccD
uVC9MJqmFwfkdg5aK7T3X+8ddzrI+oaOUJj6Az+FoV2ZoC2QbtdKVMH5dpqzH10o
+pjJ2sF1g+0wzlPQ3wA71W5YhpAXBIinh0PHWZFmgoqv4/+YVvZ92VJT7yy3Uwc1
l2oe7HyHrktIe8q4JLhbWesRnIENX1RK8ywVYpY9C7IUrwYRjLEq22E244hj1vp/
YfRGS0AUGClQJ+DhNRNfXHnuHNDjMdDu8G7Gh1nMI/sXUm2i+VXd0Y0SvmAnVgLq
pZ3gbDKZ/yT1KDf1TEbgBSYAu22EScenu7hhnmJfNi8PbyJPV3pEPadnfxuKTHww
1sIJKLNQTv2oizGQDImHRKg2icqVOvvEX0iQ4xHZ6BuMwnoMMCKXcoevVCTpdiKr
QprvtMwWnaU0f00OJXRC7OjC1MOmeE9qf32eC5DqzHT87MOvQZtIg1FoPUREZS5j
7Ozti/QfHlm2LfKb9IQy0rb/BJsT6qbfh8R4L6mpmYT/0wEjHrX75e7lDTM30/K0
0B9uj0D14nPvQNDrOVo7oVd1U1GXCyZZU7/kWkyztnv24mxDXFZv3JUSe4UDIWlM
/8clMpnSxRlwfFDt3siej6fdJVJyTKYQjHRovYkL+E9FuEH9IoINQ5UKlYPSgYek
+i+cI6Mch5D1Py0pOOECPYifyaXPC60AB5ec5/WP7yhg3BD6UJf8S9ZHOcc3PbkP
mjGg3ougm4ZBHXDcF92SyRZmtvedzNRPiGsD0zRCWbjuZ7Z1gw8/eZY5QnJtiywx
T+vq0vKLYlUHXrz1NWLlpp1BaIiRIH9jFS56OT8VrnQBu58ScYFrvnmJxLjBW6Pc
xzEn/tcRH+UtXUbbKTEq34rLf4kayCGhWi3I4r4lGPmEH1RUfCjf4wgHDoxjSQF3
dXrbj8vDyjwyXrOI/PjktLgDeYXm64DOy4nBR+Wrdcr9Q4mitUwRnKwBTpH7xAe+
Wv0lyyQidgJeEtB8mRqJawh1ScpdWXjKuhjY8Z7gtpYLnkcIdrjM9gnju1qFeqRk
4EReQjgyFwOYXtbnOryLTky+WA2mFM8z04n9pfv3iSKjo+yFAtOKqfq5qr0GGGrR
QvIGR5RP9ACVHlkAsPFk3tPvzPy/w/7X4mGLeGzWmklML7xnLQPJ2SX5DApiNx0E
kZAwhXnBt+GEWc6hquJKPaSZxo1t10Hx0uBw1u7RorSFAiy+obUCN/uZ/8dTJVjk
PK82vSDyz/2v0RbmEisAMleeP+eHO01Bz/+3MntSJIDZ8M84+JCRsJ4+9y4zgiOs
eYOpIEU6xQTBlsgHQ1D7f6YL8N8xup9+yYzGs3l5BAlCw2vq2eGdc7j7yr2CeAmr
W4TN10llBdkWixlBSnvLOzOOKKgFwYWtDCmaqsei/eqE6ENvBZ+0IX5/cpp5TYza
TWR9R/JKeqW4UMMIC9JzIstQOQ3Ic/hwqusxx4fNg/x5afRQ6c+4iqqs8f1GecA+
Q2EKTjqeWnuEdzHTSXGiqOAa/9NkfBD+OnL0IsesMDZMNCFXVhV4ZwKcISSdIx26
WeeM7u2SOH2JCj4xnHcvO4bA5EVEqMy4O3V9S+1dptXUo5/fZnZG/txHWdhkT6ZC
HFM8qUmRHFkiiLq+r/8ZPdzUzy880ftlJYt2xtWu5oRAAGJ3Vv+WiaTFnFxA8ikp
mgym6XGFvhArO4OSW5h0mcRXlHeRgy5K+k5LVFMAzjFR14SEsSr/lWq2i+bkldO/
TMAkL4HpzsJsz7izf/Rsov7z+j5LC7OhmPCvy3Up2LeIR+GU/ZWWKmCA3XrvkU5a
yM2OxUv/+1Wwyrh01jVTTA==
`protect END_PROTECTED
