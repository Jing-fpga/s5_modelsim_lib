`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kaIA2yyEXcaap5O2T8T3rZM6pb5CzuYzWAd+HRrh0fJulCGvO+7So9EjVu3dC5uV
E4EWtUZvBNM4MDg9HPC/uoGY6hUFHvH0GMt70N6/fHK6P/74OFWUtKWw4WfO6AeS
HX4ucjVvdvzf6xSxhC8DJjzp9FQ12IXQlXuLmMeQfJFp4kGGU0usPGF3quLRzDvm
PNtSN6x1BOrlJdmt5mEXy5n06wTmobWJd4fIF2OA7fsRWnMTSCetm1oQaQabItmI
hnMwUAer1ceiGUXNLxo+m4Hu39FojH/2oMRhyEIt+XND4WRh7760Hgrh8A8uNcMv
QqPzkpYQjpQQ6Zgt5Rkc2bU0cfTvvMcgI3mbc7NIqxn4UdeuZm+856SPnw/NDBx9
z7aybPuFw71D0p2JS4uuYXWAn2fE7FDzpcnj6LDIkVivcoWipEikDb4xfuVi5gLA
6Iemw/3s46uRZE8VPr1fmjD+PbsE4aZCu2riPVqvKWOMN1RAPpUFjPDoktXXIdjs
957m38m2wpSI9Sf4vQEfth4Witks82ed/7np4opuHMyiFgaHm686mCAr2xk+GLpf
MWalA0tjZH7Q06gnkzfTDFO28WmjVe3e1sMQ/AUzhPSM2pznteabe0/mDv6mh1ux
5HBp/5f9xGEj9Jh8ebfF8tzIWEAGNkhl1xCoXGGs1vvWmJ+1qoCiSW283G7Supku
fYAjFCC11gPRwOBshqIWjSR4mW9w/vgfV8thdm8uYEKCRmudpjUBmgUij+uivoMJ
z7V6hvaeqHTikDhRQAJ04T9cNtgcBCIRsDA/Gx6Wo7JGRLotv2MIO8fOuCL+uQ5f
0w6x47K9AbWYJx+Ug779nqkfXin+iBk5/orTqNixuLZcaqJipbBajhkMQLPsDUBX
KIjPrGp+WYrkV3Cb9w5dWeO9ErujAVR61VsugJ0T+IvgUTzcQHMBWDPCEej5RKy8
`protect END_PROTECTED
