`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J4WYDfXuJaaNJP5J9fRqB5BKmPoqb3sFaor2pBLxoJijzzjdvMmmd+OGYCauCwZ2
XN7MUC2oLE4Rf2w0vuqn5+dg9dFZVz8bCfC1SY3hnbfh97/wLqbQycY4t5PTIdAv
xJZZLRvl8i6IelVBak+a6QwzWHJFdevQsLjNfzzACT567pN7Yj83p/gbFWZLeoOD
qzgub+K3qjmzGEBzzhutAiTO5Y9xCHJbnBflwsi70W0FJ8L1DhmadzP2Fum4yy9j
sjELEnjX6/zvQuQhwhEaAZqBUPvLfCmfUxuNbJSa6ngKvxbTawSGjycC2km2OdDg
Fer2taEVV+s/HGW4Tzo5SHxSzhhpH3vJh6SPVNqYGcBG3ZohlWFvWxZIW8TWFB1T
kOW8TD8Xix0iHg3vrAID1Moly5+3VX5NSpZKJrCE5an9L0B+OcHeRCUnmso/+zY6
idzXxC+g4A8zfc9DjTRcPbWK7QAA7frlF24HrOeIGVoH9tEuUx53dByhKvl+e3gY
3YQzahzHJ/JAqRNxhX/KvYBtQzpSMXRe+7EIf41+DvR92b1eyEolBviz7QO4e2+R
16yX4KIJMPR4vyjyyrjUbI5Sk+rObKv6eMN5/tPJiPj2uBPadBYaxHVM+H487vNU
KHWBtXxQflRbfKWc4Hd8WbUAmP5+xXyv+vqzcy8J4beE9tZCdekv5+Z3YdpmAad8
A3mR5YOb+m3AgdsIAJZ4Lx+FX5LeGntZIm88mUoiLMrS/bZbAsr2wKIIHINslHFu
y2qw7LZ92vwX/R5d/MR2gi7YHZ9fHbA5A36ykdQW3Pa7YtHsq6QqIKILbgH910Rk
9FZcPEc5C87EeKktxfnnaKThWzv9VXpHSQegGSQPuo5jDQhZMell65nYlOP/yorB
EVT4fDu1bWf/ChfG7SuROoeOa70To6ct82uuKxkdAaJjjLId18Fk1Ki27FB33BTU
eL7fVHzyetCfDjb0g8jYoTIZcQuR9slvkLEkW1eFFq6dNWaUmjzdT0675WT8keSm
Nb0+/zFu/OwexILyhxRMLGUqDWlTr7DMrpaZ0Sg1Za/qeE6NGKQSMshhMEhIEdhW
vkQRYZJvwk8weGn2c4lg/AEeiigKYSS9S427xfsrnHbMVlvJhGliT8uXaknQF9w3
fHYb7vhchFtAdHo7SwQFKddB1xtgQBeKJ1syyPiIkLJ5ZM1KSkCYpbLuJg1lGi2m
NsGVs2wzHooYX2JsWDkyGw8zwQgOKEaLY8FpSC9S+D0rhiCq83fxXZzHJz1m/hbo
8hi/sFvVEidld5fp0dduS8IFSUbI0ElTYoS/dycr55NKJgtWpEkgAo9DD+j0fDbC
u2kbuL60sJ+xjCPm86eGllxfCHMCXwlPJBLckY1WAZXtydwEt72ArfDGnOBTJo5S
5bduDXu/nMBpy74qsrffnTgZ0B/bZdPYIQT2t0/f+4c=
`protect END_PROTECTED
