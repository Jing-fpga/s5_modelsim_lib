`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
muAUeNdk2OnWIeAtz4+fQGDd5z+KLCHB/ycRjajFWrTrHsAMm7ZWw0Yvl0DizAZ2
MS/hepmfrur+iohvnvW2k3mKbqpqPycTRkpae+4hm1Axfllx/lH3TocxypvbDveU
lVBl1/8lHlxAoxEmydXHKR/zEGSItkx3Sjxdwg3plR1BF1dj/cVYe2w5RtpOTeQ/
htdIzub/LJLKchNchlnSoU8QJmXIOJQ77e9BG6cnNK2EOjeBFaGxGAgvf9yDjLxK
XpvhEidfHeoSDKk7P9+9HuvYrUJJzgrvmsF1vxTef18FZHHYecUc3sz6urTFzN2U
y7iJJwRgfKFzPW3p9ky1d3CT6NsphxDTovHrUXhdSW/5NcjzBSfcEvphvdaYR44q
I8tABAQ33ZrbgcPkjlrM6WkKlTnt58Ns/6GBHPFjUsbI9INUipOVR7lHzjybtmeP
L+55pg4vFarknTCAjmyk6yolwqG8GTBB+PcnuTYdJK4BPoBTmgbxFyEYagFUy9Bv
zBt6gxaYUIDIrR8+CULI3owTPd/KD8GkkOShomkJ5yNfrWsH0N3LEIRrnPAq69H9
7KxuVSmydwbj/7yCn9XgX2qotvX1bfGPp9LC2lrmDhiN1XM2Ol1MWtRkNWSkfct2
xzLMlHUKIPn9+83DYzKfgFLpfJYXvzLjHufun3rcZF3k5SFJD3dANhjjQd/9aLum
/svFYhSmjOZur5J+UL4hOuNqdUOKpLbYhVKCxAyVjuPcMVEKT/532Puw4HDVbVTq
4I+rWA1soTAO87fCa96TFLYwKoWPuNt6LrjrcwMFgLfEIJu2jvnfn3+iKV/gHcQ8
0SidOAXrkfID0i2f75e4VI09YgaX5lrfTrJ+ArsYVKFWxDGxJMsq+RaxVQ+hBSne
zNm13Qz8jCF6n0kshF8TlrlQ4M0NdadN+lUZepXV1sVyBVuNe1rkJFATfYscdINv
TfZoDQ4BBJq8w5TT3QG4rwK5an1ECzE3jKHAMUyu8hsdJ04HKeOgfnrHWRL/7i81
3b/ZfzdS3pJNrT8i7JJfDlBvmjwaJccLRe8DfwhVc3MayYrA+WwDzCxh88et81jL
kFq2lDgvCM1o0eVSXNFlv/tFmQH1nWdTffcoSBCskxz5EX9EXUFdJPnknTa1fdTk
GU0E+606IjwG8TjN4CAAh+ZJ87hywKOaZicsi8G/cXTuKEjDFwYc7wBOoTsUCTug
w6KWcIfs4Fq5olpBj8GB0YycMvhnm7sIk9uyFMj/soV+MM/D0hrkBG0N+I9e6pJU
BPREGpGApu5Re0nJItkdVvjrVB/z22U6PQCvTFfLLbZU7ETKMfuD+F76oju//nwW
fou7DsLjw8H7BV6Fghap4YMZcfkxR87Ifo8DW9BD2vUTKvfgN2PHEQRk5z00ISRq
PkIn/xxmuy4O4LBpMZYWlHA1Z6A9xstCyNWsaByeVWPIq4eHrS1AaQxtEF0LJDWB
wsHyTep6M/twlMgrZhBwah+vQ3mAQdRLm2ecuQs5p/3gemD872b2LkjJRMYChr/Z
RQt5pwqDqTrEY+Fhv7Zpe5Kd9qqPLBTSyH551PDGApjjKWKrjmigPI3LkoGSrIGF
KMoQEVVtI28EuC1Bmd6NgJMTGkHDXYKoY//gb7/Xycs/KTTRXO1i89cDUrR7uEQD
c17i2FLuYAhyeY+vb9WyylHIEsc+I6XycFmcmotPGBFcbgnInaG1Tz6Ql0H/uHIg
Q5S8ForFoZJLs+KGMO4woycrLPTnXutT5kbc7pbj/mbIRJnHLW1z6eb4l4TteOYk
HK70SiabDsjZHQxTGrHd6X060tRjizWGBiDXJsD38bbj+EpQztjW9AL9cZyc/BtZ
TGFeXudnVAoMLecI+sp1JOcsQcnxbAmeELpY1qLd62RTivyDpNBI7AOFUe2XalLK
Be826JmgN0RXYmgknRCI7/2zlbkNkdi4Qj+Zz90Ab8zwDjdnv9Izi0mHLyVBKlPx
lgm/RDjz1qpzBbIaCe+LyYzYECP7ayDUYD51aJC53wBsscQQPijPiCb3DlPN08Ga
F/WsoVnu4sMWI+WuStjiYDeLX102G9rua6CYxD1AjtUI5I+4l9ChkHTx58txtlZI
7uW/j5Z+YXu8fIjhlXyE11v8ArO/KLR38rR6o99q4ik8pd3Is38/2fsuz5D6bMWj
1+RO959HPBv4Bgo5sI2LFu2uFTWLmK4QeBNiXo8u+fo=
`protect END_PROTECTED
