`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
du1vVybXLQoxMy6qFNMm5tyz+/L/beC/5N1iXtLbUiIg8P+2BEigF0wnofWHAYNM
kHakL0azoqH5R/T9VSC/x7VSiCN5jWSP6f9wtmkGGTc83NPgj3ST6NVQBb3Jamwn
vTHXs95ETDlXtvEhQrKeGWHbjtiODhj2WC324TZVfkWDA4B12O0oL/G34Du9GJEP
zPCL/mWvHLd0fbNpxuAd1ZcXKjA5tItahmdMexnJrgXSR31PH0i07M4JYnvZX2e0
t0c/E8VBNlHIs5pya4OW6F1bkPIjGh6+ipdfo67NjIG8328N9shfp/9ShB4PbWnr
ltKotW/ZbnLmjV3JJmMlF8CCCycwfFrwGKereKScuIxUXq7F4+zQWIUJGiJNnQur
g6U70mQbkryRfcJ6NOWeP/FhCLItDXAd8j59BGZKqQYoUApN9X9wL8YUJA08yh3M
+S004/NBASvb2TvBMyu8FiZ6wypxPhSRze7BpT2YvfYAe7cU6S8itpDQvjQ2gSxS
DAN2ImJL+KFYxkNGZ95PS3G7sElMbFDxeWA4eD7whOrukCRDhlDZLI47BPFpcR6/
BwQMAgDRKYSVeY4c+1bqkGhTvJTES+ppmt/m7dF5kP9zMZedM33z7/f6KuRJ0+W+
eSuklOJ2UWkGydnT6AKZNxnqSA6K9b2Tyi7mXGsSjJ/2jNx8kAFnP55teAL+WZe8
mZ80Td8rX6hiYzxuy6mNfA/WVZQxZghxPuiIDjPQ0RTUeYYNuZAVNOxhJQvcxbMq
WlGO/tBHs2T5eqnMGUUnqw==
`protect END_PROTECTED
