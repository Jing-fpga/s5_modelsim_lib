`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/eeopLFHP1i/cADGlK1bPvHQz/RCYXMjHvldmV5YktfWZCaii8YWMjSHXTfobcVT
yypGjqUG9LjfM/kPAMLMpN4Ayb2oQRt9iaAY0johtJbTK25Rq/eC1V7ISb/aD4Jd
PyiIYC8ajo+GZqZJOkNZSy7ZgXcPw83eC6Yr3WqgqQbtAFGYKyUY+t2iEoLhkfMC
aUFAJ3Pw8/7O6vXwDcXJuRZcP6loCRyAV624E1NZEkEwZRcoYJfUw5LGLDc8n21+
RAyxnsQpHJ+GRiaEgiQMSlnHau23He2siMBy3QmHsbRDYEKUMtNMyP/lckLrh4Ns
qvlJ+Mi8xDhGwztCgHrHU8Ij9dLLqy3q04eGXVgxCMz2b42y6Pur5Bt03S/dJPv9
eaX4MmJcze0kFJMooeycCjMn9/iP9TfudXr2cUhzGFjPM3FAFIFHnUx+VsMZHk1v
R/uRVlvwQ50qPlOcCLY5SdeuveFunQQTL5dqm1NL4D4vrtXs6z3CnL7ICh33JVDR
Iz9RuCt5X4HZSy5BLFc/fogfpAOVv1mG/NwgIutjLE5hQmvQ0zFUZGsexFT5ghcQ
ReREKqN1y/VkckwCLWK5Bd91D6RJa/61eFciyJj9xJ9PNVz0BDegSViqRLfezD2y
Nn1JVsh9RMZDQiCGgHfXl7DvSGFKqUA+qEtXc7B1FafgSWXkgH56j0tLlIS6rsV7
hKKZyM9Lbb0FAID7UqMTMl2nY3J3snpvDhtwJeza5mHWE3hHgapHdHuDVezFeY2t
wEIYih/ZB1fgiD8fZeSZ9XsWI487JW2HITUfc0OnmV22LCucAN30ZeeUE5oE7taW
ug7BFSaXIIhELaEn4Lw5kynZ+IyppWHznofyi1jb3S7iVxAIVjS/UDe7UoMk9AZq
5HnmwEQXSXo0nAILACMtsC1lj+c3+6p+spwnNXT/R67dzjx/kqG89JOZI32/2p4S
ZJpLqouzq33yJepBe3mQfiEi6Rfah2KucuScBzaofaECrQ3ife5xvY++4J+D81o/
pIaEGrYdb7E7aiwS11pArJ74HYaWry2rjgcl2yRE8nsVm7qhr3A33d6rxLVn9lky
Irz2Y7WYHGXTNgOFT2zpL6frdZAw88huGXJjxvY0D8W4fCVsZKfKVP5TCBmSHSQ0
ouEJvLJENKEcbUYL4kYPk8gV1mhcO4ubpbnqVrfyI7TWOsunaBFIf9jYW9miT+wi
lyPLRQ83JXGgQ2GmrHq8xStWTQODhlNqPU6E4BbjEktu5+NQk6kv1knaF/bOyiad
XF4nHtOPReM3vdy6o1n8CrbFllPP5haa2l4EAFL6TvwzdfkZg9GNjZywrGzEzsF9
Oo83hS144sVTnpe7SLtFFJrOZLAeFPuNNAjDQzAhJYTQohgudWMOAcs2wERjGvmp
oQE1b4y2W5ne7V0LZT1G2/1QWp0rBxQ8WHTMEBw3xXu+vIRbbIzQFDEM3zkT0LAF
5eyUTeRhsW6zIpkyQmlAa80LIObPzB40snogEhkRNUh+hoklUJ3uybwAg+Bmivpz
2UX98kre3RxGs4e+zSsB5pQbAVhoQ2OO46wb18usYz+8om++tMG6GkgUpJIxfSsl
NbisfDrjwXK1PHMD8PwghXogiyeqoXfUlwAG6sXk4TPmvw+JaTvn0H6KCr2RLsHR
163eikEbQ3Y4V7k3seXhIxxc0rYFZD9EefBku8PxA5FCyydirbd+tz65cRmYrrYr
kIN3x1m1w3ULmBv3CRyh2CXDJ4JXd7wtSIV1DePNJrS4ENXgj9tyV73ioHJdmTWP
nbqRerdztnSUfzbN0JO2YW4JGyB+/dMTg1cNlPn0giJGASagP6q5nBkopauu1Vc7
a5fNH5z/7UHLV4P8BlxIP6YtycYzTVVMEHKUHoUDeNDjZB/NfvVBsGrnG4I7veB5
PJGXTOFiruNtYYLA5VpidhKPl1sPE5h0aRURg11E0Lpi+aEb43dzpgZTeFl9MsML
0aB9xCyhZ8fJ58EU2Y2WUVCJieGjY0c70zcJE63jr0fD6/ySX/iNgbkBT7AirVo1
SqEpNLZVw+kd/6AdRuUgriNg5k58MJSZX1u+ZuzuIZPcRcIGG1TwjxfY7n3GS1rY
j7F6bVL4dUxmsjlCZokTSqP7YSC+Wlca5G6P9RLzeFy3BKLvxdb5fVVDZG95ScOS
5E18SYk5oJO+FSY5Ka6d8BCqAB7ZDcGjPwuwwoXBDerEDUDSmXJivd1gmofQNqUQ
Vp+d27lKIbaIKIPnHDixNpXfkoON8j+yXvZWDR7mjX/bqY0tC/SwP4zdnlnABOWJ
prhLLlkHZoScV2JSuOv+Y9rhEbwMsZWpdN2QTiERJ53TIfsmwaiqrVxMJsTXAgAb
A1RllC7U8AdqGjm1+hueWhcGK+oQAaUg4bla9vSHqToN5EQ+I6leEI+nRFJ5T+WB
SqADQ7MRhu66Z4gsPfKNjYXs95BpA3zcJIl91JByZUJd2TLvXTUhbnew9HJUvGu8
G01ov8relYI43s713U3AmnaQlol2iKJHSsmVK8qQk5qa8G1ok8Yi+KENlkzavU/o
6gdG9DDUBEnhOXa3E6hegWRATOuTesK+ZnBtkiSPxltdlq6M31x9Ye5eUcC1OMft
9JywRsFoi0L3do6y56JIKYtoIwO7PVBQaa7d42jJ1Q4vS4QcHgpVK5vOh2xE90ij
gOZtE2/ioRVtTMKrfM07LLeTx1FxIgznsOIz0JhmHFfzZ0Zdc0MuhUOsXhA7xmha
NsjjRX7ryC6j8SLeT2XMDzXE5U2KZs7rjolgFMdqNBIHhvGLg1ycbPr6N6UERCGw
AVF/AjIcNrppRnQd3n/3zq2vw3fMiyTQz8czgpXG0YaB3gxXw5SvULTbfmvVBP6/
hFMsy1u7o8t6zJCdT73eEKRyag8J0grCUSwCmyp0XeoiWWBplccRWrx/BJlFKMMD
8R7Jjf7dFhvt5PUja3S0eBs8mLcvFsqMQtGgtGQUCkjfF4fuWYcUwtuQLCqof7D2
dw+FVMGgdvu4MMtE7qMoEL/PYUPxbXEWIrYG+S2nR5j2QjhZ87SynK6JJN3939ZB
gHStcMTGUl/m85Gg4iFR3SMIoGCgD6AifOwFQzPLy3WUu/gmiKkwe0FHGemWk8rb
FYbazXHYDZxe8hph+BVWNOXXzUAKbwqMR2Wq4tZLv2Osy06rHxn0mV8uz95svkHC
5aaIOrd2Vnk8thJpcVYhCM0akphtwopy4EPz9D+ODPkIdC0OVQmBeMdo4C20hvK0
+vo6qSQlt77FNb/Vqji97Pe9YIM7oBK8msjF0n/lNyGkQg3GXoRI9tVBTWkg3RgW
/YwqvIc6akwAVeouLGGvRG+PhDRvBOVSJfmrpMO/W1E1KwZePxnsc4/0sDwFcuCZ
AMkONumX3jPFiNZwDIYaJszZE1LRn+waAYCYaX23vufBB2MypgojGwJT1a9fezus
00AGldwuTtQhI7WovSFD6rFYC45CokUFVMjYvM9tGYMRa1MExlpsfkqrIHB81LAE
5Kb7RHCm/E3CwVd2xsGFhj+yc6rT3L5myAL14aubDbFPXVlz16zgrnzhyOpYpB9+
uL8NL6+I7/saF6GvMx5qYXkZ9yamLQ5wigiFUKJ5iy2hWP+J8nbK0+3hieZCmqxJ
vVv7w7M8dmqOtN2eZCNjs4fb3lhKqMxMilTfwBXfLe9Cnw42a6K7NNGMJDLqmR8L
ZK0wu21LTHJqXGlHkzQ7gUH2zgRDgEffcdIIs11hfzxmDUA8+7pXMCBkziAswnO5
TdfGZ6JF8GaEm75kswKdli1XkSI9cZySuvXOM7qOX7eK3YI93RD8I4bf1BfzU6+e
9zXzUlj2Cr9jw5XVVQYvp33sk9k9V5PPl0Gz3ZqEyF0hVOy3CWW7X1At659/YEsj
YY5Oj0REZvJfPkGcgCZ2325PVN+At9PZXWxO/MB4+IU1Jhd8qR/ChGCgxCDsI8Qz
eczG5b2eMoJ4S0HvXMTHOjIT1JS10sE9vjIRwCB2I5bmxDoqZG0utQiDq+k1xhF2
Q9qQo8ZGaL+AhnaBm46ThHMQZXetrTN6Kjf2Q0Iqu59Gj7FpJMxNch1c9xg6hjOv
xuhzXdUhPd4MHvEhJajumogshjV3A13qCXcYhiJozCROz/Zr/9WkMUejVFYIfhA3
o404r9q37OkS88Dkor+TO5To2c+fVR46ZD8O4zccqC0oNEqEPo8ZMTEjagRBGvG+
YN81h7WV8uY/2EYeWN/tilkVqpORBDE9ICMn6J/4bICFF8fKJa+LI5ls4QUpK5CE
`protect END_PROTECTED
