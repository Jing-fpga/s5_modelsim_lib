`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1zhhtT9ghTdXSyhtXnl6laSt9WstljGxWdFZnDkL1XitM9L8s9yUN2dEZpazpyXQ
YSaF0NqhygkIOZ1CVCH5Vr3T6VhoEGvsOFEC84fWr9eNsJeysjq7XdxU8h28GUKB
SNuh+0nQSlX8fkyZPBVcw8EE+SMySDI5fsbVkYGPMogtqa7St9GVlioHIXKuM8j8
z56Ggf5BQrNreV2yiQxJYwJOrdjOPVaepAuNZbKFcWbZUpQkUHvpZ/CvUGPlU5bl
MiY3Q53snXqN93Du2cAPvPPT0skrwJgL+mL2Oy9WD4R4qgS1hz5vSpvCQ8/cMJJh
MI+i9Y/MEPL3SpgZNJQ+LJV/oS86lz5nzGc3gxr9RqE+vAzexl8as1DjlQGdr7jL
Na+e3bLC4Ff7OmJQMfPMlJ8CMlhDf05iaIVy4GErM3oYOxxQF1mFNwB8mirC5tzm
hhc+SIP6kDllpAPcYjqTtaKPMCu7ktcHjEO8DDk8oOXKp2PgH2QFME4wK+6Wypu0
H/exAJPsDlnnYk/9pnGoxyHkacjOBjG7kDhtfu1OvnjT/OMDB7ExAO1qaGXBmkeY
SbO8mw1d9WNQdii0dJ7HVM3ZrV6RGLw8ehQ/bYJEx1CKT1hScb4MfD7CCKZe8VOj
lxNklIGKgxMtb5VLoaPmv+wLpMFtCr35Y+1eqaDYW7ktQhpQ3v7Th/Raibdc4HPZ
CUbtlNmyo4y1xBe1IoUKVFwI6Am/M07oGr4TIIvj2z0mKUEt0b6KBeA74NsW9pQt
inRTHsbD7JHCQVdagVSIq0W/dYLWGcJSc8n1K7aR9uFH2eHWVoZYs3NC4KTO8TEU
Bc9xHPWx2gOJ+hA/vKDzePbAobV+6uL1iUrFpxQhWU0DLR6+bXpFqaSE6tfGWp7A
Xl2S4N7hY5aMKTl6qYn3pS0VHyVCDVcYNIkBErdjYGbeC/vu5PZ9GSx2rHguhvhr
qhdU4hZuWxQSBOxgRQ08tLLlDSEHS5mP8ya1RoUwUeDe6V5nfj16E6c/98y7RerN
Dysh///yMSzJz0yOGyGt6YqC9RmgeFwN0S0xIoBkHpfiv+gMxyMq8GwNzGJL5Fm/
kExFtY+OUNCAkw/n17PnoksK2qFLPhFXVfjfP3Mx3mRFAgSC9KGE3hyyQvunezNF
KMNmRpcj4dCM/JXGCSpOrTp0gbZ5hwQY6MXpk4lodOMFcq+ORagDK62CwUwbcUqr
Jed4IOhE2d3H5hwttB9g2+gPrsaK+aRvri7UsroCZfIztq/zPZ1gTd3b1G3lBel/
V93DGrGy4U8IeKRG/iOwLpgnk31wcA3wl5/yz1WrJZ6KVh0gIDkNy8cqZgFkwe8i
4Q+EXK9WJ+0h7G7xxxkIjhXmM+zuBwMDgaEr8vfdWkizzkrAX7EN+OE2XwtpgBQl
EU4ufjzAiZlrnsZCf3vpZssmiUYVFN+STbOaSyUgteaijJ3t27D/xgOCm5LoXaiJ
HK1O+ynPpyK1/a7tku9yhpj5d7eIPOCM5SB9Z5pXWjfNNJgEECNXqngJ7fE74Kca
4s6MgARpOyNGbiXHzpWH5t2le8srw+N9hJRrENslKH7G9r42KRD9xcduKdxoATNu
Nd8WAgmbRU+310dyHgER9Biw451vcAv5DHT04cjuvJAeur88BUK7CXOZBF7ihscE
CWe21bhmmHbgFb4O8azzNhAdQdUt772Di84EnjJZjVLr2Q1TI5MIjEzCfrNzoImF
`protect END_PROTECTED
