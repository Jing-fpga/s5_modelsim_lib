`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mzVhZoEr6nCMyyUMyl9I8zksWU68KcR3fBEyHjfbgNtqIjyhb3Zk6zHfl/fcxTBo
I4RUwjJCgIqoZ3OeGMnRMM6mpPvjgzmqI98KZb5W+RCDx8mV9oduU43ehIxHplaK
byKK5ONPJmMepGeDYtUg0FYh6vRpWiV/GqTECDOPjfSd8n0xaPeINqqbwUtA0e26
ic+ois49mPPVd5K8qc5fJKowWEScU+cwT9ee88QFtC2bFS2zPF4Gu9U+2vtdrTxo
Cm1VxLwtYpe6mpzzFp0mlpjWqUGMxYsOfiqZTE6iMkXCGnZWWHaaTDiYaqoVGxFr
CZPpYwwZypO3JDshlaI/GOCKk9YfYsM0wC85RZDK9wVpHeEIkE8kO4rBVVGzdS0s
npTFDL/wyOpkgdrbZrKp4DoMY0yqBlVLQvwNQmfvrLADaWiuOXLEE9lX9yhpsjf0
daMtGbgPw4oTXvbxO5DynokYHQ4GHtyEPILyAktDJTAIM+wjIe3+xuOI1uWCyyfi
U4aed0EOKw/1zFidmCbYBWaUCq3n5voqS1CmHIUWUcM=
`protect END_PROTECTED
