`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wdw5++ox9AYCc1U/OEvgeFybZgQzWnEDl1rIAx8iIG+RcH7WY3XVd7bEa5ZIxtc2
xRr+oTiH0d2efYgaI3O0J9BcNlAQ9VR0WqdxamssKlUz6IBChVia//VHovdy2bAb
kKrw36Rf24fO2dgpg+2nfElnz1TGLPlQRrKAvcj+OEDUoXkAO3fCl7VEe43KpWd4
lGj13Sin62FULlavtiH+7uehptWhzQH2CQ6MG25l3JfEn+dkgYY9OtVpR6nOLrt/
EoJtspC+S807bGNLR7JPcf5zsH2XmpzEeVKPmoyspv9MRsRBYnY6so+ZBGdjvsIW
9Qo/AvUOHwzPgZJWLOXomOiJazulfQD4DMgm4DT84AimsX5pDB9pk2lLZJ7U7EVg
sq3VxMFbWiQEX2N6xIx6TDmOvRb6k9+uI68ckVV66V6H4gi8QRH4wMXqZ1PTrxuq
KCOT5xq017wy6vuM2xourMpsJ7XnAqA9B6d87ai5ezSzXFn7U+SvECFR1Y+AxUhu
4+tVdKUjiQ8Go9iLj2t9Gi3pkFZMC6lTlFBYuwADWZTIxcsP0tE5VK3BQfKCb583
6c5RnNq7+eTFt4l9NZsNU2MnSnouN4ycCJzpcFzqId1oPFO0XOwC5iW5Rmy41bVd
p8gi14wnzf/bw1YxjXMQtbul3SsuZQ6oU4k9vfT+po0yzPT/aYozwe9soa+WvqIZ
bWaqZ7MNUafmarn9klZ3OSzvFO1z/UfWPM4ewt3UEXF+1AH1sH5D5C7uBFggS5Fm
w46ZbRlBHYjJgT3ffEy3vHvMi8BP1YbVNqEopxS8kbSb9fukdqi5FXdBClhtI39h
b2ecCdEWfyeRodi6bimJTuSmQzGypkd1vMmNYCZw8mgAKr7Zio1LmFwh5y1PJcN5
JlxBM+zV5VUjOEwLzH4MoaaGRNShDOROk8Tst1IPA+nB4WH97Dv/TWyhJ+ZONuTE
0iYkOLVsqcolXimOEaHR0ACmsj/IyZngmANfNjBRdsnapohwjQPGetBB6QWdK80E
pof9FwHwsld/wLd18paGTGWw/7QkFIvNOZBuqqq3cM84feFtBWgBU7uHfVEfOjDB
QukDD88hKic+l9mP6SSZTACbrB+v9kENf2MxUjT6d9yDyvQoKJVgIFlMpAf71Wp3
9wv+95ZKxJ6+ifIxdvBU75pAMOCCAt5Cm9rPtWgXt74T39nFYSBiilddHGycxDTS
Du2+tCGKe/9t4e3l/jIf49NN2yAUuNOs5X+vNBxAJGwfUvuxfHR1WrlRoQc8Ev0R
9AfLoU1Di+fZ6vQY094IRRk2UZkZMYH2qTEQtUDcb2NstipoPFF2MbpG+CyGx/Oy
gaiAnd/5cKx6ReRtCLpvi0nvsxNnjVrKX2b1P+G6w8TIxDpJKPf3K3wTIZqckG9T
UJNQpEy7WfK9FpJAPW0qKyupRM/z25VO6n+t8S/y9MxOE/Pg9Ncm0oAKj6T/16yZ
05qgDS1IlGJSic9WB1kqmedVaP1E3LhvusySVTGVlhIiEVrSZ2mZsuBans7sNH3d
rLdTuE/DHB79AFTRPpPKNKa/gbsYag3Krg+fs82BMYx9o/tYSh1nZfnyetw9Nl6e
ZKZ41sQbNqBGDvbDGyvHog==
`protect END_PROTECTED
