`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lzMh8RXjYVgOVSTJjYFmfxnnVewI20V7f/78GmmrvTIj5aVi/7DdyHih0lAAzHvG
QS/1YImvh8XydWx0/8WU/Sc8UX7ZPuZoBRe1KLI0PyQgzi/56k/sav7BZ0GTmw4B
1kBD7zzAnlLunPMw1m+m1C+tOl2jGtCOMbL5Asw5sO+ca/yHrP7UFFWCXeH9V3Su
7yYvqk2nQc49e8mzI2MXzptWglXkB1QnXFSesl1KRfuVu4ubhkqUL31xhD7+N91z
8Zaghmltgz5sYdu/WqDuTDPH3GXF3zYordUdySFSmz4SOx7LYTDwrb0WF943Y3nx
46Lt6U/cSYAXV5z0aE4Vf+LQJnduVhiTnrCr3Bk44F+f5IEv88ofJdd6hdiJWUai
PcR4l+CURDjJsdsKF+8MkyOEBJuiiJxGYOvexbXF6W0uXNGxu9ydVcNz9eXe7+ms
pxyVp1N8I+ZWctXRE+7t1qQrM/8cpRjxhxOCoMUX7Nhdz3bf5kyE5JyLRRn7gOnM
ouSGQ15+MaoY3c7mbX9LbbmAT9XkdMLnEhnlb0+GN2z9DGTjsdRwsq4H55l2vobR
C4Yzj0a4iCqRkwDorkmMTOyIDbAEVJmzVy44g00mqEGqJQZ2N89zZX7HeCNJwY85
4XJcWnLiQdwXNqQSLu4S+c8YfVmF1er+uC94QXCq0zSpOzxktDYMgzAFJoAFkNFn
CpeZgxKMh+k68IfsdZu83Sk1jvuTcTglpcYTAb+3cpwdjk9PUoLKAdKNC7rgxcDI
vGno55I2Xuv6qC7xC02yCdrvyoBx269chYSiKBwhwAhceO6j1ILLabrqmZv5iAhv
mPkm0B1fF0InrEglyZVZ1obKtEjWxD4EhUaXaUdzN8Q4icaOppqRtfRsd4YTuoGd
73AmUNp4H8aPKDLvrJanuOZMk2dJJZr7dUyeNB6d2OctqeUqN196w4Kv4/Z+Rf8w
12Y+r12OnyoDJxLissQ62mEuAFpNuibA2lrkZ7t/80V6h0Mh6tAGFSzBclG88QOf
WQVX2/efvSxuUMtHxisnrbp5OU/sHnJJLdAh7ugePVHydGZtaJPT+AnQPtI31YHy
paLbHUmMhytYr9c/sKMWhiFwDaE5FCMVSB7AmPMd27F88BMWYM1pR16ZEJA6EuUF
I7GNzrWCiqkZN/mTpOu+q8apqWlJ61fQSId9fOy0aIvtaqH0IXYZyYwn8dN01JVM
31JpHx+e55+H8fku7FqEl5ZxnQFN5jKJ6mJa71RoK1ZFKC/h/aPkI7MGZp3s0msc
/DKvdonVwuC+1vw/yxpqJnb4k9wyMX6wKUzWmsw8OZIWsAbMIrVCM+UbuBiMMgDF
JA9Sm6enALqyaRA/zu3KnJiKrFFEdycaiHlnX/F8NV7pwu3CG0aBCwSMO6ijknaM
YMzdbAmGY8rDM3eTa1jCvNsuTfzV3U4AycmZvzUg3S5C9RbE9AFnPUSiRcjp9EVz
xS4LIbrboHYmYjZpAMxAfduWIvKTxR1Y/pB9eDKMnCnKldVi6GemMghkyZSLHtVx
6+Iv+K+PBTOHsyBF8QdY9ZQAEGgIZjALTkJkqVIm7VHCk9Ge1tfq2v4J3wCy6q18
aQ1bd7BKn5UufZu2RWwB4Kbv80Obi3iVihH4IGgreP247pV3fV4gUJT0roNNOtoy
ClPwLqb6s81SBLdj4+sjI88axnMhIaHnyWR5Frn24IZN37nKmR/7I3c5+JawscF2
pJ7Rdne1RuAH26Eq5270O00tBIr5rvRJrolDVuooW4MVZoGv1hKLbs14x34VqbuM
pKhSMjijeeGqhdoPT6wTPH+FUIERmSiuDKXGmJ6c6TD8z7il2N6t/W2rormoxLfW
XG9N3+uobAHtvu7l+KAvlEhkYDW9ub2PBuYfOK79iIwYPJyDwgdpp5Msir1MKQwE
aadp/VufIaj0Y06LetQUCcj492omS09Zad/QQXtUYT3yMXR56rfD+Q7YaMOhlfLg
QcpJLX6raAI0fXXmVoq5mIlF//j7LUKVdL9jIbru6KG4gOLBwyiuGRPiy2G0Ru7S
n+3Pi9BPs0cyLDSdrlpYKG1Qhmieil7CcZZkfq0Uj2y72yPBF/JUcXpfYraTd05V
JmrmqX0ak+Em/57sMHCw+/MLEfo4JLDlv4GIGb1SermfEsnt6Syc04HaGRkL35ZN
TBu5j2ofH+V9swAXQwvS9SqnsEme8RaSPiddw+P+2l/rsqsVzd5gw86GS/8jSQOB
u08/idqwdJ0LssTT5P9O/xDNfQZHA11HBClGw7fV+O/sJ3kyqNbY/yh+HNJQRJCh
6xceikAmq8Lk5TG6XMn3wIK7yvxHaixqSVo0DqIjEC0k20nYujAe/CjngcJ3BGaz
tTguyGOpvwIPqi7fd9o7bQvIrwfHHaGVxVEdknwX6Z1LQ/rCvg1RqwImavN7hBCl
jjhxaHsFkpzpNv3ndrAtl+jUFsIU6aK3w7FPhHJwo6OEMYh80npiuadNqy9mpOsf
9dio+bZ+h6uUypxwj+vQx/WxstDISxlOuE+UWTs1IDpjMAFE8hhZZ+j169PDE8Di
GTCwMl7bDOwOtBl31c1mu6XRuZFmhX5s7Q1DwImR174QrjtmFDHX9PsHekT9jRaR
2cnWkmdAxD/tmFw3gG3a3QEsp0gPPTke9YK1DRxplHfLug+uP9J39xEpnYPGXgJB
m+UObJ9MlYqKmGSi3I4FoasYUb3zZzVqVNWcHtQBe9KjQBueUvZCC12R6q691IHq
gr9RrPx1AW3igsHWgdXTEjN5dpVg654Aj/CYm302/8H+oHkftxUBW/89k6zH9PGg
kLBRz8p/RIuV3ABpM85bnT4YD8ZJrthb+Us3PM7+HlSzFyG9TlX9bwGXDHCvbVzG
6OadDgCROZ5NhYrzvool3S8HMNJsLSlC7z57ALhyTiw9lRpJAnhIk5mTPByrD8DU
/q7hN/0Ut9hY5giqrh+3pWdSD+SeRVE9R+Rmuv+Fc8snv1P4jwDhTmRiEVT22bqb
9L5UJSFv86P5BaKzpI/lIg==
`protect END_PROTECTED
