`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BAN/dya2f6ixXt7Lh+FBNj4VJBhMKnorOLrwsMsn/2MkqCLWfwp2a5jMm57eW2lm
Dzrh6q2KJrGV/gznWoRDm2jKQXo1c+OHe4k2YRTEI59GWFKQpPdNs0dSu+5m5oJy
wJ2lmNo7uaAj1E1xaQ5NZst+PfFQ2zn/YJbK6KGDmM1YC/euZaeTduyfA6cG5J6x
klNsgSjCfloI1Lf3XNGjDGHEZH8YGANkYT+qm+fJceeO+k7av+zcEHDlkpnXTkXc
nXdeivFDjk3RZ8N8NXBab4n2KBhdzw8m3s3C19iBoMxYozvmo1w0xu557q3+0vgW
xg6PkfsRxe/fUQn4Sv6JaWklHMaXZS3sJl7QHvZar4rq1G1zztpVTqbUNIjilHFF
/Tl20akOcgsISHlZaTkpFzjPSpXF5GS0FiaE2mWnZjzJrjIBZ8gjD1CltEKoUs9F
J0Bu4HpSi76KHvdrI0NcTalSV95A3CpLRcLCMzbu2iNKw4xEcmmAyV0+zFyO5W8H
Zu9Ras6mAP6HtqIJkzCfHiY/ny14jgXmhPux5AyEAOdCVXO31mbNnY8loqaBJsii
NGwdumpypDVVI20Dm4ZZKIyYkpgBv4+OfKHCzdS6VkmmZMXT2WX9+fpZuSRmrQPP
ttvI/qJ6Oku3I++pBFidwYMAB1X3WLm4ePlIia5H2UvtHSaD8nZFfWUtLXZaUXJB
OAr0u1eCbEvN5O7qzb2v8wjlyxGy5kByLMJlIStdu0KSdwEeolkdbqgDqmstYF5D
slRe3X46DMZlAFxreS8rT2ZaG5WF4jwUHMBfK7c63kAjXTyxVehZbV5l4WRGpkG6
f3I9b08Icgj79jiwBwoXOrMYKwJuWUk/71NjQNkjW1rahOenBa+xvJ9RUrYqtifD
HUByUIwix2OMZEC/I9hSWUpI4eD5wRw+lJxks7g8RAB/N+KT2eNZfenINcVFYZ4g
1DTB23deFxQHFCELqJCi0IYnCUWH+Lwd6srDEXc7C+8109ZLKsGP30dTkW/4Wxsw
0U7/qXuzsbXJ5rTjzGT9MAd588RJP8PABUiXZ7KCacup9hJqDPajs11lxUdduMcW
fVoz/bat3BHDzHCQI+eC1YEqsZeUHmrGG8/+ZkGluDOvpdNvM3vhTzGDq0bY9KQ1
9rslOI9qf0zfQOex7S7mq/teuNlJZC3ZrgytAsHWVnIPE4y532MpQiEojaFb9KXH
is1dyVWiOplcfBDIu2Y2GC40vuXTLHH4iahI/vH1eWy7DzdMuFfijKHJGd4PLLQE
fzTFFk8DHfYkeHGZFmtAXna+/ROx6zfzbAhrLgpWTZEQN0LL67j1Vv6SipDPT7m3
FLKY0YLMIak5FA3r1IR6lxUcM7HtxK4mw79QpcvaOR0636u0sna8x1sf8owMlm1y
YyxUiGJw/ih5J75BKU612SRLbV1PHi8M9jkJATXeyNfPe5cMDCEEo6BwimcQACRz
fO4sFDev7ywlbaDlQVunxWYHMOlD6ij1ipkrIfgrY89tfmIjPm3QbUFCR6igbWvB
bikPoc+OuH+D0s/0fBB8SZGC9+eqV9zHJ0UeebBTA5t6iZtgTSJE29nTiAneKKWc
T93yC9JVa+L0q+L32aejnNKm3JVbrELRY56ztmqxXu7fW6F72ijxYelDfIHBcxBt
jQH3BSPxpYqH+8YZOSgt08k/vfG8zKTmSmEWoEUIIBT/620G+SZ945u60Yv/uX5n
fnhPWPYXv//n1HLtIY6Ol9UiN5jKHTLnuVxeGJS9ikf0rasToK3udiJtYs9mkyj8
BIeOfTghbQ3vSaI/2KucToKAHlbJuVCwjvbUG8gb6QADdKYTjFvbHt2BnG0MEGqP
wZCo2HHXbrJBZZ7TV1ldP0sBbOh2Jjcmoq6OZsdNuV1CvC3By6AjL4SRKM4uAQFR
isdQagc9kStTfGWGlHH6M+Lb9f8SDAA/BHbBjWTgBDEK8yJ3AdkciNh+Q+U+8v4K
2H3xaC6/qd1FCNkOIhlOupNIsgg1/JkUwVv5eUvcIW+J8/QxYrqL0hpgJg9DVzY2
VeK2nIvO592Fq7tbxRMCBRvH9rjjeNopewjVgTaNkqGbe6TCmoeHrdzvr/NGiz/G
ElFRtRJVPwBc2ULBxvlrjnKF8+lEH+LOyTzEmtXePMH3ZrYzJXpjKF0V+NdqqleP
+cpmQQkSgmgXXw0lK57cyKnxi6ux+PKYhidYlzHlRQK/WvRFZfLBU5YUOC7H7XYr
pwmcr1yUHa5xjGoRkQUCGL2I/tJZQMyPS4PyOFG5obnLvZl3ZcL9QmFw86Dgwc5O
DPyWtVsgfZXLINc2GvkqFxgT/4dK+fSfYorj0AYPHcKyUg7bfUFRnFkXDg6Dr8wV
vbudYOXc8Sm1oDRD6DBobTyTpuUh1eNCR1Lx4Vqn33SUV0MU0Bq+XOstgolt1xzz
W5pZ3hBoRR6nT4B3JKb6jubeYARvnZp2i9JD7ZziAFQfgdLWDClgfTd8SnOaoPK4
UAE4SrpR6Q1AWE4aAnLX5xr9SZvthjxcQDG5zKjl8NK5OcKj20K5ZFN+BzRYT+Tn
oeVXx/E2hYQzc47B4v/pYQIXEqPthEOOTO4afPUj+kAbqdyxqKpzGETJKD18BgqL
OvohP4AZ3fIm9jPZ26S7lwyRRHrmGVa8uNMEWC+pwbo+d/W33+0o4SfuN3ye8WSX
/I6SRkPKMrntO2XDhJCiyjgle9+UOMz5tpf9sl8t0lQpOrzTeTi7wv22inLf8V6P
tZLpARdhIssS64U2gO+g93/09DerH7mCHJ/4OHk8pSKDnUOMybo8GJFv+eqq43vc
bRF6WMbdsQ6OfpEA+PHBqbqvDpKCWCi4UTRa1FG3LGQVFDBx0JgjT4R07Fl0fmbN
zI/Sbdt9tv/c9I93+HFrTH+dBc4acblxW92a7M7iHL+plIGM8qxUe0y1MZcjupwX
G/fvYJwF8NaltLiY2GxWtfMBxTVq3MbwqoYRvPrpIvzY21msY+yq7y9lHPFEjVA7
Q1VUKgytP85Z3Zk1rUa2OUwumqxwLHog7RjaSQF8RSdtbqp9Ky61zFviTpZMSL1q
xLLe39+GhdLqofhKuMQ1DIWaeG1bgZgdPLpjtEMQRfI0TH2rzq+qau7oeuq57gYV
4ZemZLqKT+cLfM92M7ualR4envJ+HBHVu4vqek4nMu9CcNy/ZakB9+Gkir6AJwSl
8g16yP8dA4JUtXSMqOsJkjYuGAGyyLwqxaEljNJSO4vQTS2pGV31+oiZUpCjIChG
6+z4vd4Ivk/XBV0bqpUk0k2UUO/0vGhWLMEGRs5EEoyPMw4VySNCiTmFjScT45qo
bzp08f6nUfzgxbd5iyp30AKSzQXgztfYC5O9pWItaBgcK+XsHpMdqdUYrHaQhLev
WsYWiEQbatX1lU1W/M+qWxDWbWiSvvDJyrigS6ie8GXfew/KN2Zb8sc+zpDBfLvC
aN1VkxAkSWGOqOXL/SvCW/21I7GGRIp61838Jjml759ISuh1YHO809Nm5EjS+4Kv
GVw7qEtY2Q9orE2mwzrrhOCeZGPGTLmTmqNpjMqzXha6b9tUsZhFt3L5+LVb/lDl
i1ikoymzGopDH7IS7WIDf6yr6x5RZhNLm6L1PKCvLHXPDSH+0FjnRcRj/g6R49TY
XLE0O+NtI4AIe91U1MIW7WbB5/x4Az4stydgWSh8PBllElde7YpyfMOz5CWh7zO6
EZmRmasrKKrGVYV73bVazgiQemUX0qfdCtrDxYLmETySLYCprok3EL22Duxmh8wI
Ivg9MNRfJsbaEWA/Y1pX8P5PfzounTTbeeUtjDuCPxk8u/pThvnzfkLjNx5z/u1K
e1uiHbygkZiH3SS39wniJ3zbrtCEU4fMWIUlx4DlRVyACasCv6nGpsI9gQJRFjg1
j9e3julO28sl89KCqvLFz01UcXY0pq42y3Y4KvY3aQxpCoZ34bvwhVFtGUNRX/j+
uj+NuMKrNCWdXN9zZy65qH2Hc/xfCfE5HNkz4Hq0FnKoRyldZl3+OdwcTbhqS45E
w1AdCBRS58utrntEwxikjpyU4GUsdOi/Naf9AerVV1UM2Ws95qoa6KBExpleCsKU
mxdcnEMf9/UvCwwKrplf0p4vswUrttgs51LnXNDMFbHAq+Vw6wdFDp0TzKc395FZ
hKyvC0kp3LFBXH2LyPoJmP16DhdHT2IjDjoLrw2gYwsC7V12acfhuU8E0UHMdL5d
m3DT/MGojIidLaJWvD2r52EF5ErEUmqUthbh27Fk69Ay4h0yIkWnFh5JoZKg2KAC
oEqC4+mYNtbP+olEnCRyAIXtkjaqUNGW4iNalMEW2j1f1HWnS3lhoXKhC3sHClpZ
r/euFDOFvqwJBdCMUFDVwKsx0XBJ1b9DOsDcG0Wxw3PYBLTouzK4Ril8DbiVqc1n
hd/z3DG98Iv/EjlWY7D6/O5+YInDN4J7728GNGtpv00tv4WYfVFh3KMfgUOY8zV/
iPgjxUBshBeKXL13qJSRahLZAdc8l0ixH7fuvb4M2oTDL2vBDpFL3+76z5G9PRKp
WDkEAzvGPyPJx/jXpSO2tQ5hwkwZhva6ZJzTLygc3sqyKjf8T7BNW5CQvideO7b/
6lckMXJJlEeLYynhlJl0uyQkiamJU+1wcZdnS8s46lWjm9eLKcAr46exS6FQHo09
e0pHZ4fhs6zuZ6aWuzQPJjeGfz9EVZIqXbb4D9w/R6ZwNZ7vZYZL1IzOAqhR0s8g
XQYTlvypEJEulAvJNrPkWQ==
`protect END_PROTECTED
