`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6HVl6qfkAQhO7Ieeb/Q+QCAxqeULT9hYo1zk3PQl80H4vbjq7A6seAAYDvt6Eab2
TeeMvs5VQCkVktRaONAh8/xm2yyARuk0FslUFiBt3PGjVXcg20xk/292txQaNdlY
3kguYuL7DiffanXh1Sjd4hjgUJML57Wn2GOXciDWs6WP5LaDmY7U9fa2JWCfOVQZ
PUIt6GOFO6jhf0NL9FmIHPIyFoIpk8grRNK8pwScRmu8Be4hMx+fDWYDt0EEpmGb
ZllCYbimowCka1ke2soA4kwLwKWVj1DvxoBguHYg2QgMorVD1SydUn+x7OFwWtbj
BgxFpkC9kyQeAzN+sRAQ9a9mwL1Xhi+1FMN6vuJQM/FBzfi7T1ULazxJ10GKkz2Q
E3AHsOlHRWlme+mEIFeupdSA3acx604AitkyaYXXDzj1OoDE3uxobyQxUPx1TTLU
wstDJ2mGz6CyR8M9U3Yt2Gri1+dwLuXupCBq0Mg1XUXIIY4+ej4Xmm9dy1S/ipt8
IMixmEXTMGSKqfhUNIu0evfKGEBQ1kYXXktG85deC94UnTwNBmBLBOwmEKEiF0r+
F1ivjcmJK7zgw3rW/nyHbPCW3qK15aMHIq6+fYcucRcIE+FCXBVUVVavq4Mi6L5C
KtexKi+mEH+z2ej3nEJOnfmQrDluZSEXm9EJOtOaTRztnzZ7jiQtj8ftUNXtfiTD
/KVPmPsnyF12B9rHcKb+aTUaOs1U/kqzi1ooC0YK0UQxahm4DkfuiEPMZOQVBXIh
IDH+cu3wm/DNSuUVPI8VOtovmTcuTaojESfKXUqaCwQoUVHK5N3/kztRoNbeiCZn
0ULWeSh3RT1YSwJFDFNVyFBnMlHZBTsGbxtSn7Ze9l3XhknTTSapjG43TW1HVDrB
K7xjWFL5cr2m6/RxMaiX5C58JO5NJEuOZVEV5tRyovL2iTK6uW7WjLRa72tJWWFx
rOUc9aQVDrcNDakYSECF5ObGA5yld5l3+mdyruka8UfGbOybEZUVn+HMMBcrQYhe
Emw7hdRMIH97CVeL/aldYt9yRe38/6PAGJ+P5Pat9Im7bSkEPf+MhItxs6dmu3n3
Ug3ordcNj15vR3ceir3X7EpYOHFqF6RccKyKueZHeTuxQOGykwbTK23F4ceckjtm
ut/1VVeW327V2XMoMGbil1FkQo18A9Ixy1vTJe6znZQkGCLCFZKNjPWEheKkDH9x
aB87JthTPkkOarsPzFy/cRSWbLNorGNk4fb+AxSV2hHNeUvC2VSnO/c+pu9JTYuM
Dl2Dhl3vZVmXZlwPq5g6JRJOaGzYDM+wEVajQ7n9KY2uvTtgDOvVAvnZA0pfYiX4
NKL30KM8aR24xLpcaKKY2ts4jtXP2uQOghnP4f7ROldUYgQf4053ll9eXasFLMs8
SxkfcsWazoIZdGbJgDSsSg==
`protect END_PROTECTED
