`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A2nzAE0vyLnlFt24FnmrEVC4qYva/Hrz2dyX3WiTUyY2pK0+Klhggsbx56FfkV8H
zQ3yXbU840Oa8CqwzdQ58mO7bo/nXOPkj3+nSlmFrUgS7/WILUVCTYCE37vTZULh
yk5dxEC2cR5TJbtoO5ftGYsRRGxsPSozyz3BQxhtWebIPDSLdNLhEjAnJol+6AnH
Sa4mMDBpOy9ErTaptL7MgQ4k24TYAkwn83Ark25b9UcW/qsc6SU6Sc60bH3TWqMn
AXMjcRD3lOTSXsOllZJiOENVAAdmEiWGRbWQMl7y6+lfeKOvtJlMyOkkE1zXe5zM
KxsNjyYI2uyj7PdJUnNxQDqjOLqoXwL++jN7Sik8oCyqWiNfT1HwN1CL0iMvp/Yk
`protect END_PROTECTED
