`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sznFdxW8KZWc1q5A8AHd03DMLP14sjPCivDibo7YO5K124W0f1Dz6UlEjNxfKiy9
oSP9fpHpmwPcYeaXzO4xD84ykPm+nelk60pSjiXSTJf7indnBTiWN4X6baqPLjy4
Lg/gR4lZADLS048sKB4b8mrU5WopPj1pHsHKjfQRCyTCBLlq7wt5bMJawsbZHXjt
AU3m8vpZNt4ZEk2rtgXRG7BB5W9DSMcPAJskiNZ6TSDDrdD5X0+5HyuJKOPz/SsR
LFvd31fsSc8/eaUZwQw47ttp0Gny0cgvWA/+zbBwggARivFc1wPE4fRyr1+BfKsU
gNUPpFhy9E1L74MHvh5/dXbLpCOWEttdd8DjrcboqC1Hch8bPH1chENCeD4+RyyY
PKismGX83ToV7YsEXcOY8rUKrIow7eI/G9Ag/fLhZDzku300sHwD+q1cuKimU/rS
QBLOL6oq7K/yQj9+XT4wq7ALYF70efZDMWXnmHKS7gZsREn31Ae38W9NGWsKUT43
glTkai2maS3wjtYc/oXZ0YdpF6nWFK67s6tIL1j6ZGhBdfsKUuVxhjlZSPXKNygM
T9+O5EYGYZMEFOanWL/fQk9u0LIqOCJz/DqzM2+FJ7K7WXfPfWJV27Hni+K8MmvJ
`protect END_PROTECTED
