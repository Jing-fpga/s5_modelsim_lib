`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jaWF0vX8a28XvD22O0azrH1IYmB99zfuLxNg4WYGdxRWhN0kzTDPkHjNQFkj868I
ynV0xufdiPhso1dcwoL54gq2Ks3XTEQv5hxf3GZXR1zS7rDSRaHR8jKpHO5OM+fe
Q5fivObzqxZyjCrR+CQqFBlK1wG9/nEDIweFei8EmnMSzXPjI0mphGPbUMqP2YH7
jJxsQvc44DTbGAKqkO2xb/a4ceMHP9HKhe7C5ZVtkJr1iTRstw5BLXYd0jAdXC6x
NJe2rfU97ikD8brhsvpuez9hH1+QgzwObtFjEQf/zZceTQE5gTllyhjyQg7DR7T7
inauG8MzdwUyrcPff9g/8cJxv9Tb9PDeO3u8pXg0wIr56HCMhQF3ZFcZzsaFAS6M
35aCy0nqrqQfIyq1JR9v7SPbJlQphh7gh2TAZI4fi18vMNxa3Lklekn79Qf48+Iv
Jwts2hESgjBlTMt1oMX+yWzx92N292op815GMo5RuiijLF9I/AkvtcpGCp+znKb+
BtEkZJKzJj3B6zIjGV14EC9aMxTANYLvi11RfIwRS302ln4lvx5JFeY9UozF7LIz
6/8I0mDNlVN9F2CUfYG3utTw1Y7PpURWWxSaCtKO+Ijj55AMST+X6NuSRfCZjOMQ
g4tfseKwFoCXxhou05xGVdODtfkbVrr5qTXSEwb+37DOjB3kK3MRim8ZARKY/mSJ
KPQDuI5Z/zz0nJvD+GJviB/xKdElXB526pSkvRVLC8C+OuJIUB1tlrLUPBcHnfnQ
vFeFfLQ+Efjc9l/W/VocNspPyMinkJoqeeNi4gRWZPV94OTFUyZ4OUrEmHUhHgxi
n2ujBwfrII9noFR7D7uQlkC5flNapuJik+PgapnR8t3klC+wNi+EG3RXoqmHxX9B
SI2PqpgmwuF+6cwlqrMWMoJzrppzmR57ZnTXqcLQBi6idgx/kDZsUCFm9pWs3g+6
ZxRxOWezyZhXuFaagfbX/pnpZCK74pjH2fv6pj5UlSaHWcV9Pgh89FmFL/bcbrgk
W/56sh8tLSoxbgdWyxoWGkM6O5019ZGwUpCPNpmuqJMbr0CC/2IGDNzp/LuiyEGH
advyJfq9BE1O1EvY4S9T4Yhw+B9NwOVsV1BUt157IJQ7FNM7Dwyv/g7Hb6XhP+VQ
RM/Oyn5h56bQM/fjBBH0d9ybkmBovXOykAURi0gQmHqPJqM7r15+6UBQNbjw5XLd
rrFtumLPMxssH0CEOCo7ML2wwDyqdRrAMg7DKOIRpzJLrMViQ0HRyXNWToF3/as8
Qkv32+qgHn2pjaC1NGNBdVyz7pHzG3AmLbjcV3niAS8ZCLCdbsqaq/wGEbU9ftWM
sC6UnTdWQg5hQnhjl9KrOiu5jtBaBdECfWPvuDZMXOmCoV6TKTEOBspOkZGEh9wX
n1CDbhN63Ck90BkEotCvnZRSAmPG1fX5pxAm/b5k4B8Ae4YmeaodMaLA8m6YhLKD
4xU9jX46c4fnbA7bawzaQ50DHS0HiWR3c+x49y2rAdVIQugga/AvDxuL0c6WNrNs
JnudUkSaM3v2AJTdqYNmDNufuVeBYcKTnBBrpkDAaIWGwmLYg3+9+cDGFpTQCb49
foYlgXbOj59qF8JTWx+wEFyYmEk+iVE2h5HY+TWQ6VdRLPEvb5j5odiZ9AUKtav8
dxLpDixWECPN+y/92EI4hQOeA4WSLCbQsfZ9Oxrrg95+JN/XmFwPc+WWqoGWftYT
CL14ppKFgs8He+07cQLGx4JdBLDIpRthT1owoPGmXy0n/N13xsKn7SI0A2nbH8X6
r6LVfFCJzSc1KK7ZOufc5QrOMuFWheERGclS/ktqsXPVdmdZVYfZMX1LaRi0QS2I
q1KWJPPI/UDB4oQEw4n5FldWxNoauzb7zld9yNR5ekKsxK9orHkxMPiaaCnaD2/f
md0s73ypYAHu7ZxsDip7WWzWXD512hDKD1IO4P7lsyqEj1PZiA3XuGseOVHj0gB5
aaIuZffyu0+vWPh1YO155LIzgG26eyfGBZUjWfBZ35g1lWkx3NINmZqv7d1vYgaa
4RPxpMZUHRXZADwMtORm4BOJZCu9wkFltutgQ/V4rky8LoiWWpg/Yg6TlSq4SdLV
nXxEQnDmb5z/rtTWaUq+OaDAc9mfsT9jITNfSlav+pD/uWTjod+lHUB9K85iasy/
TmSKWBIsSfbq5QY+AUUtFUatLMfZlNBL8b9ucKs70mYXndEmzT1oDdP+1J+UfVda
U63lzUEIw1cyd9Cdry4ozxWkyPTa2zZSwoJdUV0V/yFR+TF9z76U7aTduNrfbiaq
Ej2RSYfrmIqJLNMuRRQoNKJUDECM+kbJXsx92guWgkKfWKGWwFXrfn4B4tZhlqPL
IAdrHrYvZXAd8DQtRfyB65k9kRynTtT5eHwrWwoKZRSZDRF2k4IIzS2vHs+UIhxq
7MGV5aP9jGOhC0ifdHVI/mqswLWOsLETUHpmo1le7lXR3TDK5jYTM2GPF7WGqiRt
P2ICS82Bh164T1YegYR5Hg9iuBcDXqSG2JUTTgEVZorcsqzlCZ8KufwwFj97oApR
nK6GdmGqN85/Ln2OJcKqQ+AqHrhiQ6RmZiqB6Ao67w0c5EgX8DkMte/AnyayQsj0
/usdIfDE6VXMhvhDLysCp3QlZd5OY89IfuJPD0/ggSFQ74oostwPeDjO41bm05GK
mS2nBut1PlOMaAnUFimskIeD4vpqclArVNJxjwTmMBVqxY4HpLG14q/oBDTx0HXs
L+8W14nOrSHGlm5gZs0uZmOPot7Oqrek5wr349SH+4oDZVJ+NHxyoU6+ILf84X8G
D4TEnjCPvzdcF4t/eoDzvV9fdmUcVQL8zxjqu5LVqJRdlKialmsBvCuv7lsZ20w8
0HbSbhN/Q4MpsypzgVPfQh1hVSj7fCgheUa4QTn4PfyK3d8pu8/8htwA1v5o/lNq
i7ShkR3WnkVkNGQZL6ViXq0mbHZ2AOLhmOonPngO2dqHS8T/4uiWA7Qq3koEz1DO
A+ZUbnW9Kj0Pm5buvNUPmx6j92sf+v0LwTGw6s8s4kk4Cjo3Oc05GtRlajrL0v/J
LBVBt5rOnEQTm18gHc+++3pJN8dcOMkGUDnEuUBeNAX0lzm/7IdWoXl92Bn6SIXN
1JlGx0tBA8Mb27QGi5XzjO+E1WrZcuLrlfgB21nuBZGSEbmdSHQB8s/4nm0MDZbJ
JLdQg6z9cyNTgBxybYPvV+TCwQonJIIAWGOo+hu+8RmyldjEbHhVvbg/1rtrX+a1
+Babtv9ijlE16nTWYQVRGKuurJT/H6BsgscAH3HQsvY8AMFf03D8671Qv17wB2r5
JELM+wyJWOguN88WegZVHOtnjN5aZ9whygSJl24UmyRA0YLZaFIMUrMHCVg3CVG8
xBVXa+dajQb3j8lkRI9D3gUjp0+8snxM5ay44aW/ALmoyc7qGY/Bn76x62380j9G
P1t4S7rg8BNexPuCtFFnbazuPVAyn9f8BhJBvb0uolqD98fmtv8/lYeYnZbnlhtv
FrTkZYZKo92+ooXnxb03CUYtz0zeYT0z27g2UeRO0EQYN1iKIvxoc67GxOPgJOUG
kZRbTLjEOT20svNEmbgLKDM0XFrH3l14Zy2bpAr/8yA3qxDXjvxyf7z8S4UZtEI2
ApmJ0i+5dOSN8SWqXPbO8z/OWYnPs4qUGYG1z1zs4/ghTe+2KVlLTGazIfnhZ3rY
CYNJZOjjBTV/ZJFlYGdkxob+9Jya7LKija6y/h9FzdjcITUZdD1gQzHw4vc6JxGO
oFM/T0qOLjDodEt5HajJNan/glAVyaXiww2YWqPSBvHJbLhRVx49kQKkIP2Jly5v
yZxeldN9XjD1oejdG9rEkw==
`protect END_PROTECTED
