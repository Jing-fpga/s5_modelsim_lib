`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B/DOxGKWIMfGE0cwO9Z0tbiJpPzM+AfjnjnpUhdsMar+KW/fIo6MYJxZ1AAUqcCQ
MxJTughYdwq0RGS4xFOqUxwPgq1QvKVXnNiUlSOX+L3wayRrA0youSJ6fhGdSzjz
7xyWZCdEVDETmagMLiuQQZs7METSe/+k5cGXXGMClz0WfpJhLnsLmgyCSyNSQk1z
TrKYX4GphKqMqMrLyYvK/DWlzS8Tfef2/KT1UYprAAxwTVb2zGMnwM3ozmNitRXe
lUcKgGFVZzkfn3yz/4t3PY6zbrkvQRVig9uTuVvzi3r8gCr1WjQABXse6QZ65n0t
jfS5CRxWKNetUaPJpKoJIFFAwa12ZyJHxxLfsiHoELrwsERF/b/5ruTjztlDzDaW
X5Ub71ETEFLCZUK5gyc8XaB6rEaojnZbi0SLW4Guii4c1D2f3ieE6f9jJRAEjTZO
P3u+O3/fsL+7EH9td1kJxHUZUfxba7vfjBnfA27M6ccGQCaxd/+vuAcKZfE8rGYh
S2QER9mn0ixmAbLAe0glDnFi5By4PTQZ0iTY0TmWuzjzDC+Nc4mwcFiNkOnNnszc
JRUcGspzC/bOf8DjnvPu9blKEC06QUxOP/cM1EXzSbzZw52U5VDcir86lmB2VJfm
RmwLNyNC5GWUwI+iG3mxexbQDRkSrMtpscjZDta0Sg8bJh/+XQwtDvlB5NBGIsVF
q9vBsXWHW0pUdP0v4cgznPnGWbsokdUAwAbHTTnl++2gTTA9OH2/BsxW4plVf84E
aIwxpJ7F2OhBe9je+hVr8TxIJ1oQQzpnF2ESNB/9baUR+Fj8PIjsVGk/40loXJY5
ueir9zCPKIlh91y68rBEN1ZiRZzObmc87MAP85SbZXkPmKS/nvONvdGBMWLSiZz1
xuxfyWhwTyZV95y5EBpUoDbct1RFQDwhW05T/ocPwJu4rJzYFHjICF7wuiqsohxw
5+XcQwc3gWSxuBZIZrajwthUT5o4OYge65oxgKFmBD1MXwRYkgVV6J+hGwSOKBbm
F2lmAXXhy4Sa24plcmAOjWESgeE2lphvTh73RMbwsoIXxeVE+r7hmGYPqZNF+crw
ZiYIIeJKH+lN5g9Ojp+q/cmbZZpeeIEoxJjyIgnDrmmF40eqPo62+kB/hPqzIkI+
py8BG2snM6wKR3+66olh5gUKDqkShcIU3ZqS+ZVVAUXvDmolvmj6mXGdV5S/B44N
t7jCKksd/d2I8z4Ewc7G1lrXdXVmoXOJo8cEVHTaJDjAw3LuImiEm/Ay4jGArCXu
Mxl79IlUcK2jHtnwlxeAWBwPxLUQZuzG9aUycHp+eQ/uzi4IRyLg2GXbpB71uiS5
IUHHzEP2OEMUbO8H2h1qkYV5985i00696FU5NFCLvHcGdNbnZUQ6Jn0V/Nmx7TXQ
n5yQH3oP8oRHGprO1S3QY9JGw1EkETKLKXB2F07wLJ4ra6Ai3FXs9WbgKHPMGIEK
WSkrjSuyy8UIOqnXKs/+o7qHrg20i/QAutQ+c3iV91MACeGMZUF84841D0KIrTa+
KE49CB0K3STUAsoY6p75CGaX/5EgaDNH21XJ5vYN/kRTKhOEPNGOMp/EGuslv4b2
ajrPCUzTLgrLrJCmOIKO8JRNccvbwOAwL69k3MUDSI7k10t5er/dwkjgjtaoF03N
9uAMSSG7o53b1+tEvpXCzTs8g3qzt1XjXXAEuGklQQ0J+kQjNvtycTbwtiHdjgl8
huMu7czoZMJc1tmLUpu9BtIZWaqH45+C1URN8t2E0FkMvMHklD7G02be7HiGct95
AMk1XM0e1LxhLT4XV9sPCxKHnbId6QPsgPPJ5dDw282ZnVTmuPKZVt9KeHkRp3kZ
FtM+hu1K40u6q0P8DP3kYNfqfvZeBidgCqhDagIuSmj6PYnTqDI+b31/IuIIU65S
ZAM99ppI5m2KIxvoY++4uqaVI6zU0nZ4SK6wNd4hYCJ59kb5otRK+Ut008rcHc87
yPmcYNhnGhqL7+Xhh4wJ7cD0Efq7z+lh3DdFVk0V4XGdd1ycEh+XxDccQ6GQ8uH/
4dvPCMAkX4biTTQnB96qAPa4shqiqCDSjIOtUjD7PSK3ykePNZU5aBRQ64ClWrWx
SCoSyUPJlD7o45U3CBBsceGVGKM8Qr0PGhXiR8eDCcQTZn9TNRc+hph0a2v7cqoD
gNmvPFgDMJbGzJNMtRelKQNklrth0Gjd2hRNbrBb5OK6Kiq1qs/6jHegO5Npm6Ff
6ILv9ZQ4eonPzq7w7H9mhazA7vF8elmSmHQ/dPp29WQUL+FZiVIz3vQKfZbIiFsN
KjIU6xKh+anRm+cWum1QOE/ggYlLr2LjQrNXdxwhN9SpoPdVIp2hvJySJaRM7wIy
NI6eGNRUfd69KNNGf8VCUnAPXpg/vDPgYbgeREEX/gSA1hmmY76a3DsHkxTfQ9aC
JMZZ7gs8yWIeQemqO+YWRodPBR9CYgsUOIGNYhv4MW6a1gLCX+o21m0La/fY/1CX
W+goVcKawioL7irvQ50K+QHgy6EGw4aOP69EPSrUDjRezHf9ZTOMxmxM+0rDrO9W
cdeVbtBHZb5z627qg9ltHf/lIwUq6SJhx4ZJBHAKJeWR9TiHCwd5JA2edjbpMRKb
XK1x3ZVl3uxRNZI55Bns08cje44qcSUYwIYRxhxQgDEB7kURga/1Hz/LTLPskZvc
y8YKmFeGdIARyVARboieOv/VubctvfzsaINNkMcdkTPN47ex1JxeGieW4DXxa2YS
csrmUM3n2tYvU0IIzU9R0w==
`protect END_PROTECTED
