`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sXHwL3VpmKP8fRxeKP6AfPS9uAq6bGgrDTIUWf2VIwBD+xAUMuHm6bI9KXuhUlVh
IXU33zBsurTTlsK+Irm6G3MoVwCKP8RHKGYAG4YqX8MX71p86osbyuT7L8smegVI
xPllDyMUSvUkMK3xTCRLkrYLNRJLFNutr4wxRMx8ofXcD0YrrvscuBa/lD7k5C/9
FX4tr/5hgEmxAaYWcQIdTtYI58yrbZ7tUfR8wsu3HTsc0jHAGZ7hXr5vY6JytGmo
etjatj++EshhyQzmKp6WkCo7N2QvPTXmp3BUOgDZ4cIuYSvDZS1Jto0k9suXJF0A
hPblCLbNMcbHQ+/59dRR1yOmBAn+EPMoB/SFViBBFrViVVJMOwo/G2luLwgIEr7n
AClFlXkQXSikS5I+P3p+xNrd/Z6PqQXQbroJFRJrP7S4oozLGwQ69hl28Pkp9YLL
d9rhXgajUETtjhtevAho10yUopvTA/m/3FGn4eru5IGyyrRlz4USP6gIjLaNlw8c
Nk3wLfOLo+HjtRtrzH0Nr9oXeR3lvmv8VxqxqlC0pP7X5S2fVNwX7v/RlmSCUTwA
wD9Z0GDb3SLXsOlMiXPGF6sP/pHJerMKEI+07yDlqVlRbRcilmSKhsxsxXB58YWH
zaScZ4yffLsPGR7AQ5dPI+47rwx087fom6ZwByzev6cOtxSXOsVWMT7hKPmiTCYV
W57oX1YDTGMfYUQVlE+LNnx5ymk/payz3lCT2JY24zHirsVOcfIHfhZ/e5F2VjC/
XZ44RpdmGSby3iiusCrMuJGtu+6y58vLtNq/7JGg+SlnPylV7mc35lGsWj2Ig0wP
093o93X61hSxmFTS4O7dGBYiicfzTCkgSneupkjwehoFvByLjaBdWP34m+c6N4eY
88QypQhr2l8q9mnhLREBvkJhBY1uwsvLKfh9R0OKuAIR3lWm0kZKU0L9mYczIPFo
jMhDfW3DvIXRvBEQA5dGHuX8IFLpP4b+y+OlAU5kAJ0dQE4pxGCqZHoMa05KCCqP
Df6HI1qc19bBbbXYy+rOI2tVXslmcaZv4WDI1G2qcuRuZrV0mkGUOOJpBTjEPUTH
N6vZskmIus3iYSBMigr5tUKh9SruJY0TL6WgFznh4oqF1QjsA2oxwdb6o06B1JgR
PmhHA1enS9FIPym3oPRc9/Ts2QYn41/XCRqpk4kJ9g8UuRMdunwaYOVp/qst7lv1
we9L/tqO3K7y1D9FPvJ0S4UzGeg4So4NLiGmcUYyShMM0U76/qVql9QNRXQXZEhM
Kd37/1PAEq5DESWSGdD5KV47QTpxHr3e1tb54lDC7JxTxTmEcipZZtNeLEEl6rWe
dsGGD9r8cOwzu7ODfk+VNGYwgFkuzjTrQGOCgbAq5pDR/zBEEEQe9rOepH9+BVqF
7/GU0+Ff9oiAuePFIWo/xh6xyKPrs4m0Ode1ub/jQmOwmBL7p+C6NCv8kVW2q7fA
pHqoXxsomDfEHFu4pLoByA==
`protect END_PROTECTED
