`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NLS9W+NXCo60PthiuR67vcqs4OHDhbZNVgnFZWdsFax6nzTo2ths+X5f/sE6ZeEO
AlsOt6gIqxiaUWpEu9Pdlj9TRYe/yaeW1H0lGVXg+BCd25xMxq1c+RimsYRdwV93
xlJGvEQvaOf7TLxMQQ6UctpXZtaBkFPRhv5UmszF+OAc87v+fqpe1dhH03/bxve1
jA0uPaBBmJIFAPsAsaWXvI7zhaEp6L2hNPN6JMMpYnUQz+3lHQsw/SvCFilWbsQ8
F5ZqCA8diRkizOGck6dqKrP1lQLdeBEh01WYaqTo7J9PACNTfXjyQr9QKYDe4Mm8
z3p6FsIqADLwIC8vLDMvIs/gUgefb/HiVcKj5eGrcw1tUHxw7J1lDrbfm13Som4d
DdqX+rVRwtxA1RxT6dVQGCP+1f6gJ47v2EzqVkIgEilK5NixNmRHxR9+DDFAMn6I
O0qJiRSAJovIMHwsyj8JWQEw+IJxIqvo6EV7N4Sxrjbb9nYsxZDUFgKSZmjUm2lr
SUmCb3ybPMGfdWiQsTl5Kr66guUo2/5ebm2mCZdJUam25EPHp1UKWfcJ2Kd60iJA
59GOPh1/o7khb22GKn2RL3DcazvHtlqruB6jsEFkYyAZL4tDY97wquOBWp6ZaYyr
qabG9tGltnbCxEe4FUsmtCtap/+5KD4qAu4sYX3Vb7Cu7iF+iI6RrSo2loJ47Qeb
fjkqC614zmEDNobuiLp8AO+SUuvxd3q53DkCzjmebDHRB4HYiMkVBMwfAzcDCRk9
+synIbdQT7R9NL824/+box3Ezk2EU04Ldpi9vixUHvb4ZFRiY2jPbTHjYncYoe4T
oiJNiyKvBkyXQ982y+UoFuvFhnuVIuuMOvHvdEUKID+9RV1kXhJX3r7B1+dtoBIo
XHTeCsDj8hfJH8Z9XSBul2uI6yFbKjiNBRUCJ8AAcN6Z9OyMv+C15q4FezuMo2rR
gz00LD4dtSpOTXQr7y0Xkpms2G85WfqPAZIHwBoucOdNdhHedY/YG/c3nKj3pDSR
Oillv2LMRdb9zGp1+oX8fHqgzUHWNvSFOBLh0zG499qZls9gzaEAoUzfTv94Yixn
zPnN3kc1xXh8tMXvlWLtMp2gjywgP2bltcX423iEpfMnmHqlrZAZIXt4v/4HxTsp
rIGeeKcp2m436aW1njjP15Oxg3tzTRVCdAwrV1tVc/8ehZt0W3yV8HI6IDgiEH3z
6tL2VXhurltCaRMg4ZMiEr7kN9oXScDUBMUQZ3838Tc0Nnex1zifZfx44A3aDOaW
KUs6C0z2NUyk7/QZJt4GrlOvYKWUrnqRaz4j3l5CMa+IrGEDp3PK74a0QC3ZPcjp
gtHhqa53sgSX1fHf65lpjkgh3CbbZgmk5rxlnhXcB0qUOnAgi/pcC7JiHzJtZu4b
TwpXG78GzX3JVdxHX2RP6qio/0LEOI9X8nzfqSqw5bPnZYX3w1IxZcPPdlrnaKl8
nWVKcirNpkKNE4+78tpxZDv8xGumtlKBGihZ7PqoyoM5ihkXhIK7clNtAC9of1c7
nuDd3h/K28P8FHAtmKAes+QOBMjqhX26ACxGuHiUYt3HhXxsB4To5QRSHswix5q2
s4PXyf81bSY34t4xOW657XgR2JFmMqDQyUg/KbW9oKZJassjdXipmOk2TdcWn8Mc
Q5SUpuHqlgzlBPoYvnQDehOONfSXdQFij3urf8y2vVX3WbJc4SVk3HJs2Ot9nxSM
aAmBh9bHuDC1338vcoIbXmzdSHflqNOFSWOcj3DRuwuLm1V5/imoJECtXft6ZhLs
GFKWcoTyP7w+JtGC/iBl+05W/2bvE+S45tSoFbKnn+d34HgpTTfAkPY4K4/pixQ0
gFsbFlmSWShngv6nYLZ/4JhcMaoT7hUE+EJtovjEd0V+8JRQUJqn0dOlCy1bMHvK
gXkjbsit9KZTlWA/YfViCq4WR3TBH6aVtqzVzzmLiSE7Q6YFvDMuyfuqDAop75+C
76KcHLBuwg2cL+/5MBX35xa5tlCdDpdzDSdjszaKORGpPa0fxIhUfHlQT2J5vgLI
pcHSjE/OZwxrUlqASJtrkqaarw823Kc0EgZj6fziwu8QvX71A2e48vnCXHJaNGYm
gvwWuSnRYc+mBczoULhH0NKEzMIaEpvUHlVVqWMMO6GEek+g92JXFMXVjt2Apl5n
ePOSJVlJjQ2PxpxaK+RG5WOdFErPHFhSc5c4gfO7N1MhfbdImn6BVf162Oqu91CK
UaoVYS1TgA0V4CyG3javQhnRxqNoM27xZBZ3/CG0dDM1QXzwPIZ165yN6CqO2VCD
4aUQkxkA8ycTCbrhdV4xzDpijXF4LBj8edlREWLQ02vhTOYddYyLfzS+Lbp/nr2K
gAGAu3Bp91tcZG1fOnAkjvDDhoLLe6FHv8ROSZNIs86bI4G8AvHYVo5KcVnvicio
UtoSDGj0KwDSoGemHPjyt5Pv6TeHg7MF5T9mINrkUMQ6xokbO2xF22nbYRiPVF7S
VPLEnejYrBtYcJV0rfkeuGO/x9mSX6CzrpQftzGIEuR3ANh8KruhtcnUDDDoY1Dh
xEXo/xTDTO0y52tPPMhKj976wP6G3UahIHGFO88OEVOUW9w+MRahRte4Abx+Nj5j
68wBc9RORC2PodJjwA5YRfDO94yD4MhjFCQxKUR8vpsuAmDC1/ZtQWLKBa9sHCch
L1sgEIfFeaHZz3o0gDIIBQxEutdC2T4xn9OICVKmyqXWo5x+UL/8qRF26fYBCyvO
PyxLahU2V6cdeZIstj2YYH9Im3dkbrlIDt3YEIzC/LrY61qoDOD5R2gUJbIkQyUf
IMRkf6xAFGlWdrUH6TNkUJKzgVUgwVsyKXsYIBwTLBoLw5IP4OdGXMClSiW9Pf6v
MEDhj58kEsdVVD9iokBY1w==
`protect END_PROTECTED
