`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V05FjiPFwsOcH7/N1tYVopgD9Fb1wsihGmAg7nQbzAqY74wSphD3ahyip0T57GUS
YEfHiRBMRHc/sL55eK3DfgmRvw8rKOoH4uLwSERCJAcYlHWrytyB71u5uPYgXWyr
MvLfYAshE4N1JV4V+o04ZBs0BQN+GupFg6VdQv94o9614GSybT/xc0wKQMP6nbhg
b5jO7j4zUQdysJ9apUqwE3tUhxPILqxEjiCDMmKGmHDc6z5kjPEurRZJOqI4+vij
+EfClARCsQWTwFHhYDWIxdZ4oPeTdsyC6GoUTDUSXoyjFZ+lojVzkL9IYFIOZv2E
uTnwn0DDdkE4FpdPKXS/5Vk3MGVQLSUQET5KO7O/mnKdTaCHSXFAF/ipZG2JYdkn
EJ4+WAtym6Ku8tNWSlLrA6GGw4+ivVO7gfRwP7cdsC1F3s0ny9w4KGmfSue6hU0e
YNX4It7Y1js1wNvlBvNqi/rSkQExREtX0o7uZo8vJWSZ6bksuqGhAd8myGnbJWgn
UaEb/S0Db4t8XaCGRQV88EQ61Tm3gkmGx6vGgqyT4Yav8+m3fkhTkp7bHfjigssD
xn0lQxLt5J5GJEInVgSApx8Lc8YTbeBlmkPWy9QMAakXK7LYOIJ+71pmlxI/RzIY
Dcy4bKlRU/UU5qmlM6IZoW0v5jmU0R985XDiTfE0X7a3kjYTOyuvEHW9XZd8TVb4
TnroKGLdh//KT4za1QndIEvK/7p4cgw0OEJLB0TNQWD2XaleBTis5mL8s/Yy+2e8
LcGigLMtTKe6DslEssjBN7k7Amsw7Hx4hTMxn+7kZf/pMGKXn6SSFZwTe+QypKb4
Iw+6ZEO1Vo9RVF6S8dTXWsiX0vx1rp6qE1dG1Gbe7MPuAXUXe8F/byYpUUcByzjS
UIlu77CteZtTW4Rwc78vQEl7T3KRQZVEEVHWkxzz/wgrRgb03YqKSMlKmyL55sVx
WhPxXqSK4WqXNtsXxIQMaZ/3HihujLGthDwgO1AJXigHP5KQDLA9evgXFZ2vr8Ya
Cfk7Y2mwEs6zDJnp4bGVlPRTvjpUYYXejHSeRDtMu1znTqIz8VEl/rAtaNFF5w9Y
ukhkiPVsAwm3sxLPx4BnMcBYfpsCrDhxW1+rfqX475zAoOmmiuJeZYnSeK5yPXn1
JtguuE3gY15fhOueOnvfBTJmRTIWMxITmVeDPedOqK1rAbnqmbiiCBZzFG3wxpet
JZqbdnMuD4sayRQMIlRxjZoTWjZpVfcXsJ9wL9sHd5lVJC4bmOWzm123Z9VIkUqM
8ckKsQt5mA5dDrnn45m+/84GtXtOqk82iwMF/HCmjiEWzh3Eg8MV7+HB5cD19ZkH
3CoUWcYZ/UPMv+ImSgB/Kw6WmAIXzIV3wWIWk+RIX77Z0ZS2Y6pOY2axYj914bmT
HPLdKpMJ75zn0sTN28Tpfrj6wZHGEAOMDIgiKYtl3uzc4FrW068WBB0tC72rE+S6
Q5yhZNaF03su1C9D/0guHWqBzWnC8C8iQ+Iv0Vw/ZqtN34HO9HvSyiR8JWhtsd7P
iY5zhiZHqKDM8AGiFArOPVb8+R41lxoJR2vv3nX5Op8fPutH4WcJV9zT/QEwBxBa
0x4Bx1S+HVfPZVvOfnq9KxKSNjPOGSVcOWL/jWGaiLh8ItvsKmPQyw+rZsvhVf8Y
SFL0EkWAzwATwljajPjgizwVOLnjSziBXAdlmOq+cr63GDmXC7ftxXRq5iHnuqFY
LNPzOIkPVC/x+YAj2BeXc0yPmstBG9WQPSatyGNhWzAaqmXS1JhBbm+pZWFQc5ed
8PoDgRE/IzxsG7iVk91Zwd6KBlZ6EnaJVfYbFc7XQuY9zHYWTPEJaFV7TQqXKjh7
IAPDczdFK2xGp+hTvr8zeh+79O9EoL+TbpsPHMYG7N6O2UdRPtKhw3ugC1bi2pFh
MZcoOQNsHrh/wnI7nbIq6BjyE5hxF/A7nYv0w3JoRWZkVO+Swl4uNOKJdi/PYUGs
kmpzN5KAGeTZAJx9fNjl1jU/YgytB/3cVqBwXQ6SM08kKna0bqi+QsOY/IEcQm03
Pn1f7xcEZEVh44EZG7UMxtrDh84tawlOct3daH1NsnFYQm+ckT387HNiX39aRonj
WOugrQwkLU1CO0WcxKP9pxyVuLStKJX8li5S5oLpoeh9dl9VRRmiW6ZkMzke9XNL
M48BoiUSw1Wkhp29YDOksXnxE+04y4M73EEoqFb/6xgg2KpPZTn/IZfZybQGwBOo
WdZvxRRbRMPYdlHyC2dMQ4dotJw5H/ivTceuJ0D4UMplL+xhJoU5vB1ugl2GNR61
2Yr6ZGDCRk4NEP5nPaNg/v6TbKIL+DgXH5YCSwueorCUvY5goNK8zZkGueBfm3SE
/urApeupKtnwLgpt4YSIKDjXTuzscr0SGTf0PR6KhoysJ8uHDdMLn37Xq9aoEP/V
d0rEoMPmV+YkkdGb7Z0B+tE96SqmKtZWkaH21bM8FvZzbnRpfRsa9YSOjJJqNXoy
cvXxEcHlSkhdcGFJzaCvXcDBdPxOBamNez2h7fs0PKKsS8zjArWRV3x7o1/QjS52
6+Cl9QhlzRYYH0A+LTiYz2bsaZC0+m+fUNG+YIynERRhr31xgNfI8X25+WtNrOvD
yRzxP/lf2pPrgKfq0dCkUaZifRd9MgpHjEv9yYny5BJ2iuD0jANnCmeQnPA0iwfQ
8ZCAejigGOrKcDdK57Zc5GQ8yHoAfiRTEa2MLLX2j4ApPPH0s2pIp7AHn2voQC4/
/EY7JV5fMV7twEnQh/52wUkYb6v8kxCCKIxxKWkw+n4ICWW4g4tqTBWa4vo+zV5c
gEExEgx/u5C692dpvjvxYteWadhctXUyTDRAWoMADoKHIn1P9cWtHN6PQDYqRfHZ
0ZplWBsvMQ4S9sy8nosRqFhwXeDbwPHFJ/TqNqxjejMFAZRN1AD6Or2JbDRw2T3b
fRjWolcj+ZufHM8MREL8AGd1Daf2kdMbTD1AoCJQtpHFEgUZsrHZJMWZGyNi69EI
XJg0kgJ+ZvosFz4nAzFHzaaUbqfigRJpjhh/rJX28aks6YQFs9cIgloqjgTK6d2w
DsZ9DUKBFZ0ivk2N3a4zbJIQ8aFFe1672NW+3FgN/05v1exJzH2u3sWG2QxfmB5a
eqE3oVyucWZ5H0wV89QieIBYIYkFFVcTecNbw+mqKM0pYDi415vGhrhmzrWhQOx5
ovthp9SR34XBYDeIv/gxlfxpsMLeq4chXq3xSLbx+3gtHEJliGx7pGOSTGhGY7dl
e7KZEGTbrVjvSIfnD06xkaJ4Dc1djDlIqphhvOoZWD1V09XcKYpYQ4qmCR/H2Y+s
PvrhaJAiFyoOnGY3AtQOFMa3u0MPMqDLAYaxEHbXXmIReexDqpuodYATOGuYSs+o
ajQZELVTuJNZK4Rupvcr8FBydfK6GRAo1pJJh6KHCPJKGGAtBHn4JmJv29ibqvDZ
35w8Xs/TV90sMH5cbsjPHS9zUny9GxlGqNQ9VdMeuTD4/JK0LiWM2evE76LYK479
XneZLMfdTUzRdwjQcu8XyfiCMVRXTQbnaUosj7iLtna+u9PwBAd+ONeKLFpq58uE
JEpg013m/FnuNxCmrxPEM/g6Uw9GRKPAW6LnitdQRUCYqDYRrs4HJZ/HM7D8mh+R
dMz3dkkbo99Hm5UlJu1uSIig2S/RL9MWbcXwBMUPpcCACzmbHs8qS89NtKIwGnnq
oJWBmUsDSaSWLmn6q46iz4LOmmEHSrNWJyD+vy2YzqxU5yuL7cL4ntgyZ3KTm82j
Y/TTcmCGOAecl8U6MA+caDFKrnXE2+3olvgA2e3vYB7/JiBRk4JEqU5UAi7Kiszw
rLHv1OmMvmHRX0pvFs5lrg==
`protect END_PROTECTED
