`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yS7oey72MoQBQXEmftBVu1fAqTLWshozQZCbiT6CJotSyfXhZEeXJj2KChLEuYC5
+BhgsZA0w9r96BuGvSIsyiobkilq7SRcuQJRQOsrPM+j9Ouo3oHEtWcwQj5nwLxM
8L50ynTnnTVLngrdj3RqZMRfpibzjS8DJzFGffaenEgEnPduxGhro2Ola5KAnddM
4c2zmXOrpWTkK/euXKPd1tEWyEWzd0MUo0FdrQ612CNifyoCpaFwerSGW18MZYn5
No/jrFjxE056NyLMEQjg6WVwScJgpBSn2mB+Iz06eksQ8kQzywNGnZdtIZUyeZhK
mmJFEW8iTpt0Vk46r2A+Pl5HCTBX2sZIkkCsmLs9tBnFWj0BAV4tjeb8zt3RAH6L
SAeqXuXByqT0dWSD7uy3zXjqloYQOUZKXuVkH0yRaF7GC9wmeCMp+3cQNLVpgMTc
0SkgGalC280Qshn1n+uf6pJ74abXmE5urub2LQqQvxF7QXw6vphHPXHR3ynKnQXp
l+KpA7czSGijkdGso5j199UtjJLeDvaVLprXpMi5U1l6T/BHwhonreUR1u5LYEq8
KM3DjsPNI25hHXJKB2gaDAK0rdgOlBNDpL0Pkqekh5Ss4ug6DzZS6xv5FzRvNQ1c
Cx/jkIj1OeuMDiYDV1uNANGZTXFp2IgAEKvzmjvegtce2oNqLsfMfSe5bSAIJMP9
L1d1RNpJHdU4tvDW7ymCp+kd3TwvW7wGY6SUNuYvj3lTzPbCh0jWnwwYLai8VDVd
XafNVGkIqjgmt8hlleEtS4UqziVnmC2jP2vjGgrJX6c3lPK/3NYsgJyt5GgQcP2G
Mv5U1G34J5eUsvQlWZf2z0CZ9LOkWqN64AZ3dsNTl5T8cIr7wYE1kJKhbD+3w2dB
n6cKDkdKhh1QMlx4eqb9awgPmbBwzFm7/wFsy8n8LepwWi+tZCanTwj8sWQK5usx
ENXRaxl2fzdOjKjLpzbwxBI6jISBxwlt1yKYzKEwzrFLh1zD5rAhUMduSwpVUYI8
CeErC9tjmrzEJxKk1Fwgv+ADTpyscO8WNy5c+War0f+dK28TbWXEqcSK6yHhFBCE
uTQkhgYof9keoMhs9Vfrol2BY5U9+L7e4FVj/qX3hcrtwztPAEnIZqPWTKwe2356
yZO1K/d7HnR4MzkyrpLQ35NyPtz9VnQ1m3y/Z08/nlYGh7PnwpuWPq3vi2iuahIj
ucIqShzoMXxc75jkmLxRDQS42t3/Lqhp819EvqdNEiuGoriqVGyBbAd/uFMAMLBr
GsK1Ska8aIyyDUHul4IlAVEqPsuCB6UYaPh9Tr20HkiMJ+aDlitWZ34Y6Sl8jlYI
pF7e08VahGzl4796I6/0yfrea/d0M7nxgvJEbsG3Nd1p6N50NBHjPvvFZh/e5iI+
RHC6STsdk+YBqqd6KXWoGjm1t7D47fkJNzK6SGwKPZstI6hwzo3J29udScE+4dBC
wobZYmFvmkpnMd2/S17kX8/NNpwNu6sjiAjmprLclU5M08MWfsMvYX33owpRos8S
ORFzF7B/GkaSJ5klbZ2giMW2uXTQZ4Enc5pJOZQD2gAP1j2qvdmhWuUgGqcM1WoZ
URS3u53ceuHwD4Y6nuSmDXZNWPopJ6sl2RoFqLU8Nyd6Zao1fPaRMvBasf6dmbzo
VXVUkLX5NICkMp1EQAxk1iEAelyxGwOjSs3CynmwiXke6ocM7Thsn2SaoqsTsDR6
EowPU1uGkWcqrXnC7Y3XW8aPR9FtqUmxdS4wn5AVDK3DO4k/2ZD2wprXMEuDrOGs
QDCpkC5v18YG+InSoI8xyd+BTaX4N+xfDcZG8mL+q/iHq5HMGxEUA7m16IfELDhc
OItlPXSUK7UaHl7S07xf9cUKdw3yDpPShnd9SLGDltzYGCW2UamNUIXVZ1lLYCGf
IPSzdddOXL2J+CMtlrVTA7VirwbQo8WrHnT5177rsOg9qChLIyyRlgU/aqkgv/z+
Cg33LKzy33K7TzQEtbVcdUoVaTejA7aDW3ZabSorGwgbJssR2aqhDt1sHoCpqLjO
uIQfuC8aA0AWu0qKnh2WJr0WQHSXDa3ixsCBj/E1UEDBkXWxbcEKbVJsX7E0ryTD
DeUSAVwoJUAoRkT3KikYxBczrRjZQe1v9wN8GI17NfY0JRTy/HyEq9DfWV2Tej/S
w06kbVkBjsCwmZc/ALyBMx72iQA5li9kmGgUt5pffrJlS+hBAB3LE4F/+zEJbJGK
IGZoc8gylJGX6TwByqfrETAfkCVpGKsuN/XQaR/6Q5nIv5zkDyk8I5sDDhQwBsAT
zlqJnzrElCErSWfKDdcfgsHMmMcSyuZgqqMMwVW8o0amcJ9OIGUvCE37z72Tf98D
RBhGoLczkp5JyRoD6w/qz2HPWwHf8OHcQz6ts5jaEXGaaCWKB9YSxB/RiQK5B5gC
`protect END_PROTECTED
