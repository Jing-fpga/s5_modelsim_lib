`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2659jBSEKHVNrAXQbiVidOm9KT9rbSbN4Fird5SmkUsgCQGGTQXLI/dxhvPTuVTM
8i5V3mooI8cHyvWPqfzjwv3dF/oi6wsm9oVA5R0/YCt/f6ZtdamWo3oDQUQ30hoS
xvWJ2DzoZAUFtqG1il87oVsptFeOfH7TY4Wx2AH2uPZTBJvxsneZBh4ogI3c0rJN
jA5nwCvQ2OMV7Y4UqmvaVftCCPKb3MUfexcQ0Gu6K3xncxn9MmrB2I8wif9jkFjk
WpEWXVMLSR3XmWm2q9YkBUWnWHdXFy4ItjX1VDPDUoSsnar61f+Yih0fFXAmuT5q
AOL7WA4vj/ha8E+BBeukbKygUvOCkB405daT4BGh47aC0vHxPv1Ejm+/DdIRzip8
`protect END_PROTECTED
