`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RpyFhRdqgaETfSdbEnohixalU/mf8PqF8y658OcgQJvZAhsa3/rVhJISzBAWlXfW
w0E0Qoj2kkPQFgfhn2RuxYwBAWEVtmJdJ3QIL1Z61/xxppvEytsBYoEZYw99EPbs
WU5uTZgAjpzufaKJ4Kz0FFl3htVyk9X5qQEzDLXEzQkopA8imZW4hAxyyH+GMSXg
27XSc9VBespskZO/tp+eg65HwoE4BG6sMsf5wPbR5/muBsu/jG+sh/izbJHBbZKE
J7OrXgGADETQImfF8vzcLj/Mk3nLu1yEVX1LSNfy6RC2vPwhjcBtWVMR0GTEAEsZ
JqHkbV9ioewzY9qHCD/b6dTytRANKXCi7Zq8Ff1X3LyC0JkVML6jnFrYimJK/zWS
w06UTW/lqmTlqefqGir2AAy/Q9kZFFS8g275/PEJaPT3MdMs3aMv2dEN5NT7wJi3
b7Y24UmlQ1lMTrXFsPESLrjfFju/GazAdvrmfHWXHoOjqyY6rL2O7gpfW8k95OnE
T/2guGgwYICurk1IBuqbdoyfukzRdvHq6KUR/OETAVITLZ8sWuLzfJXxb7FEKD5G
lOhjdvMSOz+oyhQN5OcDhNl3d2Zp/zg5UdwJA07xnzhmTzq97xhjS5CV37ygz0Di
sLJLKGHxB5VOc7W2eRjYPY7VBjNmxcrlGQGyZGWmzp0XtiA3dP+dA/59v7Bt/Ngj
7vZkFnSbtB3t6lT6QwNKSEJTEB5ozAQ0774965K8yBcoj/OAV09w4TNY1IbLUuLT
TJJRi82U+2bIDLJAPqOnC3s35PcojnLFODd0XmUO62jMWC4sPY8b5Wx4yerJGfaC
uuAoUZaHktAcDwEnsGh50g==
`protect END_PROTECTED
