`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JEDdy+tdRpbK9w/qDeR2RL3aiCAKcFaDoVNrxSJTkyIqpdAM1DhkPHkUD8W6og73
WtQOciIL3cYnVmfNRpYwZXS9CiRMf7FZW1w2ZcoCJopoLkz3gu/GqBELI2GA6xhl
R+D1ef2f7SZiCyxGbp35dTPwqVxwlm778Ru0M+L1yu/GzmJs6ykpUscfhjcekouV
MNEl0PCuEJcUiV+Ym2O5+0R2UAsktbrZ34f5b6WSo3HPDfZBzOXRBMBew2Hv3ijg
fO0eTiTL2iVHSzk4tu1L7lcYe5740uBnjNJ0dizip+ZmQEe+A20QecqNslu6mCp/
fsB0PI2TCXOsE2aBgzs94cWgLhBSc5n6GM5ZkI3Y0IqdKtoajCGZOUmh+ICEyh7L
0Ce2/7LQ8WYASU8c+AjPXRW49XHeMCPiersfaKkLLT/7JhdWT//AKbZaWkm7vhqu
lVbRWs5s8WOsmHcXUrJie7+/y3fPtsPcwYnIU8LjVWhsfnUywVmC0GjRp4CAwCfO
ZTggxVAOdieqfK2BcqnJd0qEw2Wta6cVrc4+3RA2mJJeUb3nxTZHkkbxnWjwGscD
wTH+wAlOaDf5hpZpIB7BNbY5itbbIK2s0n6Xc2PRUxOQfAzrAhUePEyiXjFFFHaz
q5Er/rYELooj5lHCCUMN9gHOnFXZa+72pzeaQwdOYUzGQsYbgflOsd6DE7jsaKz8
LCLWiEitdpigOc3NjBjI8z99Y68LDoKTpcO437iE07vKN3gEc5eEv3mbazsI0nLj
hKR7MaEd27Kww2cm8oWcuLySIIfvsm3scA182a5sWnrfmZh6nWek2p7jowdjNDWT
QR/l0QIJUR7sPnYP8/5al0O2hTydDV5J/mvOp6nC6CLFoyCQVM2XzPIC+PH8Om71
LwzG0ojyKc1tSeTK9z4FZJI4nBxQZSZhNVE0RXcYH4CjjyJBP6RLI4Ntn9Zow+IT
IaWBNK2ra3CijoB/xlwlMUWIZ2u1ysExedipbmMfag2XapcC4zuWW2pZAw32fkjt
/wNvn+GZQuuA4hR/wI4sAUBsmaFF+mf6GreLwdzgbwmwL+CoyVDnyb0MDzdtWi0o
125EqAUJPDfSgxYVv7j7ibYLA5hElXzqVr5PreqrCuVYj3uvhRKtQNr6ZMxi3D35
+2hC4aPGytQZAzhA75kEtkImtf1KAMOhf25mrddllRtZUpf8Z8qu5XnVBDIUxhPF
s5e7I9PunS7IeC9QYXV2lLq0ObVHOw2MeOcYL8MMR4VaY58DWujNIgfzeL97Cq9W
DC2jKKuBzasRvy4g+hdxlNAXs54Vg8US0Atz5a3dqf0vwPnfDhuZIz3aSR6xcxmO
F5Z0RA45WEdtUv+ut4UwSyyYPUUq0CjUgik5kFF4tN7sZbx/piebHL6WSjcN/NP3
SU1yOghp7rb71SmPYVZBBWc1XSIpUNdci0I8PtvQZ4bXOmJj36FKjSQt77urXuVs
XIxG4Da3SjTWSFzravQUqtyCttDPgyVPbUnWy/z52XAFr3/1kOwpR0s4jlZEXNzq
95iZOVq9IhbVsXof7ul3GNbmj55Z79XtyDN/51p3ce669hFRkmTNVOnq5qGjL4A1
9vCYzGIhXT1TfXdUn98I/8q8sDJ9NtAs8eK5KxLxEaNZhXCzdkOYYby2eWm3SEjl
JAygK1G1Oo3FYZtH0yZSBR1m5nscqtgIj6uXzldA9Xj6u/D4K4Uj3G+ggm/wN8lq
UwTQXRKgUXpMZRgvxxqt1ngbpUilF92+6gAZa0rVzA/fMMcYT4Iz/DSVDfl7FFf7
uU+zqMvi6l9tgbMyin5LYc1VtVz+KjIHH1NXTLN3+2wKrhjmm1yLWmkeRjbxI+ko
uuMhya8a2lukhm1+1bUQ949LDHnHOM+3KJR6jHxOcBqrF2EejZ8xX+d8LS8cQwq6
QssWi5fJrBXSQ8Cedc7IOsh3MYP0mjckHwqs5/9xCzDtWb1/t8aiEn3Oqx/NYPTx
ba0AaFpmX8XY+uV+YI1k5iA98bknA/+8oeKXeoBWwRBhiu9/FnAKeABoZti8mllu
tSpI1jw58EvrVZBnfLLY+8axyIyQlVugg9JQh6JC/VVbD5ji5HVgyvY1JqtP9lza
hVOJ0IKMA4TNs9OvKQpWFspE8QbT7HExGTi+BDi0cd2Ju1uv6+7jFkzEvBEUl8wl
/3LzYd2rOlbZ5+7KsWYFIw4YJL+McH/BXqgnU+Eu8FYBlhmq0vBsxBEG4BtRvdfS
G0A2SiqXtVJt3eS/GWJw3Q==
`protect END_PROTECTED
