`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BDtWryYpLzr6IhEm19/g591I0n/FhXlgEfzvvAK9xBW6nLnel5gtTr4x4O4qQ7eB
aQb/GqZCBtCQ8GfeDCvPFsTs06Dvc+5WMpdq0k8HwP6lSEvscGWw9uebshvqs845
AuBQYkOLUb/sYspv05nKwCLkDwLbpESiOd4eFmbpIBTKopyKFTziRwfe67fUpI0r
/XM4NYtWDAnePnn24onSL5iSpp0L21lxsyOsyppDnBmyqUI58UlUg4fZA/65X+/X
T6FfD4hxd+MTFVejHsv3jSvDDQeJCO3PsMiIiSslgUOhyeLQHWMQ+gmekeqYvbO9
U2tS92nMeFd2vX6o13VZPGBj7WiqPrmtEzaeqZ85R1sB1VX1ZnRbtyR/s+NImdnx
+XQjdQ9GI0bcqFj+FnpwcwBbgOBWpdl75XxmqHiKdT2/SC8xdT/R1HEI+Ks2kVkg
rP+96NCQ1d9mECsIzToKsoQgK9qFGSN0E2gpXLtjOna1io9dUrAx+JS+rD0Be77Z
czXtmcfBBUJuWxdkVZopv7aDTvl332oTyKsVpFw7TooayKtFGClCRIb8+L6pJf0O
7SvaFtJsQaxmL4hG/LXsJHjG8Js0DttyH/3kfGRqi9WsV4lGYWn4hPAQSiPgcocq
hFF3SYSLsVvh+y3PMrqWtRFXmXFbnh6G1oo7X4zt4OEgdS5+2t3u0eHUvphWaDlB
fjQbLLIbbLcpWXfEF10H+A==
`protect END_PROTECTED
