`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
seRYb7K9upxzA3PSjpNAj4sPWdCPhDSYu6TlqJmzwdvuWIzsHw0natdnytnR4MVW
T5dRRsb5qxAKHjKOiN6b9RlVqGPIIq5Pzu0NYZ55m5hzBQNOrCBlxAbFjxAYvqQi
wNb671o6sUttLkq/7Nxut74nw1g7F5GpHhzFZVkc5j7/kBys2VaUCZSydXslYi0B
ay2UK1LjkldKSOfP4657G1WTjHWzmUOPg6Qg7YS/KrPBo4+17VBzURVvbmt71/dU
VkQhfbDoxtfO7BAGIkrtkP17gwrTmpLzympj8qaIXcneVGbi0T7zc+abnbSli2h5
fzaHSPOpaODUy8yqF5RwO23vcMUVc8HPV2tomnkd0qhxwNmpypfqVSqPpfuwu6/S
JAJB0us6Tnsq3FrKhV/570oA5G3s3Ydqgy7ugPljFhWAiCHHXii/oRJd3U+G7SAD
8UoLoVMv2M/yt8XGg6RnzLoiDzpF7I5wgHymAabuCgaYnbqpPHkebylKRXHpLb9I
OKuzLALOmAIKLTkYYlj6qiiipV+HbJIac0Dag8vunEKtF3bpp/6pCg0HDuJFKgQN
tErvNKlfUps9iW/hXMhO8T2H1+S2vDGApGohikjYtP42Ke/dbRSYEulDYIT+MuRv
1in6JhlydSoLNfCje3vQ3NXCKLHQ5qe+n52yNn7+n1aum6/m06VNJgEmkwGkIF8R
zjTeA3LWOFr2BJFSGxRhLheQLKoRT8QCbLFALbSI6Z4tIqPRjB2Jo0vuWMw6jTn1
eJGM+VORgzstyO/Qo2VsT3tP9iCoqk+Ih1nrk6Vwjm62Mj6rP2vXMHw2BgAuZQ9Y
`protect END_PROTECTED
