`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GQb+PbCAPU5XAF5DxbUwzHcYD5Lq/CCndWkRBBSr4Ajswnq6MpXREcif9Tc8B/2i
UIQxq8Np4RmF8uPcPBYD0WUqHCJiDopjdhlmGg53I3FfIQoJJ13uTkSGFKHyLuE7
cVYuLS9FeWY5PjP5CGU5Nqicl1nINJ9fw3l8Hz6EuCbasRCm4WoGBlSoi2QEUk0u
DOSscyFTC8Lc8SoH8HS1WzcfouufTxqrh/mhu19kGX6I6gp+M1j6z0ujCBsm3bwX
xUOwDfZF6KE0jsUT42jStIz5QqDDuS/b0yiasWdLJEBnp4KDxQg0xyqSEz4JMGHO
nhCSqFkmwJkp+/AQ1R2+wJnEY7i8dTLtRq9mObg+sR/UYf4k7wkJpbhrVVMz7rje
V78nmNpEnlN4mhAqBi/Y59JfM1gb0XqnFF1B6o2eTXJZMGKuZCQTu+w3nUV+CiRM
x222KkPHV2bverz+PpYdDR+XwiwZlWGZOAusw5WWEXaMIDW4kFKptbEEqnmPQrxk
MJVjz8zLXNGvugNxeT8vzoAqktMiDoJuNt0Gis1dAuNXHNrCSbmU56E+m8A67wUH
Q9f00Hc/5JSKzyIPFR6Cn/nBW5xeLc48Px/S+ElTk86wm4iGIgJrjShDRUpWReIX
8rd4vFF2Vmud2nm8c2Pyry0Ew+oCCXqmrQBvJ4hfwCRI3Tv1kj46g7tjauE0+j7N
ncguBQhiFp7eNTiF+C25mIi/L5N3kvXC51VSMyufuItYeTCBzeUKS4Uw6XxBoKm9
BWr1PrL8yBN9ss/uN1g5GBcAa1F6AadYGP3CIRgHuzpf1ALDOzi2eSnLf/43Bu6g
l5wVEm2dfek4CYNBnW8o7DfS3pMbjHESdgz8bRtbmKt/OBl2W3jTVAv3aZdesTUN
lxYSZ/kw4rUw9zeZWlhZ6zMbtOh1yP8z0uSpdvFPYstb5exYOm1BijgKfHbcvt6J
D9yu6R/cnwQWdeaz6eZRrn8UrZgZNcCamtgIih/CpAIK+h8RDv34EJZ5NAu617El
vLfwCyNYz2sGCQOS6aiXRRDJIrIT3LwjpItmEtulCgy+Nd8WWr+iK1wEgvdO1/RN
BzhMv4VJkx/i+h/BPyq5bjOX/Y59AjKnYE5qEGbOml6AGMUSgpKRqzk62GMAg75J
tZ0aqWxGWDJy8r9eGu/IBAx6wwBEVzNW45tGJp5D2BKl7PpITL7p/nF5dSZQxq1+
huazvqVlo8GL/fuG5PAzQfwb/B4/jgOOjrSBVtLUFc0vQqT+c7G9jALYu7Lnluuk
ImwKk1Zwf7CcM+AMd5vGODTOje+Yp3a7pluJwdMlCvJth6NVVlTI7+GV+aQu3uYz
fWGnGFkO9M407o2t+9FJqxAFXQ4rndKWJoT/DYZoh1BgAzEavDF8hN6MIghEELTn
Jq+Xnl/36NHgkYOq+0fD+d4ICRv5/weeYpJfwMiKKmpkWJH/HXVDJb2bNMC5dY9C
lJ8Du+UW8pWJ89EeO6k/uT4ikigS01uiT+Ib1HCJ+vPwIGIdgwXw2QeNzrtjEJTT
VuFCOHMzCEyiREXJFuvwXHHuVJwiQNDDMW9FBfOlFeBdxyikcEABukP+mLSq1OxE
ROYu+zY7iUaCDbf+iCGN9hzBrIqrj0Vp7lF9TYp8aXTldKBiGKGWmb6lNzsEoBE1
GuUqsOyZSjVpiAYOiVKaP7ysUegnRIe+F7P2Y7dsFYnqAsgdn95r0xqygQAIQsgQ
TGEwjDq8PHspHgkGLDHVCqceExQZpETMNol7JasSKbMpxHpHm81QabfLIHaZEesT
brve3Y6+dLcrWs/mDPi7wTw8NMrajI2WRisKgzhM/TAfM/z574qTclBb0Z6o/47z
tfBUSDK2mpAfxUeUWTN0uxWxfyFSimVO8NDUQIdUjmtR1tD4Jo2A+ZqPj3M8a2de
01jCUQ82BfTddzS95n1ApgSgDcbBC0D+SB5UPnM7rA4Qk+DRggOEhTVSo5Q++o5G
99KHGT0lpipvW1BQPuff5qMxdmZhn1uXTKkJ3X6H7lG2XD2h6lkeMerK+zkZurTy
Pr/OSvureQZnVnMH90nF/sxhmrijcyJ1fr7RvAHbEVyfz7raFrRWBJYfNeRCL9gX
sLXf/k4Uhmuh/r7k+GxQFgOuIbza3NqjpQp4XUvH8em9IQ0kCzG+WVSZg6N5q9cZ
I5XzfbtjtVSyzoXot8Tjton5E7ZY50imPvVxC4RF2+oZtLbD/nOTBas5MSRxer+h
41SVW1lwys0CmAIPGoqEqcVSHz+D8hwTHW2Gmb+s3CzHKxVw+ChhqAvESYFQgLdZ
bn6usAJAQfJ5X4qgJW4ut92PX+2r+zcXmBzUzaCwhUpeEkZ0IqLlQqXojmVl5kP0
bErtizZ9YzoHF8Ko3pX/lq3ZGp2eJEYTzROsjF+V705k1DBBL2tWP2qZP0SlUc6p
jMqMiuDbVd48ezV9/RxaukegAdhihvk5gJz0jnE4Gi82CiWEAdc1bdI5rMLqzkhg
rq26q8IFQckCmtH4xf6xn9y0XpNZDbcgZO4qP/8RmKzunOM6ovP9U9xeok1z+4jt
gASuLJl/V6zewxE4l5hSw8YYTptfGRUpGk+aXq8tNjgs+bXPnbfDO6sqf9EXoZpE
V8GHGvJLPnb+xGOyOoTxO3mweBHF1y4D7w9VUuijN//EcIBtuTEuNLgCqyA2jTC/
g57zqauR1HT58rr8SOPo8vIXCWULM8T9enPog3tnq7vz7F1shRvmEw5BBAOawXQK
A4gGsjEwqKCX+uR44SKs0H+6wELio5g3kaOHByzdCFOqv19Fd08C5Z/rNrzXhaDD
1QxEI5HekD2/qsHyJ4cL8MR0xduWC0MNTLYuYH/FGoosfBemyUlTJtXUmdbYd8pS
lW4+jFAr0XA1hBXWdyYfHPh2XL8ij7z5sweARHX+/6eOm/Z1e2yLGjHlWmH4nocj
F34hG4WdKD45OvZ2jbUPIwUQkRhnSD14tGTGG88nSusQEUBQrL/Em2s1MAZd2UbM
lvU8V13q1wf2h4ydNMT4RVmadNZyHYLa7tgRy8ftpG2SoHmXtxhbyq+aZ82QJl5u
FfVTLyuPLRWjOVRp/bjsC1NPoF0OEb/sZ5geC4fM691d+3KV+IspbpYzcmqfxFI5
kQ/OsZs8dekku19IElB6TdoWhEVk+t2oK6rfTp+RNDzs4PE7vqPfKR3EMY4qWKLf
30RuYbEbAZxk25SunhM9RmJiO8KEJSPY9vzh/nPeFQY4TcdeNItc8iDyqqlSfi9k
VHpkm3O7ez/dLyFPWbyUzcI9L7oVrdB/NCtaoy3ZW3RrtfD8X+vMGqlsCTrrWiS3
DkwTQjI/MlAcOfNJPE47WWkpc814IWzav3z6A6FkedVm/GWIQJS9L7HWof1hfiP7
QkK+IpaCed4Y2wXoUk8tSYDnFsK9WjZUScp9eEljQxTk8RhbaECy/4xNFV6XoIaI
3KqVK1k3sedpkXfo/YyQNOQbpDF5A89Ho+BWL+/YPx+OFlGxeMvclE9rHhsIJONk
FncDO+LTMghGjTIWEvxXsfZ6h06wdTpWonQPy5SyadwS+Xedilq6j90kumorUnzq
RBD1kZVByfl06HrzJyT4SuHoUegv8wu6g0bmnQUOqWLwuqlTNykToLz23XswJMvb
lFBqmj4kJQhP2JtZivuQVukkkGmIihjfFm80+M0hYZ56bQoEBo664OMsNn3bxPsH
aRFGl3Npzk/kM4gY4F2+UCbTGZUVTuNALQcOMc2ovIbxiOLoXLORDC1jLErfW0ou
xXWiG9f7nxKP6canFMbFkMxlB10M2Kz+hGgwx1ncNnpWN8v/szeOFEav8P+p/r1C
gRvctFec6B6BUh2Gu9lwaQrOZm0CInd9LNDdxDtlrGuV7UbbK1HXx+rhfUWEPjju
ucBhLtWyrByNFwOT2lyy6MEx03BggpMXnjZsXFefEk+KRDgccDIpokDH8ui5AzaN
qAv8KR+yyPz7jfYC26M29N4LRT688Hete4jEMJTGET3IBDyl5GrkwkOLIVLFoTod
0wnSGWbI8RWXSkAYGu0TULe69F3V5ofTtQ4/hsH0YN0A5N9OWMLrxMo+fnIdvBWV
LBZAetU5J8MSpkYgGGyQu5RXXcKbjWw6XFU5kN54Djdlcv/mQvXC8NEwXDQYWsZk
Ul/uyYQ4RJpGHjwOZyheCQ3wCPpJrv0zvGFDv2EskB4bUrFuXE+TbPFRr/bH7N+1
2HsWhGFgjatbBp/R2fChLbOXRMu9KybTaq3qo7oOC1R2Utxe+YRcnzfowIjO7EZz
KoJa7ZFL5iwO+O0oZXa4yHRjEin1eHHQ8IUfF4RWHzS/eCOfttjGOuR0GZwB1XXc
mFzrCFaZx8we60ItKzD/EqpKX0t5O3vVp/5Mx0h/wLcxGTxDmo+ZF8/h6MaHMxuv
reYO6RY5ai0vf0vMTfs5e3LLo2x49kp8pDsKplt4u8BTrdMCxAugFLEdZymFDuy/
taf3BO5j2CetIDxCNwRaO+PcWh+zuRiF+HPonYZedPO0yvAu/zu94JWcevR99QUQ
WOEL/Proc0gpq4NoFA7ORsgZnZA6bZ/vGJKyeA42FfR8LxrG1hSEY7ogq83Wl6li
P1bT3soqWpi1rBSLLAWwwi/SJd+II/16QpI3od4iEIJLkZd6qvS6Xr5A7iSA/O4O
K7ROgX4mixC+kxhqVi7PbNRrZb1k7Y8MP5CnHgQwvK6ull+fhNzIGvaLOBc1uGpr
1f9mVf/YYPt8LGa903QGAEU4L850fKAwKxqGjerChVs=
`protect END_PROTECTED
