`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v2QUmCo4pv68wE8Iab54BB+aEK0ealDdpH/Y/90XmdvsIEP5aepl7hZuV9uA/dnZ
2mWIc3rsyEk9S5Sj0R5lE41EyLf5nlCyiHa8rBcfPUMxNTgG2Nq+poeMSu4/2sQP
uMvBicDM1hCPNxhVNuCQWMexu0Dxmi6glGCV7HcUhMhjfFa7+aDmpwzmYz2OrSMl
55LzFBI1RkmxYDdIP7cUmVQCMiu/hjsorCGkFCebaImOKjZymB9IdsUz+65f2TnA
Gnv1cLJ+lRSXO8sQK4W0gfrS8FbPuFVEVtGkcG1PHqw03a0UGuENvaByCd6IX5gY
PuVLRIkbaCI9O6GOpHylUkLG1EBgfmS1d1o83hR74hQYfX3EjsGjzdnt/MwpM3xg
FLqvIKPLFIKoMiSj9WWqlz4hZtBGwbuOStvL/TL0RqZ8CrhubBf7yDbbNgfAfmlT
7FXUNeEgnnemkGT/0TP303HnFoGnbBbmU1L+HznNpQ8mZ6RBWDvXEqTXf3AEtAPv
tRkvYmTs477xcUySbD6Cp6W9ZlucAyVmNLKW5ikhfIkaOWJV6B6OHE7OlnFeZZdd
JOYdEvSBIg1maL2FzXtFXLSu+MlnmHpAaUGOd8D4X+nUlv6bVuIc8Paj6/fLxXR0
vffS/61Jc/0rT4dhyHp7w5gO5Kn2QfPPSyxQb94QOZazFZ0Gxt8Y4bBK5+HXC9gl
xfs2pC9eZD4pJt0yEEz7xcXyzb6pT25Jk5xnLfi/6f7v5svK2e96gwjwnJv1C88m
wk7q82sytgSMvxlMx5xfLCkbI98n/uer7MZXTa311lMzg4h6M23p+19EYwfLWqyw
OKrEYd+MkHdcYlTC4KWEXqLlOL+jU8bQkT2xxFBPNsBGp3LmHO0MEPqDPH2/+FCd
/lCMQ/eiBAgjTI1OSMWoTw7oXHnREzVy248omnrQxuEKjPIzre9thgT7OJqZOO+C
A/k1hao8vQESNVsNqya8poef7dm1LeuY3HdNIaFx059Sv2dqQZG7i1p/fIO/rrVs
zKLgHwoypO9cKItxBWvuMr6eAsUb6JJ3TB01yNdpzZI=
`protect END_PROTECTED
