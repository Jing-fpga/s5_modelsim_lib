`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ZB7DJ1VGjHoDOpfc3Iga46DsAKfX5Z/Ep7xuYCuqcczZUY0YqDWepjnjPF3pV8y
Gp9Y2cpmEZflr/TLRjnio/URefLA2LrDYrhPRgk3JuN0ZbspnLXuMDUhgkf+162R
gGNqBDTg3GVHugDcl+cRmpLiOqqWhcYrTsA0O2anvm+j1/qo9F33UA/ZhenIbomJ
F4BzDUs0duIo4I6QTXRBqbXMyM5nX+0+jgJSYdH5hGuFXyuZZ8TN6IAcf1xtyjXc
ngUUTmNyTK53rJej5P5uLyJDzberEsVMe3m5frmKToP/oTwp9edwc6pvg+Ttb5MY
PFQZ1Ydhuv0kaMMbAGCuw4jHW4K+mhS0Owhyj25xwDjlq08XPKHUPjUVc6EwQ2/Y
OM8qPKoEgfME9AFqMWENAEooaNyc4ZFZHrx53G+JLyhKPqME5b255uMz/ujLB56n
XdzDpawdIroeHfMtTklHkl7zKse/XUwWuqfaQqQgrM7RYEtfikf9mJlwhULezdQG
vIhcV8SC6rK6wgLO81H/JAoA3lECZw25Dem02G/0/4cAK15ilcwzpRnPneest5Ou
NmXCjL3nnHdEFd4E9Da7zO6LO5niy248kqtBEIw/qkWID/E3r/0uvXehr2uSOxUS
VJ3V2jr3wRGsLckHbKjQVtrqMQ2xPUaxvp+MjZBhezDboJeT2CjOL4HYnyON4ZKa
hNFAjvqLIjLh4pT6N+tWTUwluuLXe7KIBd1+fWxrU+S2+NfxhZE+oanJZdQj8PN8
K07/pn/82Y7VQ/YIrnuBYN8qzamyzgScFZAqT4IifrXveTiAfl2S3SD06x9ea85M
w22PU5TeSj8KN1IKdlQhjbwgXSaAvZN271wLi5M6YlwNnoe6vGGHZPWUnAjzUs+n
KNCnCPC3Ehc2HbggbVkwY8S4IjYogqE5ySymryzJ/fZmzMWngLoUI0749ZNJ+Ds5
jyNeA4B0RzCeOiBCEM4Rj4SX1nHZGv7iAxUJbrW4AGI6R+s0JMtfenlQnhrkcZCm
Q1gFu56UBta/LCsNM84ieMzJNwq9uLZ2/LNa98zTHQAqKqZGzUuvjMLRZkJ5giWF
vtArnudPC06Jt27FGoJTKy7BGjDD5AE6J74pAJbfYP/3DND5ruTMGPtp+d+4URKj
EdHA+sHSL2DUSsCDuDR+6hCba1hFAUg105wyuIEZhvjJ0K3GjluQ2R6q/8TazkNX
9FjaETwwoMzCpcWgWWybFnDbwmqLzyoEDGk+M4jFcLw+fns5ysIu521+JCd5MczU
4tVwWsZngqIn+EaOkEOhAExtQJUh/4gJvKxEQtFHVipr3EeMAcTrwiS/1BNJK+5W
1voboVDb8cANLHbrTRdKkDbq2PFxDPD8RKmRmNH/OTrc6MqlTf2odA0sO9vCVpHm
9cPpbMcDi0yfW5DHA2Kn+Dyq59W8eYfUR5bGeinbxuPUkpW45uT3YSmwBOAQhTUd
sQ/EIdoEmuKC4/03IToTXZ+6zXDfy5vZHiP++8y4Xmut+E9ydvfL34xV+mO7F6O3
3rnVyl+aujxslnD1ku4mL1srGrFHe/E8dMpViE0ky4tz42KfmI/XZF1vwJi2Ekuw
EqPu2Cg5xpFg2jk90C92Xrr/vnV8nHz767XBbZCqteSVhXV6DsFu0aF0YAgYDvTw
N68b8SwSkZGl6Jh8FMo7A8jb1StI4C8eyLh/6RshGAf5FnotlxnZjRXimCM7RJLZ
k3iJ8y2f3JoC/F4sEvWuCADSurAHBbvwjg0aFTYiV6gZaUezMxXDT5nMY1tPkFi/
8TMaCEj/OtGrc7oZYKkxbvjW4d6sPDexjFgW2/BdycEBS3g05fvrFaKdw32Q7t+u
+gRvVtvC1cbxpg3tcDMvVdalQZzJFlxutBbjUyNFpuk=
`protect END_PROTECTED
