`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dzFLL6vq/ebuSvIKPsujM4S1wYZZ/4jyLEUmkaSxHr0iUuQ5pfAwMUw+23xS+Jk9
NzZPZlARCR4bGYmfEB/v/sPe3farHk2QUdDPVNNdgCkuELoFGLvcTPm1jgvzfcxs
DZQv5sB7UGsB3+mt1r9LHgcKBrPamQ3hGvn7hKJjuCGZfx+gT7iDzS8Joa7qfc7I
TlKD0o97YS60e2EMAp7Y0lGb4fDG7ig5b2ALPY35PYFSP1DcrEboMWHxopg/S1Xa
YproyQ8KDUiyi2Pfed9b4NxLj3CSB36pmCehH0YMoHxQni9MaSYCTg3bC6lWPWdI
DN0r68+ksek9TUEvFYurqwqGyjsS8rC3Ecnk+NYCKzzBBnOXNXbEoA5O43kg4PVd
/KwKuBnw5KE7s65ai3/Q+hbnOjAof2G2adrbgcQ403GE6hOtBYOPa4k9glWGBnQC
`protect END_PROTECTED
