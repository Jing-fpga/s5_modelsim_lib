`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XPRMXaum+5E0Cnbr7B9V7xuRD7cM+P41yvnvC4eVF2vgPvv/SeUqkSZqADih97C3
R0ySvgZaVS/LEwF6ZbE1P4ETXFBLDIC0tNY1nOiEZK6OdTX6pstJ9U1fAQN+cq7h
CCv2gHG+wkxeoM3+262sqRpPzAZ/COVS24rb24tsP60MD4YUvA8rIwRfx5GQUaDN
A93UcjJl8LDxyFk+/DyN+00wv3Ri9fpTGLsAIF+LgsANCVh471M9ERauv3R9rLD7
lMGbgkLeT1+hbEMjPQlP4kJl5bvxShE+OXRXv2IgwkhK/zE/Wr7I0HqR4UABtz4h
CVNJFPKPMOH6C6gsHfGV9gqJg3tqmSKnfA/AQ0bHAULh1prgqm/QqPFfnu1FfsXx
0RCDuFybQhGdcX3BDJuwNG3ceQa2V28Rv8dEIphJowBoTtVSVdXrv5gtAbUEzkaN
Xa7xg98hoY7uS9NPYdYUkwnImj+w+E61m9ntwXMscx0RQeMNYlbryZgUXUMh4UGz
i29P/wsJeFPJXUrlNCFsz1qmJuE1P/7qmZ8kSMn7qRb9Ew3uIC9NKDyNf19+855I
wNSpUEyZtq08j3lFldCv88I8y6m426+2bzm+28MdmkAEP8Cu89qGGQuN2yWfmGJA
ydNavzrhlmAp6LW+9RwJY0Q5gcTyenmDGOwUv/Y7SMlafWYoRs1acEwe609jbWpI
grXwJmvRlt+Ldhl70yMwcJWqDdfGk206p6jI4eDNk6HgPjbnZtfcQK/RTXXKF3J+
GhxRUTqsq0LPNZQJ+G6QH/8y+uHxBo94E+A1bs8FVjumhfAlDJ4elYE0+Sxc5zf7
zwZNWq0mLSxfcW9IImlKv1EAG1Fe4z2UqxoVrxtYsp+xF+J0z38vD7NgR3u0a7u4
vCZWuxVI1bqYyI8wZ/07wzZzU2SpX3VsGwhdVtcQ+qkWS0SIYBk63hncRSgR4o8s
5eXID5l3et7fQgz37t7HHQ==
`protect END_PROTECTED
