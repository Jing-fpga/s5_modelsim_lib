`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ppx9kdVjHoxLYaNSoY/nboBU7fjVvvuEBMid5D5QFmE2RQjdW4qJn/J7aAPqhlqN
Wjw7JfuCwG6IkMTXVj6VLf38Y+53McXvOuSNQ5+2RwRz/JOI/l91hm8rLUCkH3zo
HjWc4SwSoM6SQcc6pDH/8bbDUUkqqhuANEzFRedlcv21EXNj6C8ycmure8TtnUad
8p1koRGyWxLNZPxdJb5JNu+404A5psc6Nh25WI2klxmP1xSQ6R+ZimzbaCTrH/iY
yZRCRsVLYa13Rv4bDmRBPsC1cawA7oTclJsm47TQVaua1nw2B6QvPlh6otDVj142
6t1k3iVxgfSujE78fDAVJj6hEcDfL2VThCQqwO3+MUAPtuJWRj3zLcfWclIGUi5o
YEke+1qReE8Ir3gAXn0FYasH6d2SHML80GOFSmyBbnAiwoEa70GLyNnBAy3ppX1o
O7lCgdXAAxwg70cS1tdcfWe7fp/DlxBhuhDpOwC26+u4wmXLegwZL6mG28Xk5UiH
l27LMVslGNF6tz9C9PSEXc4KcjTnLOlhw0hrZsIZ0Qk7kkllE3kavY65R39fovud
cgCGKjAFI09ZVXzlE3xr7YcxW84hCNEKf46u22RKJmxqs0UnG9+0qa04ugo+sMBw
oarOKKWq+xCa5+KzB2MrQHSMvUxlKKelV3zrUbiMX41fmKYwdeyRedgwVLHPtNX8
lT16hz1fcQcrneX1HkyLJ0PiMiu4atw6Cmzr3Tk1PqUhpemw4Uw6hGrzqvXtGUtN
tt7U24LBasAGuH0HtTmyw0+nRMqiIChfnAIUtD6aY6z/FfuRbJTKWq7ycvuDNaS3
5nKIxbX72icBq5SLZta+onsJ+QA22MMk/taYZFPdXaIjPi5PdFyNKfEG3M3hP7ws
YWwjdsBQYxTw+A6FEc3VdGGypuVwYjIzpw0iyWszDZw4+yVVTLtY4yVWQ7ZZUdZ7
ME8y3WWGACA8VmaUckCu7qWL47wInNiFJJPpRhQucdju3okVeSEKhYfmgUAxtfgF
7xSrlGeYf4Rxp2csdzRFXQ0be/HTkj7PUxQiCgGIAnLF0FHe2KE9Pd7TNAS95CBD
O87yvK2n0o1HKpSPZwyi9A6VF4M37pXK4wpk93oUj3A6tc38q7ibEG+Hg7kEyKy8
lBE/Av0xK+SoBEUi1yhqXOL2AWwA7EHGevL4OuUkbSwAUzpDW2EHtoJwi0snWNgo
107CM+7s55HMwLLex6xwIONfuKhH7ifeLbPdBPVmxIU0jlDiRf0Jox3gP0HGqY2L
r3ENd0MunmNkdGGR22zBo2tr1h9gSIBgW6q9n+t0Y1etx+RW5yJZsVSS4N7FrdqJ
hCaauLhxAkMIAeqjB5FWqSCJPagcHf52R7BYIsu32p49UnctX7dXA8U04CXtLJjf
oQI0Mk8laTCAgWDGALJoK6yPZjRVyobns5y25X8xlZoWH9cvGxQ/EtaSlKOCln0I
dLFFnnrNajlAQKJvyhDSpKoNO8RJqP6F7QVvzlooHxyOQCKbQHUlYrRS4Uq0hz73
bIqY396j7rUbu5kfVmCIMpXv373jtEInbDNidwcuHB84DOGqg/MjuZn4PQjcoJ2D
6WH6zKTyslwJD28L0P9BPNFWtI0MnmfHUSDU/tUIlGVkvOgCnfK/LJPHLW+YzzTH
YwfrIwUzkHkLbAmn07NN3GdIfk5iowLB3GZPt7qeuHUoy0f+GKG+DoYWt0kUpdBS
gRVbyVQFRtU2KSy0CXwEwjqnMDU5jkV4laqo9DmW4D9ab7JTTjpGw53JQuGTKUFQ
abvfv1Mmoyke3/tiZ8Qu197GmA+JxNDZA8wc/jKkERQTMgsA3f1Qt4mY7e0pRZLL
Htn9MRtmeTcX3rmva/SoFrpI+F8vfjWJUIHh6/B1KY13SQgiGvZ2rQ5e4N5n+z6e
PspQgYCjTEsalkGY3AyXwHjPU/Fc003+CUgoHmK9bL3ISSbHuRdonowWcBI3Tuc5
DU4laL9O/6KAJYm8v/tWDEYhyzaCDgwGjHCrgqhXYuvqLeSzRl7n9T1rv9nsskxK
FPxm/B4wURvZVOgA2vVcAFc0CPuw7xuvV6HoUO0WAJsgJTQW4nh5TGYpKqXOhbn6
cPlcrVAy3ahpOdQJ6UKBipXEHTHm4v4e9UQYRLGbt9XMamF5mkSfXLTqoD0b3JSg
0m6+f2lSqa5IUfUsJpApJNYT8Eu9Kb0uct+hAsNFgG+o7YVsAIzi7dL/eGk8MUSR
auPkX8dAiAnzP0nnPW8xt0Pps4+jvxV49+hGFlD8KPCXa8+qzUssgVXDs5+3UmzL
gkjdJvTkbaDkIj4lsdSuEF81P25hm0VdOZnaJLpSslQ+wDK1HgXxTtIWOwc7HeCU
4MdNeubfOlmYFC8mWSbrY3XhFt4XfkqN3ytOTTdQ8HfAkjUVYpsTLzUrr3Ej+YmO
Le3LB2C2C3xfuiaoCa4kCGMqeVMghSBpsSiNj5sebBVaRmYbgndJV7uABtVlJX8b
Yjuln9TCTfl6FgJwk1kdg7w8KVThIwTSp83Z2Nmia0b7VajNYwktKSCcarOac7+n
oycnxMBJyW7bf8rZxyzINgMiMTMtMbf008euxf1TwxRQcxlmAjZySC20chk6wB0q
PLWGndGjndSNWWZmz5ZsffIVhTyW5ZemBu20m7iZYpGlaPe0Q6E08EdPHR/2FpLd
grHXTtpam8qcZQdxCQlo1+UeRw9TDUmX9DpqEJVr5d1j/qmwAQp7iIJw+ttzHI5l
vxAkS1mHo/Sy6WTyjSwfirbjINQHS/mHH0qM1o3zH6OqDLn71Ynm3Z9LlUQzWAk0
V691AzEYLW0fS6sxwtEZx5LO1X3cjqClxMSNMLktxrPFfMEUjPJXhFcHOrJx8HGr
3Hk3GzDaEei2Yn1J7kztwxluca8Oo0/mSTmKnyYUSKpjYLm2UIOUPLoMIsvrHTnJ
BZ0xYQ2lqY40z0Fe7uTn32gmq0hvBEWuaPTUtrkZSSatE9wBgsa6mqOmDMksvDAu
sKj0i86YIiPku8DqWo1wJK7mrZwOqN7DjlsHNsniXV+J063KCFtnAmaJGiZDxfE0
mjultQxf89beXql41WEnRk9dgofZ0U+oTotQjMq12n6TIM/2JmEXZJJCw1QlUOPu
+wB6bW385o/LTU8XArQaup6xSpqUpwpFgM2K7vrS9qPiD5Zk56x+qtDjgqbNyj5h
GLMArERaslSww6fKbDE6daO7602POSchyyyVFbuscZ9ouAjFSKdm1JEHArmYMkLd
WTurD3SCUkhCM8DaoI/iHFdmwz1NRZGMLVN1vkyjKZDcznZpctzUexXHA9iv5L3G
vcBQpnpXg6fPIlht6nKjVVMxfxCgKb8U4miGgRD84xBn4aSf4Y/6UkaNcmn5QtT3
10S+/6y8OpvgPWLeeBvyzFxSBBUCBmxf2DuCwtZZrLVkYcjT5JAOhbHdx/kTzxwL
vyrf2ddIVpqPmzdkakjcXkhHgePImXFug5mfnLwJYXxHHtsjn936+Pv6copvUss3
ru4+OdHDyk1cjsizJJY0XSFoFuat8XQKgugiFbvt8oVaUDd93kBegLysrxCJ4CfE
qsedzN15XI1ee+NZz7a53sWM2cvAlke4Ue7ym30GgYg/CK8qcKva8e8KhhOr/3mT
Zo/YSmIqLyqwLudgTKIbGpZPu1PVL8xdj/yXw7zy3JioXprzhUv6DVILVbkW0+mz
ZdZ2urfgUGBRGjeUqaQ26gqXmoZVpMitt9ueEDdD/4NwLS6L5p61qYWe1ERdPo4z
q50BTcpD7axII4b5WO0ECz9vLwuQjANbRhwIvXaGFNBzzUViSHjhe9zm6evzCXtj
6lc70tSOVFSErcBImCy8bejdzD0hE8GcVbPX4NCHw+bxqphg5sjM//s4A8wgc0Ij
h69nRJWPY8GvU/82S1QfVj95ocw2HU/ayeqsxuDsyTM/CNK3LcQjDwaXyTMATfO3
RTwucNWBsttiMzA++PuHtIKTSyA6zV1Fob97KA96yCrqZZ5zhz5F9cxVhJ9rAHZ6
DymfxVoti+Emz6nAYMra+qXQRTt0oNmi7fB8z8JMHuDfi44N6VZnqruluGzyKAKU
5Ey0dooeczaPj4TqVe23gG0hAn+MMdEngW5fMeXPvwxotgJYIkH9V0eD2kAhY+Pu
3TaEBS4SAv6U9tIwQpSJtp/5+4nhn5OgOxlgkl+/XXT8aVEEjLmCP7rt0ykCbrTK
reuZaA7lRHX3xSYIVXQof6cLmVuRfQuVoEBxld/Jtv27ma8Onm7xeO8c16lEN1BW
BAfCzqUjLbDb0Z7DLHcP9ToJDWvHbzz0JZXRUALl9GqasG+N1J+Sadtn0XggMXXL
fKsV/HZNnVsifyEobzA1VY5JAhiorcXs2WUmz+A3+pWgUtO6h/3qELyrF2uz/0nG
9YUuBOP0nmtINrsvZnBIDw7JOXEA7HxczjdCUxF12hKeme+XDxVasOdhHeEc3bf9
BgBd18GYD7Fj75KzzTXcYjRu5FV5rclNnwQTA8ByzTPIZ65ceDuh6TdrXeV/k/DZ
ffwr66SNuHqtgo2yft0tbPOTqaFjUrMCqwTqIxgiOKPABw+5I1ZlkiNtYVhulVmI
7XM6LCXCZYrLnDfxK0cNEUeKfjHzxtIk6B6PG+v5WDc=
`protect END_PROTECTED
