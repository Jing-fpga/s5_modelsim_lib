`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2vapkBr4jTGjbz8cy6FxA5d0Wvxb9UTnL4T9ndw6RjaXL/wk9xDmLj7E9lfigTBt
UKEOAu5yb1AqTpu6nyTwt+TywKHTIkJ/yITwcUvPVlutaMtAej5/aGBkQ578gW8b
aawJg5xAXpsiJfB9vsERgIZcFN0NMtHzH6+ffUmB+PTHGyipUC+IRxQF9zBvUev0
XlJ6ghnjA003pROy24lIj04oTAaP4lVLpkis/YRFYc6yu7/WQSZpLFMJWN5ozv2g
vvo/IHbvuvxskTT6Ym14O31EqegZ1W7LfvmG1/rTBxGWaeU9C5JfoX5qBMaIUw1a
/LZgvRPxBuTv3oC8FEQKbY74cwz4Tf37ZsCN17/zzmZGKOtFA+PYp1TIWOzHNgIA
BbyUvPH17Vhw4Td4y71ZsmNOJbvp2V3PflY811RK50kD9tlBAlFkaCi3hgC2YzGf
eBRhA5fEIlFB+CqoOdJd60k/p03rRkG7ODOFXdeThmoFRGfEtRLs3Sz0m8j6owCK
qGOhZikXLFxqN3kY6huBKDNLyQx3k+QtIj5Mn61Wf7S4yEBytY/ZcT8GgSLrqqhI
6m/8xql+KuFEgVHLfCs+qHkEX8XX+Hd7eWuhq7RVMIjDkqqjfgoiZYxi7lYBt3bu
zhATk8KNM3xdeVFNrie+L7hze4RMabYtkYt6AZPpBdKUMtMp4jdKB53cFKbBvGCx
WK1FTu8LbAAAkW8CbpN9/pAVK9oIWxoxTvDW9TyoIoLf/4heaaQGsefwIHjdkpXN
SgU+gt0Kc+SRr2V0YzowsdKPDVCXQN1bQgo+qhUUJbJzjsi+56iokq8dkxbyneSa
CGrZGQLCHrbacGDgMRyqPirJw8JoLnAoYkzDZD0GrdOB9bEoWCb9FErTHB2suLez
xnO+dYPafkf3hquaOhWLhoMrpwqS4Gz0KUjGPD1umOHV+JA4iGRkn/B62nRyyI1W
Z/uxZZX9rqenTgH8SYeF7Hjkt0Qd6i9M5UaQSSY2W746aFwbeEWEch1Udxjv+wq3
nZsjcv4z14XBBH0wLMA5Gg==
`protect END_PROTECTED
