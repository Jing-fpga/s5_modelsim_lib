`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cHLz1XrIJ9mRuhaSIkVInFaiOOrx5ooe9iyrIl7OmIHgeZ098BUkO11kbRasvPI7
GVimtQlQFC8VBaRHK1+65Gy6D9lSt7p6ACOewF7qLgAVj7ixuE7XlIHPVk1BD3ja
pSxjsgJhcS8YigiAIGv4uj+G8r1wGt3JoejcodYjS6D4n18ccCXXO1528s0tRHt6
FuIoLct8c08YthkSP/59oNmdvAP4ZzrWMclo1y28l4hoVQ3ukyVJOZPYJ/TxoUWj
eFwR64bPZQfL2U37PLqSKmbvtJSPetn0HSRkuEbrj7beqjjIDYgTcP6ZeSTfyrpc
+2yeFLahi3tu/tkmZClU2VVie/Yv48VaXr4E7brr0CbOQCY2f8AZrn1wjEy1JQ+I
fYa15aucY04jJr69alsoztNzGwuiFrJGcwNn8mdtlCYUL8ZBxg/h5lhR6FJzL9qy
jd7jRxsV5iqF2uWjsTzth726CLRGgsjisiQSfWUvsyjHg7XwCbqmxy+P2SMs+R9Y
IJf7G6mZWv6Mgg8HscbqMqA3D0+FHLBpIq2md2GXTU8tMec4tgpjM1VmNqLq1X9a
0ryQlnZVMCDYijjIg9L984uh5qng2GcIdJ90Dmj4vU5LACaKVSZLW5wY5mdrJIjM
LN//+AM01gi1sgFsOhgIXVlo4AtauSrZUMByhXz1TZXZsv/Ta3z5ydrDYIjhU4oq
Ah/6EXyvX2zijMoaK4m4CoaXq/Y2MPCsiwWYyg2FtaVuj4I8qYf0R0Uzsar48eoq
LKXzdn+o+Yp5/Xm7gKJVBgt9eY5V1trWcaqcUNMlzME1ZfLdX0uk/lhbkOIYcQWu
saCeu6AfymIrHRMxXemV+gaMnkHmJI+5xL0/x51D2HouPOEX2uOQ8eCjBD7MjEEO
OFmxTZc9WKkqlLEKaJh6iqYYEp0wpIG6OzSprK99fz4CfS63m2kpeQJcBVJgan+I
PKCrH/2Nlqum2yj2U15opIW3p4l8gOMoMiRdq+5YJ/dRfGym9lLGp6YrMBhEs5dV
cbcdIaQmYUATx/Ly6pmRC5bp/nzTezbW9CCB3EkeT47GBBYtOO88aZFA5JEKnkte
esVazwSIo8gjN4Pz2f/4pwZ/mIUuHKdbC56CTBGtTkF1YPTPxXOX6brA2R30lzMe
817WjDv3rTvHwgRnB8ySGuuNUssW41vEdDFbNje964zwNo5lihzCfORHZO6gIn2r
ObSBu+jUEf4A2bMznDBuI+IiLOePdDHzYuxjlfse5l+v237QNDjOkcB/tRkSczNk
i6Qg6kemUK5BGYC/hIRVV6xg66WP5XTfk9DoC59Ummp7Xf6RbzU8Ivu9LXUdnuku
4tdd7+ZZ/1SxCF9L1Ma7QLYrq5w8vkAxZhxHiMDhGFdBB2aqUYFtFBGAioG0X1pR
hNTilWUkmgTfer8NJg7NZxJIhJceC8dZD1IvbwaWLrVIt8Dd3aT2zHGB8Rvgr3db
SRqRed+9309FC2UXbdPtmNBC/Rku7/aWd3wElmav0GTkTkfL6ebsmyLQV3Yh4/RP
twWB5CXBXyBkniLrEzhyjgC1nfm3G+7RRrMYrw9Lf8uyIGff4fvJitiwxdBdMpjK
XrTUKg59NR+wmjo8PqYNkV5FXmN3baTiiXvZGNjFyprXvT8jx5xs7vKvHdHFDRXX
j7A9KE2J7+/Hz7R4+wiPNMGCgxF18/8y4CGftFvUjawvnTjuuCnlFJvZ0RPg4Je4
0PSUP64SHtu2Xa07pLSe+94ndhLCJ5k33QXb+NYUefOnL0+mGbJj7w5D00Yt7t4R
Lmykez4zJ+uPK0zkPwWKrrWgVCCFYiePun4OGvzZtE++DejHOMvMb+WKpxNuaLz5
H2UxbhxSiqQkjG7CoAKI6s2sIuJr7MTEs2hcGVvMucBJdR2h0H6p0JAUKLSecIM1
ng1LA25rC00rOQYb7NqEzSUk8IqEgtgd1oOq6xQJO3px3MRZGdGw69HuPUrGwzWx
hPV2BDOCXs6JJp4903/ge76cxsC7TKZoDo5JBmR2wY3YtrIdsvBbZhcLswoFgpVp
U7IEHy3oNwXgwjYG4sOqwy8SK8qwpe/H8hbORIYfjqdC7Pm5C2Pq56TzFY0dgQHu
MgbISg6ZJEnVVKFpwRWmkSbFk3AOSjnOlZ+nHPPzyUfPEMVa5y7nHTknDA2RuEIc
ngILfAPj4iPMhS2Dj+JARcLcXqrgSjGvcWy8RVrBLoJDA60sIOqtP+vVb9INrEvh
S0uqY4Qx7sk+Vy1K4GjOLdAeBFxiGaZjeci9cec2ZfMk8zXX6jaZ4nMtfxzE13tI
739qtmqIz931o3G06o17egI0iYjI6L2x5RT1e9B5ydlfP/FXVDI6wtaisdXEhgCe
4HgqlHynNPSAADl1DLhVy6BLZvC89n9PcMPfHJDjunMqw017fSWiypth3MfhQvGm
LJdQfcBObLiewHLPnCl8MYjCp7CmbBN+CLjv61MZUdoxvZR3JmTbz11Lu2gIoLI8
VPETUW0FpEQcAgLcLCP6twanImctBHBgeU+vy9QsWgcGdA0dhu6LTQtG7QNaTNKH
DZtV/cxdQ+65/HtydM5x3xc31OwNHtqAd/aXKq9gqLZG2UyB7/wdUqO2UXdM0o75
7v5R2CPg0bBW/Tnxiw4Q/mjWReTJ2c3TsQ5M5OZ1d7ymzbssB/KLgNiLfWqXldC2
NB6QGAUgv0vQq1O6y2JLDvlghQ2EznWt0eYgJjRsxlsSj7Sf3mKE6ys6TxxM6KDA
T1SmPTJe55+DnGhCIscXND5J9W9ueHweBz7cNmJsahN5ySr5MRuIUdNMjHTfEmy1
RABNsHa3yyMqsMqIqiq+en3R+ZSAoLwBAgyqZEq64PLwx79NfNz/CtiQgLiTZ9oE
RJYsuqHUw5d/bL0GmeMrn3gEdspjw+UFBWAHUp/KQaWxQgye2kVGZYqAGpmdYeXQ
afwluYmQ5MD1LjknDag/XY/0SuvE5q/MrVm+agLwI9ywgvqeM/7JMKidWM3sXniC
ele8Oeu4cZrSlMLvfHxEJIHCgOSUtSv5MohY5L3AAkZtY31wCCVrYo2r/8tEs6Bt
d+waTBKZrnx0YS4otZIMTuzzDlfR5t8xp4LbbHlcgV9AGVXQdmq2UTF9wJyszhZo
9MtLVM57XCE1Td2bgJkE1CaqQ346FO343/maf+jE4/joEil+Zks+vS2y5V2E1WMD
hjDTs5PYx6O2FrRyJEP0Yj0KTj3Tdijp49ovyHvNXONsQwtJy0bIzsOukHqLvbFj
19fUIUIsKmNzB6cMd7Cov1WJkTQ+2VVDFkSkG8gH6l6U0zgKMDj8ZB6uL+sDgPMz
O62N/ioGxwQvch+2o+8Z1ogrdj41ulm9cZaq9Gd8DkOjRCeVt5E/bPczNsGcVoP8
7i3UAjh81vyI+X27JtZUqMaGVQrULHhNVTkoCOgZ5c+3xMvPC1J7/epQfpmavjwI
sl9wU8js/UlPq11Pzq5Cyxl7cL+54Q+NhdMYdf+FDgk+0YExO0IztH8FG8GZCBBl
WthdkMlUW4LBKlzZfhwcYajs9Z0YhDjluhLCu+O7xHPiFW5n++GSOfc8roCAB8gy
V/yAPkSvriN09/rOUlJcU4IfisXoMfrmWg4YXmQSI9kiEUbk2p9tvSvGcF72WR4w
DdIaSl/LqpVG5LHU/dOiASE1OPcccn13QPl1xPFATISLsp6dYIcuXphNpCbGbkgQ
Z/LSjn8QT9FXsLhgoczx5GBORzwgMqSetLRd9wow/0bxS+fQMVg2WR4edrOcvXtI
cGXrUhQ3DnkjqL5zY9YYjpPM92lX0BoYGWN9qBA1N+0mgWVE+QZyOcssK7sy6h8N
E5gavg0DPOMzZx4X/LMb/HyAbOqeEon1+l0bVPycMdDaL9mwJpcrSyPCYuElrLQg
uzAiJrs778Tc4Dmznkjz/TpHgtJ7ZL9cAnoKvKVpt1L2MivC0fnhFLpsA8CFmOP0
yjNZKoSX+THpmmIyLn72wnVXyJqV7fgRf0Kt6Z7Op8RNg1b5vXCtJw8n4xzV2kF5
k/9Zwnt0Wr0F0cHYXGYQ3DUUMPE3eXm0ECkZK1iD7tvCmjLGN/O6qQLZmJeE3DGx
alypPtIhJ2YCBhvxuv8ayw3fqhyJ1UaJjuxh8/kvd+ItlfIHFuygVVW2DiuRJZ2C
Z8rfVqgL0JTABN573bBEu6xNYcdT0ARk9zZIKqKWPke+KF1c8ycIneTNWPZ3fEOC
lgHz3SsNvNUW5EVicG5rWqFIo1qCwJK8LzIlCzTV0h0POkT/7C8NileiKgebojjF
yjsEYTczzBg1hNgorxS8Xh/grvlgE9CB/1kCO2zHg7CAltrv1bxca6h7dwSwArZR
73tMtDz3OvQXgJxDQAoPstNgiylNd59L0PD5PYUSXcIlxG+NJWZM1PSAseSWVjef
KIqTFEL6ZK24F+Sg1nkr8osz5PsGz/LwGVLbGQBhBan4ZUC3Y1qNEvXbLlDOhU3M
a0PPZoY31vtw68Es88x8iKwkoByu5lCqi8LdbaHp1UUcLbyXy2QaV8AcSBRx/ofJ
f+ldB5NQFozKg4jCWOdNncQwGUYs3ZXzqreFAcNDDqLhalwVm+sNDBqft0DJh0YU
8gEAUpBb4qjg4zLrsOSG1QoSEp+oT9PRIe2fYWcnG15VU16PF+S//9xmyf1VvaE5
Lk6CnutZG3hkxL6/17wrKd3Y8avS7WnkeU9hZK2vJ8up1xrbtHZspPpG/MVJlvVL
ixlUjbnCAum8Kvrno4Q3osSdouwDhGFb9py8hqDWtZXg3e2ZJTMPwkaD+D7H0b4Z
0Fh6JxW1y6/kKARn36ooLoAHkwYDY7NUopWphfHWQ9H/8EFrwygeb9pgmF+UqHWL
yz+/bLp2OhZMDWarzwpGzj9hRk10/mJ3WH7R1K4QSJMWtpUqvpDudse8zxP+z1ch
hne6xMPBHlp1Ht+hZGUGzGdNrudugrPPg4YhPa05vZ56ocBrcPs+fWfW0X0xJY5j
TqQxmpToIrilr+M5na4PT/+bxLEU7BWf0F3UbZpw2JRKz/K3O+Ycif+EzkvGPEJl
l4kwEUt+hNKZAG3UfmWi4nZuy0ES7YwwFyeeQ5zFZlPTjOJic6vQIr+AyAx6HqVY
txfZ7c7ouo76MrnHYhZeyviZJxn4sCxNgaXh5Zw9lfAyc7rSGx+IgJ+wlNeYg/cB
MfZiyr39k2arnWyGtpa0OVzCzocNej41EakvhfOG0ARgFd5M8y7Rfv3MnuMOhkiG
CjeNC3vzGRFHm8xtpF5TBrJTva1GP9K/DnNBvY09d1LJlDuELDvA5R1SR4cbK5FJ
dQlGw2BIHUxmKdHjOECZko7e0i8inCcjyu4J3N1WX1JfULvKLnnog9uhdO2W8/zl
yW8GoCONnXIrsbzpUwaJVzntaBp0ko2nrt2okeReXFcLR0wsT2DLm6Ogc3YWb59u
eliZuURnwr4NH7TVZ00nPNMw1v1BH85hLM+I314G2ZPd/cF3V8aqDIUZWjy39v56
q6lurQ9ai4XoUvDAawv+8pOrI+kvueKT9K097Rneibr74EDOJfMDG+ln6RqDvYSj
vTXuR7yKrUOjnvZNF7AJuiOYzc2WjKtrV267S845WrMcX9HVme+UV2PoJNGKQAGq
P7sHwYt/AcFsGQvqUFEnOwtFHBrSih8P9jevaSmZxPMReUr9cI/9lk1sC04Qs+K+
agxzvCEVp8wq6bejui7zarQ03WMH68ddkT7qbwDgHRepPqt2waQ6P42xU6Kzzn1w
gEVC8vYLk3wD1s6ae3H8RQ/G9KS4WG590EkZbj03Kl+pRLGAwA10MjZUB0rWQuYX
Wim9OZzC6bw/0bnuSUqSZDAyEi9xzkfV/Q7wj56W4i1rMVFIcKMNXjwAwDHrJqUS
vg1917219NtEVYnJUyqKuQqSnde05hNnuvNWKrXDai/0yXPsvmz1HJyBymxuV7gR
NtCxDKK5LDB7pBJ7kicT50+4LtEM+jEKkBz5TawzsvmkqDJU3LGQX4M+cj1T84TV
hFQldEaoImK4mJkuMCetQm4goq7IOjzeB8sTae+BNW61pgoBpMPYyPoYq8R4l/kT
6bCqtJMmzcqlx94TbwTRlS1C6qlRjeH0h5l2rVnjYiKqgtpifrdb/e5x+7C4LaKE
ZXOqx54AGyHTyxokoNFuFDW12pseDCxt2NFqm/VFFMXYAjnaMxENTw0J+6p1NXd0
CyssavDQWSCjHZy04QNyhou7v13CvdI/muDRsrOTAWK2GtQVART6za7jcJN+v5Me
ZWcW6eKKBvT7YGVsNnl4FM5IkigHNgFjQn3Y+gozK8xbT80WhpWU76/Gz1pqkc5N
4IsuKlekEAsYFCWGYi2Um7qALY6aVTxRVDQpK249bKVIOFzjCPZtrIH74/liuwtd
ES6S+H6bXquV66oTlqmpVrqA+6ycqdk2WldbuvqYlFQyp6H/vT4XLdCQwWdySKeq
VHJbRf2pPp3jBfQti/jMlkWJRWozmMnrZRhzVilnHEizODL3uSGEQ+pM7NqzogIM
IwS4/L5YctU+eWYfmYuXiJh+COLrjuQeVNCyR65O1L2404F1/cQRysfaA3PQR7t4
CQ6jmCeS6heX7v/EvlfF2H3KswZH4BoWYaK9LT/PFm3EFdTqmpWpVqWbOHEzF3Lp
+gDYM7w9px5HWIyiP9q4Kjqkg8kjHfcZdk8B0QoFCPhroRnZyGEjACeU2vOamBWQ
C81K4SyB2dgOiNLuDbUA6MDuzI+3GxrmU+iQc6pmggas72p1+RCMryTdfmvnjQNt
29F9YRw8jW8pkIidW/hfM3W0h1gEPtwTMkenQSsLRlov/q0gCKjm4kzUnTKqtV6L
QbrEtrCvtijA6Vc/EEDayjuGpxFPRlx7P8F241zuZtLPh3xMN9yDS4kUPJPpf0zy
VdHWWed5wHqHEua+C41aAM0V/tS3v3v4KHZ7FhdB4MgsoYm/HydSwnWea303JiP3
4HTxtss/Y9YeqiguS+UKqkGPlSE1l/L/z/s5Bb6h1Pjq28N0QeN1/Tsxvi6MKT0t
GxcYSTEytJIE4BEvPKIu86f9Q47Xy+9zB74xhwGkcQV4bOaQRH05SmX2w2NoWcUH
yg8/NpYM5OhEKA4Guh7tRRbid+7rKKUGeNgyFp24GilYzNzTVPsXHZxA0kOAsVUe
uSuwvye3fcINwQhy7NReCplWNUTVCmul7gxytBayt+PK1Ja65Jdq2c3gSGal1MT6
uLJwPy5MIOin46ujmdg5JWZReWvsjJoCC/XWVRvgWRpKgM88HmfjdK98uSUDVxd3
PrmfaM3u+iOgfPNwZzMPB234wd5nLi7X4rWPzOo1ZCH0h8Qqfwem84yKaB9kwsrV
CiL5Ko3r+sOX+RSmEdR8ya+iaQdeQkF2ZF/O9gi/nT8vdjwDEDWfuuEtXHi/xxHW
vDBU4bwAvZ0lrbwdsCTmRrfZfSKUyHQiC2XrtCf+kxjYPN/N4T4xq7I4f2aKTF+L
qRAyJVu4PkiuCc97oHgbiZ5RqwZt19FBCOQrEq2W6EoKSLW3cR6u5yBUKOSSclMT
N2NUqf3V6Q78FGqxtFNZRF7b+g9nHN3CaETlPkFC0F0bKSfSDywNCpK1L9aPOfn9
C5u0bAwYZeBij9zzhfqc9g7DI5t/OARYl3EpTApcE5G/fS594fZ4CooXLNSb28i/
o+SGuhRwlTK5nIonvVVKtEOepeuWcVwl/v69lZ7VsEOZdv4+czysNNQEJy72a9bW
pVarJ0p77gImD7SeCL6DWwyeuZj+iieFoDE9w6PPBC7UlRpNryFhFAAc9cz0Lqic
+fuGFJ+Fz0tRfiKAnTgVFRI5vK1zPa7pW7VNtw4kPy9vtvyL8hYWxoqtq8BnBd3X
neZqe42VtjrwZbtv4cTptpzlkyn7DHjnvpxg2fZ0pAp1iLkKmn8g//fDcSiwbUz2
RxN4KaqZ631kcPes2DFUMK6m27Vg1X6XERTSVYb57q2E7MpLIDcUprMmVYiXbcy2
ZPzs5bGV/oDg3Yuc+71vtdBbXNAuw/V3N7YdkK/Pn3G9S5ThtaCsEJuthr9G85wE
ZzQbDeSHQoOT62DVMfUsZPRaG0RfaTRyN1CXIXvE8PScCSFcQqLVHSlWPRYEHS7Z
jOz68P4aTgRug/Fm1vcPC5UEiXVhb2FVt8e/GnQ/PJgQ7m4YWRN4Cep372xcXM5J
3XJseepcKsT35+f04tM+ew/82voqPKJx6MyJ3yIyLEW/GUVBJ4BxXOeEjzWViMwY
RWXN+6OOHn6wKEa1y5KUWc5eZQftz8A4S+zskNNZsvqM5QUNfvFttzvIUGdMaMUG
9DduFItzNk/20pngmGi+Fu+WIKW0H/K4Km1EtdB7ZmWh2U6EGHqNZwSITT8YVGgW
AUnwHcsPqNgHA9L1wF5nVCUBNLW+/x51UQ/F9G8fJBFmy65S4fmwo+7Rse/2vM9l
5l0oF5GndVHyynss10L0tGxstVG+sUQ9+374gPgbyGTpbvPN+vkK+2eWQlwNYVfr
c1fDhzWD5UEbCte1YPQtfe3Tmi5BMzV//Bj0qpYGAl/kjpKabZxr/juKOXlctYT8
iOcM6EhOYrV9yYGI4wq23YZESrwJqjdm5j46zW5jRVSkoslNb2b1YfE5Iz5vrAwb
RP77ARl8WqgySbj4b/w1G5bC/Ydxm0bS6Rl+jHcMDVs4+JqPmsL68S0Osp5e9E7/
srMMPSab42jvbak1fbvnLITQ6gj+PZgOwPH6mRdN6/FHR0pcVT3VmNb6XDBynk8q
hDcMiUICbjxv4pKL5BXlNnE4bqVUkpEK3ir9t5WFxSCGxbFx0Q95pejwLa6hCdC6
G1rVKTnuUfluKT0y7r5qEs6c26Yo8VZRm8kErtOnPWofNOqtshOTaFcXKjibXQGl
3PGHgGYHqE4MkGlNPmTfFrKEoejuc2TSH+YiZyf1P2l64LYKwSlT5I1Cr2zi2Udc
AOGogsk5wpow+HXX6/Iy29KkJbsKoibAUhvnKm6FsSpfzRRpM/MErZh8cvMZygP6
Cwx/Su2Kb9Yv0LR4iMja/bInBYGUYfxDUjMDGEeI0aGjLt/nfx/y4ifvAHg9z64q
VvdmhHq20XS8rM0q3X9wvCDVCW8jSyO4N58bmTaA1sCEE0tysjKJGoD6Cf+JyyGx
Y7LltYUCBnTGfz0KrBLYjR/JlrHL6afF4donIEaUi0FumYGkrTJKgeX9dH7FZl9q
gOJ3DEvr4BlxRst4wmRpZ09luPkn9ZtNz8u6nOuYThHUcCvjCMjaxqvQUhHkCWpf
HfMBd/+K0iaXQ1akBeEYvD7MCWQCxJJiD2QLUbul0oDseuoh65EcnE9auIny6rQ2
RAZYZcxNGGmxX57mnNuyOWRSDIZOad32g/lwILxsBoUoY6AWMLOLaZh3HGcio/tP
M2OJI+oqWYLKcUCMNUBW6PxJ5HOtHuzO4e3dmf0J0N/xk2nu5s5mKYRRZbJGIOYk
Pa0SWRJO238g9rj46Yr5XDaZIuWPscR4GOYTeMTdJSeHwzF7rS5lQ0tUevpkP84r
PdueMvOeGuF1w3iVwrMm7rSvV5cczl4MtpU8brNDAIRdl1Ql18Ab3E2kZw/vfjV+
lJfxKFE0xnmtSdubq3mAdAmzm3skefD5vDAjW+vUjwFpWvaDlr0tkSupXR6aeAcr
BrooDTkVYWvSkQ+J+KRn2eGJF4XkjecCUPyrK9PPeKrps5A4AcSxlHb/68n0wf2u
6rFpKsOm4rfS6wyBe93aAFkrWop3+z/5YKVk0/o3JyY72MfHjyo7pGKhkPXomUSc
wdmZi4r22BLivw1VhGWPvj0hWLHTtAN9buliZu9y5wcnnBN6WldqyzfTiVOI4KIX
dcZx8en885SScZg90s9rM+j/cqFE0xy4ZjPfsEMXO3G+ubTwnXq0bL3o+BqHxrkb
EYOzJf+G8n+oGKu/5LvTMvXWkVf1EQVMOJnfg7gwA9xDz9ybkPbf0qv4PRumaJEo
4BK3EQ22VKSJXrVNcR6zdk44y3mbmq315iEEMynuOVcUuDiMjK8Sbo6LJ2vfxbOL
CTHnK2S12CDeuQLxPV9JzjRDbtxcdo0Xu/FeGw0VQ3/h/kAFRKCamWppaKMJP64U
MMVg2CF/ITA5LmK9eyXT7Afkp26fxFr3IkIJSUTcvUHQ15LvGfkNqC0EE9viNub9
hn4DgtpxvtNGUaxTqYXS4Bszq7xQBuHAey9pSgZLc81B4ezOOLL3TXY3AW67pm6T
8zBd0lK9b2chz5nRY7mNWbX51HqoA1AovO0bfNCYUQbr7v6WbXUTHCB6UJA/4SXl
tWYfIRrloPtYOmGxayi/mMWDlJ+Za+4cFb31xU3xkLqdEDNnTpNvAaG6bxtaCv4y
Axy3hc20fviBJTGbYLMnm8bFW+95QfeEJr3kGIo0o9ta3J2NP+/gWvTZgtanKdaP
TtqCZIvZmVUOmcEqZGqLBEl94MIqpTn93+txC9GDvMRJq2n8hB/ZyIfYinu5OvL/
Ay8Z7kXejLLHYHjSR0Bkj5qPTjHgN+uqlBv1dpyt+KCwtfFw5vOz26KIvfGoJmoP
RFkdmPLnSbZwJSJ0ZvjoNEXg6cxQYb+A5fFhHSQ9vDvCdOtya5ShDGzvojG3X0d5
v1E0nR8E8RICuEmNu0efNazL+7v0laftZhq05JMfUCIDcJELBt9Qbdv4fLf3rzkz
kM2+hh/jsEyQAMTZNaY7qOQ7G3v6yv0LV12gkkMyH/2OuWmWN7H7WqDSWFOAJaxy
la5Hn5Rf75UghW/Pnp8HzTwkHYZkss7mzme5VCDMSWbwXeK1N7ZpFHAL+lygCBsx
et/Wu1mvw+u0gJ+a0AEpuZ0QOc6L9KlQ1u47UW0fz6N8dC8iQ5I3TUttw1d0HVYD
5u7K5CP+lksRmcHWWypOAJftWNbX8/xUpk/O5zN/6I42q0+Jzbb9gBVTJqXyBM5Z
/S0Zwstle6FHgTarlktdL8jv+ptkSd5ye5KUYZAruQLb7A6iEVkEyL+FdYkyQZYJ
8rNYbFCbphQINmQ1+HZhuBn6aJj4JTU2pZ3ssft8y0OCaXM52YIzY1bmd7dA5VOv
etNj4p6Ecuy2xiGnTFQwl85Yw0MAhhiJ6XnO7jsUOYuAnYgtMGlBTGaotTyHTJcs
MnSMCR5Qdh3/9a1yBzkPr1FHyeB1M8A0PwsVw+EIIKkJkHfiP3RpHbrPNDcOhoRc
E0DK8v+L/sWgE8okDRoZ6H9+lh5lAISqgwaFBvpQ7/mrW2SN/2GItj8l23IqpmT2
FNXINRPOLDUErgP3ufscmTG4Iq7MClLgf14/alQ44vCuy/g/JUwiuczhkFS6sREA
NrDUF1OrdNx0RbGjvfzuxZs/eVX1+P8lX/CyCf7C+yCEafANwzF4F9biMwQNlQZo
I3zIPWsdVyCSGPD+FMWjS3jWcJIL3HaJYA5rynZc4Cb+8U9ngPJq+40WrHiD2Hhj
8IpUsCtd1zTQFd0hTZD/5jDnUpKl6y37m+tcj3kxMT3Bs0LBdtMOU5u89MzpzZjq
5IlgPIeTvypccAmkqex4Tzao1aW7D57Kh+SRq//CqLmm+M5Xz4fzzfTCAMv0sfvv
ekfeF69gKvp/BXcAtf26Rs9ODilxOipi5pk4NRvAyz8Sw/5eNm7NtsQ7B6Lg7blf
sNXsu41EnXfg47w2GXFISSSeSrglEl7s6mwNOrm+mar7Lg+dA8AEiljJiqjNXbET
QSbynzYbmW0wbwezRh4pyhF2HksxJDeK7nDz2/AdnYoUZWrAjx/QomZlGBIFexHg
lQs8j0GBqP5tgYNchFTMNxUg9F7zggG8d1lvIEg/xkqJOB8WokC4MSBRBNm7BxLd
qvIO+tVXb3MoQ0Rlg7qQvLw6JnUOV3GCOlkids8kOvsPlugZTNcjYIMNFnwko0oR
dbhtl1o5mmKjbBEwkmdPqAnG8DPrJjNoE1fNsDGnObpCwCApGThNv8Teo3u2yK7g
Jo54ryjZ5H7FbgaxhGm3RRC2kcYQMtzlAqtUrCVvGffZ3mhB/N2if9lZFTOs70V4
Do0zWGB86PyOnyvJfb6HXivV2mfP/lR6kJfvx3HO0tTtnmu4lHfgEljNmL8vBwnX
rYBMccU9W4wQit8UUaf0t7s2bW07f/WNtX2OLPGje4seQMmX0hf5yScGjkrxMuMF
oFX/6VMNKqABRXWlerUh6AT2IDNWcmMjOhBDB4yIBrQfTOy73euW8xQLuHGZtR12
n1oemmMJLgxb9jAJ74F0bUaR+cvO+4UOyEc0ZwUoZqw3qXC104m2LA0I8TICBGRw
f/FE5TUdvof8Bm7nVwe13KQ2yqc3Ji+NLBk3vsP7MDsf5Zjzvj4xk50hyJFp9BkH
2l5vLqRBDjcrujGqxM9yq07vP3aL0FMxMRH8V4Ble726FhW84aE2JtVyPn7RNEtx
99R3LsBVgEuS1oYrTbBpHuw6oR4u8929xAEbU1mFYlil7I8XNH6UId7ZP3nChlq+
Kh0dYxgXt+qwyEkZbRNoH2BXk7W3FWFsFjxw+fAoZZdz/5Xl/HBlAXuUc0fsV+MW
ohKRbttYfVm0yzvQYEzj7A5q7LWXVcR5mH6qcpU6VfOIpJTmbyqdYI5P0tYm41bo
DoL9zLpBXR5pwu8smJQ1HpC5sFQB884yf1qeuIKpOSuVtl+4BpmVTrfTFzc5b/QF
6Fp9+ZiDFqABDmUXdRbfHagaVlE6gqPw8qSA5+FFyfdyF84Bhwx60EFJ8PLRt7yO
Hzd+pdx1TUUrqk6GVHMGjGwduwRwtZKEGbg3TxB76NIRz16c/dLTgMqoLZN8wweB
`protect END_PROTECTED
