`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lU/omgPch2wEjt+61OOwOXCawRuDLsxTNSHpU2oe0Hv2eRkF8nCINHmQN+RTnIw+
Vzrgib594dznGdSa4yeAr4CdcOmO/Jb9XOvInzSbo3cGqaOUjPdKkcgOev1ipgr5
Wf1o3b9i91ufyNskajfkoP5EIX8U+YPKxtp9BlQKSHGm/jUcYtE8A1uwQJLL7gOa
imG4W3Lk0LLGanxy39gJujELPAXpFbY/2MzTGY6A7kpT8CLncVRUy7i8FaZue9H+
94cvT20eMbDjBAfr5KVLVZTsm+tH0qol8cWkGQj1BNInk31OpTWUGSBDmvvenndP
biIcWRa4awbHBmowv3Lauexm7o1LIbmT0I92W9flCf3rh8HvS8Sh6LpQbfSuCB6z
IZsZdTvF28si7o2JAQZSux33SCXvd0pRmLwP1nyGJRDIvck3hYQ9faVtv/03/sgM
AaOBMV0Aw5uRHBzm1Cqu4WkGExJIHnSMiGYrWze7IioP5totmzP85lmv7pjJrKMd
Vo8eRVtPadOfpkEs78AWKcZ2OAcUvAlRC/XomD0+c47Myn69ahzGGe/11oA+vQGu
oloXxLWygQtYeOK1bbBVAAQl4O6X2kwTEbVuxJgRZ46BnjlqfuCXoDMVU8QsVrnv
40TB8BjzUf6jQFiGPfq6w0ChtCJiYvCivs18MW3TM75isly1YtEr1cdAdcBG0dRU
jK+ir4ii9iHZ6qWfIXoGhzHocDRhj47GoqHZnb6w56wUJZyM3JXse9Tz+QFLPaL7
v+DjixzW3a8FyROv7iXtrAOMbMo6y+G4/V9gmPMVYhP5P+nsLL5wD4tXNxsS/Oy2
mWsQCy3uDwghaIIXBO9JypcZ19gvZ4IYhmoqwesR/bg4S5ZTMwGXIaplwCww9vZZ
8AvBXatgumStU0tovIjGZr3f5iP+o+xXcs29voPTViaW/+FdC/PJKMRxuW/XfIWz
pgFI/GCcYpXvRLZOzHXpiN3xh3ZZXXME5R3Hw9nkIX2nZ/0aJ2cPo3a7lJvnYOj9
J4Kma/qgDVatyw5zqdnFgf1GeyzngK/7TSc0BTTHUp5u5tdMI2+lbouqCJ1SECCg
U5hfQ3Wa1HB7q3j97e3cz+Z/0EtxYvbjUix0uewxoMsQhAY8b0wRQ6vuuOOYr6bw
3dtvick3SLGlQLlti8Ib+4l43SB8ve3/dS2I/VQVDzYunGRHxlbgwOrKR8X85irl
H/4vEJwemsDwHxozeYDBPZaIT4PRCmJRaQkJ/vxLZXNpmL6/Pbbb7KN6+KNkvOcA
vpBiAvImGng1PqRPys5umuSx31dGN1wMgwD1ciZhFAbVEq9tWnHhfzBmS2fFlU83
VL2SLnQDB9cI7MYY7B2J6PVRELFOOgpxzDmYqo/h/VuiGdyEI2Vo+enBWCoP4PIQ
AlX891f2F0PuroS3hU8q2SC1TWgA3WWE7Zxt4qF6M2c6t/wwY/JwzCOMuGTwTz0s
WLMZVClDt8eWRPWf8fgz447v9hZHIIGfnKHTBq+kDN/tJoKVY7SR5UQNfC/nYfKV
B+ji4GGUDrDOpnvLPbInyV+oaMoLljj1j6v+Ii4c/fxi2Hs//1EmxvuEnD72VOzK
uHplHjb7O50UGrWZVJcFBT1tl3jOFvSF2YiOBRpfwMyLmRSzIcICynFQMPfL2E9X
xbUVnOV2hSGLEiWo2KbgLSAM+LSAXH086ScPfEE/E9Vai3lHCZomTG6MyYabT2gG
Bn0L8r/aiHvy1qnqLZTU307UKxhIbrwtdpWavZfYuyY=
`protect END_PROTECTED
