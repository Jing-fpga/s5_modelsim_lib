`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qko2G6KnrnbtpPTfEGsL7VWXMFF4K+6C8ULvTpfo0vfOYrZqSlfKl6hjdHhGfUdR
9Nx3Dr0oWtttsX0lyu7uqaNk+n2Yxg6qdegez+Yw/qCec5lNVGhNl3dXmOtIGhqx
tDQe0sKGLXN38L9J1a/pWdwIaJsOzMFmvPnbUnnQ/znR9NQJxFtHGGzjnONKbyKe
rVbDAB5n6tt+Ivzk7QLfEyemD+fnzE/a7ZgxMsW7Zb/fOk4PqPb7iUv28BSeqOyg
s8/98Gl74KwdoO9z5HyJ0WFOybX9j9xyKSC5EncSRZVlEuvaU21ZzBBvX55u2NSL
+thPfHyA1jTh7yttz3sQacq3SNL0R3sO+k04v5ofICsd464zxNpd1O20Q0f2DctU
NHtv5haFOBHp643hYV0QXVDJQR9cdUSRA0L2Bo28qqeb4N1BsyQG0ayzy49IzcQC
TxDwqK1UuBMBzMSI1/UCx+9Ate21u8Arc3pqJfUvscEvq+JJyoF/egpQzSbQR9gg
6yjNFNz7rQsnKvRnSLeJ1rW4FQbUqWXVSlNaTrzvUOQvyBicQNmMAcl0/axtB/MB
Whk/sr6WcDBjOIj1vSdG7YQ3RO6WQNcD6teWobSUFACP+jq08fmQIt2HFMr9pA9w
z/HbzKKubQjZYS81sjAUHv6VSapVmr7iZZcwCBC0dNYe5fzIf3uw7vkjdT3QNnKp
aliiJZj/nieupnRpXOYVRmD6Q9wwxTR/Z5NXyJxTwU3t6HIUAEOKysL8BlbrfoR6
DJh3fKgd6vEGWWItpCG4b9qZxwSLJWK8J7gEpaBDmGGn1T/EUhIaYfyLiifW2rwP
GLUX+G6mVRhqlaEsOSviSD9m4Nhd6wMHGGwwy+TpvnukKztObnI6x6qYaTj0dwJm
xVWvyhSkdXoiYh6qOj4t7g1mhsA5ylWyt7PEOebVNQmzprv36GwTCH8bIGjCR0Js
fdh/usppgH0uxTVBGUk3cd1UrRHqnh1n+rls2JUsbIHtnUtfi3tJRp5GFPU+N/GV
Yq0mprdeRcXWfjG41y2dMmXTb9pwwkxG69+Q7YZk9qkZwnd//8Qj+Iykb/N59mpL
omc9Gsl/j8y4uYP43SCilv+2y2XVAwBC2QQf5pACnyt4i6gBpwozHMuV6dYfcIq9
EBhhfuxgfaEj99Bw0TxaiD3Ocv/m6GO5wMF1/8xM1F0uyUkmeVFUtAEjCj2ux4AL
S8ONXIQ3oQzlSrERF8xc5vABQuncTYppmCz/++F+78wvJybbi2asFkoqhaQMuMnd
gYXVc9mORz43W83nPc0b0CdCGfJIjyGkyZiNZLDO5fZQaD87slNC5Q0zuOoDecVd
74tTT4RkK5Vw+yDPjzh1GsUpJKqc5sB3SsQu7Ik8D5uXDL17crXkvPFjZ2FqHyl7
cMTSQdOg3fHnUTGEy2GoUq6EwHwAoKRhW428MjT6APXG/hJiZ54a9ZWhikS6gNTy
EpVt5NOhavHMCArImpljcUIJe7mY8fSOZ9Kgl8VqkVNCKsUr0p+o73k5sU7NiFyQ
MyGuDklksd+fAMPtA8BVEnDM+kwD9A+KywxbJuigz9/RAa8GBSfWNzA9CVXl8tz+
J82PnZ+gLkwJX5/QZEvIz6mYaRpQaEa6vF9J5hms7Gv+7qIruCz4h5V5u+B+HJkY
SAhHt/wxQfFd+LnTwMpU6P+u3Dlw+moKsrJmblaz2YxFfEq5WMieufdnbijpyfTh
V7TPTEz5bmVVCIwc47UlYL5ZZzZIx9g7pOhSQkh0AMYEVIydQJqGxialcBOxRhh2
806eyEhv+pSqr7W387hLqLMVU3JqKgo6G7Y40oUaYy/ywiMgM/FK0Q/B9RRmNwny
tKpseDHvvDNaKDQp6itXOCBQ9r/lbqiowCtAa/fAJaoU8pPqNYP00ozkqU1Mave2
VOuZD7/Yw1Z6Z31GFvOWZOGFxmjun/gVBn/UIiz1uQ77lRugwwMfbswI5bx/3U4q
NmCuZMMAbQxfVkGtgJJy319ZbK/fkZy5ztpUpe+7RKwnwewBLJQ896dqODr4UMN1
vooEJ9oVrR/xdspQBqGfQ9MGHHZwvVm2sAw3hGO493nlzr/dzVwPgEufUMl4l/cS
f0cg8KH0tC0gUrIwx9Qj6jw03eBNMIn/g1hsPvwjW9s=
`protect END_PROTECTED
