`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d2zoX/c8EjWymDzD8RlFzOLYpXZfckuOQNDc7yx8HxQeQTklO31gS1SxhuSdOUa6
4P1wX1+vsd3EaLXBFD2TCE+c8e5qQShXiMrjmyYZM9ErJzGN2FMfhinhj5/5WgbH
6g6nk5a+uFb8g8CnWrlO1nfiPxh9+F2Lrzkj5T1GSKiYvMGSLM9OrvDvZqSRN9cT
6Flq/bBu2oNilfaiA00sDAmiXi/V+L8A79iId0BldEIW8mKWVSI3PDAmu0lGbU3v
OsuybOTigAu/7QENRI+5sBWPC5+1vmwvuG4bz/X48cpCvxpLc1hzf6U2FZZNzKHe
SFXxXE2umr8FRG4iSyhVR9/lC4x3/CsDnFyNh0NG4pBKFatKWcKvHX1+tmeoz6Lg
w/dMJnaGn9vhyEnAZiUi1R7284hy65pHK9qEwVNfTW6wKPeZsAGxZz6+jNKGpdpa
8l3Hvav2Z3PLCbjMiaiwTxhCmbEOW05D2jMvb4ubt1PEaX/z5aFjFmXzCMJ6wXt3
IOG0OMdBv6deFrec0YfnKpXrrpO5L1DCgjMcNqpfjcckGH7DhUazFt+UL4fVGzxU
rGTbMlxvq+3Qw2jrlQxHxnRJuKeMfUVAAJqkxG1LFUj3aaymZybEz4m1reRXKXE6
vCKbY8vr/dbg+1TIingRU5HIDUL8MtllQJ29CD5PIrp/kjPQYe/7rwWkdaUVVMVe
81Jz7qjMN04WObh4i1Cp4FbrseLAOiHA8mqZ+l+xS8X391T7uBfoSP6HvR1mfi3y
u7aKU9YLnnniMZYhtV45o2tO38R9H8+CRG+px6Izd6vCZPwsUsauGXxuK+9SsJiW
bJpcxPlgiq1Q9MM5bloyqxAF6MfGo+PEdcSJFdI6mX4781RsoJ5WUBWFQWv3ilkC
fEKxkZaYyDNOGtAf5OGWhi0VdmqSbTlJMbkIbBwlgtW8w4r2be7J+5gBzND0VNu+
5pjnMitI3hqrBXpTUYJUOrrLgZ1inKYZP4PbGxK9irFcunE/3qp1Wk9P3Eo6Rfuy
N+EOGsAfLQGtgSmCWZ85/jaqXlBlarpOP3ROCL4LaP7ZE7tqR+pkeKEPJ2GJU0sl
sGu6MRkVg55SQL5aG4ApXntTbyh39bnDkQal+FIm4S85zIei50eliabl5rk4CTW7
zv4iTCU7Rnk9qjjD4uEUsbLNTAgy1MbDleh76mw+8CDzlWTMSDms8dHIlVcXybYn
s+tH8opnJa19FwE3iH0kYEACx7dWgpVx6SYcUWwuYYviT7t4UfiGQZ0/1r0optJa
IB9pKsYshBw2ZcxC7G9GEpfXrVj4Y51M1V63SEw7xgkfAjC8TQU5Tj/PTsbiiW/W
OOgD0G+UIgM1HYHJINiz6dp4e/mj6heiBihwhsym6Kl+jW0gIFjmutZsY+rSWvtq
GexLJxYJCyLa19cJP1yl1e+mRumHo/uMuFuUIxfeNztJMdjiKVgmSBO9YVv6WgOi
GM0m8IPoSh/zbcLD/F7k+6pat8x74Oip+ifsJOgRWXXp5nC0AIKPMGmShjxUR8lg
5ZIHdoXjx83WfwF8RmBlDEKAW9zHNcRd7X7gO3GwUKZAz5X+7PDDWVZsnLaSbj9w
8y+93pvTDzMYkWimCqOn8RHH+SceXfcwE2tb5eIUcJEC741SwZP7FRreOPbPiHtJ
CT8aJ0jTq0ol7ZP0Kpk1V/XRwns6RPZQiU+LIxuk+yZdS7au3CDyVPjp7j2o3nnd
PGrueGXfuiKOm/CampcsEN1t3qa8Wae/DfkJTYevWhZ+GC0mh6Zfaqm7MywMhzLH
ijt9QaFGErGQWbo4a6Kz2JHHknJwPZPIzXTxge0NP92yQuxFO1JtxmjvE5vCaCy1
+TOxrmxlUCYNBKtCixDeqXcqQ5M3VP/6iTQ37Z6lxJ6oWZFcjNfjVGZK6k+f3Sak
fkTgJayrzgpThvVBoy2412yziT18IfiFcZ9hX4fmkKabIGA272bWVjqBDh+Q9q0N
hlBDVTUnGVwhTXSrujpdI+/Oji93Xg8p1nEzwRAk1U9ThXbSpM61g659cXYsxacr
vnGosEh5az+qaomRyvuWs7xaFC5hNk62MKtx+Q5P9Mv1/XydggnVBgh4DorbAj5x
kl+G4XqqjMDJRVlaiSfd0rYCvfm97/4E+znyVQRP7ObG5R1RQlFKLtAs9wgydBRn
+XBaJisK9TjQyUQi91qJDxpcH/Z/ps3+bbiEoigw0siMKYxDXw2XV+ZWL7xyRTgN
YhmhF5YQbgrkkVnT58G/sJQ7C0pPr/KgBhnS36WhseNs1iQj61D31WJ8iowtogyq
Ob2hqg/KP2/NCG/BmUkGoKby/OK3633xcl4K72vSlxpWMH3Yls5iFVM86/hAkgyw
aN8e7s4M36g66vVnpNodblBPJ4/swEpiY0t4K77WL3y6hbbez5EGfb47dbywl+or
Av/ORxBU5DahgZ3ziHgF1w/Zv+t2vb3bAiJ6k2FW/WbYJVyVu0Fuh4pcH5/Am/eC
Ha+jW4MugDBp2duJl7McFXBfnKtkjYbFgEJwY9azThbuI2YbYY5zv+MXkAr58S8T
aGXT8AzsUXzG8C3IYELEJo8QpDCHpMQGoX3H975zmqZ/4StmNNIH/KqowNNcXlvQ
MPE0/S5NrJk6wEp3fkNMraiAICwmqfIj62+Av3CA6jNXSjw7JtMNKXjKrCgKXpDn
D3kk3DTnaqFIv0TpeUNqhq6E5gpCnRi5oK2XjGNGSmtymStdC5hy6NrdE+w72cri
3skcG/MjilDgpDaI2G/fUcqMSqJ6GI6cpBezdq6tO5SUt2GzxjtdnvRoC/RYbzW0
wNwD9xB8J8XSlrQ1HG0mhcI6kynPuFdXiZ9G0SlYfF8a0yjz/O0UnkjeGUQMc9oP
4QKwOp9q1iNVTp7aJJXm9NJssfhi5F59OVyfppC8sDTuNhVn71piLvK5u8K6wTR6
rmpk1amsnCc8Ahq5zeMGB97seUnUEw2uErv6Nj6nGaPdh8Ol8MCauuUTqZKUexeq
zjsGr0wM2/WdLvO8PLiP+iR25VEOrWy7iRM35VtXBq1trTwDq1kGFu+1A+W6woG3
mHjdsv2gr5R0R2bmMWJbOFCwZ+Kn9TSqyX5Uy50rRpMvsm3dCci8vgd/rCmoZiSH
9Pr7JRecKuvPhGW5gbTIWeCxZMikKbQ3rW6P9+ESjsgk9a+H4MTlrtL7Ovx3vyu4
Vshnp4kbwrbXShfSdQCGva+Z/WKTVm7cIZhpbpivexcTtCz8sNyHobAuxuYvm/m9
Mqs0CCnoYkuTMwiw9J1amC2T5jcMECOEqrKE73xOTqJ78vocOEgD1CsVqvRDp7Ke
QiDB/WzKHAuXQdIx2kitOQf91o1r+bznbVK40keKcVfrQFps8Qu8HQa+MCRnfQ8l
oISMGvK3m9zH9JUk6Ea7F9h0A3JwQdBFC/V+mcb8LUv3XMvhun4Gd8blYxJI6kbw
`protect END_PROTECTED
