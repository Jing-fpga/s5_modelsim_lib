`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hlFE/lZOBG7Cqhv+9N8xLfg0cRqaaKuSviww202+MB10N48P0XR2jDd7xRpeEYeM
dFHKJ37OoWjr4Q8kTGSTOBq5MphbNh7dgmeHMfEqg5NJNneUsiZmp7UA01RpAw+o
h8XR9rDGEb4Iquqdhaht5+xzalfkyv/OsssVPwEbypa4/CZuRrqrZOQBUVQ/6UCT
hBnh6WSkSVR7+gacJ4cyeiGE5xghrE/eaz2Vp+M8WJYe6w2nzKw+kb9YeWazxbKf
QWwkPraRF81CjG2qbjkL3INLhegx43ETgpCOHKodK6it+ZPpo0klb5wiSv/mXQvH
ilBiRPUWCwv2SHgcxpeM23wtBnhcERg7FW8Yh63FndTnvUmZ3LxLi3rfjgxdHmJc
f/mrVvfAnJYXiGUgt/AewXZarsFqI3MQny1inpjE/kbZl+sRRUW3/lVB0qX5U61Z
W5Pskzjck7BdfXSDX7zqn8vG2j0mP9xSEo9SJE7lMAZr40LV9ICPN4UVhEVDZcXD
OqfkzKFSNuax7WEufNsN2DbftSuongQCA9YCFEk4MTpqZL67UtTqESEaKARIrMjt
20EcvA4MSPZ/eaMiFVRUv3+LzYz9PuZgjlh1eDvzQOy2HW0DRT9kyoxym8KMT7b6
7lQqis4jWo2G6Wao6d6kuvz3E6Gq+F1zaDeSUC3XoFrqMk/u6QrL7gugN2J4aJpF
X0NSnC3B0S4xGtOyyjyUF0fuZR6NR945YtXd8st4S+klF07Ccgm+Vgtj9xaQ9xCE
cyB07tgX+92lH6otnDdDCSxaNmvvXM6ktX/zALIKMUZ+R82gac8/+faoCC2U9rOc
VqH7/KmFpb5+U8yxIet2GhUplP6lxwbrUzYj38Imo1MwHvv6vTdKCDymegOP1fQa
`protect END_PROTECTED
