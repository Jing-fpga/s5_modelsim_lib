`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sBVUT0Raf7T1keX7WqRaqIaCn/dvao9/UbYcf6uGsaBd3Dqcs/lTrOEHJY4XZ0UG
56SkihA1lvXlQ+WHwtzybajqhFbl6c/Hv8KXFBRB1pH6XKfqWYu2zhDPnunZ8/Nh
xQTV8XlW9x9ZiHLqzwI15Wy9SdOY71JUpRTh2JxvbWYnI023vF1WshVwpf3ld1eO
0k23sv0aGy2WZ08doRFRPzDEwxcAKyiFWrg//qINyZBJQnOtlOOZLiR67rUWjoAl
cWjZOqlYen0eJK7BsVM+HdLCDHGeQP/fLDzODggp+HArXQa8m2bT0EBsBIZlsfKq
TgjdW9sj/PQ1ypcx82nZ2G8If5wTCBSlJHX/8SH3O0iUOMRari0gIAzmnETtDGBw
WIuqC6eu2A9oWn/p1plavpFJPy6U3GWnEp345DBr9xFRW/paWo3pITxqoj9BG77/
j5qv58togvJ9+Efh9RbDMSTnoGlTv2MATuBxaxvDvrZ4CD0F3QSash394lOYopOC
C2K4zes7qNJ3UlWHiMqcGYn+D4ufRcYXt+wAZeLdRR1oo0l7bAwL/qH2F8qqJsOY
ydy9H1b5viT17QuVYFnBjgfvMwUXrnkkOyswSKrESObYLvxyumrfTjoyCa4zhuPU
T0SRN7r7vKxMgenNJ/7Yihr+w+gLdkfvsJBgs7RU92DymK70ctMi/F0XcAHGISLn
tltVhNKgs2r5Z6nGBh6UaXC2YZO9vF8bud3AET7F2ZjCm4j4icak4rtXxPsjyOV3
nutppoprKq3sBMqO0PRHh4uB8DjTgxC7+xjhT9soSYM=
`protect END_PROTECTED
