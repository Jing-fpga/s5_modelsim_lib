`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CVPBXN68iXQh/JhN7mZnoyLeubEOzkxc3WYG9WjkRhsW3/3gn3sUNGKDFzznrJAL
0s5Yr8TiNDsmJI0GivopR/lFq9nyL/qF+ZxQw/afSyP+doS5jPWRMxMfO1+/49ul
5eOo038ON28x2tKHNXRLfs4Lp1GCNkltFlW2zW29H+jjM+u/0sG14lqJ4Xq3oToZ
5EArYTQPAn55+BTWmFehIQHlp63mR/tFTvfXnl8z1tEV9kZC4vEQwK3L8YNBUeg+
ozwW2v4AG6kUUG5tQ7rgHdLHZZC+gpPbo74ofh+0WBXbiHLgL8upWBlcX9oeMwFA
ooyMsIKnkBTEDJZLVMqWl/8eYGcekhwTsB/qikJJvW05/drQ1MCOOz2Du/3W6dnw
jdQcG09IHaM4wYeFBBXWkPh05lrHEfwuW1Cct2ZD+1iT62WXUKm2JjvYhOsaFVB+
`protect END_PROTECTED
