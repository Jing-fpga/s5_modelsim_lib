`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zrNrw7IyXIEntcby7M+4AX5/XKNwPPX6BdNsvJT4anVpyP7H1bldyuX+HI/1SSMy
CygLy8r81/ENetm4oXvProLmJ5BOe5usmSgu7euMX2S1MvTBpbw0ZfkUAmLkx+Ql
uCfHI2PSzLcrHYoAxuS5tPwrkVmZ8zb3lAuT+NXNk9hqEHt5ZNatWZHYIfWBciic
EX6ztUzD+qo2sMfGnXmNe6y0H9LZf46H78l1n7LQ4Hoooe4hjHb3VTWfTw2VHu8b
N0NOJfh1H6DIxVa+DpFCn4YKrkEkIREajecb0TYOtpSyU89PAdi26zZSN0llCKno
XwbKc5o4zUDRoznfEwnlZKP3L4ksWPem+V4lQAfjKk9QYDz8hjTVdrgr50jqcoH8
AMxLWjnZ0Oolsal+dhtzXEGYrf4wGXTqdgOzZblHQ1IhDvuTKdIqKjbkSdrlDcTo
AxKxjBYl0pZiPfpZneR0U2qYOGiUEEka1ERqA6WoNpejxzXxtos9Rxc4dik1t5l9
P9BOrru9O+M+yRN89lDpQn6qZc2Pn9BVihk1qdvyvollVhp1YoWh3k6y+mZyl9+r
C/0TkmPjcl5eARe7xVoxaUfsH28AbTiQAH6TUQ42AoaLIOd7BWxrHSV4+YIqAmlG
FQ+PxyuJ/jnqx29tACjqBp+4PYgAsPFdUluf7HsEQ1xeeRpIIeqlSTBGcBM6y3Cy
aINeKqFA29BHIrldVIu9yZfv+rdFo4LRs4tc2pOAGI1LxniTvRayFNNWBWObpibo
Gp8QjzaqTkxdeZdx3+zwasmtfTDAIlZsG8ID8x4cqY3yX+FMr5sbV5FvMGJ3gm8T
vDI+JtR1XQeohFwMXE4q9SZIAukAZcOPpL12nk9bz8yZ96Yw2is2BIhLLTm4ZYkE
asCVAozKdi6kiuJ4UsQi3U2i5J7yEUPiIxSpZhX60Z+20C+gfPR5gdJ3+Cszwrb+
MBJqEv58HFeLp4/OcPNH1UEHEGArzdMr/57fPLjkIKQjwqRw/BaGNm2RZ1bqXP8S
1hkyiFLcJb0WUY+lgrikMymRoNat32tsCCzW92cSX/YBs9JK73mVxaMPS1K1P1KZ
p4T+sCeNu1BlzrmK8R2uao/3Jn+7Z19szWh33XeidFsMyaMhXRAWw4VOie6R6GXR
jFL98NkIm/hJ8exzzGF+msE6T0Y6ydjGqHLS3jh6s3c21MXiU2DULi24i8pfflc3
1DQmOv4aTT/w5XK3fuWv8NwA959VRMLxNuVrOxSfph2lciJlPZRJJR9/i1wUbM57
TiNQEWaDKdbGulWFiwe/qSQ+FrBZHYWit+YUiKqcZxGoTTgGwPXuPGjRng7+2UgG
iRAnJQicsaWgVECYE89/1ikxsF6DWrGFMdQDE7DZM0Kev58NFfOTy+VJojvfgtYN
ynF4WZToneqv5DH6d1lPqSVQOt/MVLIPzA+F8SA/lzRat2FwWrzfyrpwN59v/vKE
LETWA7pC8fwWlz8wkCeGvb6FWeyMMr2fjS+yU8+l197XiL60ljtuHTj/tHfc8qlq
88uYzPjrr36Pw4QJuyMC8PdMgzbV00umWi0JAbcFNfyOPiyQPV2KB1AnI27qMrU3
/DRwC5gMEKlickeJ/V8iY+U1B8Gl49HiZCbmsf7BtUAmuwdgIk625jtEBDUZ+0th
UiExCHyBdAse9dXEQablaRS44tMZQ4RjZ2ccQMunN25GFwQM+lNswIbU07w5tofr
sVkBpwgyzsG9bXRGSTquFHfoSYWsS9MGU3x1NpwZGh+nPPtgT3b7HDloA+5RR6nJ
j3osafDFbL6+IFXSniGNZTNKbBccycf1kx8flIDIf6m4mo7P6pLCn8BLgRgOeayV
Hkf+RZOOSsnHOcONQq1eZRym7fT6jYTl+sq7XR9mtoG1fXLTMv5J1dCjr23CQcBe
m5Cuas6igMPDfRKi6CXNm5pTV47ZRB6pwJonXSYehAZjv8LoeshF8R1u99CEurUQ
vY1eqm8q9k3vPw5WJjJargxTElJCxYIYsN1i2y02cxZrWfay2QXKRdDcZlNv/BSR
tkcx+Dr2LmRMNocAAk6RWOIkYZJmvcC20Y8eC5uU+kNcVsva+jiAaWl9DhWRp5BC
R3wtF459sdJO8KbkHQA5eWhCR7pMHePPSpPq2j9YWKjgYKx3mPhDMsO4JY+5ecvf
MdlG7j3ckgwhmHdvkhS+xE6ntoKwRwp1M2N/SPlc+rXtIib8ohGgUZCEIAJ7P9Vq
X60IirFRGQRtBObDhhJCip3HcPmdrqPeRFV1Qp8RJWpGyxz8dHjAGlru5KLgpBS4
jZT+iM8Dx3xdwUjHrGypMR0x6Oasv4JiHk/tiA17Wgke1nz6CV6paoxpNz0wGQHU
lpuHgRPyq9V13AaKtUm1+ibC1LM8mCDWiyj2iN47FAewSGUIvC6NiAjlS4Uaw2Lu
QKMbK4DgVx41glbu9jR4nfkx9sMmngr7XLB0bQQ9MtSH46FQzQqdN8x2TNpZsKou
Z/YK61G8nyHfU2Vq6I7ahOf04bZWEWyDNA6wn5bOKH25qqWxbIPFpb+4VllLSU4o
UfvRppE1UIFi2oX1Ok0R119GNgjXIXpDkXC4qQyg81Uvac70GM0FwgfMt+NTMOAn
cERxS7l0qTwXTinbrF+N2nA7gBZlrWZQNrjrPHLntKvBxIq6Aw59Xdu6I2VIucGw
oRoIsPGV98k6i+42mBG4OMI3kLWN0mMl5O7QYBKkllxQQjWWcfL4JJdSzbB30QW1
soDOMiW4H7+1tat/gu4WY1pPiqag59CZE6wIECbDsgs220h48vozrjG+zRU0behG
JPoHkhT5EyZRT4TeYBtnFvsQeO5x1j44/x6PPiBOXSElL3ZIi9PMqSnZHenPaCOD
NqhXkpMtQBv4Q0kr3Vds+L7irYUl4GFUuIJL9n7HHq8MPIPCOy8sFXuMyLY8vhU5
aLhkn2NXxIW4rybGzzzF1ceuH+vEbyClz+NGq9Y3vwitB9BNxbk75iha8JUnzhdp
7Gd6GxGxErhMJfb2mABS8HHTlH9U0/atqKC0AbH4PDgGLvxKe/xxIMH62/LGf4ov
2GUUY9aVxH4dfvgm1RU0JTtH2+NnaTro+vnpNvvdEDGzW96G9egfRmcNbk59T1N5
8lTcuE8YuEfp9Ren6o3RJiP2G0rYHkPSRzJvhg67Flj9wRNfMHvZQHkdKKTsb/zx
GG37Ue1WvfUBI2UmBqefzy/rj0hWcCZtOhuBp2IAN/z/sLI3ncgiLFehztSq04Jt
yGZoqC5kQIhHYZpan9EkRbp7NzWRRO0fUCfhGjnduwXRSdj+ab6+O+OavJ921YyK
sy/oWsCbJOHnwTWKqzKii1djODLEz8GCnpeQMDmM/S3b/jbewQLKT2e834Km1kAC
KYbcYhBUv+CK5BDwHIJhkGCZhr3I716Klm6VTW/j03Jr2vGGs+Lt1vn7v/4ONerT
dsJRZ4/1b4xeBw8HXrEVULnjEhbTw0AstNuLs+aknouLYNhJPvBVGN+GsABqBWGT
GMcMhFClI8JE6eTbcZjqPxTtCbzPjh/I8iHdofZ969bc0O0DrNbJMhEdeSaDwV50
7oaCfZRcckgTqu6B4FCywzwr1TUuctyKzod1IHHdXxyS4nE5e40YESuzxkkBf42i
eWWV4KsWM8D9LrZ+TMdxJwJSDVXiCd6PbBY0SDZCyXNPHEuJuvblvcLUK7dgAv+0
SLEES3YQb6VcBTtpTqw+J8j/qiLPLHXFk9aY2Mow1zzWJ6rJRt5lB3vQFGFvPKhZ
g4a7g2HAF77mRb3LbG0UV9nfE3xjGKxUtrG3ZwGqb1qhf+/YkYC4uj3HW7TXwXSH
/U4f0x1UYsKfQSdXFSgTqVREImX8Yo/R2fYxYR0Y4pgq/rSl/y3n5Kx5UAM4C/fg
7Ml+h/q2NbK3bz3tEbLHMdZcHIrtwYutPN5g0db/K6k5/dILKIO8GBs8ydVLhRYE
ZgHKqVWHANoMZXQbY/CqJ0jxbZb1QocZWysfdcYZ4ldGE7AGy1+wajBxFF2MpLQN
MfFQ6h0msGxr3Cr1IKSEiUv1IJ9abZwp1cVDdLrgp+y4Usok/Rkp2iAoPIj4yIoO
ziMC/oqDCPZjuXin9HuayyzTAqL+nwG9Ip12HJd97uqZQwf3owlv8ppK+dBLBh3O
cC+F7IxpvzeykTydgaABYPyH8Hgnf/UGUEBgtJHuCNjUJD+VOYR4vIcAlFA5k4Jn
H/rvbD1H7CBWkN8opRTSsqmZ0qdZ5pDVQB7SMF28iZBa3VhVuGCGFcpkZG2BVCTF
f/5OHUgg/u9UDiPEuRybNT+yLUdB2ZkYwc+GJL4dbLOMIZMHh9T59tSRnaugUEEY
sXaoM+6Kjf4w+5dwL3qrw+w3iajNitr6wDhl44qo2geq7fy48O/0hwTV4ErM5Mkd
B617THoXZGgU1ZSHjbpLX0qELtfoO6vIEotYH6Uyp6EGPB1EsuaJAjsFMDzoXZzU
0gNrbC+pfRaVEN4YPuz9A0R5eTOCJWRb8y+tKE0p/ly40wgrSWGN/67Gr5+kbBV0
C/YzIGbDyp3woxvzomzCq5gguBBAUWE31DREIej/58jo6qjHFjIXzJLK8Gbfuw+f
rUO7PyKl59bnrlzZR2jRghn8SawGgw553cCbarm9vjPoi5c16JqYWV3vJ848dSiG
DQ3fhafcjYjEoCY5w2aZJ98b9t6It4i4mVarzxCQoW8=
`protect END_PROTECTED
