`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Et4wZqsBybfXlC5P5SIQFtf4Po6QnxI2CUaj2bG5EGQJTSAEnmKG3p2aS7TrXCK0
LF1m8RQQigCNfkBSvtNkVVS2oI/gEYsROTdNVh28/S4w1P6hzhj9cAry/937wm1u
HnB1Xs1dMNIYhhxoz7sceuynhc9V6aw9Maq9yN4RSHLWMTRjsw62eW8nkjvlOK9C
IPifMZfUxTPNZWGFsMO8tDOzbLnVKqWYwX5m6L/9pkW/h5ioZrYhUqvfv2Yf1N6L
kAcVgc5PHIXfMzn0AsrAm0mydcryDAZvc4vBeW7WWQVmVqDvBUuymfSG9Lr5byfU
yQ1f5urbIwPUPEpNAVssvHW8TOoRc8MyNvK2pA90mh4Wzu7A69ln7mA38UP5oUh9
H9daSlO4mucPB4OhMrl/qlEL9+T4yVGCvn6mdjQ38P1wqBJRW721Z3BCauqe3M6k
Ji23/bxBrIX2T9+b4yoV0tRFXafU1gAmxJBkbxXR1lc5o7dPJyV2k+UycdwTr/VQ
uG16b5hn7UbuEQs0KvfdGlahrsPV6Du8n14K0PJTFE905uJERjBt4cmyWXr9ma57
hhwvrbzeRY2NjVRLJjDtwm3N9EBbcxN5Tz65pzfPALqGSpMG4AMvMXxH/TbPPw+h
c7siDwgtQDFYKGMxXH0o0wubBm6ETFojFaPQLiBLQBRqpoVoUy1cn/TzxrpQfvSw
9or/Ps7aIKb7L+HjkRFYuMRVizZNyysSrIHdb302y+cbO5OJB52YHh/Bz9JnDRrU
zdjVw2hHdYdROKODGWaeuInvmNx+5GZ6NpPSa6x74ZEegE9Gqrl6jCsy1tyGtgMe
jF07cMpjPbIZ57idkHL9D/Wlp1J+FZ00QfcktHQCzIzgawyluLReTj2/bYeoHP0P
BDhUD93GPGGK08Og+0FVgXwJ1yAVNiKen/F2PLsgd0x8Iz2/kPhW/ln3kePkecbw
747GcqA/E1IbRiyN2morKOVPkZ6ADKSdpv2Rv680M1lKyJobBvTRVVQ2JzbYAWtn
BCFahLgLganX0/f4HeTv8OlL6hrwD32nCgAKOqCjQzbGlfRYvGXX6Kxl+SPyoNsO
qcOD4/zuzzpuyHNs/Kvo1TuVc/1jVi3A7qpb8RQVpT8DE3PRxi2kPBHu14RPxoQC
pKnU/KHQsW2adZfM2m43dDdQBc4RazUDEnSkV4vLWu5S1BPz2Vx+hgMVh+3wnAOZ
mgujWeEWkSi9pa+6z/xysSeXgj0n4U/bIzfW9DmD9HqsBIOk1Tpqewpj0DmFXdTI
76bK0GBPiynYhhYcx+K2yBvrfqsZNLHo5raoyXHUhfp/Yrwn6qeYxmt1i0t3n6HB
PG8sFTRpp0yaEBPnA0dg0dNNCyZRm2XWvZa5Hbx7ImQPXlObBgnxpgP1boRdr5nx
aBaYS1Y1Bc+Nl9kV6wgvjYn+8jrxVZiYO56BnS2ttOmfsFUI4jmS0c9mK+8aUyHU
THaVee07u+5nvxhjLyOMr92Pm9FAuzKaUg6x6KDkB1ySwAdPuvYQwY8koA5ejNGV
Ar67lgtjJ0CyykepOpaiIk/CG1S7FhoQ7skcN++sKYzJVdX/FOIi8iKmQHn8EF5r
LX1r3DffS5PiX1sUedRiVbbzlV6PSi2DxGbclBJ88M+750kfyGsb+kkb7cWpimJI
i3MrmeoTV3hOGOdyMYBEQSUmFfQwjd+mmFae9RTW67rqnNISAB6Bq6pVadrcwMFp
Vco/2lXE2VIKtN6HqBXbx6KiR1doNQYBd7uKeyv2B+oIT/6EhLmg6IuOk0c4xXsd
/4emZEpNu/UOND9ZErJ/OLPb+WtwkMTkoYTBYNyR8Zi80YaR1qq3ad6X3Y+MDOyF
BEmgp5x67qsPacz8YGjygh+mGa5lffq8R/5kwsMCwdqwy3gvYTCkDx8U220PVzFS
GMBGZ3FW5kLQBg2SMdb+gzOf9aoNAqDfMRMFqS9gMVgCYgwNcB3vYwqf3Hs1XxhT
`protect END_PROTECTED
