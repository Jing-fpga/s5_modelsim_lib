`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yzg+xhbtn5iEu0K3u1oTaWryDZNkijdhHCClrKCP1H3Ddm4CNwzpPldUNiJm+O/C
nxgO3U11wqi2+CR+rwhvQC1OAuVk2XQlzsoOJ2jjfIUsWzZmJzQ+5AXnwLytLkXs
Q7MzX0o13OJ9lIOz/M6FT14NDbZrVfQxzsQoMyjUWlbCLHjJM3hy/d1kmxJsTd82
5gI563bVFh1Mtt99rKE/PcQnKC3owMpuw6a7rjUQQvbb+fQoMgPO90QR9ya/itTr
iX8FnuBTN7+NMYmiQtYO6QM4567jiJ8YEf/C4v9ftG0Eo9eRdTi6KA91fFHVnne/
HGeWZNzHkE1v2GGBU/zy8miwrIeefS67hcXAdvv/D3Ed33FV+U5KyZqUkXYwFDvk
McRJWOr/4r5ZRfIOO3ffqd9+w288aN9ApuiwxEpZzDwuUeH6yXiWCOVhOFfu8mfj
H3vxalsRDwPutWS31HWG/1oTaBvx+eKUfKLnoBIJrjBsfC6y3x2DjTMOzzfh/4z3
aGBIu2K2Qq4LuClrqsf3ZLfdPAW6j56ZgxXQ10MwZrLKryfDiXxiejUx55rq6/TR
HPMFoIF+Z6rpzWHggsd7q2nhp54lOIGOp8e92yXUSK26NEml5OowjMqLcaP8m2M8
49++vfTEiuiHAaKKdVX5wOUpA/tpDoRHf3Cjdj+YLGRbo5W+gAKXpwU0V12PudOQ
XjT8QUu58uGvEN4CNjsTdKMZ4+7bDUTpgzhVrxPl4MuWSBeHLIx9Bw+JqsACAu8b
91GmhnojY9A3rrzRNmSfjMyUSSwUuDc6zpetRHG/1KH0MpssiYI/+06bSj+M+9GC
Cfk6aCp68m2eDsXVPSsaKjwmlyjQf4LuHgHh7apRGGcq4B/Cmae9H6HrHJAMv7S7
2DigiUS6doGgza6R7P73fYHtCR2/2K7GV4jIai4NjeKzS2ZMykzm12spTcpf0yJS
/VGCkVAmn1pw3TsVQD6ap5zcjyrpWulaADSgH7cxPKwXdZN56jtEolUNb3CH9YO0
r4JPt0OnhA9MEtWV7qYZ08Zhvx3pfIwaPpXs8k84HkW8wzPJRugkJXKh3LxC05HM
VCJZTYbuY4PFuGkmPubXZDNIIZ7e4FapGMPS6t5cdnDBJX3vIP0+Bkywn0GyJD8I
OtUu96O/ykzApNWPu8PebmpkvcKAOm626uxRAICOLE8+tv4lqTK2TjGdbQlKnKJx
2egDj35TQaKnUCQlZ+SDs9whqIMhPy5dJbyBDzbuCt2oAMwJlPnjQikiXxGnvP1t
e5y+GMVSiIxwMtSdMGNZT3n7wS7FAixXl3Psfg23O1jMkNlFOsxc6TQoWOYSQ7KX
ha7bU1Vw1VIw6DYaPD0/qEYyXAMUtu9ExX8Tz+x9YZQasoKuYXc5iQ/PuzpgE/Nj
lA7rPY6tBeXmijG0gTjCzl5XWTLspyd33eMxkQCAiUyezu6QqxWUNOjzeqnbzE+x
3RGNyKvzlHr0MZOnJLguh/hwEF6BKog1IHiIphpL9eurRxvgPmSSTehQvR5CvgCJ
2oveuyf8EACux2eZy3PucuVIIA8dMwn5CAyFue0lbj6CW5DwNBNqUMRhG+SMJc5E
79uKYjl8A0Dw1sp4smEPH1rQSowIxP+V2fSX69lpPgGlMsIxqOKGK2FV5dXRcZaS
9t4Qy7cu5q/KZVrpIKYGaTOEgibluCQU+GNnbFR6UcBz8zWRmfs7VyisOeGlUz9u
YeeBxjM0D3UVh4urRt2FFCfc+7PX/FPlbLratYFNnk+eTmjYC+VVMHVL9Qq/OLlk
pGPdQP995rqxfgA4jEgKP1sENokAFVJGZnwDHL+3wDN7ArJSV40ZdZG2XT2fhvEx
QhhZmps/9guwh4J1HfA8+1UDTAJ8gNdCHY1CCvkOs1p97fqa/J2fywnOMwV12nkf
xz6R51TWO/+Fr4X4aceYKvf6XPFYPskHbnrAWZDDk2PZki+qNKxTpPhOI9pW8CYQ
Sf5J2yrd79MT0xNtZo9McNBzNbpm8fTgV3Rd+y2KKCjCcSbaQA8K546PDzNlJPaA
4pZ7WLUMmbCc2O5JPo24zOI76HT49JkxdVEUHyI53LI2L2iPBQab1IL/vnQeFYch
ulhmiYMdQOE7YsodPSMmOjE6jF7rMewCVkOAyy7R/2ZY5ctNwLKehBN0s7KmQYws
AsQzBZlXcqNBWw4MM02s9q3B9uPv/PKpsCCXLRYsNWLvVF1EH2nfziEm7USq83Va
3P9eGiRmm/e851/LF+JBirw+CMZlGi+Mwrr4cQrVkU7THrkqsfYSp1F+ikIAm/M4
gNqXA5SuAEvFX8M3p4tWpCMAyit2UmbJoYrg4X2WkyvQ+jqVmlMF5QAks0w/6WL9
mVxLx/cLEtUMp6Mw0EGliUDpNnCQAVXKUo4Q14hI5iuMFWaguo1FBsvDiUcu1kxb
fi7H2mvsXIdSOvJZoR62DQ==
`protect END_PROTECTED
