`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dTv+MAeqIE0o8rV2S72Rz/F88n7++t+AC5L17/LQlJKCrIU8oA0ZBSalX7GafQ/j
svGre6JPYj96ebRHvpbd8l1/WPAvLwA7CFeAUntjAzCHPIOxCvfNUE44mi3/UI93
sawPblir2IBLCIdEJo62uuRs5Sb+MaRHrANyLofaAfeqn3p5VVJJXTyvpERe1idz
sVvqahoh4JK7eohcW6Sofo4svFycCh+yFKzvV6oLdShQKqJw2yX+A29M/iAZkSrX
qmbcp0DWyKX4dRo80m21l+twY6bLFLgSmdva9uAMpZdxt+h4rJyos8MZVGlHo7ks
vUIEW7uApPzA9V2Ei42K4k5umSrjibuFqVojqOAP2REqt8akNPllCrO8Hijizwn3
LTb8AtDYPItoaf9bwk2VqavGL8/TOTJsWlpY/gey4Mm61ff2T93EEuKbp+hQo7eE
DCUYLDZVkITU9eF2W1sb7CtysAZjDrp31vSqZ32XHnlhL5Q8p/kiwvo9oR1pEK6o
ItpNAAG6RtJ0nhe2SuunpV0S+xAmql5qpWELcYZ05z4=
`protect END_PROTECTED
