`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O9Bm+eexHNY83cTSKQQndH7wu8zqMZW8FSqJZ+iKPBDXOUOajF9zA3FfSyJtXXuy
GjcuUbVv3GfABQBaeO5Yk48vBu4TKMs3JgtY8jysh602eIQrwlR2LH7iQRMWra1R
vXQQQlECW0SxtFBrgIGFJQz383v00rLrA4wsFIhpWw7zO2Zg5Cu7bjX8K9ZeMG3J
qY0r40nu69TWgK32SdkbcZLhbYSxAYGovSmuGyp8/nOFJzdUaTIIPThw5duDaDNB
vHQoy3hhUvLazMYWF4gPAQXgeCClu1HRnhmRGanKJ9+XLjtTI/nw95jeOLJHgFqJ
dxGWlJaVUwro/CtyTK+jwm8E0om1r9Lka6IVw8PvFIHs+6owWwmbfnQKd6LIFAZc
ISE6Ym1wZ9Pglc4rxpoRRDS2y7mh81vFVzx1DCh8VXDIbZQpG7Lj2JDg4z2jf75U
9An60YZZawDkX7nwzbvGP3MjiISzgPWsZW5hYjNVIgcRJHM76g/HtLIqjmzUHTNo
yCZG1SvcekOXsfZu5S3UCabzyNa+qoxXCrGGg0Bju/bA3J1eSZork3uSYd7c8jiN
Pa8ACiBwgWuC118Jk33w4LbxkVepqEDt38E3L4ZaAgxxfC5/Op7WBNaX58ZXwrY5
LrHl0r87GpovXifXsKBQjkJ2ZTKOcxmi+CrjiuYC1bOzj4CqGPOQ30OOYSqQtO/W
ikmNrqj7aGSgUwjWIZ36KrfYs+/a6pX0G03XPsWmHeuPcE89VyBcju4yiuN/bCLp
jLIW0SpTZJ34F4cGO4KgVj2/Pbs2A79p6r7EDaRdlZ6+9ZXScdNJ8/tKo0ug9Ybk
E/BH2VdRMB79tMJ/zWCNqM/IV2yqTgHwreyEMBZvXah57PkqJJbfCzYdf0w9dWB9
E8tuggg9y01hNO6QagEIyckzYgRFwGnlWzhHXzXuSBguhDyLeCSgdTXzVGaI1ijX
2FzxAJwdFSZsxzOGzHaX18HcvCSKdBGoqzkTAM2Ubbqh+U330GKme4y0C3t/SlDL
zcIBOTfXVpfrkKUeAsaGDSGvjpkx1TXd+d9mxpjgML6pxsQrFovxE2wCficM4pj7
EcR1Z3dDTMiJyv6Rbv4MX1LJWELOAKEV19NbsKxHzxQ2VTK2pCuBeSXmAPkYgd5l
W/0Xc42p/akqLWuVaPr5AZ99w5/UFFfnAHc5KbQJbfuGDmf1ZUVQha9OAhmAibdf
l4HTw5Hl8K2Vk7TOG6StGOVonVdh+Fu7fBiQKi3z0+nI5avHRwi7uTjUc8o+cg/+
D6+GzYy5mpZ+7RKs3cmvu/k8yiKxpccj+3BDL7kZ84dsqNXC310pmC/a2780dG5c
MuTuMvAJEcqVnls76Kx1x2pgT3Zj2tdZHgc+8vnT25S+dr16qravL9gKUBaON0iL
Mux7N1fU86++jE9j3mme5Kg9TYXApiUwBKkZ6cqJj9FvWGKueg6VDpBvNqm6gGiI
16J0cy1W9oZrb4rcVK8WU1rZnlUizaKgikNF0ciZmMeoIedIR0KGugaK+cQK8e9D
Jpit4FbvKeCeD6KK8TghojfZuNwpj4Y07SNDqmYyeLH8Anl4vSV2QhuNGHhn7Y8A
rmsphrRJgq7GbzaWgKoT2HSSjUr+8MkgHosyJQL/JqHSYYhiu02grcsKKlBab8Pj
PtAkUVw6D6KEbUvgdksYc4j5CbK4nHIk73fbcoQV7YgxQ9FOGY4lS01CysevGhr2
I+OuLOfRC2Sdo/yJrmF+oh33vBkTCj60CFCKBLyPg8z/0JjSPdj6xSwqrgCR8x57
koWwPQUTNMGrYQwxAdgwsFDDr/IZCfQxH4H5E6eGYibuZQQ5akRzIyouFUldVJUE
mpSU+Gjv3g6zVziHpKpjBpv44h0eDoec3us9oYiDnRfpG9V2ZvPEcb9A5MUJaPYp
GaMPi9aTorOvoSQAoXkceDofUIXBlPPjD4mkJdq7E4Mr3XsS9rWbkbco2NzI9R4d
XizgKLSguR3oK5Fri4M8k8MlAtFleDR2XSHFKHNrvFyT8AYZX1TaYyeGWZ4ytkMp
HkuIUy+j09/qn3IeW9lXBz8OOLm7DrlMCZjGHv7yZJ3KGNo60du+2ZEsSb2aT7XY
hrVICAF1LxgbUlfqParu0DGTawDWfg+mfIAGWHobiVA7r0YKfiWy70PLnGICT0iQ
4+tGsQWMNXUUKlkFeqOah9k21ZQc680dahby+/BGNPhMBM5NY8hTA6YIUc2JxOyO
3u5wJQe8yJG1Uubqn0OtON5QsUfitLiNfMP+nYh2eYS26sLZhX6K43bl+tMejrFt
yPnfvPQEMqVQlrmBfibJKbPu5lG1KIl5UIvYXdGPLOyQws00mtJ1Omq/zwquuzAE
CN2h0O8vT3mVeb5WBPQ+zvZmEJgMYThM+DqtlEcubXqYO4oZkV9XH4G4SLUFJxTf
Mdbk2Xi1Bm4JA/KO+VFw5kVoJ81ouvHZA9M0lkidxp2vr8umTI9/Ue0ZyJgXwPUq
yqN+MlaajAi1MTsJIqDC5bEkvBX+29s7BIkYQT13ZOGO5sjPFGiQ5ivdIEWleorC
y2ikNqwp4FS6DKiINHXJ1kt8jEgmCKEfjIhanB8cLoIafs4rZJgNFULG5gkUedFq
JVO/XA1kQ/kCuTu2ceu28MWxfDDpKzX3QIHI6Dh/3puu/YQba5hCbyhNX7LNLgfH
8XHDKcFwl4X73HAFFc6jw3MgeN17LeOqChdgGujdfkG7AW8Uo/eHCVwgo8wQLLzA
n0PZGm7v0p1pEoXEPyo3ag3oLzuhRHYx7djdiT6ZSwznGu9PxAELP2VTaNNotEcC
//ZgoxHj3SeCEDHyn2Q4QrHjS+Cev4Sf86glI8Xc3ksV4t7Fe0/Vr6yXTr7A0mN5
LC83j2Lm6t2MiQS5J6zCnhIODZ+JwPr6oaXGtpsiSEzyVhAusAxhTivRDx/ss9Q0
bBXGGMm4BShB5BPzR5Zwppx1vqhVEnfxE8tB4Ua1XoeHPKiDsiOO/Txvcf336syx
bltu/q0DxEPEFEaikSU1C4qr22IYSTyEmzFT+JRutjNgwMXBBblyOVtZzrFkmzce
+A5sP1LVHHxSoamv+BnCY2XGTCwkRS/SYaoJ5OAstlEVNYM5zxheje/hjHhFw6Lx
OpSsB9M/9msd3VL9axvWg4rDpB0TJTg45U2/18IPlUyGL8nWIFgoLiDhmZu3pmd8
FBstNejoDC0WcWY0ILq0K1QvZ2goQpTxhe4gIw7NTpDnwPzocjLmHX03QOvJyv5s
XuHtX7w9UpZXNuEGc2ZwtQM8xFuiOY1K7jDuKlcAyY6TNBrcCQhCH4TaVnIbaxir
Agezxrxl54HlJomy3xtv772tb0hpnchDqqumy6+n8AerTvHwVwZDEz/4EYhgQnE7
BiDNtnh+DOwUnYmSjVARc7ByMCDZc80VHATftG+hb6E/tjxWOgKUpJBdRA5yVZHr
9dhfD4DILiHjcsJA0bAA/I0PqyfJjLKM3Kpk+MeA0jeu3/Vs58iOSeSQjPxybglj
9Amv5HhtspYzX/w/8LqODABs6wmvpgYeleQPM7nkSLcZKbf8I0EZlyR3VrrqpOwN
EF+X6NC4emNZUapItIMRAbIZKW+pyuj95v8GkjykYow11n5/XIG1ckzLT853t0EH
BLZ/iWGZr5t9G34sUvExAZwv5ZevrfKHeqyEkXP3PzHScIS0MsCXdn566jsUKJZ2
XmMS5RtKt3T3ClzkStrRjDaT4FX2y9IAN7JkmcVZCuWoNjKwku43J6rGV2XdqFKy
UFJyLHgbtitxmyzbdbjnXpHlgR4xbosOPXxClEAAdkQA3yYEUVyIVutD6nPmi/rK
PIKEQjTLtGucE6KcvUlKDCHb3j9GclfOgCmDQUVviVZWIi+6qVc/+ppjXNgdYcWl
40TiRsf+xXCQVAYNnm/oUOHI8IPaT4Oj6K7eTesOIuCPQwrU11C9uiH0pBbMKZnn
pRywelGXbUJLe85bDfZy0MYs3TqULIMv4ygOFLkto/+7Dw0egbzBvRRyObe+QP5x
HAe+UC9p1JqwT3cKojUrcGCwrS14NZprqJBr5HGAXPupPcTBQ+biNQLXztMmVLc5
q/vE4xuJjNwIwKHwUn/AtE1QiTtMMe5+xlEnXj6cfI/TKo56od6kHC0xdosRjA26
zj+3ZcxQLISHToKkZcmjiCHTo7G6K6Id/AzbvZXuDIwjLL1dKYAly4HTD/27OMry
Qa9dl+Jw3xhCE3WyloM9r4OHrwwL3FWoOLoGDqw3hjZaPm+MFbjp5Z3H1Bl48Tl+
WhpBQsJ2MjhbPpT2XcWIipQfgMAOM5t0noTM9eBRw+S47HsFdiOEiU27aYzAh4lu
h2+swfkIoRZeL75S7fZHwvhOS2J9nTwRDI58CAuS0i5yMZk4BAormEX0tqPAZFmn
YqawEpEI/tSph+pVCYfzf1Gw/7D2CwXU4UMJpxDYXK8wPRbxfHdGhpYRZ+FkmhvY
HudvZrx5CSW8b3rB7Dz4edPY7N89HV+tQDbjIEze2HKqnuT2aHSYb1cvFYKbE8UI
iwFRjpGK6RgY88EwEHvVN2SkrQQJ0Z2mxiuxNZd3exRg+8n7hSbka+cQ23fpbqEk
c0e1nfpVpLRs0uuoR4Tc3ByGcoklV5E66zSyVPo1Qnn0ADk14viYiYtK2490s26B
7We/Lgn0/4HbK1DB2GvFsuPpPS1oDeA/df8SnU6iNyFWUhK67/YTcnoRUQ4Aiyok
+/dOtMnfPJGPcXTqtnc5767FR5niz4zyOAvPAeXnSdUiRcfzqjttuqTGCiGnUVNu
VYSMwNKGRnRn7RXNkqjbTR8EJ323TxnH9mAkRHfpcM+aRHZeDA4iBz+bu65aaKgv
zAB3DJN6kCiMQXNmEZbNpfFiSs5MdfacIWrhzGuvcpphtvkH7lsk6ShzbM+ReONE
jeilxka+2ECy7zQq34y66mcyl1eWIi2wo00XmDZR3fmXk1Lum+lVpfWjaa+lRh+Z
Ut+/sB4kNXvlgoejiCr3LTJpAbWJJpMePBqUKK/rh8iJ5rPgBeEXkX3+AcNNvL5I
N3zPq+HGNxnajl/Vcgyjh6CoOKJlNo/n1iVxebOYrmD5XTF6y4zNl4msIRB3BpJ2
42nBfGcxwxcEqc8vx04gs3EycflCQPSMP8GVFOgBSFmVleF1dCfU5CQGfHBBYw10
9j5DQaha3slPU5zmsJHGalkoitlQZ92AMKlr4d0bfTbOsW/8K5DMoWBJWRIVOOII
zI0MqyEaN0bgtbL9SC+B+l8WLjb1FmO1Ywj2HDDpbAwNbCUHHs4XZuyeTUHjs6Ni
dYqVYv3DuQtxt8L+4a6HgfYImfnNrYRUGJoJt+rmo5zQwP4/bSaSmrFcm5s1qmEg
ANyEzx0LEZstu65z5RAdRnZKkyngzYISOLhcKzOlwtWgpvCxh9hHeVqMN0P244de
DM4tgD/V2i3J1He2J7OCW95nL8+L2LgSZchcR87xF8DszqDm9cGtfAmOyBe7Xek/
HnrWlHmdFU9ZE1pi+A4bHC0gDbLobhRItLYXatrFlfl+uFQq6y3w/mP0Jc6SZ0PV
TfHppWZER8RIlQeuoMGLa5qOrJPLy62+eyfJA8HfxGBsUb6/p8PbxNmCnWznxyRd
Xn4Zs5yhsqmnL/LEqG8+He1s8NR+zMusTfRRZg8OaYdHL6NuYQQCjZIo0ijjAzPu
PJ3+sGbyav7te3GhaYgcGyyb2UkWtkEsyXVFXaFD8DNAQDFuwHVw2epHhhInvRcm
f3Tof6jDoAiCXfRs/CB+mbGtFQpoi51iqaiX9y4ZS/N/Gjn/PwRT2JnY1isZ0BsA
kYheb9gqfJL7PFwFJmvbdvndznKwZba4bwo4yXl9KfvEigyx3NR0C7aCdaCAUPEs
w8l2VM69z71nt39oSTMvBVhEO1i2T9ix6C3t86X2ODzxgPN5dGIXRHI4YmBiS6Er
QPHLeEHCfoQExIA1jGBT8sB7HbNeSTbJzQ8TG+OYvXNgHKtnIy7WHMYCYzJ2jtqi
YUTP9mza2/sB70d+m7TXrM4zmCvmKrrsabtXCX/ktTeVIJ28IjMeRglDgIHtGqwZ
gxzyXFF8kEmaJaeE6i2LwoyBS1in8/ukgTtSWgvdC7qLYXkMujJJ+SKkLnx0viuc
LG0VVLVA67RfjQP+5K3VDfXZebhLDPbaavSuHxo+3EPHRI+4yezcaWE+DWQeNXKP
3g9NQ3SGDtiLl2rMWi/9EoqiUDBwXGUGAcwXYS6DFwuBuPRpMh4uxTjeSMqWubo+
eLIb+v5tWrZA3eRlYjnrpv/tJA52y2EeMwXjlj/ew3VekmJ2e2gXvV+3zQILLCks
tciveDqOuYgKs0IhDWPkIztWXk4ENwQ4DkYqlAE7txHiHYg+xfcy8uGs/x2RmA0+
UWNFARTHQ9Vj75yRWAYVci/s1q3Ivxmfyon24i9izcRcmyHktHwJHBmz7hYjXXlw
ZHH1PRiDKVpHPE7+BW4mKVzyo/lxYDSTKTvgIu6+IOOkel21pfU8VUjToEir4H0R
tj2eZL7lgu7siadhMTaBTFCNJ2J0wbhwn6ibNGJy8GJkyYFpkHlAEkNGfgaVksrm
f5GbjtuohgohTHv2OdwRW3etkRY2z6k9RyETL4Ex/1g1MEaK8TD9Ci85ZAHPN6+O
ZkDx0yPmTJ465xiIcI5RIOAYuGb+1bYfBFttL8g7dxojkHN9zZYExWD6qY0eNZjK
SaCJeVdd9f4l42zpxOFG81JHsdKBi3KM/mzKsBQKVrDaKbpdzSg1pSOigdBho1JY
mwAUOjz9/dRvVluRKWUIV0AjRHh/yJG2J67k2P8nru15q0XbFP43R7ynXVi54o4F
rRt+wPUp6hOQFnYGi48nd+lRqQihT0N7bRc9ldqRKiU81tI0XEYJ5/XeGX4SzK39
I612oc2KOYeUtpK+Si7Kzte9+EPwobe1bJmJimbke/OCbuDsFyXirX+fcVsZEkoi
L86NQKbQkvBKehh54Dml9l8F4SQY0A0nGB+Tdx3kxBtEV9Fb67g9urRTugrzIHwY
3kFcYnS9eWsoTWsAR3tVaTFLdQAnQoUQNtUSI0BBG7edrnO6XQXh7ufippAb3v/1
hrPs7rl0Ok4KAPvdbAc9QjgVzBXpNO1QXcqn4aXXIvJZJJd5OYgmgCCasqNmFmcX
w9nb/9A0jsPRFn0pW4IvQrRWF8JfflmhMuSYlFqBSkqAke9+oPka+7cE/ACgM/EK
LG7BdP4TWwWdmRbLePDRkI8AIBKLDElhaVjOzOZzHMt3GptxtwhQscA2pfSHICNw
qpzOXKNfCxFHEHLU1+eiIvZ40NyHmAjZbRm1gK79ZJGBp38UyjoHMwuWYLJUNIMp
D0VLlUdyxnQbxcoVQISj8oCbmIQDLa0XU3iet2GNQnAn1L0eaqqvS7Fxgt2/qZJo
2mfhP8fMmQPT295MUfrCx3XrN0hF2jD0uMGcq3zAW0lrIhohxQREg98Za/44C03E
v0UFyLnLZd0Y1+cyM1g6i3J9vKBp4Lpl7fpOS2WpXMLr+IlS+YZDx5ZG4Sk6IZPk
hrvAcpvGNpMgxBcECWR6q1PfOJu87K9Qda6sUeAsNEoEBbWc4lkpuI3ZXVQrgLAn
nEclLrvIMIGnDMZGrqBDENkc+5KbpduqgEGe1lE1Yey3k3yFDWFs5JBUTl/7WAfz
oxSO/8jKyG3mwgtvvE4ukZNPWGUKb9uFU6pUDGc6bZPDMzmadanVHmtTqPQd3iaV
zkhm9+D9MgIyA7J6xYapP3HPxKnSVVs2DG20GwKl0nNpffEP5Um3txgHyebea+kt
g4bli/wavzREo5E1a1GtoBWWxz0JihqqvKJyiFDR583T+ZnKuBsRU4OHOHEVhAP1
7qjBSwx24tuKyg0KaClsVHJQGyvHLqsAkd9iEph3NM8qrFPKegx37f7YSSTr8Uco
z2PHHOz3oqy07RirFt8A2m/yvp1sIzViHKEQ81YorDNvHVjaMmYrwWBim6ZOHFjE
3d53MTXMbAQ3LBgGu2fL+3Jqh4wfjzqoBYFjkgsieLBX4Q0UbFjwReTeRTL7WOyG
b5N92yW2lAxwWinMWCAjXsuf3p9GyI/WOcFk/8mz2LXFCOWEArdpq7uRR1vA1k3l
L7KRfrWrCEJw0wGX2oZ+r7ZpRsaoAh62qjqsPIhgZzpF8jteenIDfMoEVGob62wN
hCGQcuEV8kX3RaFrWJ8GU6f9etE5uHSxWGp4TG5Egg5wGByT6ZdGaHs+uKyMYIhC
8iBvZd5hOG0L5TXFLFM7uDLKo0dg3rh3g0xMTqZX+6a40hZQgYl80YjWUnl7nwRw
2kabqyNrgJpNiaiHCFu75Hp0bM109Y5qegJygfhSgJlIUz9EdbpGqtJADkbcrnRM
SySORVBiQLymjYamyQN4IOtc12pBAOq+237o5FFX1SOYse6l+tijz/KDKTk0+cn7
AYMJKBiIz+mYxXB5enEezEiYKdrdywfzG3XQtowR0x48SqT7Us6APH2QLz/RiNdf
aubQ7DF9td0hmMEsfWtnykkUrE8oMr5V3n/zX/wge2eESPNxLn6IL5A7MaNkFrBs
1FQyQU6KGXnFm/so2PG6IAW+mDtr4xLAibsMjr1wRN6Lrl0/CkcPqMOl8RYdHkB3
GwQCXTCi88YYCbZTKnxc7sJOXeqSkSFjSEjVOA0x0IpuBE8ussPMXKOWtHZX5Rzz
baubdbDhrOotQO4K18mdkZ0gw4xKYCMPQI1gtLnRkRG7d/MaBbWIfGHaChw5A3Jw
OJZBqPO6Y/kU2zepYP61zNFrJhLo8av5NmHPeCCJOvLoUF3jnATm+oKbch2IrXxb
+tqId8eEZdUuKXrFl+tdkV7MFw+xqyWdu4jRQYonIK+A1S3Yu5pUdONVp5kVjQ8j
ciwuN/2Kty3xqJ8/fp8hE9gAw2jw1xr4KU3EwnIPuS93ClclRQfucWfO+ZadhtUR
oMgtC6IHV8o+m2C1yrJB61uvqgUC9hKNaj0/jnu68rdv0mvcyWNlQ0GI/clXwU4N
kePvTuVx2y0xLsfWyH2bywluvVuhGQdmq8NwgWdZU0ZFnms3eGyjP5oYgS510Hpz
`protect END_PROTECTED
