`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6qNJ62rY8I6EFl4rIS568QDYzrnlJzbanGgDmn8RDW9nz8iefxeHT2QSAN3KpNXr
U8CShBcsQpWlDqSPhqIcCugZAvBPIGz0RX64/vuDDaIkTmCIKLWBIVMTXRXSSuwI
1mve5mR/SNUtD4YSoJkXSxlfvilixrfDBMhhNMDYoBs6Oq8xiLQDJX7SzAAGzQlr
DZchRq5qR/2B44+W0vyXxc48L2M1j21r5t2i1QtPdo7tTdniRj4yBj5yiYpioFuL
2/xTRmVyeTGiZntH95kArpxNXMqOrQSnePmDUJN5xn5TRgnzGrMiu18KmV/duS/n
OL5uKS2gtmT645z/IH6JilQjs0gK2HRDLfX25RTIiA/kkkZnAxyk7DQJEgQI7zHm
30v/Q/aIhp/ciG/SOR3VxooEQVG+YTKAaQ/CKVW+eADUdBpWE+vDOO8MFx9wue1O
e1xjgMvLG0/yJHLVufFtrVedV1EJ+RVWmlhuJqeiyDC8VLw2XeXGHxCUJ7ANIuQ9
lrgB5J3/GfYLMAAvdtGkubkeMYfJT7RUUf5AThBoXguF5WCBH1aosDXr291z2m1q
OTrrX0LeHp2KHqDYnd85MlFT3OD8rqcCiY6HuEEtYrhFQeAhxE5wc+hHwDKhCc7f
7PS+O2bvYFomf36fa3ST6q2shbZ+Mz5Jpt9MqwxOOTzibeHLL8YGFXxmpDcw3al7
/z0RNwjAI+KE7Q5GTAhhR7d32b0EmFJFtal/jRL/dbYFI/baRAuVGZemxURnqF96
NElxSAjEgI8hV59c8lcX0GaAGW52HyjrH9XY5dv+bzxVFl2YEptcF5zGM+lLZNl5
LKh4DEEAAf2O3CdyR7LxOhLhT8vv1qAP8ja9OKLMHaeJn5NvZ0qtCWPKzngconE1
ELPf9HZEu+Sdz7ANWLS/1t4e2qHnSiN/mL/yoPQYspTPupxkkcJY/uAPSIQT9eOT
FESDIj1Z461LXBUIa1DZseF1l6IhdsoQ+FhdGDE4rx1M4X1q3JIcSc86sRjYP21t
s1lIPDVhUQc+cq8Gvs/xRTE/dMJBxj6RLVg/hGF5s68NNCpebs+ve5eRlTw6Fobd
aKMT7MvJ+1PQwRxs8Zx0tJ4wpyJCsN1gibAFg+YYXGYu1yjaRzHkPVksSJ5KPMIF
MCcDwE9Hx0EDCvSwOsi3sApbrx9aHSoEu5CPAkbMcxQxaSpmar3GkaAxp0VLu4zc
95/hFuk67Yl0NEdxLGL51XlxUqdZ7ByK7z2OpA7SF3uFS1iwPIvZw7Xsev8OOXMz
wfTHkZEQZy2ppInkXTQB2MnWkcRwIgYbAlOSw+yk6DFAYXFGDn0chyjzNHm2VJm7
taLf1x+yMckz600gLK0mnHdAXyNCWsMQeI96pnIPsQZNSKydwOEKySRP4s4nNjyF
KSIFTJRekPCsdaIgp7Ab06fjL/arkQvEJ04xeKlYLKGLelfbpdQrEf1PBQHhci1V
o8Pbp0hErlfE9ZaKv9LsTiboFS4Mu6B8zwvPbaaC1sZb0RGRO/4VCXD0+vdLAYza
sv+kSfvPK9MGVpKlXIZNkWvkKdFMU0Kds8KtNc1xY3NlHA5ykrhb8/80+YwMOKbN
gKB2IsDayGt94ng13YR2qqjAGvOxXoMHwnGmPqsD9BZDaJzKSiDir+sK0U+kCPdc
vUimxeBHsokYueMXTUlVdXOA3RvVnod7TdXI97HvNgbCbzQyXZKRvZ+u4u51AHAC
epLXilhe/32uTzbap+hjFvXvvf0KUl2/FUUgfsSU1iKP2u9Ib/rzyYyV4b7HhjhX
VXz2A/EHkzxxCVnZnUHvdVIezFQPA7lfCPV1dJd1Lu02Z14qlKUiV5JKd2OOOeKL
zjoex2EVu8wAAPCBQvZ/q4heALszGqe89EnH+ufIa/y9We1o346D03apTJjSiNiM
89bJ+vBBajTa0uvcUAQ1v8XErF5zK+1Iy2I879UHwRT8NFQA24KRXZKSIEpJerco
Rv+bgjOBvH0vITCC3FvMSOA6x5iQ1nNwDmD7pzzSGqvmYsMBVssb+sWB0N7paQ5k
WTD1xMZlwnBoqY8ieSOaSY1Mzz7jgF+L3DnvRXUnyrguiWcNIc1pp+oYms/Rp94N
uqGDP0JjHMX5cpgO1WGGBJ7EgV3/9K4TadlS+9IerCrEBqFGh5IQ9wcI5r/1XkBq
bjPFiGCYMHuspi45t5EpZxwtSSy0W+WOKYc4jar1D6vzNk70ePeg7wcFpNUgKRSM
TJGzOvaFXt+FGdGdDdDtB1+RB9OSiUj4geNFGEnty4VAq5RjM7ThlFlkXyqJiyC1
g0EMzgiFe9OdGNVQZv30k1KR+ZW+6XDusBK7krabTHwRFYVqUgLvgT3aW01BfJZN
jDXwq6vtiE1CyJzDIp9QXAK0MTCK60VxkCLwJBh0FhMl34be+ufP0O8K39jZsRn6
BA4HJcz2ubFAWqzRL+yo6JfQLVU7LZ2YD8N/qqqHnCXWzZ02k+MDZGHX0XBkZKwH
ZcquUk5XJXGYAV9dwInfSHATg9Bb/oVL2BeHPuXbCEc=
`protect END_PROTECTED
