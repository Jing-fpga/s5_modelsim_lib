`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XoqgzbbcAUyBZYSj6hcGu9TzCIL3tOoSzLYNu0THy99c3OBuN+FWVZuLsWStWvWW
OFYyMiocJOdXPAfDkM6CDhedMGzQD4UKTVgtZt8Bch152tO+GT0jeRMUCg5YZiie
I2W4tkZQiyJW4jMvI7pprV6tzooYxBrD3TJcsyq5OggLGmHj2TSxjC0uBtfmxYSU
nSwni75zVfau31t65X1CVowOqbuHB91yWd2pHg3QHrpklDKtkavPPsB0X6SCtKGB
MqeypkpmrS0dsmZ9seP8eTWgbtM7qaDlcA0220sLIYAFQeTMWVMcQqhuEXfq/fil
f0u+dpYZhNFHfayQSjF/+bncdewA73WvixW+g9GrOXJeADG1OA0Ms3aLKwRStLjJ
UKtsIRSpGiHsa1pNxMADVfclxUVudtbGAiSjhV6BVE1z6cjr/JQSvSEfJmR6/7NI
+WYmjPTIj+491FRRi1LDKGZNTt4McJMBkKZc2idS54rIr8HNB/zKUM5aOTtTQmeY
`protect END_PROTECTED
