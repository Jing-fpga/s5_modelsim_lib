`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wMeXgQ3SpGCJkFmCxOjhJwxkgxD6Gm2pB0XRdaMJ95qdjxwSHFNPxx7ttJ/CmgVj
Lx5yD+Un7CAnCeooQQkvmakYJJnZO3u5C+BOl9wWM0lNXPUovDks46kActWlgWS3
D1ANTxmTx1muCmgTBYewNnmu2miu8tltvq/Nc4tWDhFOzKjmUNNlMs2mrWS+LBSm
W5ofMNdcfezJSAnIH6n9DYfX3SEdNDZ7ifNfKu8OFvYBFULOgP7/00MXsJQOSxto
q8JldseguAV4GMgCqVmEuI1fsjPl1/vzLiG7Co7drSWXDNrS6nLxUxgZjC/8mRRm
KKuhm77gPtM1TWOMUjBFCedUcL/PfklTiDUF/gvJZPP9ww2mAm1i/IKHDI0hnbqh
zUYah5hMupgE6/8YAQvGJWeIdzikX0GHQo4CpKF8uWBi+Xcv8BSu86E/awl5sgb7
v9CqvYMlRRXcAz0QSk6FoY8R+3x2QAhfmUOJS5sMy2Q8h7okxyt37DXUEg1JED1A
GfNlcaUQuC/joGrZK7WaPmw1IWJNwUZQzIBtq1H0YnS+uDh23fzQsMT0K7Vo2bVv
EQ+CY0K3bEzThpCLfxkbanuBZil30BuxVQ6mOaQBjDGKAWeDVq822Pg5BEfFSR6W
+hObRPiBUCrHPZsBhX3jB233DJvTGy2qmxoFaKFAvjbOlr9MxIjfhNuPjsiIPe3C
fRcUbv9XstB9GNZodxsXnlCtE9K2CmMd9OnTtYzQLimnaeZz4kApfqGGzloKhkzx
5yMt7tVBT0lTctO1DlHPeeFBU8MUPteqpdewIjslLgDv5H/nuwjj/FcgwRz0TaL2
v5B0eL+US00kjMDuO+qsi9ffiQODIwnMJj49BWLEH0sFd5dEfGqUIf6JoLYBsoi9
QfKsKQUURj8TyyIGlYDfAFy4e8YX2ewGY8smdWAANr9OY9gvIzf8IzhUjSTpznk3
XrOt3zb5bj+iLwYvQJTtySTmgptMwEO8BDsHXQRVdHi1MLWu/liH26Qfk1Cdgp3I
/oAC5aGpZKmT5DQE65o2fkA7Lh1Vlg3It2HYHMhUrS56oiU4qPpJ53q1MtWsvR5R
YE8adTiIVSfz4XntaNnC/NbDwf0XOKFPH+kaR1yE8XWKPIpteAiyj7KkGUMs0LZV
8SD/8DVTxARzPqj8imIuslIiK4K81h7Qi5gVal7OcXnpug0hTHy6aMIpR/+AJHaO
A+RURF2L0p2WXT26TD4BA9TxS5SaZ5U99DtDueoEYFi+oUowR4613NgUjX/xGUio
nDfntxu7nUiJNtb9l0mXEn+Os73TUKYAao3elLitkWYx8js4IupocLNaqDQDhfRN
33+8CA+kW/Vb6fcj7x+/O5hFrDHiG0p2ZEXM2z9/voZ9yb3HO81fJyh4ylhaU6Gk
PUDikrmYfBFsiYkWrJOfdJIxTOIzq/G+8poH3g4XK6T9p7Pabm58+UEbbW4HK4hT
kfGfO3kVke7MpCMLh+MrdqZlEdMPm3a6DoBLJRD6aAPMONwNpWnTnH2vncn/k4BX
R1vBAOjf5JG9xJI9gTEBvTQKyoYu7yJA+B7bFGyJihmRKwoxB94HabqDk3IQLyD2
NY8satVe5IjkMCr2tvPs3bO/NYi6uHOKGZgsvi5yacfmCXUba1158JuJRHyiv+Eb
lkeG6kQene+IjGfVrlaSFnZ/cbGD5x6u5JGnwJ0mSG0p9Fa/zeO6l3zENsECeTSi
SbL6VeYLo9Go9ueVYDb3FXVh6GHSLD/9U1kElTTjF5Nc1lhHkJjMPtF4/QkL5YEP
uBIT6INjuAWbC1AmRqTnOEWscioAi7ScIRqqaJB2P2dhyKEByXFBNXAgBC15UHpL
8LZ4Tb3eGL5C1AZhALJygOUDAaRLowSdMF67lfvvrowBzxFF2foOCMMIw7uk4ECe
5+sV315k7x2UitrKiYkGXsVxjuyb0NRXcZ/kAv4S/dvreMh778IF7t7Nga+2nPqh
HZOxK1LBP5m4cpt6krYLOICbyruFA0R5eUTByv/3G8TWfp5qnCqECUILxZXabKOK
4nbaGQr0t44Cv6wiNrRtoyACA/3XUaoAZsf2jXcdwzZAPP0HQdWDC3o0Gd0YyqmR
VutLWnwTW+Ye0nA0pbOPuKS9IaFA8CH1XVMrXZWV6KCj+HpqLSphn4Pwc7Wr1MKV
SU2m2/3CAWFhni2F2LH39NOiYU/rFh5rHZBcK1/5jUkZh6XbXAuWYS5qjgdUGZR9
VsJAYOuctrDdD8Dkl0mVfPmtn/4H+RX4vIb2fk0q3xok6HTwRd6J9ts+2I/ct66+
MGnZL6Mj9Cf6KlO7Yq+5Z00RWEjPxj33EATyrg4GV3OwLf0nzp65QfvAvrEeOpye
knWrJGAY5mKKICU926BaYLdIbAnEirbRO6KSvks8jcSoDTUWIwZb0ZnqSDJ5SE3E
0A22JUkBl4Ski763kwy7JdOpQ8jFdXaK3xrGGJ+hvWKLChBiuwh4mShNBr4CtH8m
pUnlT5h98CuQNxNbCBrgtwTxtMfM/cChZag9q5s3BO4PiH1mk6Hu8rv96xEbCKWM
8WZ+aV7M6TEPsGimXwrGadljrvb2xnifIbnsgHaxomzkZ1D+bJEHXRtT9Du8M/ck
41W7RgOB8AiTrRlqfnrkCHUiymYtGvv6aKGsneJoVmCYRz7R+Pm0t+2zzoH6LEQ2
btMR3zNRhhmNzmx0XGg2UjXQ99ysvZbrAOdmpzLQrWGQE4ACfU+RgBIVjzotddTB
M6jMsgampHPFcndrVK0kPea4ID2RJ/J+Of3wEvaG19INBqIMpnMbT/0kk1YKTQB0
pj+9YCJrQgt3xmj1TpaYmBDyx6Rj92Y1Uj0NHc9h10wEty8H9AA5TBPb2Uk7SE5u
Q+5rFxHK5SJcBI+TBs11mdgPpDeaX2dU1JTi2dwPRyc/1ltfEphHcKyflc9NmWok
OcLn+BZGTY2XABXOqUyrfdTYJI3o2AEi4iupiMdOPZYKXpQa7kQWAPz6pd726B0E
/6cbVrvmNwC9qRB+z4vml7n54M5269Xkoq+vo5s1qqlZ00/B4KYro7WCijdL3ezV
DhcReqk1sqalk2mxERILZ0vIhIKKKQQn9VWRc99Urgolu5/ceW18DaxXSqrIpw+o
pRDf3WPabzqBzVJdptrc9RPtbI1BfWuylAtTT2TqkgUEOAnXMlvZGPfSjS9sc8SA
AQWexUfzZa1Bum6ltWvxlhJ36Sc1Dlu3nWaJFTesbEZabElb1Odyj7ydD7axkRPy
SMlTm/OaqarrHeyRyEoVoWeZ79DSqpQLKGXAbdXm+mPe/XM2kcl5IBIndj41qhzm
U08CsWJzmGstR8DCCLH3C5JH3dhKlG8r3zgXJ/e8rdvJjoXjr5g/pWMTx/KuYa9T
Wj+of0zeuCbiRYn3tqvXvpiQaGVdQSB7cxk5JkXMeIs74s4cxri8eh1yptT97exO
ka0YkV29+iQk8ybYFmviK/AIWzadA+eTbTIcEUoQq9YyJHjTRg0GxIr76q6Lrc2a
xB/eLLnps94cg53hfaiuHU25OFORx3/B8uHq2kvVoM1dLtxXSEH1t9EYCGRsM3IO
vaQwkpnC3YIId+EsnJ1bAgAeDZuuMO2UhbrAoObp58MZ4+ZtOcCQJmLx5bStcBXJ
tE8YqhUoLtxqOfme17Sf7DIHjbeq6e792AUI6wQNZC3oqTI/cBWp5SPcbFlQUTKx
2/jZf+1YDQy04+lzIAh3jiUXp42vwkhp//fEfoEvncwqCJ3KzoVlTXnfDZzjI2ly
T9iBtzKQz6s7/O7t0vBvkWl7p+ycKd2OgFhgGX/1oCYrYR2J36446r8ppU7bH+3l
39V+OPrif6hV1x/Rijh+N2qEOy6ue/feDQmCefPthVf77J3rPzssOLhK2stR2N80
WnuP3371JZUD49TdD/NgKoUqpzeL7kk9gPargwOQ9rce1y4N5wvlLUHQAPxl/l/I
F4yZdN1IrxFWA6077bzpFZlcgjN1Kkz7jAWEpZTHNP2rXxIOt82napFXK4tapJbs
k4npOZAL3obPZliBz5yh5AlI98N2h+ShojBPZguDe4oIHAwKHXbATn8s/4+LcKei
7ccUYevXVJEufU2QSFMDo/d6bTfdBLnZMlj+WqPMRmzIgoRalX+cp0G3o/B0XYoq
2dqXMX5OhcDN5V+6/VzSXnRPSg3BVU/8Ze/DSAPXtqNY82EBcgWIf2UZciADoGC+
rCUtJHr8i14l2ILVq7qoRcYFCGAQCyqFBeXB8wGvEA5DsdbBvtHimkzeSsUBWaS2
YPvw/Fk21M5/b5oG56JPbdWMnqwLedDEs7m+8782LAPFpRLWpsHd3lYrfJIAr3Oy
OVlo4aHpriu1pB+R/WJdBlftfMVTXIPPIiNHMha87v8irvrnI/XaHlNaV3OMPKMy
st5NsPzR4X3aMUzMm0h02LHogCGsWUH6wC2YfVQPZQvlEXyPUL0MXfr3gUSwqQCn
I3At0idMhC5lNBr0Gf3cZwBL540509K2kAlHoUlLhEan0AeVYKEkrcFQ/+RsizlL
7WnbHBHU3BMDC099F65wCMzApRBAzOpD+YOZUsltfg1mgYkuAOgte4C6iYi+ZpOc
p0QTKkboWLtj6m+ZLGi1L139y50VtDxNrPlwWRC7wMo=
`protect END_PROTECTED
