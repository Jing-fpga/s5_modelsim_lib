`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tFfh++czIbjrnCBTNv89FAux9I8GUZVoREhfzT0pT1WjDw+A5mWe713+zHz9uXbs
tfzLIVa/DqQImRjN3Jahi7gf3r9sSHkI9BL+d+Yvzw1a07TZZsF+h8LGeZB7yxYl
c8QFo99tWlLcDpZiruzgEgLCqTiKlVFqq0JpTAzDaQEditbqkm6gKHkQTNK+ws6V
xS9IAR0XVllzvdmG7XeO5PyjkKkm64HMDu0GkQYhAtgUMU5Ley/dXWoLiV6nSgFO
de+jXp7XzbVJBcNKUtrMNW1+ycj4XlL79uPDPYTPSi8FlUCqy4vAZtPJKa2N48fv
WFrJ3HqKPhqwI1i9nX/bIgkixgaj2qMFg6nG1i8uncEb/AAcwniAgvbpsRGPu0BT
lDIcs3u7rpX/W5xwL8xR+78AG2AZRJJdJSZUAaqRnbzT2n27Rqa5iEEPPmrB5JUD
Knq8BPFrFBjPGedDYQM4Bgo+msCnPCYAX5nNYMsiwaemX5pdrEzThbzW+j2P7P49
7QR6YuBrkPN9Cc7nt5JUvC3rxucguyIdRlAIa40HrH0WRWnVteDD7TshrPnL1u5K
iZqeQ7E7NjNNUM4idQVJRwstxBO/nAiDGUyzLhUBPtqwOcAdkoke04Q8ZLDcaFqh
zBnIK5mYKFP67on/aMqqUtIcf5a0p7A2zyRkYXuVxUeoreGJIYAsNKiEeGimwKbX
FRDNbYXW3zEzGyvRzpLwqovYONtcRgaptY0dDCcVl2NncCi+bnOWnm1XWGg8HZ+J
uRewIbmbrw0w36Y296p2b/SXevqqPkBgX0ozauzMkzmbqJs/JEWI6i4L2oXctrmK
7iD6yu4C6V5S7HFPginMsRMbdH5du7oh8E0M+yVORp9nwq7xpcrBYGHmN95yztw/
K6Y6lz9BybgI9ihyXCMKNqp0AhZlfga6TCe8zCePIdaZGi7d6G6Z9/pgiyJAnWLh
2xUuq+nfc627bk7AHeKLV+0EbrV62BhMWMa2M9IX6F1K3jW7ldVuioZIUCz5UZ9o
RoZsSVVjIeAVQntGUgt4Rv0L6zLrtdNOIIUilTPKVCUm7dv5m44ojMk/d2qsE/r1
EmZoADR2+equSa/If8ZWEoXRJbxF4jiL1wd81M7XtFZDL57wD5W6NpxnEVRFbp87
ZBsdcpIwHTMQW4ZVYzxixYP18kvn56jjLCCzfKnfK9JAn+koQVexHKW5UVnKlEOr
ylTqdvuIezATHMu52JoKq5dpPmCjCynKoAoRMtdALl3TYjj/7t9MjzghnILDdHH5
BDxh/2dfMHB8JCbF8Sf1rvK4FHafjepl4hS/Jmv9rF2LIg52wB2XCAv76cNAY+XV
Tly0OVIRIOlfgf2sGuqtLOk6CbCENTQ/yVaEtDkiMTU71s04dQuCgPsXGia/Ok4D
p/Q5QPaRBAtfbETV8vveI67JWF0jJ9UkdQzNMlr294237CCFh430kgAg6IBkkCpU
52np0VvlLH+PCKUw/EqcmNRErekx19lOOJrfhuKO0DUyv2HJsEYteV/hzbxGezHr
MBm/iIm+SbLWZK7FVi+sSlOy1YVIUVH0t/1qaXQ51vcD3eqUhpT9QM68ye+sj/9v
+favDMoM1VOSH4qRICjCOCgD3o3vIrP+FcCkYQ1XWvShZ+kVdOEThGrvSqosz4x0
/5r2zjzBje45otvnwiR8ZpyhHdnFAiYdztxe3GYakUOQbYl39J2dVf0mFgEoF8us
43iyW6EOyQNyWM8EtkusQf3aJHi1a6AsKLDoJftrFubjpmR92k8G9oU9Qwvm8jbw
dHCUpnm5Ar5OAkciD8sMvMEJIPjlueZi6SKQT1Arp09Cth70d25/k1Op+MXbHvwW
uj1nH4OTZB0nZelML77+TL+W1RuNMaev60JBpO1w1t6By3FNICbNM6VBOV3WDEUk
s5rXOeVJdqYSBcT/6YketRj7sgSHhkoBFtbwnbaRTwJOgH+wYYPVA6sy6H3Kti6t
gow0o05hA/uMQUdtzDx+fwC4/ybdvl+z/w9KMGCPD1yd4rysQHbPq81pyI/PvqFc
EdqUccdNhc2W2GFNmdY/eHESmnHoKu7l4NvqX+Co0iCEQGDEB9Ws87c9Gm7fQJ6h
FoXU5MAuM/6MMYaboLGxe6QRurE/1X46GWEXR2+a0/xRlEEwvDPqGHt7WsqpW0Ov
/A9WM0fHfJKeexKQWYAHt3hkThdONtrfaCC6K4cLSPnxQUbs30SeAaeQzfl8yx55
k4rAZAWLjiRUcY8FWtb7weLXYAHYEorIQ+Q1jh8K3z7QI655N3QHGTmKcaUsX41o
q/H6LWCS5HrnGt4wGm9yZw9hIYps7W4SALjTN31+72xsCkKXy8Vn2uy+shoh/P6Q
8sIx5m9tk6SuvBi+x4SLW7yykl953XmmjB9KJQ5MDvsUd7m8s66HY/OMlpdSooZA
5buo67ryXLiKP2oMOnNrhLF36QMULt0LJaGpMUKPB+FUZjgEr5mRrh62q9AjL89X
3TeQRn5qyeTSap7Mt2DPs6DWPs5A6bo8QWca/ZnzhpaPK04H5fxij59SKlXUw41r
DJYZMBn1CvC3ypJFGmntdaaW3jT1ROn6cNUGuhBU7Glt1fod4Tlr2yGr2Hb6j7UE
Ic8UxercCh30xcazyyWN8fBOCdmBNM9mlwaDqMdCVq3sFprsuYzU/DddSsR1obPh
`protect END_PROTECTED
