`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SJkPAEv/6U1ajyjIv/ycKtEcrD0HY3Lw9auXNzTPtXc8J0HqcZinQAe9qVhGKwMR
EPNw7V+f8R99rIwkHlg9ViC80XOgvedMUm+iDlY8/8YolqEZGOYlKjuStF4SIMbi
JGmIFNyfR+bGQsU3qet8jmije4LZwTZA66QBeOjqyBTXLh+pDtCItH5qTLRL5Yoq
3NaslLApAESpTQPiIq4fazXaLlKcUBH3842BKFGM0sk23W0zf8zD3gaPDdtcPzOP
VbtdqnXsDcvCFy5qn++siXepWaZI+Sv899HUX1Tu9fA+zATvi6NM6JfmEcB0QHPp
RnjmSrt/HRWxa3amBhs+iitb2bgk/p7uYD10WMoAGmgsPaPMBmOjb0RF3+XVmiXK
ETUGJUlla6E+n8v7JUD12RSlvHH+jPnF74SQ2YFzZdrQkPnFlsvNA6NxV1KIcQLi
7e+MTZZlhcLzjZwDs2sixK+3aFjVSjKbJESnXZifk9yaFawFbtOTeJcMCgo25Spg
sUl7XQD4NhxBGyV64YCADew4sWikpiEn16BCFlqntQVLVgo+3Xz4ZsR7qAWxplQz
AOceNNQ+SkOAeK+bsQ32aE5M0vUFDS1e6/tXzMy9d1NxU1DVgIsATGxqNx/QTBne
uvLrSx5ZZ802NFJhWnfQiixYzlWj8qxDwLlqdjojOMESqlO0IivA8s1Nh286wYzD
IOjd28JB5sw7CfcZxfsyUzMUxIFnFelYD9xd+NTA3S/jM4viS1YTnmBCYFPB6k+v
CJCBaUnxRSs7IUMOC/ENu93H8kzCWzfy7SBtDc/jfepOm5ewIYRusbQOyiafn435
ZBgW7w89AcamV70jzzrZbeoiUGl3RrsSlo6tLzwUu3s/7q431hhnomgrJEam84rT
kUbyxVO33WJsGecaQ2aTL6lYu80j5Da5PBNg5FNuVIzslyUTGDqxtupbV6OTxB5P
BJuTJaHzQAngX8LKLWTvYSpscin12gPT2H+86uBl4vTe9FYfpzLLhU/Ka1PrjW98
V+ni4ga9ARb+qV7EQUqkYMwf4RAQ3quBxOCmltN5euelJ+O5zDlqNQL3CZa7Y8pz
LqS/pV+od9sw1u+kANinEpig1AJZsJK7CCz/Zxp9j/6PFPW/kx3F5QfDUZmC9ZP1
jlIh9iX1EUy9BWd1la+/VhQtuO194vDJHRrDkbWik2vbqxNObRBmcgTFCX/FSnrT
fTEiBS4PJlWrnpsAIu0pxHJ/nShkdOC6xTm9CjK9/7RxnaxuB/89x+IhEFWq+xz9
+hccK+OcQLv+/WIevLAshL1gr4npjCwaLqNou66WCIaY3k1eDvA47yC0f6GdmzQk
T+tmj7iNFkCGx/lY+cADuYwRKtgyg3kRVMioCaB2OqFvLfVL8nAPcS70D6OZk+gF
FkXbQ2e/oU0F6pjEroSn3WiHH0KmDvo9uLm2pxzl6BivBGQLlkGnKe/Ctn49TPUh
K5/QXYu8IxhlmpjDKPlAwSDhr1BfUqJ2KIx1dWFOkd/ObGq3s5DwdmiC6XaHm/qx
upyzGMpCCB5WSUKl7vES+ubT9/QTA/nclhJ4plKl1n0=
`protect END_PROTECTED
