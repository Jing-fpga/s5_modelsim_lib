`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lgGNMhLQqc5wu4kypqxbpZ2qtQXR6ISSoTW62URrD9PjqTRS5Dlv9FDa0veJU8Jq
NwmJ0PTnbfGZhQfKYZejtniTKbrePaAHRUgukFq9VDrtaBbo/MEqylZzB5br0r3u
TrNgXAc9aTwCj5qiKEw79ztRr7e4VXjS98nzIFAd4FeK48QIfR9HnEvd3IRhS0/g
HkPJBIuRRU8tC2JJz7/yPlaiyGPzOHdr+/MIcb1R3bQW6fLaMVqdtkWuUfoUy31W
ITCGUr7zOjg//9s8jzjPk5L5DEKaoyMNDkT5w4MDeqGia+fNfkTfTmP7yxklAusw
eMI1XUYR/tFqHIcVeiSs8LB9o+Z9Od3d8iV2yJeMIvNECRB9LveBg+GnZhrlFKeq
s6FubKLyf9N83YYtHRNM1rq3yl8Lv6IgAwYcuUoJQXrzK+H8eJGDF8RsNd/Gq7F5
/fN0zqEBqL6+L9Ipp4pcPhnyxduvTVLPnirESnN2/BZCwPLHDnrLFKOnBNoaZRRU
XCvrpkThoZ26EvyrYwyzO0i2Wc5jgDx1G7RnMFuYch4P0cn73ZZrAvk8dK4j5gJV
j/ZVeU77yBvL1n8HRK0bk52s5rs03KUniPuQqiklmcPglwnEqEX6Zvpk3SNcCdvi
FQJPzl9wm8S2y+5eMqiQGcezrxh/q3nxhtGLTuTHTCbYcTLgC2PyCwNOQibYj+4G
5/EV3gYpv5Pb32ygAjDISUuhubxgDe5rDK4FpgT1Ztg9nsp23qt2M6kJt43TREVT
4r+llGfA0icrDvKSh64dfRN4mIeoNpkqksVUMPK1WE2iuyAeVXMSsEtLCiR7QGYF
vpGQigDr/X7yUhIapbjJPXL0RZu28dEiwQE8+rD9zFJetb2lpJ8klv1ZFDQ6TOsB
56VsG1Dd3ATc2bl8J9l+RQHg4QqlmH+5tZIA8252owPU4UbWLxeFdgaNE8bwYeow
LxVV/7R6bL1ivRgzEVe9faDBIE7W21dAyJCBIMdUELKX+ml+F0NRPR/+jYhfhXzb
rWEGGPw0tuHGyIIw+pw5vdU4wTbD1NIFZsN7CIM8ilafT2R6XUYj9+9uzEJHWZRF
aAZ0EmNAAA4f6ynJLwEzUcspzxKQ/ma6tg+8lZOliU9v66e1JzEF4CSPh9P5ikYv
MidUdlxT5KWPh9+HTKZags49linqusKotHC2Atb3P9dvbb8p4sD1foHq4g0F89/Z
`protect END_PROTECTED
