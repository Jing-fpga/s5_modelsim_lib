`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j0VYYHfVIdfE7Gb6Y88lZvajLfQaGxpE4AIP/SzxyvQF9SrqRmdMLrJE24ENqIhZ
nbVaTVPI4+WBOQOut46iSvtGeObisFQBQdgxQC7u7WqmKRVJVQVRM8KmyLkxo9jO
skejID/QyuqaWubNlcIGhh9CiY3qjM/FcgMHndCwTx4fySmk6NPtzR/fyKqHlHNu
UvInVG+RgU1gMlC6UnBPjYGQyqrivSuJIdI9WC0yagE1yLR81hG1iqmmehVhgfU8
6phVqb6mGCwP3g6z9SC3zUlU1UB+bpP8mgc+zkSjmaMdFEYp8oaFkfBnQiz3IocQ
JVSkVsRFmV35+OykyUN1uhsO3myZ64fioGf0oUr2jrXYMl9PIFL+3liL2pXAVDOs
zRZKLg2DdgdpQPG3fZ04xkDRImFOeLPjr/wZ2gBh9QE3Oz4wTSbF5k5r+WUmmqQy
t01aMcD2CnLFRv1mu3oaqQ7KYBreJN10k9Crjy953N+zja1ijS8WBxWdfxW7dAVQ
4zaH+Ly0vMVpQ6Ynb/hR+Q==
`protect END_PROTECTED
