`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RY3YnbOFXQdcHowP9Ei+lvgAUgO2DaazAXGM7yzPQbs6+rbHufjy5uPN8SJqRsXs
dFS82w4V6wT1w2DDDpvSxl8+sSlc2qu8W552/xXvQ+xazFk/ueF1VFD1B+ZXYyi/
1Z7gEtENyGkCwRRvUiFTGSSMY9joUZsrfz1UVAhoyu08NT+cMAphh+LDg5om3y/g
UGsCYIAIC7VYL5AaAyIGje+jrGhoQZ2+lQmJCP2cu2zU+7eG3bxCriL214dnQ+Cr
dw6YgnwPLAwqvmjmA/OxSICjj25MJ2thHxJdPry5UnbZkF7xbKtvhm33b5qZvxiC
HEsRGFi7bQbjtKR8DGIxEUK1kTY+4RgoNR+7TV++HmK39SKbNE8qk6h8WjGGqayX
T7CXgA5IouzaWN55HiO+pQ2ixOGwaHik9MVjboo7OwIT30TnhAhIhYrxjSTeNfUY
w46ss/ReX8xfb66FftP6Pqzt2QsNcEgVZB52RKbYzZ5gUbdvw1zjjLRZLF8wdBsb
T1diInhplXltjA/LPtp4mK71PZj0MufRCsYnEAKBoXuaqnizMDxMkFMRof2bCX2Q
RjhnB5c9SVZljuD9D7ubPCPsqLjo4bwx3QXvt8d0io8fEM5pa9kfXuCKtk6RTkKV
o1FhNW4v+OFP9HRHjapKMipQPchq93qmaZ3DBx6cxpO3f+kYI4NrQ3Zjk66P4m/W
k3e8yMo8Y3Qcml0ADfJCsusNZbRBtmdTvg+IoPHlOx4zMEKtZTAooGkbJn+9kD6b
RGihGi9Azvlk7cgknqTyQVNDBf/VRZGJXLPiIp4ks2n10e9NFFVFiXjfnxE8XF4Q
vhxvrjjTqO3Vs9ZxzXp7a3DnO93eBQpNkS08kxpvuoTfaNdr3osHpZm55hwKyFrz
wibpux39CU/QOlUstTKDg5kiuNloUm8Z3as/C1l+8FYrr4brx0m4mtHX9Aq9Hk6O
9VBV3lggIYWo6tEWUkDKIrTtcAZvDZva6eqgsK0cqAy0xwAgi/kNTftuOvHiJfWc
NYV7IQkxJyWUE6Hn41tt2/ncyW7rK2eYDqQVUxtVhRkKSgauf3bSqm2DeC5n7avp
FexCWspZfZ3yww1mOKJ8ioxwuuu2kqiLAUrCoxIdD+racDIS1qSv3+pDcZj+ZRfD
5HEWsJt3oeyPrTjwBIOp/B1UL9ktjSuYeJL366/pQy2m8PwZxf9sAlkShEg4LXpP
G1s+2tROouQO+ib+jakgo6dCBhd0VlmRoD2FBdvpxxpTflljsyHKklAzQPQFi3Uj
tKLi2kUaAhb/nCAbWgxDkl0dfwqlHZ5icRlWel9cVLgJ16aMZuP6Hit3a1ljRxcW
BnqqItmzoTF3QsyKNTyJU+OY95qlmJRANDfQw4SqEjs7E9ooA+dxl1iX8gpRZ4u1
1ee328Qm7A+PX0bEGqOaO89ynk6ux1C1sFR8WHPK+ck32tO49hLzmAVX7AEQRgLG
RjQwq1hfAoBXi1QSwpOWOY82DOcvmud1SIVkCVE0+RbqZQlMElEHCULcoxWYIX/y
W3FQR/z1grbBZd4zPALkCTO4xmlmejhDdJ3L3HUi6ma+ar1lKI5Y5KsV178a2ixR
cu4P3igY+6LdUwiOdWzVUTxBOYSOGyWd7GcrSUF0i9/gx1Ha3nyePqDjQLLeNjFC
EXCimj5jyLGEvCr9bwcOD+GweF/ffAmZredcJrRCwTbfaJp5ew1F53bMbbHN+Cp7
0VV7AWW4X95z92cub7JPJ9eRZ7CIn4ffLwk0PSwbG0Ne+SyRKykWX9AAqpqlMKDF
qfi8TuorXbdK8Ms2Ivecaqi1tZbKx3w0EW6Ti/i79mjuf2XFPfM8csWBkfC5tfP0
nBoxSw5cCGF90y11Wm5/uH1UhpcML8TaEktZMrL1Z4PpvH/YqWNXi5BNtfpZrDqO
icysJxlYMYFFAlYmKudUxVlEU56JRqBgMfVsW1Kxsipyg1JzrnnV5x8Gh7Th63Z5
JXKNBXXEDCNfGaTrESEAuboDHBmkosdQZT80SvwOUiLhtDArA+sbIteHf1cKx6mI
Djr6TpR182txhjwa9KYvziVGGszx2l2k3zVLXQ/1ZNc=
`protect END_PROTECTED
