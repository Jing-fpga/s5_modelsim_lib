`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WZfACQiR6HvW3X9UZd8Dbc1I/u5G28M0leWBFexn0n4RP8beW9xDww8T9COb2itb
ZsBJSt1kUXfAmzn2Iw56z9qHqkSl8pkzjD94WavRxZsZVGbfu6j9QaZXR8VDty8Q
6q67pSbiv6Je3w8m2tdK91D2H1HBxgpHA3LFPuteyX8a/DIB0fOQKWHhV2wCCLBD
oxWXBbTnAJpUwylbPkgcu9/p8n0pMRbpIEY21mJUddUHfx2p8Lrp518N4sr7vqc0
5Y5YnsfP3oTWAUcMBHAIW3cF7uBJqhNAKFeiZCCg/DmR/xano5XDzNwtzKsyepl7
W931FplwA09z7f4DGAhXduOQCLOJqMcsYwADguc5vEk3m113WcT1Jwz7VKuh0E6Z
/aTNtnoy1CV5I52qo6jenZpV9rYVhJEWcNIZy0LIPNmKHxkf3Yy6XJ9VBJD0+bGI
inyr8q+w+EOjPyXJIIgWK+v6jzM//4s1yvW5YaMXEZfMG/sPTAhA6selbbkjPDW4
9ooz7OiyqOKsFbzJJOseTRw0/BMkPwLfPH63lwbXYvgXQfmixshhvAdEYmVdXYfm
CNtalyB78yU4syLLIHgwlCKT1dRfhUWi3IkqXxBa38N4T3Oxe8bV4Z31K18BQc3x
/odTbNVifYISkdsOUmvZq+ql5nIKl5dC48MOA8SDhLd1nzSGLkwMFxSPP1TfnEQC
7AiUTwivW9UQh5WtkCPaVnfbbYPktWkJVlY1dNJh8tvqWcmnZMrquCkWk0Wb9Re8
MxUCztSem6usihs2XohoZxeibIEKelvjjtpuW1mTUpurzwnxW3j+bSpA4XvA0KhB
y2zSjdprjts1AMy6rCq7bPa9tOSfr7hrxtxfaTRX99A5x02E+4BWew/p941pDwZg
wa64GHzuLgMTngJDonWV+lqLxsRBarJSSzixtW6rz6NilgU1m9F60cIUo3WAm9zt
lvnh6PUdf2Al4PlSR9wzEd7SLLCVki2GejVYhO5NCkYelew5cIIqC4/G9xMFSzQh
xdR131GgEkPhWvDblHU2cl1qQaZQ/zvGtGeyi0+dQbq/UgpvLaUn33Toooh79LDA
wHfyNMNsjxLPAEnaIRw+NblnmGagL34jDJtGKWVw3vYvFb6TgjX7n/QnTF65QbCj
Q2z/UuYI6eI9NOa2PBIv7PwWQpq8NvNHjbYX0mv411g7qayd4+7ogFmM6gyeowWc
mnMBJE8y5YjePD18erZJX15RXbyF+PyAKpOwFuL5BYuvK8v6U6Lli8DOXuOuONu0
fpSi4uZQlL3HqDR01j2rwa+shL6GbCxBEIcG3jI7tVQHpb25Lv0056UxepD84vcf
I2QVnAfzBzoABvCM9ZjiTO/FJKJwoofO9Y+/6S88iyfT2jGM9qhJODotDNBFSS7l
xwQMCGhcAcMKOCpCkWmZpJAPhxBGmjF8o6GhFzeNH4qZ5IRc17QVheW11WA4Qil0
8ocrCp0cacNSJAXJ5iv85CRLbBgvPnuA/nWL8twplFwC2ft9nVsXeBRgxAhrCleG
1DMWJyHmr1WpjATQkDdlqA3FcJNNnLoKKzNT0YHaH+GjScMY9eYL6ivuAuC6JHp3
nxu3PK4jK2kFlK9rF1IBxdSzZWLFw9m+TffOa0Mmmin1q+oX2+0JIbfmD0dMOs/h
l2qxNf/azX8pcT+Ni8sFkT7q40joRg6na7piafk9qWkhjrbya5FfgrCYOdE3hMbJ
68Hgtz7+iDmJA16JQ3pz81al4HSN1RIxv8Hmge+pmReCA/Uv9Q4UWUKynRAFg/Ye
yYJ6UvIKoD6/zs2SLE+kcVdh8uTz5otlrNXzJK0u+i3VEpPhhPa8HM9BCa1poAao
6KgHxLJAs87JrK6I0HXcs9UYcltXUGakPKHxb0+80/DLpOuWhKtuiKw52Z+vBiOO
xtNW3bnvknrwlz+DG1izg5jgo4kYHOntxL31GnMsSyrM19tsMtlsZy+YWn36ky0H
Bjx2MSvziqeGN7DDjTJVOVCE9zxe+TZhE+HLoop8TukZ0yuclQFqm2Y+sh4Y5cAM
Sw4+Mx6A7JoDIVrNRcj0/jXJ3gA/LLXTO8c7zivkMp115K/4556UnV+bLf786zGP
vICvLWnswpWYUFteVgBGWT657k4oqDU8e5GAxWTqLg0VHJgui3n5kQ6aGv8v+/+M
M9haJ4WAINiTjZxauG3t2yTfzxoyzISjR4AFbX9OMVr69HHYZ3fIcpi05DJVmb7C
07Az0x8+8epCC2Yblk9LoG6Ja8mYcs6Mp7u8a8uzROXb8ndB0al7I0h0wNuh+h9B
dFgCjCx8l5QGG1E4wdnYG6R02eLdp406Hwpnn/4h6nD7wVGpLiDcmNHKUvB9FcNQ
SfC3e3yrtrz7r4Nv+Z/3t9fnGHr+kbt1/Soi36IDoCwNpi3ePLI9N0Nxpbo0DYWP
qSKysTEXl+TEiNz8E4V1XG0fVQhKHf/KMfd+cZ+r01kNSesvH1WUH+ZErmXbDIFb
7Aj5cXGIiPAI7phq73ysqDxwb4+UMsfkdCB60ye2d75wEX9A17CFwpGoWyCbg8rU
rdSriEdt8/7+k4oXxxovVOZhVu7ueMsYs081P+y/wsoBofZyR3/IWF4Kd0oP4MgR
jjDe/lnpN6HT9+J0ek//TYyQI4IO/h4VmFzaWt3LuNNkDKo5x3zT9MFQTxDxrhpY
mzAkcQ7Y64U8x+ZT/3tge97bwkE1Ns9yJLVnWCzfmkGUlJgdpPGEfNlroWBT+XhW
wsz1VJzpxJyDgSQwfOVp1mDENfGubKWBkcEYj8g6q5G5nIdzYXMTJS6HlVMNlHQR
zIt0m7yHvn0r08KtPtUf1FW6n6hfkmM+ej31p9Y3eQgR2X14eKx3DpcI7paYo/Y0
9j50pU7kPBxYH8wKqTb+73FiOGjPf6rAIyE3VlC5x+VdLKPjaMRwAQOKij8R1zdq
xC3hfHYSl3CYL3dxPupgM2CRsFIfelFSuTeC71toNhYvnlOAtmJ7ICWmq9SDSHkt
l6hsA3ydRvlupJds5nSkDRVetONnWZLmvQup2yc62yV5W30CC5dFgcHWBdai9GDu
MCyFDQtqXkq8dt8Fh1sPp7BQHOQZ6RWv3UA2Rgn15gNBEXfyaxCkiHnotB94V9+h
g5HdkrRUtukjLWZaa0gzDcAWIC+/5w+ivf7l5Dru1ljIhQnBbYfjAxujn3T0ON1E
VPbwZ1AKG+ngDPsustq2BWYWvhazOSG4gU4YflxGDX1zf+UNY7MMjfWzmiSV8vkM
c/FcxTvFxtfCzZGgOfRkO67dn8jLJx7OfZa5FZUvE3Lj0ba+dsdzRmEeKDaBNMtn
34Wi+/2JpvECZemaXPfAgZKeMUHN3R6qHn90x8Yj+12WJ1j6AG4BYv4LEujBL1g0
aONwMJgHFta+z8u0wAF7ahKgyKW288pSAaGVEtlg9HLE1/CEYF79FsYpQsu9RGjh
dBb668/dL3yfi8152sQOJqaMvHB7zkdeTvaaAupO4US0J9FGkRbEZ4niVD5zykXO
+Ox8DaI0ewzuKYbyF03K4+AG0B/EvHypdCecPRR+uNWBK17GflCVvYu3bUbzWjSz
06h2m3KbLm3+n0yyGuagaUo6Mu3IhwN9RwGSQt5W5ifr0UrYvODHLTVaE13vV1zP
OMo7+n95Go6kJ5uMBDYa/Ba3qL9dj1bMtfa+XYwifdgfb8X4ux+eCFIxOsBOBgSb
LdHh25Wx1q78WPiJ1d/SUss2WQlyvO/Va9CHVI99ZAwcaMQFs1lfRujf89+z0gI3
Urbvj4QnKuEvHR792k3ExDWqdKSeQFGmH+0I9JLfn9vXh4WEgire80bdl0y34t6Y
ZiurPPeqfYLTEPdUp0NZJAGybEG9/rAeBm2NfJsCyaRPQc58JBFnmvDwrt5uDIe1
FNRsAyTFJbFuSc64iRCpjr1xntuooAiNLGw/Z9W529RyzKCcy/3kc/ynt6HwiUzz
KwHlLmL5wwOxp/E+f8Uq97ncCuvD2LEJDCcgtQPVSkGoFCFdCfp3pcrB6Y9jv1iG
7GUO7sgYu0MVkcBjSZeU6vZ+00fQT6zcB6N6+6GFX4AX6z/VSSTQtQFttkVaX7lQ
roKAxXtzvhE0iOUZUp3ZsovxPhsBSZgBU6ict4ywk6vlXPkXWNy+xz5ZCmPxefby
t/cZ7Y01qoyHR8R0yWy/oEuAU30fG/P6R5PA/S9YpAv3EEjtj+mxJzia+eRcxFaF
1PC5v9SIlluLtBfqx3kX+Rw0BC675dyP4cXFsSu2gE2hN5xFRgsDUxAFL1gt/Sc8
0mvSe1bfM2mhaOHQq3SWzcfwDGo68bG/M0c7XSvQkZJflziTPXkqI9XTZLo5EtA9
19duxtJdtqnnod5KzTfNPvAaBIlow9+/o5vP55bLQOVLOEHR2queIB0QrSpN8gBp
2FDxexoX2dxStkkJETcsQBLlnvEszveyCiSu2r4rSuHtqv7AStwMDCg/7R4bjlvB
ExID1KvfaXO/pklCTC5jZtC+ujJ3bgE2+iy8wDARXJAKj4L+5M4joAsOcwSnz2J1
yZvBbG8bBiEz1oaMSdefWwyTi7jnB1x/UVy/RFgQAjcKGFhxAzBONpFvK6B36SQL
fs0d53soKjA9d5rxFMnFlGxCf5abhn2e5J3PMJiWW+jjGdGMr472jWmZ8m+DddJC
Ap4vXEDuWDlMP0rxDZvEqaOZk+HXgoG2ZBUrONhV7uJl5rZfx3wylhFT29m6BFdc
nG0sdzYKDFHlf/ArbaBbVR35YmsyZ1fxyKEISaglYeV1W+eh1GOlymMK6582JxgG
xMhwlz68kPO6lbEGLvgNJQZ94dX9iUFEntSH5EuPq3ueB/xp0jVEYeXfDKOHZMRX
U6sumTgoazimDxIfWSXtIdZzGsl3iTh8wxA3+axpyuBTGe74drvF62EF7Co2CiCi
NHofwIFA1A9mMI7A0O9/+M0hMGidg6CjeEpOfDqmH8mXT/BM/WZmK1cr+Sd0p/c/
Blv857Cl2Kd2WoY4hFa+td/I03lvkSz+NylGk/rbFR6d0sA6jj0enq0TcKdJjM7G
bg3xKITaf/lM1EDZhX2jrToozK3SFGcpZxLsclP+oT2zj9a23si/QEsjgmoa7VMc
ZPOIf3ykghgxLcwjqEXTWniklkiX1R73N17DpiFI8rfIslS2CBZK7bvrsPrwCkgS
kRQF/9Zbmppg3h2/42d1oorwUn7i8QJ+wPCWiCW1RipJPWtWI3HX0AG/YtVjVLmw
mr8vaZ7IZy1tXd4L2mYdVFcdVVAug8s3TfYW3sz1Q/QoUVHK4t9qgYxObMrNn4ZH
8cUkRiXgVAQek1VLhhf4yMvwWnE25dtkiz3NRrzZREBnCQXWeblWJTiw2URdvlrm
7bd+nD/UwKrF7MUOOQIojDv/dU+zFdSIF1vDBcHyPhXhC+LElRL6uPgwJ1qdijZi
AekQsqjTsC+oH8S55NR6UajFn3OGc1GsDc5sWc+ZzoI=
`protect END_PROTECTED
