`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WrUhbiG/961Cwc9NWZ2+znpHGZY6JtTP9xSpKzaz3Mtgz7BMDcUY2S/JoA2ENWpa
f9yEYg2khQKxSqw50IGcTnJ4OQ0XFBpcyLSGBb477ZcEuxKp6dFWzjwEBPUyDr+0
t5Pbtfj3Kit/+nv8dBN9r2bGZlU0KFjjoCASa2rANMDMjqrxcD4zlM+KTVQapXnI
tRNsfiynSDte/362MBSSr3beplUKMlkK/c9ANalOVn60ZMCjcT7bOrZ7M0k5c1kM
HkvrcTc/pjMc0JoY/YAHjPpjyK1iY1dyYGgd6KzxV2aM8z3mzSpETlymVXCjH9jo
7RnKnrM6HSb7BFRiIlBG+L4BdMKv3UdNgP0BsYt+B69keqzztGGVCwUl8sbdjKXD
WYjGeURzOGMfbsQk03KSS7mxrnzDL8UzPQkZtmTLPp0BqM8OOvsG0XYw+Yq5070B
Yu7s41X/wemjxpjPduwIwcf0cPcoS30LYPw6AvYqfEd/1H6DqiaL3XgQkDPVD1Ck
hIVYxVUy5QyEYF7WNyqTk9o1cd0tOuRZJDOOjb1BI4Y1HU91SZdXsowV/onrorEN
nywkAUTTKRbMaCrfYwiMgWNF+B/nf2Esc+AujJJnJAkkxqk6vLDT3WH+gFWrKe58
bTNjJIav/aUD3ZC0o1T90ya6lF1Pt8AFRegby/8dESuzKQFSDCfdUFMdtcH3Z6bZ
KL1dz8Teffh+5PRBr16SLynsneB1s6RnhqKNGMuf1E9xxyFgiJBskGIdl2fjk9T1
B4Vej7YyLpNBNnxmcRZDUsEY3pLTKpztk7HvX572TWs=
`protect END_PROTECTED
