`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6JneaAh3hzKh6v9wQ61w8WdDDS0igeBvtX9bZ4Td1ThnaRHRIfVoZznNML/YoFAq
5WCJ63cnRNgt4koXZCa+cXJcD5sddEHBTD1PM2WEkkDWbdw7sr64TdsqeH+Xg1v8
ex/LWGEo2LXtpqE+lMkIUvJMiprnZeugo94UesgNbki86tIMBb9kxZ/WxgI1pXoy
SLRVLn7t07BRi2M2Wutvz44kYMo4h523nlfWiBbI58ekpFBvAgU8YiGhkYi3unCO
xUalEGzCU9tvt5J8r8xAmpeXK5yDDN7oWIvo1WvyLCOLKbz9JzVSuqusuFis+VGP
D6IdOcnL/Gvh4ecqJ20EQr5OKH555XVCy2BuZQyYgjmJiYM4AFf9DblSVxz6KKia
O/+XfXnPOPaNDU//NaaSRzxXEwkb0Y1HTDWE+dpFeqJQj8dpooAMm8Cughvsnz6H
`protect END_PROTECTED
