`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x3lemTn0J/HW2tPHgUDXLcN1FT7mUyPPoR5D1JaL1kdQr8zdQzetgUOPS5xUp2Kp
3iCfPcSoPbLeY0uBZ7q1a0e3hJBfPtXG+QkL5lpAJzBvIQ18GcXfEc1PmhNiTtyV
NN3W73/ofLgiUFtVhjYcT2TCxQYyP57+JaTNjA/DLGqaW03AcwElpEmKq5i7jjH4
li9AroKGcinWmh/kSchlHyJy3RbGVkyg7PjpAcx1lyPdgqcgDE5Mk6o3IO7wV/mq
S5UiARFFBonHgorTfTm4brR0X0v3qeOANMr9uypwU3e/JtMP4jHmS4E4Hmutj3JI
POXWc74Zlw8tbnf6PAq8UXUzZFymInkIyGrVXHm/emJn5ZDEnPq+DKCFHAXHNODE
k9l+n9K9Z+hYF6OgiljlH3skUAH/JWg1pggAlLFjRwd3nN9yCVXJuD59BX7MypCW
UTlEH4GpUpPefaePZ4OdSHCmYNcGfWeb8K1Ew4hJ1e9lJki+TGbIoYtFjnU8ZEki
cp/wtVVCedz+JFEYT8NLySGuMRK7b3EgbTA00U6f5Ie8czfh3iSlHhdWmS50XOpB
xuSWtZT9yg2BCuH6s14dTYZ8E4fj/gmKCZ8q9Z9CuqpjlsX4duFoP10ENTU1R2kv
ngLsj0lHX3GZVV+kaOxYhsY4TAHgiFwgFxgoHbcfRHbk0m6ks5tzJx19uPPpaLQv
P87y2ghSmcFf91lJNW8vqf5PExHIdM/2tFh121G27VlttlpV2T0gFVkJPEOaTUiG
tWK/CGBfYt1ES4u2o7tSmCVc6r65PHXavH0lfVasaEiMwxfqknjPi6n/Z/n4JWNn
vMChSFb3Iay17Qi69wDvdncPxsreBHVMVDtahFot2Vs8Ch28U9lQrwViaU0cvZXh
s87UaH76ffLXPPt81DWptZQDxmVwZ2H7fTffKkwGaH0f0HM+A6al10zkUHBm68W5
BTfK0d7LYuDHnQPG/HfImB5BAkzVbMYaRkyxJpBFsLw8BJ6CD6pMdP02jZc6vgzz
1K437LoMzQShkvowZ3CHmqHf9Qqrkv3SiSs1VEjF7rzsnL/OxBlmHwI9tn2dx0rE
N9V8LHV1jDaeWPxo3CieAFHL99cNgMulUvpwRFPEQbTc5BXtNN1wUFApDlFvBr/8
FGW/0h05jbRMc9ooulBDS5Yoz2hTXUrsFPG0r9rsmUj8nHLe7TeXVdJx2TyLs7FQ
8klxy0iHwjlBKXNIQALe1kW4eVN8VqX3uaddJfPPBevIZUtKe0sQxoST78fQVdql
msmeS7MboGIx+6abDFgtufVcDboy/toIb2hMFg/CH5Cz9QlPDzeUmi4iUaQM70Qo
64UHOMkdw+IWCmQsTgbIqe6kN6kTFKkobB1A7q3DHfu2fmaHIX03gj3sHoePib5q
wSFs/lWeg3tfRxC1CTu+l4PtEAMGmPU79faZeHwBlUzrh+M2I/vcETk2DTGV6FEr
`protect END_PROTECTED
