`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ora47qhirNmOR9UKHa81JbEs80UE3G5kpq5Pw0mY9QjqYStbt3Sp7tVmfApIvM7N
e7ftahG55gk81CSU4zIHTWiUr7Dqka0pgrsg3Tcr9YXKkfLlLEjTRaq/JBUH7hPJ
LcAHyRG0Ip9hg5kkQ2jpC0SqZq9gYECCSayoXgDNhJyE0JXtr7bih1XaD92g/+pX
tyDPWY4cP7MAK2tQN8leZEY59uMOCBUzgjB8uAEGOB7DwbdAbHaCpfFCFXKbxqld
9Vd1b/o+ywMSBJ9tzcMCTR4689s3JkqJeLBmoGs958064jfQAxgw0Eng4we0pOHi
we8/kn+3MdfBd5dOwTbFowynZ/XakmebKAXi3wV3zNqt8A062HSkJApFon4/mrmB
eBrsNFT68H9rbTQf1GVn9UexGsepyNoixSuI42CrLO9610VJ++uVoxoblovkJkts
pe1Spm6hmRY97kCPud1wIYL1qBmh257oMKTcXEctZ+QQvfcLIpdD/riaO0HK6PXu
1MJpnD9ZPLltCRl0jk0PYIPJDzNlkThaN7uZfVxJwV8GNIIQ45J77AJOVujcehux
R+25b2zTGWCGlAo+HeQ4xSAfEssAxMKbRfLlb0RUWlm71kgjkyrSKbEOQKIB6aBz
0AMNRrIRppkpWgBTBymOqrE95XPOn3RBB6wmObuYgg3b2C7/BqIRpMDAg8fnGqeW
5Y7KCY0HjPJJqHfpMhxNSvZ2h1Vyc8Lelrd71UosV+2fK5k63gQ+mJGPqw5aNCbO
y1EzSbV1PR1hG8TzCDkUaYk9SE4qFBdp1qhmq6W2qQKFfxItzh9hSf2xrvKrOkON
5h1nTE/BjpPPCjdmjZZtFpmfibxay0SgPE7cADdwHYBsnpRDavGIlnTzK6fKFDR8
jjJkPtgwhaRN2/NJxEWea/99WhmU4RX9/CuNZJkgP3Eaueiy44p+wAPqa5mag6aY
EHN2YdzRkJiWLrAPL53ap2UYeIsbXWORWA8uY4GCv9L+rNhquN/R9ZinVDEx3wqj
m5M7Su3RML2Dst5UWyn8nx8hxglLMq4WR9PFToTPfXmJldzYjasH8woO5D8hxd1p
4++bRA/BD3P5j7dxPdCT65uXLttVaWJ3lgj9xbr5UoHkhllG3i9aNxx2ME3lnEYB
qedYvL2zvVH8hGc1krsXu6WrzQNikBL7iCN/E5U88xLz9FYYide1V4T8ERVhRBKE
KR1JbAFixjoqcoSi2d4yoeoAxpzoHwv38a/tya2udIMcJ5uZBxQksNC2NHJaHOt7
GaoAfm2HD5DWCVo1GNzv9xNRNJF5WuLNODHcQs9D1Etn3MB8EyMQTm6now1/ZKd7
CWZYNXrceU4FMA5FWLtwx694QRDKKKanM7snxxWu9h9VtosuqXEj8Va2lCKV7hgm
XLXlcTD493GrZoEv6eaVfXWeqQhf2vlQQpNIYCkKR4HGTf+Ix+rHVt1WhyvvQlPb
y0BYNRiOPdcLvBlpnGgE6K8s8G9nHgn/MWYvO8CtrLfffq+2r/nuLyQGNkw6VPoV
AduCZbTVnccfkV0ZMPlqJ7kyLgcwLEcMaQZTeBhQIj4kRoePkiFhMKcNJn0hu+x9
30gIXBkWRrVQRWy8/o3G8PjfaHRcRlH6Mk5ZfILuwjgR1Jcp5bukT28omPM53ncm
PYszN0LpE23EtzKiYKrLZpN6ijjxeVwcxNY0h1s/DUQnLbUFjtl2bMupuSw+r4v5
KdaXuiuWuJrnZKGMlkw0rTqJE3Pd0QEgcg0SRleSY0Zsyasu67JssQjKE2c2FG+E
0xYFfCsZABJs0OYaf6aihf070fCaNhGJUYkiaFgl3bZJJo/3GRsHLyvxwHny26pv
TLV4RlB2ID+xaWt0vWDVscr1eviJ8FRgWcPKohySXV6hvZ6L8ZqA3MV1zhIkKF4W
0eh/ton4R7a+H1wfIRuPq5GBMRa/yTwLR0JVOVd6bEOGhgs28eH1iT4r9Iqsfj06
hYQeKmrv9wH5WC6sKzQbhzkPFFFCXmNgVHB5OiWXA6AmTRyojeuf9Pccx09MDWnD
F+zSeDcxpeU8B0cuWexluek6IhLx+0zKV8yevsveN199ocR/zbnT1SmkdGiZ9kLz
0QiTJhpzYaWjz/8qiFPrpRUKPv5pPFq1yQ/dJAo2H0sBYQKn10kjOBYqDLlpSUs9
SwS6iddd/K2VAVzs33ZBUV2BeqhcjODFzOjCiXig8ARbht7hX4PNXJQMdlEI4iFh
dLCDbr4/VuYgR12XaKrjJazEJdVuEwYLvLsiOAy3QWLlO8VF0ikp/HyL0MkZW681
huwGuxOxUmRZqq+99wGt7u8IAtfgomLcS96cX2QaIg1B2RH2uiEgHH6ZpHkphF0K
KuJF/TexCsaxfYA4uZDuj8J7QeG6ZZg5RWkY38ncHPPoK3cPP3hdwoHzgz9MYpnB
p6SxxzBvhcAwx65oMRzmef2NQ8LovUZ5qq2KE+CBgan1YpR9zSrx1GfInaSgJh1q
ACmhkO5mrtgXxrjAARbMO3mDYUdwAbyNxfeoUlgcE/YQvRcUaqpd02nU4huIzRT8
ejL3Yp2lS9L1g3Tf8LVatvqsQ2XYntInZpgTqKwsa3iH32BnbF8gOxNxQLVxM9BU
20a0ysfCKGVovfFi7L4zEp4ezdXDzjaaXyZBUgU+9mtVFAURi5DucFPYzj5PBUYE
JdCEm1QG/qjEdF9pUgioQi0lTxSinvJHt9eAupeJueBQFV0TtZa+gGCyDtKS9LqR
XsaVYu5Lj91OKBHfgXSc3QeUJVyBNacAgDOWX5K6J73oi6xcrNd3NBkqyT3x8URZ
nBMHffepnwFluqgmI/Xl4A==
`protect END_PROTECTED
