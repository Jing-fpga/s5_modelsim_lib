`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qnyUJtqMTs4myVMrXxOlJH5k3HfE1zjSlbAvJCa2jvC10FiDw9mwM3x+bU35E1Uy
oYUwWoZm5E9rzP+yCZLQzBqtcGuylwONgJ8Dv943INIi64SVCfTK+Hoiw4xXIKrS
18ZSooCF/oW78u5pKdbQjhg2WD9KqtuAKHsYPnGuStdkDyaoT4AFlOIUg3xt8tQO
3xw54eJkle0aDQbVQh99OqMp+safXEHdgJruAF0OWxP7fc1/UaCy3TN1HxRmCMUO
sjJpC7g+mcMiZPQfG4PVaDFcOmhN1WY5rK5fVGtGO+Yqw6IpB1F1Q52QE2d5fhRR
gt9mXqLzheRD6jkadSBHhvsMb9lApfqRX5voYhNLGSj8Otura6yxOVeVf2TPuHRA
iDGwnlx1gg6GqaKBDFvmdyQg+ePYx304UOGBpM6NlynoJX5N8i9vwTBawk5c8CBJ
z0aOtG/d9jbcCznP/pR3Sdg+ErUeW5H7OAdJxdnlUHIo12sLHeJI/8+u4nivF8gu
KgDNpJHEUXAkt216EEpjVg==
`protect END_PROTECTED
