library verilog;
use verilog.vl_types.all;
entity stratixv_hssi_rx_pld_pcs_interface is
    generic(
        user_base_address: integer := 0;
        data_source     : string  := "pld";
        is_10g_0ppm     : string  := "false";
        avmm_group_channel_index: integer := 0;
        selectpcs       : string  := "eight_g_pcs";
        use_default_base_address: string  := "true";
        is_8g_0ppm      : string  := "false";
        silicon_rev     : string  := "reve"
    );
    port(
        asynchdatain    : out    vl_logic_vector(0 downto 0);
        avmmaddress     : in     vl_logic_vector(10 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        blockselect     : out    vl_logic_vector(0 downto 0);
        clockinfrom10gpcs: in     vl_logic_vector(0 downto 0);
        clockinfrom8gpcs: in     vl_logic_vector(0 downto 0);
        datainfrom10gpcs: in     vl_logic_vector(63 downto 0);
        datainfrom8gpcs : in     vl_logic_vector(63 downto 0);
        dataouttopld    : out    vl_logic_vector(63 downto 0);
        emsipenablediocsrrdydly: in     vl_logic_vector(0 downto 0);
        emsiprxclkin    : in     vl_logic_vector(2 downto 0);
        emsiprxclkout   : out    vl_logic_vector(2 downto 0);
        emsiprxin       : in     vl_logic_vector(19 downto 0);
        emsiprxout      : out    vl_logic_vector(128 downto 0);
        emsiprxspecialin: in     vl_logic_vector(12 downto 0);
        emsiprxspecialout: out    vl_logic_vector(15 downto 0);
        pcs10grxalignclr: out    vl_logic_vector(0 downto 0);
        pcs10grxalignen : out    vl_logic_vector(0 downto 0);
        pcs10grxalignval: in     vl_logic_vector(0 downto 0);
        pcs10grxbitslip : out    vl_logic_vector(0 downto 0);
        pcs10grxblklock : in     vl_logic_vector(0 downto 0);
        pcs10grxclrbercount: out    vl_logic_vector(0 downto 0);
        pcs10grxclrerrblkcnt: out    vl_logic_vector(0 downto 0);
        pcs10grxcontrol : in     vl_logic_vector(9 downto 0);
        pcs10grxcrc32err: in     vl_logic_vector(0 downto 0);
        pcs10grxdatavalid: in     vl_logic_vector(0 downto 0);
        pcs10grxdiagerr : in     vl_logic_vector(0 downto 0);
        pcs10grxdiagstatus: in     vl_logic_vector(1 downto 0);
        pcs10grxdispclr : out    vl_logic_vector(0 downto 0);
        pcs10grxempty   : in     vl_logic_vector(0 downto 0);
        pcs10grxfifodel : in     vl_logic_vector(0 downto 0);
        pcs10grxfifoinsert: in     vl_logic_vector(0 downto 0);
        pcs10grxframelock: in     vl_logic_vector(0 downto 0);
        pcs10grxhiber   : in     vl_logic_vector(0 downto 0);
        pcs10grxmfrmerr : in     vl_logic_vector(0 downto 0);
        pcs10grxoflwerr : in     vl_logic_vector(0 downto 0);
        pcs10grxpempty  : in     vl_logic_vector(0 downto 0);
        pcs10grxpfull   : in     vl_logic_vector(0 downto 0);
        pcs10grxpldclk  : out    vl_logic_vector(0 downto 0);
        pcs10grxpldrstn : out    vl_logic_vector(0 downto 0);
        pcs10grxprbserr : in     vl_logic_vector(0 downto 0);
        pcs10grxprbserrclr: out    vl_logic_vector(0 downto 0);
        pcs10grxpyldins : in     vl_logic_vector(0 downto 0);
        pcs10grxrden    : out    vl_logic_vector(0 downto 0);
        pcs10grxrdnegsts: in     vl_logic_vector(0 downto 0);
        pcs10grxrdpossts: in     vl_logic_vector(0 downto 0);
        pcs10grxrxframe : in     vl_logic_vector(0 downto 0);
        pcs10grxscrmerr : in     vl_logic_vector(0 downto 0);
        pcs10grxsherr   : in     vl_logic_vector(0 downto 0);
        pcs10grxskiperr : in     vl_logic_vector(0 downto 0);
        pcs10grxskipins : in     vl_logic_vector(0 downto 0);
        pcs10grxsyncerr : in     vl_logic_vector(0 downto 0);
        pcs8ga1a2k1k2flag: in     vl_logic_vector(3 downto 0);
        pcs8ga1a2size   : out    vl_logic_vector(0 downto 0);
        pcs8galignstatus: in     vl_logic_vector(0 downto 0);
        pcs8gbistdone   : in     vl_logic_vector(0 downto 0);
        pcs8gbisterr    : in     vl_logic_vector(0 downto 0);
        pcs8gbitlocreven: out    vl_logic_vector(0 downto 0);
        pcs8gbitslip    : out    vl_logic_vector(0 downto 0);
        pcs8gbyteordflag: in     vl_logic_vector(0 downto 0);
        pcs8gbytereven  : out    vl_logic_vector(0 downto 0);
        pcs8gbytordpld  : out    vl_logic_vector(0 downto 0);
        pcs8gcmpfifourst: out    vl_logic_vector(0 downto 0);
        pcs8gemptyrmf   : in     vl_logic_vector(0 downto 0);
        pcs8gemptyrx    : in     vl_logic_vector(0 downto 0);
        pcs8gencdt      : out    vl_logic_vector(0 downto 0);
        pcs8gfullrmf    : in     vl_logic_vector(0 downto 0);
        pcs8gfullrx     : in     vl_logic_vector(0 downto 0);
        pcs8gphfifourstrx: out    vl_logic_vector(0 downto 0);
        pcs8gphystatus  : in     vl_logic_vector(0 downto 0);
        pcs8gpldrxclk   : out    vl_logic_vector(0 downto 0);
        pcs8gpolinvrx   : out    vl_logic_vector(0 downto 0);
        pcs8grdenablermf: out    vl_logic_vector(0 downto 0);
        pcs8grdenablerx : out    vl_logic_vector(0 downto 0);
        pcs8grlvlt      : in     vl_logic_vector(0 downto 0);
        pcs8grxblkstart : in     vl_logic_vector(3 downto 0);
        pcs8grxdatavalid: in     vl_logic_vector(3 downto 0);
        pcs8grxelecidle : in     vl_logic_vector(0 downto 0);
        pcs8grxstatus   : in     vl_logic_vector(2 downto 0);
        pcs8grxsynchdr  : in     vl_logic_vector(1 downto 0);
        pcs8grxurstpcs  : out    vl_logic_vector(0 downto 0);
        pcs8grxvalid    : in     vl_logic_vector(0 downto 0);
        pcs8gsignaldetectout: in     vl_logic_vector(0 downto 0);
        pcs8gsyncsmenoutput: out    vl_logic_vector(0 downto 0);
        pcs8gwaboundary : in     vl_logic_vector(4 downto 0);
        pcs8gwrdisablerx: out    vl_logic_vector(0 downto 0);
        pcs8gwrenablermf: out    vl_logic_vector(0 downto 0);
        pcsgen3rxrst    : out    vl_logic_vector(0 downto 0);
        pcsgen3rxrstn   : out    vl_logic_vector(0 downto 0);
        pcsgen3rxupdatefc: out    vl_logic_vector(0 downto 0);
        pcsgen3syncsmen : out    vl_logic_vector(0 downto 0);
        pld10grxalignclr: in     vl_logic_vector(0 downto 0);
        pld10grxalignen : in     vl_logic_vector(0 downto 0);
        pld10grxalignval: out    vl_logic_vector(0 downto 0);
        pld10grxbitslip : in     vl_logic_vector(0 downto 0);
        pld10grxblklock : out    vl_logic_vector(0 downto 0);
        pld10grxclkout  : out    vl_logic_vector(0 downto 0);
        pld10grxclrbercount: in     vl_logic_vector(0 downto 0);
        pld10grxclrerrblkcnt: in     vl_logic_vector(0 downto 0);
        pld10grxcontrol : out    vl_logic_vector(9 downto 0);
        pld10grxcrc32err: out    vl_logic_vector(0 downto 0);
        pld10grxdatavalid: out    vl_logic_vector(0 downto 0);
        pld10grxdiagerr : out    vl_logic_vector(0 downto 0);
        pld10grxdiagstatus: out    vl_logic_vector(1 downto 0);
        pld10grxdispclr : in     vl_logic_vector(0 downto 0);
        pld10grxempty   : out    vl_logic_vector(0 downto 0);
        pld10grxfifodel : out    vl_logic_vector(0 downto 0);
        pld10grxfifoinsert: out    vl_logic_vector(0 downto 0);
        pld10grxframelock: out    vl_logic_vector(0 downto 0);
        pld10grxhiber   : out    vl_logic_vector(0 downto 0);
        pld10grxmfrmerr : out    vl_logic_vector(0 downto 0);
        pld10grxoflwerr : out    vl_logic_vector(0 downto 0);
        pld10grxpempty  : out    vl_logic_vector(0 downto 0);
        pld10grxpfull   : out    vl_logic_vector(0 downto 0);
        pld10grxpldclk  : in     vl_logic_vector(0 downto 0);
        pld10grxpldrstn : in     vl_logic_vector(0 downto 0);
        pld10grxprbserr : out    vl_logic_vector(0 downto 0);
        pld10grxprbserrclr: in     vl_logic_vector(0 downto 0);
        pld10grxpyldins : out    vl_logic_vector(0 downto 0);
        pld10grxrden    : in     vl_logic_vector(0 downto 0);
        pld10grxrdnegsts: out    vl_logic_vector(0 downto 0);
        pld10grxrdpossts: out    vl_logic_vector(0 downto 0);
        pld10grxrxframe : out    vl_logic_vector(0 downto 0);
        pld10grxscrmerr : out    vl_logic_vector(0 downto 0);
        pld10grxsherr   : out    vl_logic_vector(0 downto 0);
        pld10grxskiperr : out    vl_logic_vector(0 downto 0);
        pld10grxskipins : out    vl_logic_vector(0 downto 0);
        pld10grxsyncerr : out    vl_logic_vector(0 downto 0);
        pld8ga1a2k1k2flag: out    vl_logic_vector(3 downto 0);
        pld8ga1a2size   : in     vl_logic_vector(0 downto 0);
        pld8galignstatus: out    vl_logic_vector(0 downto 0);
        pld8gbistdone   : out    vl_logic_vector(0 downto 0);
        pld8gbisterr    : out    vl_logic_vector(0 downto 0);
        pld8gbitlocreven: in     vl_logic_vector(0 downto 0);
        pld8gbitslip    : in     vl_logic_vector(0 downto 0);
        pld8gbyteordflag: out    vl_logic_vector(0 downto 0);
        pld8gbytereven  : in     vl_logic_vector(0 downto 0);
        pld8gbytordpld  : in     vl_logic_vector(0 downto 0);
        pld8gcmpfifourstn: in     vl_logic_vector(0 downto 0);
        pld8gemptyrmf   : out    vl_logic_vector(0 downto 0);
        pld8gemptyrx    : out    vl_logic_vector(0 downto 0);
        pld8gencdt      : in     vl_logic_vector(0 downto 0);
        pld8gfullrmf    : out    vl_logic_vector(0 downto 0);
        pld8gfullrx     : out    vl_logic_vector(0 downto 0);
        pld8gphfifourstrxn: in     vl_logic_vector(0 downto 0);
        pld8gpldrxclk   : in     vl_logic_vector(0 downto 0);
        pld8gpolinvrx   : in     vl_logic_vector(0 downto 0);
        pld8grdenablermf: in     vl_logic_vector(0 downto 0);
        pld8grdenablerx : in     vl_logic_vector(0 downto 0);
        pld8grlvlt      : out    vl_logic_vector(0 downto 0);
        pld8grxblkstart : out    vl_logic_vector(3 downto 0);
        pld8grxclkout   : out    vl_logic_vector(0 downto 0);
        pld8grxdatavalid: out    vl_logic_vector(3 downto 0);
        pld8grxsynchdr  : out    vl_logic_vector(1 downto 0);
        pld8grxurstpcsn : in     vl_logic_vector(0 downto 0);
        pld8gsignaldetectout: out    vl_logic_vector(0 downto 0);
        pld8gsyncsmeninput: in     vl_logic_vector(0 downto 0);
        pld8gwaboundary : out    vl_logic_vector(4 downto 0);
        pld8gwrdisablerx: in     vl_logic_vector(0 downto 0);
        pld8gwrenablermf: in     vl_logic_vector(0 downto 0);
        pldclkdiv33txorrx: out    vl_logic_vector(0 downto 0);
        pldgen3rxrstn   : in     vl_logic_vector(0 downto 0);
        pldgen3rxupdatefc: in     vl_logic_vector(0 downto 0);
        pldrxclkslipin  : in     vl_logic_vector(0 downto 0);
        pldrxclkslipout : out    vl_logic_vector(0 downto 0);
        pldrxiqclkout   : out    vl_logic_vector(0 downto 0);
        pldrxpmarstbin  : in     vl_logic_vector(0 downto 0);
        pldrxpmarstbout : out    vl_logic_vector(0 downto 0);
        pmaclkdiv33txorrx: in     vl_logic_vector(0 downto 0);
        pmarxplllock    : in     vl_logic_vector(0 downto 0);
        reset           : out    vl_logic_vector(0 downto 0);
        rstsel          : in     vl_logic_vector(0 downto 0);
        usrrstsel       : in     vl_logic_vector(0 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of user_base_address : constant is 1;
    attribute mti_svvh_generic_type of data_source : constant is 1;
    attribute mti_svvh_generic_type of is_10g_0ppm : constant is 1;
    attribute mti_svvh_generic_type of avmm_group_channel_index : constant is 1;
    attribute mti_svvh_generic_type of selectpcs : constant is 1;
    attribute mti_svvh_generic_type of use_default_base_address : constant is 1;
    attribute mti_svvh_generic_type of is_8g_0ppm : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
end stratixv_hssi_rx_pld_pcs_interface;
