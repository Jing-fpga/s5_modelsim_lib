`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ql4GCqId/5wkrp1Yrkb5GshvaaBplm4zmibPgAVDx0bG8RqG1K4jbn/5mX9mk8p6
g4I95m7nk2QZD8bh6pK/RTQAfo3fqPiJgPo/e8VfyzcJ+XpslVZcivd5zhQIYVGT
pH2W40nKQkGqTfsCdXxH1bL8wkPjamnzLWqDT8XkoDNMc4wsYkZG93s+vUH6nwGH
FeuWkni5WHtIlLjIjTy5FyaL+sNlCqyz7AX0pG9TugvnFCqPRrc9H0jLTHeV23+d
zNDZNRR6jYt1f16KEhYfstDxAkVJXHG/Erx99XuHu/Jh2YLSmxPfjkOw7b5XiQBH
yEeHKDK/tEARdYAsZmgg+2+mX5G5TglOdcB7cC8XQ7WJFRWxPLnR47tYTWk2VRC3
ZAITuxijlLIgAicQEgOixVm0mJDtZN4AOxmZnQrq2v6EFq0YH2Tu9uf6qee0cEbd
Oi1ENKfWvtYj1bQ8Pj5Aot2tplc4T0ZKOnGoi15/KAUrrXAn2SFkH+NVbCKzi/dw
Z4lJ1xySghTl8kvuHUQAng==
`protect END_PROTECTED
