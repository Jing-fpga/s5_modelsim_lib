`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XEo6nA9J18oUnSoZxowfcZFGkJgl+tELYF7f3FsxzutHlEXTaT+PvbVMu5f1zdX6
JS4kFWLDERoE4kOBPppxtturiCz0gnFsGKR0g0/wvDJ/2GzsrTp6TyJo6UmjjtAF
XuGhGsolnIChqf5ZLY8mAIL4mweO5f2SPHKAF8l5t69ByfUIYThIGomyyWcU1Hjp
BwgjsrYAH/eMBrh04q2aS4YVO94B9Bvybz7WNYe8rbLLjIO6N+3j2Xw9rAJ1GFIo
D1Vky9/PSQyu7+A6voNx9iVs2y2zDVQKMg3T6CDPVDj7p+TGUiKWpa1GFxHT6dZT
63r3MkKsulRISctZjm/QlyoTCebBeO6XTmVb9N6oWrPHjXpR0YJeqFJbHi1SsQ6C
skPo5M9G1cqFYuBqCE6NWXmyJttB1L2glcre7IyjpAu996cab+q0JgXOiEAMaNVa
rRO9E4PzKsnlRB4LQ3kHUigDlYt9HQ1PvPEGJFH+oJFXkGiXPMOJdR2O99rON4If
zq9apYKogl4ZyLtuC/JZEtmMeLbVTu41/FVnTQjAT0osRMOO1mhOaNwc2/mZq1PC
8q4n1YHEduLnIB7cG6ukqp7qEWeLQ2htQUgpssbQwqlpse8WbmIZmZC1Xk9fS/zd
UeN83m0T4fy+urLYPZLMUNS7hWD1rVIBUHSpxyQn9MBpOFP9Cslbko7nbDNnSzNm
4YFMXNObL9BKZRd5SUs3HKqRFScEErXjebu/9I/pM09AE7Jqji7SeSOXI3jX/EaZ
FYRUp+Ttyc2SaTLtEnQVkct4zHvIn2nmBXzuzkFFoAzXhvxS0tdj/dqHNtGWA70S
x/grzg+N7BMZ4rIxtifVaJ7D5TbHuAfm1tEEL9FYeJabBbQnPkhmZrTXYD95scXx
HLPUIO8RuxoLUvViL7nqJRijcLM3BaJPNIbMJ2/YoQMYc9CfRPK6PDRXtAE4EeM0
rXWpMYDegnb2Ux8VwRiHL5R+nanWivmXe5gktKp2rdR9u7dWo6ntiJ8J0r+r+6b4
G2n6gyJxbez9QMvzp0MDVdd1b9tktaAl39YSTjXQmejEfko52eqlmYls1rcWFNT7
tvbkkZ+CgBwkaN2qSw6pZd9DTEPAPkh2gIxRH0gU6OF4AT+BcK0BOGYgU9Jp2jvv
zTeoQOgvBDh3oHOvA06b8KhtsQ1wT7ZBMkNFRZx0RcyJmtYok14UT7qy0qVBftmJ
yPysuOklhERTtiIZSNog1TtoN60PCjFLRtsv5db803myE279lEmEC2C1lS8yY/Vs
AbU20+w5DnXqX7SZY5tyid8yxsdJYYLSEfkIFr5ZhiwNt2iCKRcNomBmZdy6kdp9
K5n7/ENzhXISc9OGpdmN9HCu+/QP1ItGTGRc51g17KU2WP1KxSffIb2ptwfXyarn
rlbQO7k5c2Pmu4Xey8hEmOpTNx1CDdQI7yEH8SY/d0JpjzXVxr3udN1VsljYsVrz
eP+PKb52Cx5g2zMQ8/HQrARTlnVFsIxVzWtbFX5qPnuroU6cnUvhkDTwTlRGgyaW
TRohFUyMdjNCOl6KmxCiuHdoPAdzEG4/ReGrpcA3e0AO/PrMYQJBm672Llxxp85F
xEsC/vPRl8gEwIupQB833Opz7LieJae9A2iy8mwhDfPR4pnMTfNk7BSUYaaRfvsN
tWwnIauqgbTw+YtzBxT/CzX73Ye8ypi1HJ5o/AQb+pFM6xlpAfMo0+I2lXIUHZDK
cjho2tvxirCP+txbK41GPEfpUbGScsD1iCkulvfNnGsUXXx6SAq1BAfnqopcZABs
AMsvjJ7jsKkL4zL+0LFbRkAAvWkpqemG8Fp44rd4VkBIHWw+mIEf49GFIDuSVT7m
hdyit9TDdCvRKp/As3vRT0a+8WGyKnfWqnNiS3wg+/lRDKnfxBOI+UNEoXkJOQnt
bOmfQmDfEDV6ey1++SFDmOKrIp0hUnjf/rKCEvpA53NZgB15vUqehkoM3pN+IN5k
LqGPl2XB2ypjLpdqcoEgGgxDilSwV5xTulxq/9K13kwJBDVXWvH0CYKntT3VGWA3
ZT3GSFX0/aYmQ1+4ymbI8/Q4pU27C7DwBsGzBxHddjNUpKY0bULnxnU/3cGEiv1w
1IVf7MAbI2UdiKd/CGwMcM1LAUvLlwF9ciGc4hzVAdL//4z4v/GRKrM8zmuDeYzx
Zq36/BslBJOsm/kH3LZa7PLSLWTEHf/0+RmJEcDslQVVbp27pUixREEY+IQb03pu
JHxYxKfEaWU8iMtNYUXvsfpEjdvEB/bWXVfNp/IOoTNx/Qj3a8Jjp5hFCNmUStU+
cPs/jFuuQ8eSSh2cyJ30Dqeh16TaqoQ0hZ3tFR+FTP0VhXfj0ULXMKtQIGmC4HtL
dc22It3/6CBwu4ci/VAwGpjWvn3E+wc3OzUy/HBbDzNL2QlG4bHvNHNHMTQ2Mo5k
97SXhZNtC+XksL7+tKIR4NJNaR67PI0rCjx11/Q3P3gsziC/cbkff1ASM9WEv7ma
iwY/5tFOuXTfn6tptLD0eehXqH/7tb3YsCUV69fJ9nsO+ccpKQrmQ0PpcktFLBDi
C7Snt02/y1bFLDW5UVM2sSKF3+SnTSPsaF8yYn1Kk+Zp+GEAlhqn9g38PoQuttFs
JciM3Z41TycH6Q7MHP3r+kXwlYENwR0Ywyz+10lrD5DFRM86jAazEWGoWY1cwEIk
+q5wa6ubAIF147FGY96PPTAoZGHWZ9kGml5Q0YuAZaGs9K2WKGvpDHZEr+1HVp2n
Dqu/jyhSKjVmgqyVZ593oYJ7RFRCDq195B4rh2xdM3N3kR3pBZ/buZFvSVr8DsE1
z40iyhzSAI44lA9Yg5/1OMBLC0xM0ktaymlE1nkarPK4yEm/iikwliWQRS+N4Vfy
VlN/8kr5QC0a/lBI6NUP13z8OUMZCYYYvdCwPzMMSJcVCVyY+TZOJMzmKGvK3X+M
rZzNXZo7PpRDRgOP8+BBrQ==
`protect END_PROTECTED
