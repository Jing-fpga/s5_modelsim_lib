`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FxgZm/fCqEhBeNEDMmusYi1kNBGuVlw1mpL1bLiGbwN5W2hoU++9Sp0sdXN+dqZI
TsRjJMQ0f/B9+K0RbNolaP+BzfZsYjWhxCrbj9fzuusHNiExzdNDVKZtx5GLbFIJ
mqo3z3KIHNw6lWO94wc3rZa8SYCWmbkiKhzwUKGbsNTzri5qek9/53pVsV33eYvc
k7XQl/lu4XvVLprpv54hlGiQrTn5MuNR3X/VczET9Acwa1C+HKZgBo2jH8sHp2UN
rvHxwmSsgH7zlDAdqXv2fiZVTyxu1FUB0ftZ2myxuE8r4DoesizeZDKHSYX6TzzK
q5dkPPtuaolpVTpP4pzTfrizkbHxT22hHagIxXv0ECRfOl2a3tN6ZIFTnQO+qTX9
WZd6sh4tNW4q5N7nS367BRyzBNgUAk8kioeAy8FPXY2qrwFi+ni9PqZMHV2/kNnX
Rok1iEn/W0IRjxOXBpgWuYwVSD/Zh92yF2q2z+vyX0tB+cSNJRy6n1kv9f9UDEWZ
WKHjXvS3wDvkxD1ImAP7vsELrJhF28rsWOQQzfZ3lIb+nGAetkABqZhvQk9E/VuC
CIHsTkdAgymrdLhB0XoyFVy2mBe7rHr8wuvdZTKJ4MB+2h7mP4SgtOz48LAM7z+y
BKdT9FEFQ7OUmu79dqUOOsxO/ggpI74pIlMs0/mKIurG89wY2ZKgGpPeEKnO/F1H
qmvtI0jiy+Dq3arehCp5DbyoCBWDTTNhaNCMzEFIAXXiC43kNsufbvf+N9Xxt7zV
lhqL9S5MsVdz1UDTtpXtCzc++wtkKqWF4jwj4zJ4Zr4JdTl6Jf6cZ5gwGgAEa6+K
M6NB6LJpmuIKCPxveUbSBg==
`protect END_PROTECTED
