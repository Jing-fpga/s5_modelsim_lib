`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ODgHoYtONUF/0AyvdxKehHAWwxmzRi9Q4JW0CMBO3KyRadVCPhUL7zK9P7GM9i7
cZ4f2OdKbUy/dOJr4Qz51lpizKrdrfOapKu8JAyVELrz4TvefUu1aqHyEq5f7OhJ
i1rDBNKm6UdQKBegEmjZp69Rl43PC1142GnKikaftDOro5vc8Qmu0YWwrW2qZAVe
STOK5M76CCvWnrcjt1VaB8TFJ+588YMmNfwmJluoAmUp0xsP0n6vQAt5CCUBkBj+
ahad2Uv4UfiFVuWDkckQqcGKlwJ4drSZITNbqNPzR5utXxYoqrcZK91IrOKhXCIZ
K2x91GgIcdcUt2jNgvDXMUDE3TfvawkJVOorcfyS0dMHfUqcFJP8fwjHANPGn78U
9omTWCekBpPXmKBKthnAgVH9aQ0mN4teB6KEDLsCX7H30x3vuKh8v2Wvs8+KAnlJ
eX8d3ZDz+zx9LBFpFA9a3kucbYoHjlAULTE5n6hGESYUZEl45zq/wAKFyqwBCRAe
lZSLc23SHdymOZVMW0BqVITolaVjJXwTEWTEHjcx1UFfxMKBgbEXqcd0AhoyLG9B
YWTNb/xfWp3zRYn5L45kZZYESfAMYyHWwOIpTYQQRXTpqKRGX1Tw/3JtNlbglWoW
LpkKehnzskisrLmm6Wv4T6TbBmOxf3eKOhhrKf2+0aUtKL+PgObrTWOtYM4Dz0b1
sKYsHrE5q0/XP38qNunLa6Cvb2l0A6EAIqYABM4Tbb8GxClYEJ4YqrraUQCQSra3
Ykt7isgcU7JzZeZOuBjpBKzSkpY8LiK+HrFpEMzp5+T9FaQbhMGX/LNm0JUEeNzV
kwJWrntUwXsjGnnLaWzXN57yiVRJUQ5u3ZFiZFaT7gg32gejPJhyroATMWPDib6o
RKEJlNKLX7XELd0LtnRTquh24sSqTCvnA7FuNBM4xPwaigFPmOPnYB/3BpmmK5iI
sLu7s4/5m1UtFbxbmTYttSCsxi4KZrX6m+plWPHKjjBH1mYBZk2XDgDLUdY7DOxS
qG7RvdS2t4jjMnjhDOv2VdmLfWvSFey9G/gxe/csG0E4G/0k2k9Qdqc18IO+tzzk
HOIjkcTiaPOuW5/b3rux5SQMX8ztRjU4+t9urBSaQ/swfa9gx+XeRQI6ZZT/LfZX
jesyFNgthAIsa1kuZ20+gJ6LZ/P3jDup32VJG6qygujw7R8mVFhCCDe/2xzVPtjL
5u1PZ7vj+MzEMaFyJzz31WG9ToEkGJrKkZjN/18b/wFKpNR0ZT99Rn9+9xdZpy54
ogXr1/ONfCB9ByZtlG15BTOz7CmZTenZyADbjFSBWgzif8RkQkXH5+HCJmoI5A5l
wzP9mWx+Iqcv+w5JBkW2jsFj0kcwsSReAfD2bHEEtWX7ZaOUlUcERBtTsep03V0L
YF/+x8QeMF/4CWdRNjLZWMG0jnz6bNN8mE0H8LK6Bfi8Y175Xc4xLlCZHBBWVrfH
47xBLAQelQDhqoH+JjIlL/jnYlN/IRx6HKVb2ECAJvkRSaGWfuk8rvMVij2KTzaM
eSt9KRztprF6SlI758qw1pHPJhK5fnSv7rDJVtwEzrOOUsV47SDcCJH0bfxJWd1o
1eTcv4uOqSMMrmkS72Vf518876/CGUnUPDZzUyu0toKVMIG6ljwAmsQhZosixxyi
djzrHWMifZSqUD8cWVIk2uPn8HW+YZAkVRrDuv3YD3TFGwPgnn70DD6X8bxd7xcD
XrOENNHjVnhvzXH+b074n5PbbQHLc6XqCMF7zokugPioBXZYfRPRa+PiUHYVan5s
b48OKY5rO6YT5ZN0BkEz7qzLjUkuwMmi23JKsOjHnpUASrH5CsvwlpTKZBLNpvzR
8DTvfMK4/KvkVXsuZrerBC4uAVUJV3mX3o+zkVc18Ejuc7d9W76qpGmoc30LxD0F
UOg01peOA3CXibTm+k1H8EjJlrYqOm/1vxBVg3alM+8XdMywdaClyYpj7nrChgpv
YEzp4+AD4dUk2QIxKWLr4ZjSmegJ0Jbqn0hm0mY0EuT3Tvvfm9GOfDJpAFe6CZFO
QQuoe1+T3s6uno7a4O9WhzPuKlUUlyz7N9jh13BSOt05dT3V3wXUDILZj+1ssxqU
49E6wc/S+mVGxTkVLqpmKrpRUnWjXmeJlWBgyMYgI6SAe9x9A0Y6D/UNhnWXzWPd
QdtLfVZf/QyUXG+AvTluTI9LgIa2XFkKk4TzDhwFDlehmyw8TP8fKlM5A8GPubZM
JojXwlfOyKwQhpocI07v1N6PIlwpKjWcHzEuHk1mH0B3swRIDfyXPs+s8zYTgvlb
y0jWtipcUCJMScaYc0jMWM86MAqw9wmS6NaxD8au18a54GhjXgALdEYTLklV/vxH
`protect END_PROTECTED
