`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ew4sxlAjnTkfJiI/qs+AMS7DQDSdoabaoU9ff+td3QmfktjgIhbnCDiS7RFEyqHc
xUjm9SodLXvWkVdHsZTpxClFImtfNBnYGjRkLKCWydnC+pADOJiUkQEqBQVR4yi7
e6CK4cDDOnEQ5TjYqz/IGD2eaPAIeZN80BwXYO99ynxacj3wnyrp3flz0IHLuL0w
BlvMITQ7juB2iK0WNwwyCdkcf8JDW8AJpPhaIbiPEdFbWhFJZ4rXRDHHPMYnFdAk
rfI2x2NKKDKVTerunvNGawH3pOOFXctqtLZcKXF0OLiQvGvsjDLexyzplSl665C/
UDw+/OCSGihYPyfI5N3elPkM8son5cykAb7W/nk4pMnl9xFOGtrskczB6cKGO9bR
uCRr6nbCPJKBSP23SywAEFVH/Y8OTGKBRs7mQg8OGnLz6NDDHY1JoHlovP8AYxfQ
yqgsgoLN1Wrr82IZFcY0prUvmT6m6Zbmyl+pktmCrm0JHeRpJENNPBZAl6UO26Cu
QGpiSsQgkYjAfYLrvwUcMkQcm+QZ5ieYKGnvOpclzv8XRGdwhKNbPzZn2/4KKfe6
pWekqi6kc7bUJAPntNMTAAGqcb3+niXnNk/DGq+XJ+uIVkVCSIMTP165rJVG7IA/
Z0Ux/xC5TLwgB+Q1OZW9l+HlundLr43qYSGeNyjoqzBDpPrLmP9TywttIluQZuRE
LxE3gO8ZARIYdFHRz81cP6pQOifc6H8uYUkW8FfQBZMO8oM/b5REUL0Ncfn8A9sR
KseU5BQEsiujgwc8KlG2kGBBI5EOnGFQJXwWNf4Lp3TriIQPNyvQTqkQmfGVz2jj
FzSzj86F23+NRccxvP1syyPRkwBtmTA9VOuZWEivQXbHrql2opH+WFmlaMf6w+Fa
xmgUS56l5eNLJd/aTNRmmWxyx9MdDusTNWxbfclPl5zRCFIza2As89OiceYovpS7
4xpI7V3UELPxESxE3x7xivlUVbuPDsHeTiQoytZgGahdoq5aYqAJcW0kcXh6TGg3
H1tnjwLfP4SwNuc8bZP4RXDyeznCoJYfKr4bA6THzENcKtni3OSHvuauc0urO8lX
Q1CP80c66oUuWRz46fJSD0vB7VInOlNpr6bZOGJn6q8tWWnmRWwCT3b782alLzZS
+hf14cG6Bruaq5QoaowENxCLViOw97Y/Rp9SuCbZXOZRmk4Q6lCOB4K2iUBAhw2H
fW4i3M7iicoUi5cvvZ6hnzYVymucrWwVZtWs62QCWtH902ZICui/A0ZjvAQV/h/o
MZnDl19/29cYh7UwiDAhYJTVdlKbFMFquzXLJJPT8OmOJ0FwRtuZ7dgXbuRnlcZx
yP5zz83TrhEyQceS6Msf3MCsmWphfD85xS2fPT2aAkqKs6QpqoqixeFEYutQ+vHZ
ov7hyp2YX327EYNYEUfvG5MlgvIFcUXEo1hMsAtFfogHzLJLjjJF9oUOnZLu8Y9n
Ry4wbTV8NuYYdtEtJzvxlMgT3aTS3wWI2IPY5spVvAubsUkqrjGkXoUxPk+FZK9e
xJ/05Jt7zzocIohYOb/RV0AmB+v3OVagnPQY8fuVvh86vFsvfwcS3iGnZDwLI6xx
HXGC7S6id1Q82u3DhhnsN6ThL/XtA8L8GFayz0EOYVBmwbqdKOkC0EKekI/BfUAW
nBp4Zn4IfwflRvIwmx+WyBixlpv39DGP8hV5U4MRYtGjrkFwEr/t2tQL4l/qE7Hm
v5s0WCG4+tMcUCDFQg+hrcp9xRhByt1HK0O5bfRqm0zVASmR2CUufntM13n/6+uN
6sVTnhuInPb6ivG7YidwLMIMpZflKTl60MdLv8iboZx7AkJf7XjKahUczyailQ10
F507kGbeA8IGULrlGcGKRwzgTwURD81nEwX5XSxD9B03XesZ66MvjLhIV04o05fv
dektZMYnqpTD7761RtBOuhZIH1CsT6eiCOJ4N88NofTMSPfd0NXHpO53HSRBYsVJ
nclISLkAhfMjXdh36pn2qptk0LDBblsJN1BSzDZbzVsFodWe3Fi7BDBSRSw7TwcR
uee0WRrCHWjZ9AF18Il9aKbaG6TP+PlJeszza7uaiuJMXCzVagr6V05/S3VR8HD/
VgJ4M8faR6jg8o57at1E87GYZ7K+SrIDI3AY7FYRufxloV7G9VS/efEbxKuTvkxm
LZkPpFopkWJ16o5Nde6d32Vf3K9/FK39brIL0evXRkamXzU7fanpwzOeuZLz1Xps
kPokDUcTtcDoNc1ULnx9fgW4jdKJnA2IHWZV4vy2GpUxD/q6SuMwR+3F8Rl2DasX
Wgr3+ZoVFWLpF9o6VsX1zf5H/S8Eg5yTp1sqgxkwK8eUTRH7kpAMskvKzs6z16Nz
GZjRV0kmVgsJoSGA3HLdyYyTQrQzNezBZw2cXDJ1x6VVteTnG134T4FBD64KAGxr
yBzg87kWIkVO7mEx+PNEC66J02OYWl8VbV2lyLNKhT986DEiZfVaJ9qodl8Ml9R5
Bq1RPpRFP1VC0EhtEwZQHkZajiw4aIZUaDw3PfSeuaqb/tRI36ZvSVFXEDJL3Kpr
lZ8ZQ+B3AEOsoMRAMTxT4QEpipaiE2XU6Dv8K4m4/TSeCbzcWiufmkxU08/cRFNT
J5wvFbZJy7V0kYXtyc6eJbj3toKE/Gcbu8epfn7jKXnpwKKXS0moaljAvXeZ4exv
xK5A7SfzIVnFUWgRrvx1abU0uXX21ShGIl/ltGvwA6Dx/Z2aYHSdGM6YSBggDefO
f28GP4MjCJ1elp8W4LmpMPRlCMzItY/GSukgvD89/EQjLXEjBpvUq31L8/N6W2Dx
2bOkM/VYdSS7IV61DkL7ZlbbjlqXK7NFdVV+7gdHVL8gTMW3i/58hEpenIxnxNwL
nwxhHbPDOunmnrka1qooi0NOM4r5OhwEQ4nl5/q64dC8LA/hRRA4GtuWFX6+10KY
KHU9JteBl1Q3BnpDEtjYvjKieQ79lFFKxN2HWVYO7II3yj0q+D3o05uDMPOlWswD
3iVynHx4PGzI3PtehOH18YZvCwdFRowIVSRtKuD9Qt9SnJ5xcOShp9ub4TG/4kmx
1JLNzj+yWPUJkxiSNGGyjY29e2YSFr0YQIvuQsTarMKe/D+2qSTABvglfnuqeuZK
StVlmKLw+oYgMup1ibW4LG7sU8vByG8saaJiwBv5kW+TcYlm2VYgVC/9RxhA1vvK
T9wo8xMctAeRjg8Uvn8srWOmKGhq7+SA74wYlqjzker/JRx31Q9v/o7weXKP90Sa
jbPF3ZqhAJzSgn38+j6AYpNReG/2k/wekjB5VXrO/Tgvt1lCQOtUPIfAnZHCNOVb
asPKeGkiZlX+ss4rT3CyFew94rQgt6393IWfKIY63+ntkD72fXHg32a2yOtLUbsq
rVZboJ01wKhqw7P07LDVdVMAaskac9us18+dMu1seqVkz+/+advi/5nrlbab+ZDX
HWSsCsV2s+PGtzAR79RkgAFD4ycijl9aAV0FuyL/6sv6jehUcKkIvCMvhL9KRNFS
KVqz/RWxXjQqCWqDZDNgrW0wxg4KqmNiXKuI+jZ+Raj6UL3t6oNeTSo6BThvFZJK
rc0ZTaywy/ij6mluKIeLRg90yf1MPyMTWFxeDhTIptef6VnE3i41iuf/j22g36yc
1R5wpZpo5VbfIRjVz5g4I56H6PuA5kRkRdzjxuNkSZqXi8ElygGbszaHAaXvRNGD
xsgWmbuHcVLlg1VtngD+7XS7P3cFBdsfSvFsYy6omknGZWJogBnIi1TP/PsauaK5
k34TSjAiX2qcMUwXisTQp/BhFyqUNWXdBWqVu4JSpMzpViUbZGiUK4lak/nK6vLi
25DIKgIifoW1bbYoHxPZcSA8O6u12Zf5BF2vQRPM/+fT6w0waXx6MKNCEnTyiCPB
LBBWp2kNeG4PCctPgeRGBGMxI+J38/WQsYINEkR0TQU95KraJ2Kml5Aoz04bybON
Ce40JnE/4wp/O8Bn8o6JselapBcnNfamH/7HPu3KIpYaw7U1FAR9Sq1G6ujKEaVN
aEcWsS3sEBsYmxQt7H5Io/dA0GmEnTTNJn3ItzFMy9OaJun0ZhAeGi3ZDOC+oXaY
icLg2vtH3ZnXv7V9ypJdsaSr2Y1QrnBM77a1iYt4uDoNX+eJxh4j53s40ha8dD8Z
PEGLia0S7Ey8XfHCCr6O7GPj1Gh2/C41RDVZECNuIbr2EieZxZXuL56lTZEtJ3aL
DMrAt5q8FEe6Co99P5v4RgBklkr2tg1cOWHOwdW4d25RLVi1ML5IT+R8ALH2eJ4s
UxvBNhbvmrQ/SHhhrFoeEPL8vcQNeVmeQhc1v1yLT9VME3wq1GT05pS3Y3alVi59
ejBVwQj+erW23tQ/h2pSKet4Ah4zORnggHVpZq1aTZwdNHtYj8uJrXDuAtS4l07J
PHqFXCpU3iB7SLQ30ujW4bOo+6/nNta0W0ZIyC0ujUkyaMw/gbftrGIoi+QxB0ir
UmPCTSpVMME4vNC9/qcwYUKgjwn7IbX5A4+SzL0TeocLDmbEArVtOJEN/+8EPyxU
ui+5NtpVmyUlwFUq7NGP+UZasqIp7rOxVHk+okkUImJUbyEDwsINesZBRijOVEQV
LIMlJWaDrOekbqYrn0n6kvo2LbisSKlea52xlzTCNF6UCPGsR5bDR30T8MOKoQK5
75pbjhAV3jZhQG6jr+Q5w2l5zppyU1pcMhLZdIKIr9+SdzLGKQQX96FeMgqgy6cZ
9xSOJ9D2yhTO55WWd5xNmaml9LGnXF20ukTONINH67eWXXk0O8+0rIsRtgcdpRyM
aJXswcd50e+7rpzM4u12AtfY4tYd3ndLjaSTGHOwSVNypnV3snkn/Vh0IRJMdLve
5aQfPXeqATj+KPDWOR4wdvHlKYuaq2TXATLJPHRz6SsK4Di+pDl7WlBwZI4L2Ykx
pZKdrazLnpE80lSkHAjAUd+HJsD8SclrKODCx5dmhcxXINjjjBT27czTpERtG2gg
kVl5iI8IjqLbBzfhGSswzSq431+jokg+PjnvbFT2zmcaJyUPD+XZC9w17bxKEFcg
6V1X5KSsaT7sTqMLtMLNKkyKE50b5pB+TayXHsro26e3J+5X5fdzaXnEMuWaJooE
2MMVLLbRwr28k7KY9/CGOBILScQjWLagGun1EgIfyGB9ADBp2qJ6pw4ALgE7FQRA
X7JAByxRAUDKuFTuoMI0hwe3Pu3nRsZ+g7khlOdE1+PZMLOwqVbDzvQIO1lD8ojD
8oqk2Z+slbCrdrXTUj3YIUkZswO/50Y6lx8WRtdUEujaM9hmSKCkCbyysiWKQP5N
zD0LRCyp7qNcYVEmj0sOlth/i6+mnLoQ3sd4er6kztx7iIe21aDoaJdjhTMmVfBa
1FuffwHHMqHg5uAjIOX8iHdpOsi/0OjA9WMD6d20XdaAbUgoU+OgMPxfYOgcjR1V
VHpog5pPWO5a80J5DJ9l+LsMnp6X5yWRD5Zmtlmx+babDCeUaQOqJMd58PiX7j7T
u0QoOXsen2utv7avMoNvlfI89HVMWQJ/JEhp1OFABHQJ4SV2hwvuj3adKf9+naDP
SuROfEecWDA4dfoWtdubcsW4/q0aV3QC0+UCmNLeCF5JdOzkh8whVWbKNFxSTdg+
cU6eLrNXOlzIoFhS53MJyJ8vLbr9/nUGePLU1fYcV0mF06rwqFk7gKEEVLAcpPbU
96g6xSRw0eBkV4yYVven1j424qcBB9zKPaksbjO03NJgjJhTYhOw/c39xXH3LuSX
BkdteRDT8oQBixARG3AW77jUBZCdo+tp+wfb038Kk53L09x/jF4POgDxNusowDnU
4CeJPkvpbSP1XsDkB5uridZoQymKK/VRF9OvRp58FlcRKIO7cY8SMI9uJ7IOx6Tr
aks4kbwJHNc5tNWjkGFSDqQkyBSyTq/hIYo1q9xc9jDw6wI4BqH80XRdqGxd9JYX
/QTRtZ8UMxdeyLnEdXut2WFq4cbptASwnyXh5IBJjCIiHZcJuGj4ksYLKo4LRZMe
4ngaChjstY3MyeIbNSE6eqCJvRv1TEZ2qdtEsUxMaqgTs7N//lREYD4GT83Dvbm0
zuWaXAg1Yz1qIa0KDbtLBKXH5GjvxShqVKdpxYSoRwGkaRWJPjUC1yvNfHzUi/dY
q+ZnSOlX6lgSbi3j8JITkrJtGFsOkuvWM4kql5/AVzC1qLnNangT6gVMUcLQSJ57
yh/zkdg4x4sVhdVpFlsXk9VQeJhsS1atw5YWWjmzclzdvzovLc1p2sbVuhmcTw8N
TSBWxK/KUO/VXTDdXfQ5uq9+Jt7zh4YgOPk4qHbJEyE7+xMlLWJniGwhPVnlHXOH
S13Fs7hEKOa9f6nlUUiSf3BcEONGoQggtKnuIt8tQ43HqFvf1mpxt92GfI5fYfRi
3tZhmKvFLHtAGX0PQ55uLCrDckWyG1kLZt2HcRpPrn0B/yw2yGMmQd7qx8TP6l4D
TvxVUSXT+i3BkBJTGHlLebDqBw8oTBgSWgSQE+266eR6w7p+ATbIUOAbJ11pE4Yp
KclQwTTE4SxQ6iiAzEH1QDtMHao1k1KZ2lIq6AY3meaEivXJe8yeYvwjLBzfGR6j
ORJ+3SUfW6cMs7E99N14QIGFVJlMLuehA1PdltlQXM3s2MwvJcpksSZrBzNEI9L6
ANmhyi+MFz1oHyOlMUIu7Lyte/u+CHh9hOhdQ7BcRPcqtc6SYUCbI3qk90wXkCpX
F0Yt9vA+G9m0d0Te/Ci9/SN3oG25poY4nEtd+DxHjNmtn2v4Pq1ENmnaofhgdwtg
J0/ZiwZbMPwyyudODCUYO7TD/Dlm/gmoNHpcBR/+GQ96b3um/gEqsI9wtdN8QvTF
+UV6hD0CEM4BDz4g0IRLnyKTsu584v/r6voK/HSeK0R0cecJdDKoToGb8C0kJJUf
FMjd1S5XNohVVdDE3xMua8/J3O8asZWfVtafrQC0Wiad8ni/qPv46hiZgrTVtaQY
dvUfc3JSB2Gobuq5x6n+LN/EOkzsKSVNJ7x/Z+IAlV6zZ7RpWRsyRFXjhx0rtrR7
NDwoYQLk6Ohs5Jt1YvoPnqi7vgqo4be4M/jX9dCzG+ydzB9wFMYPUxX0Mrlmma6E
gAc9aBS5WNy9PHnJjNvMNCD8r1xsavcec0+jziiQKNOyF3/zGSw+lgohxGsPFSjs
9EbTj9+3J+l7ULUhFJkU8Q5eHtDQzijjYXttkkaSlNu+0EhoAgU/YeVlEYrMj1Co
itSBqdhDeZ3oL/iku5SEqDl+I28tByA534g4UeeeoOw1cT1EiOs44UpBAzUdBDgL
e6heQ1a7x0eYpJsRbJQ15IBG2DGA1pYK+auGfo/K8k6z2GE46SGr88vkVDvnlk+/
D+msvHMd5c8z7kRF2tD3328cPLag20/OA2A20kaX1ZaxWhRSdJm7FYJRSytrDh1A
aIZOHqQ2kKL7gMcJJb5dbQPay/EWK4WWuMRNN63cmltcmA+aAGRZBg7mdUklXgFU
jFBu3Yb8yV9M29BIVk4BEesx/5CzyUzLRogUCTU38QwZMC4VYqSx28RcrNfjacTV
qOttCJmwakXCcq/eLRh4tXVjK4ucpsSnkuHmlHcfPOJtGpRLdW2w5Q/zXy1nDa6k
OO0T/qoq3HuDLLj8B38Xx/bm10lLJRK9tILQWOuSq5euDMfXbM3BZRE3fcippowo
x4eD3bAUljT3WlsFIAgoqnpGg9j5wnyXG8ThXYjTBKrdhwc19j9Z0aqBpmUhthap
0cMXmoxjrNYp456P4fdDxxtqVIaT3Smg577diRhMKt8izeVQlnmpyXu4+BItYvCy
3SoFZg5vyPw09b0waIUkmd18mG+PfZuT/5XHHt67rP7Nsd6QDlhwnYrNXDC9mUZt
Q6eL0ubEBZO8X0EU9gAnJlHED0gx2R8Tm55jZHVeCqDYmkuAONmmM5YlyE43HwxG
ntwbH7eZlXntDeyhtiWqJ+mDcJPbwDsh4INV8OnemWGdR6YrKR5HRIf+1n3B/dFm
IPfgvv1xoBQu1TIH554krxS8/YHMs1mmosa5iFgVMm6OE64cK5+9THivvPasJhkJ
BIY1SB1A/eOszETIN1SS2n07/xFV5/LUy35wu+GYy7pEIB0K4pYJ5UFbDTP+fdxR
NOHbwsvyTh9NYOCLy3Dv3PooWmUxYAOO1i2lHHVsHrU9bcEHXCKnHGKjRrSwa0ou
tmquZmn27SbxGcP5dFEu29cR5McmCaEF+iwGyxaD3yepaYz5QZNNOLz/EIyn51zR
CF45V5AjyW1OXZKVJDvCLtgnMZSWVrTVhrVpPaYqnobbt8q0SEb09ADiaFCzIRrA
/uCotwsvqyV8mGXzBqnkR01ODGcxhQ5ESCGvcu+rP3doou/jY73bcvhAj0Q/EM7w
eFQPfQsqh6/1IEvvnoz1cukWq0x+rMGT0S+2N/CKGVnPbAklV8hMFrFqoGsLyf0e
5W03ssxoLf0MWoD3m8CweU7tE8b2B2d27xh1l3d2QVvNSbqkfNmRy5T9rASJuCRf
ftV3tEk00BvM1AFuuqEzGQ0Kco0yeSnIrOI2e6B7Cm1h0L0nAqeq3i38b80zp0w5
ZBTgJVVdx8e2HtK0m2Ch9roSw1YjwWLl/Gm+gcJiG1kur7x3nsRrx/Tbbxc7otL4
yOY6fFXIOrwW39LsGvV77eL8oWeRgSE8giAxBQSF8T+qxHmShGoKn/M6JmATv+vC
sZ3Yi/8uQARS7uZjZBy5tA118um5Kgvso6Nhm6tffUvNFC3yC+NWIFCpAx4Whirx
WogclHOhfWD3jDMSd++/x3m6p/GkndpxgZtjvFB2tntpwvWKl18TvKVryHvYI9zL
rWCIojTWNy8gfm+AE1uuyOtZt6+GvlvpTUim0jUDm2tmMRlLSRvMBI9g4iOL/T2A
ZTfudpxkTSPBcUIq1zer1OazKymHi0urhWdDlo6gEJ4/WtIsok814Bw+AYqc3xKn
4sowtGPDoHVCulJeQj/oFmVnn6iur7Bi/5wi1IpoDUTS1H0aNEdG9FnZbj08nBNK
QWJVlWcKoNDiFMbx3SS13n5ehIYHry0+kZF0K8hSFJ0ePkx4MzZ9wQkxi29ZNH4c
i2UBXkubeFiG2iyAew7W2KQXORoa5D7vFPKlAGb81CV1UtKikv76gJJJjYP7cacC
iyBi6YAmf2m3AsiScWSEygY2jISo1RYOksRQbskIIo+u7nSGdB3TxPExb2TNbuGx
jn4/96kNQhTLcoArQif6e6DRO5KgNsX4TAHWyg/OffyVtxZ/BRic6iR7HgYF+Jpa
m8aEHXPpYH05rZFIhYUas8+Xjp2xUgCwY3BBsGnxV5x5aajvT8F8FEH7vibrOKL1
D0HDhWFcRpSKp/NiavX/3MRAPSmq54S16vE8TRIXaO6A9McreLkIfnqQOgviUwzn
6s/mid+nwwnSPH37Ubg8wECpJo2G2PwdJpeD4k4/H1LBuVHhWAJqcTgSvoXQ/ShL
tLAzyucM7jJFz6XLQKsNJtIXEQz/Nj1CwxeaT024TfVn32mM+XUMdDUVZsUEqNWq
RYive7rbkyolzwtqXj4leDxDm3m0ebvxwELPyS+c3ngyhhv3fSK5W9MvmOlGPRgX
6xoyvGngh9aKJGQeAPNinftyq5HsmVMr+bLuIqlxIhIejkZfRfJhswky/lR9eI3T
U2EmJQZSioBY0lIIK+t2vYCcKnbK5f3QheA9y+3rDeKlEDKzxAx4/nxh64vJCBkI
G6M/aQXfpQFo4nlG7L7uRn1nEyxB6edQe28kOOIg3PCFoCO8TvSc3/xLe4lPBcc2
i0og4FHER/Qu9cXZzpBQEzIKi3adLiSMgr+/iqmdf4tXq7hxfHfpZA/2bVGLbpXn
PsVnZR1hyvrf+heNWK8Qk+gZ+0oyhQoWA2ltRrM7DiD+GeBf+RMv230creSPhvIZ
UCh9pryrkR8I9N7KdVEnfmWK51ZrlucJkSsThLhKxcBFy4H+kfeZT+WF9xZhJMi0
JKpafGFyK5iEfBH4heES/161MECSIoPBrbqCaUrLGLjiLu3lMNOEcD4nIShy45xB
rm0FjtIILCWgiuDEsn7LTkLmT2F87YnWPvqXP/+V+v/LJJLtJvm0CCzBs8Uj5mnN
8BpcbZR01prpW9WM8RISlOGfpshpUOfgGH0mPg1N0zfJhZS4eclnG5KBwbzo0bMT
+IG578ODhAZNmznSggMsZJdTNFP3FE/k+G626qIvum+yRJn9tsP1Td2Pl+sito+V
Va7OLHSD5aapA6hZtilsNI9gX46ioVYSN9MNezqPtVnGWS7Nn4y4uOnQbLGY6ENn
Pa6vbGKuB5pjNhTmD+rag9qM5DF2WQUNMViNkd99vki+ALRdT4dg+cGxdv6roUHC
ofVYP4+tOKV51YJLoV9D52IWhDSCvJr0oRRRTrgiFaywhV+xZRS1g4XqoixaSmBB
mg6bE5jMQ1MuGOvEqOSlaj1leqF3+8aIQkN/u4ykIqDIs5N5LXy8Z0j64IF0J6sy
GbEAJzbvSl5cVlZI9Z88Pg18iMfcA9SNk/HkcVevfvt0r1XkNyxWdUcOYITZWi1q
BIISPA9J4dRvXWMUqGtFzq+/X243G+A28XVW3mOzXu0Bl6bdhph0bqj26q0TVX6p
CMcuBCIZR8D2t96zhQgPZB0/+c38NyqoDOuuw43o9X4cOJmNjeedaCqg4y6+qsHo
5LhCt2n4ZdMXq/daSobflbCzmfV9LdmIaOp2OdCN3gnTG/btPFmvXjX513bYPm79
tG9PyLD/MgGQnIPkvQZ/k01+tkiT4qE/VkaHrxGnOdLjqh6sLYgVdSAHxVjzEWcq
ga1m2keDQW9bjbTE9WVLUNtftRDXdzRNc8asLkzMKIuYX4S6/iDfh7kjVtfqadAZ
FIIu9YGr2YC3O47aoZEPHWOfPTebYwMjy8IXELP2ucHOwrUv3ztpSXMKW6DiW+7o
vjGKiWHzn0v5Mq0QR4NZKp9f3rJGKMk8MBQFfFUuzpFiWcvq8sBRup2vrPibTcyB
iyPtseWR/5y9KWCbKOQjLWQWiCBE5afUaIWB/CZ2PochejZ1+5cEuHOQTe/dFIKK
ZTs8LZXGPjTopJbpiZ7lxNI8DIvddLc0uHnrKMcz9NDmt2TsqAdqgLFtjLpxLqGv
XJfm4GIdOAE0D5DM22Li8hgo1f9wt6bWHk5iNzrv5uDaj5A/fhfALs3NSn5c3QXP
w5LMtljY7qfztltN4awXBbbUKRIwgr0QkjbsOCy9MVHHgNL6VVQi2NgzmPOWYpy/
5WlkgfacDD9FafjmdkT5d8ArdHpaYwvhd+6C5iN0hgbq7cLbtqWU9AoM7td4ewW2
fRM9MLiYraCAjVbOhHYue9wBrpb7TnvBSHYotRnH+9ECyBhd2QilNwAGeTVJbqGX
K4lbWxuie2eXhv5wjKXJmUxOhTz2b4M30OxLvLcQmUvf1O1+e4eLncpbINuplxQc
7JyWwP2Gv+Vogc/daKa9q08H5dTSm3vykpet2PGr/mRcPELY6HO43qqrYQIr32tk
p9rNXsQLaC1nH1Ml/NAwUjbs6c4VApM0GNfTs8yV1xHkrTZucKEUwQVZUGkWHIoy
P3lLYG44Zl+p+hwUP+/5p9SKtm/YYyz2V4bcGLkheRv2m4EhZxZEQw4vmDp33C2J
xgNL/b+ZWtB0gTKztcD9hb8Q0kCcJ9yq2Snr/gpjT9XoQuvaP4Phq3AdQvIMk0P4
4BH3zLoaSHYuKvLk25oLOmBYgLur1OCRp2JjmNikGq5NHIic+Rl6eRKQkk4wDATv
APSg7htfmbQsdg55vv4gh9dU2dqEZCwvfGj+fw0sKoAXjJC2TQB8dnRTKLq6uyXg
UtNv28OMuFQyjRjSb8E2FwzwCGuhWag1GpsgAe1aHQ0VPkY3FHrJNNwQOJbHcRFu
wDK/u+SnA1lhQQKzxS6VsvdHbNahe0veUYJJ+j6RMg+Z4H1l1Anrc5y0G/VArTRE
m7rgVsGnPhwE+xjsN3W3EorpHlp3PT8CMRLnStsKM3+J7jI8s1vxRGpifI2V6Pbe
jXVX1n9laOsMtE54KmqmUy8FU2dDHvrDGlxLVkaVERFtXI9UEgppb6UNDZM1dbhI
rdWEPeap/8A5MAyneqyAkSZ+yeUo6j8N5ULGX2tlNf/XFjpWix677K+7QNLUXRCZ
zo1DKafcygS+P9+2vTxK6QXl0Dt9/AOmECZCjXEijlSZ1tuSMy1wni5H5dDwP37U
bY2UHoKLP2tIxATQmImZGpR8Wt8scyxOQz+ykQnVQavchzdTYl0Xhn01HXJp8Xy8
jzuISStwNAlU+Tma+Jza+3oYJinSo9OkE4EhyWe0XZn//UCp/1ODm8lsAY0SEHt8
3Lz0c2qP6sRMhzkINbrhD341MlNpCOVdPHi0cDdDHhjEYw1gRw+PRpmQGZbbP9Bk
7yztIT0fgjG5x+6o1s1DYedtamIbIj9p3fEGqw/+4Ev6bUt3C9EAQPsU9VE4tYlp
vYFx9zMmtUMy/mtKwsG1+LsRD9SBAZPrKtCZ3yNOjnXT+GHuJpDXeRrlIlTMxPxf
KOq3PA7oR4MNzo30EzWZu1B/D31N/wO73I5WxRpgUjplBrzCARXX8eDrE/A6CQRO
vQdjccU6D0X2rrn5teDJ+k9HJULMEpCSeoPidRk/kCPXWeWhQ9KW9uR1L5ed+bdA
wIq2DcISuXl6cxOwbOLUlqE4EUbrQsigP0f0Wdf3v4SuT3cREwFH95UDb0H7b06t
K22OTQrq1yOM4c6sqJrkObjet89A48bUQ88CtrZn70AlNIglS3h/SLqsU1Ava7A3
HlwQRwEAheZ63DBxa3yDFM1nA6Hr1qDgUrb7uXlPncmO2WqMHv8fdj0HQcdnq3cQ
DkSsMk2b7n+gKUWNMY2gfNKzI7CnUn/wcni5UAHUAUKMyJefl/be8nAH48rqi/ej
dimZvQ51kjQtey/eIcHlL/RbNUXcjSPb+R93VFTDHmmpydzqBmEfeV6Oot6H0Z1l
vuiscWAKIbELpdCoM39cdWCLIPrPWXdRJDdrICviIxXhdCQycAo0C/6SQgQ6K/xs
uldrjcNzxx3NoUN/BG9jdTT7Y8mEUpm0BiRz67rHrmFggtfdFNQlF/vzxWQjvkeW
BB+WwhARfyuRsVBgi5QK/jvJ3Hpnp5IoE6WPQZ2SRuqCbMhgKrHolhuuVksie46z
y4duU690JyzBFIJ1yvRTlkkJvfYVTBLU7bmkJw02B3hKtRR3zLXyGjAN6nXjZChj
yswiE6RVMBFUqTolsBnVSczXFVBgG67EFP1le0Q+mIU+/1nJxVzSbpilkbrEj1jw
lOveTN8L6fxJzqYw7F2R0/gqdv+ye+/g8RIGAr3J7Av+vIgms9+ukSBfbehkmVeW
QBa0A8xLaRW1X9jC+QwbgetwLPWZ944xVSeGNIyx2agbHRzgSycqk5tyNIrMoOwX
VJnwWGwGqT3TOIwRiUw0oR/WFl/QbCIBNeW25c3JKH9M7tKZ9GzIo7YQhphqdcyj
M9BVsyZIQoicJFSRV3+9qusTVWS3nsNtt0JnUeI/lB3lHm0dLCon1Ow43nLXD8+1
imq13a6xruZge5oy+ISkZCU7FYMTl6srEJuZ6A3g8ajEPGQ0KLbJdd24SEHXAU5T
hpL/NnrsCvemCu+o5AFad8JNJJvpcAwwDvl3yMGB7VU7QiXbFAbF5WX1Z8yViy7g
DcU6CNK/L5HqDb5CoBVBPconMFBermm+znI382sZ/Jgcu0MnxcIx66lgnDfM6qp+
4IIOTCP9m7ckW1NuWWcIcj/sv1D41tR+PW+chyRQR/GC8nlp5zoJtFCxt8ooqQJC
GXXnCfNI0WzOSXYNuKh7x+1au8uP059TUiAlKStTWxE9PCGksovz50CrBSX8AGXj
75e5Ba/FyifrLlxKlR+lcX6jfoOrmB9SAE8iHwvuAnAQBUK53EiFXPKqHvWp6Cqf
zz/rma+ci3OIZrw8x34GM2UF4nWL+BRlefEAw8QhQOnUpslkVSa1gKDCbSQ/51Od
IJs1U24KRhmlbqcMEk0GO/Aoe1ZJ4xwKuxvUot828/Eu/t8vMzHzh3Nw9szf/b/5
rcfq+ps2V0hl/cxiaWk5TIewrTNGe8U0tEM9sfbQEnSQQ1hG9VyeH5PSt7dprLA6
KZDdSyZ8jXlfK239dvnhBfvZYpm2zQLg+1K7SQEzd7LpobHp0ry58KvjnEPqZuuq
krN+l6ACzNxnzoBZbm7VKmdWFnUz3ewQRurzEPPvb3PAVVJOnQdBiI7W/LB3hxra
1tx0hlLBiyQET9uoDX52vYfC0rS2CC5Jk+pH4VYz5CbQkcHh5r+GpvmzyM3gdj65
Id+bCeOxQdMepx46ARcpKLl8jv0t7mC2BQDqHwdCgNxXDprlplqB7wpk+StIMkRW
2Q9xtplrF2acT5U/sDIyv4Ok674o39NUmKza3bUSR4ioBedryRONz5pu1gFUQqLn
dQP+jC8L1XG+zEb4vQ/BsEI4b5TeebxFcd0QZ8oOn6szwDeR0tJWDfKqLgBdYFz7
k4p6tq7UCgNqzX77w0e/WAPueAHFozUmPi3ek6Rvdf2j2dMEG9ZWRu+Y+zavEIdR
59NKDoxsERqBHTlVfMplTqh9ArpjZbUkbXx3cHnKzrihUSanvZaTZyCj8Fb6WQNl
aQhPELfWkUHN9U7l9PGh362g6IY1t/FN5Ypuvc+Et3uXD79Dm2rhAf41hrdtolMD
wiLlkEFKVjZquERLFfx5my9KwPjpmLPaFJ8itff6Puc5oGgMTmx/6JNTi5rZewat
Zqh0bRbbY82lnrsrCjRdJhBuscVnHWs/V/Huj0PSGc1K6x5WR9oEA6mvj9LOQYnH
KNPj82bTdy2gxQWXkkoPRPjMEA0Q6GGKdM2sgkgYLRESJsJXJnSSVfGnLQCMqjK/
lFKPHD8OcX+/cl6I8rfML48kny/FwD6VI2a4oYFTD3bQYPwAsg7vBUG/9UpyHo9N
HfolppCIaX4Zu7cYM27tMvP7QR6g5YrZ7ArvfuYxnVd0q+JD8eKFG21xwMtPnoif
hoMmnCXviUJ0oSR4LgC7aoeu3fnnY3KvKHfdUrICd9/rHDXPTf8a4HsGhJqqWor9
`protect END_PROTECTED
