`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jIZbfAAtdzYcwxAxBwwFkI1hQQbOhTv//zrqH4mVDDSAGNWAWrhLgl1/ONac4qXP
RDS/zhf9PS9Cs2gYEd0f40rXYnUcOk4WExe+XY1VJUTm2SqT1me+YfSAu9t+rnM7
dap/e94JS3DZMV5kNmaXjp92qjFL99ar6i049zSMFxivojf+7eDkYb2RAapMoEuy
xBmZpjfJ2jXG3Lo0nuACDZRzJm3niydfzxPCUuwwsGkV4WVAz/YoPn1ALi745ZGo
5DN5veeHPIH/xCgOANJ67entjZyxaPR2d0zaSMqgrJ6cC7EuMh0e9PHaGptNKT/Z
ei7C/iRZSuuE+d2Gg4tgyyTGyPRb76CNhKqJfiFZzFTCOErgYMRcNI7aw6V7r2ae
CtaG9R/gS+SnilVdFbqlIQxj2FF1mpcMWrYlNfHtEZrQZlMZLoXA7ygw7NKCkM3a
phLTJWtTdIeEnbnLCBms0o1M7bThPWewOQx3LPo0vSWzOdoBwXzTosBUSoWuMYp1
xuql1EIu990WVJVsH0Ray2y8bJTx6yaRAh3bJ3Tmcm7Cm1gmzbW/PJWwfnLkCSzz
8kwEO4dTLnQ1aGVr73auDJKo/syB5m6zY04bioZsxbtFicJfaQECeip2MoNaaU9J
F9PuAxtvUY8LvPrZTyMxRbg3XbNo+ugOFxRKTyA1CtJyz2P8Q3ynjhEhZcp0QNOR
ynTQtSxLCNk8JYLKQ1EsLWYF9XjFmS+20jAVgf9RQUblGClQ2Z0m5VyGX5451gL0
4xV7vJkTvcn5ppGsBfYgYVgP4Q4+UE1LkcxsBFnzk0a5OU36bduond/gT+FtJs+O
wzo9SAHHF+lhT7SmKUgxj9q3kBnDyGOY0cpMRIHBtVhqvc6k8EcBoqGd1RE9TOJu
lYWs8ISdzKKRPndD+LL5TpcXdxV5kvPoA2XrxWgTT0qJ0vurNoYPRZo04yDPvKNi
pxAI5Yu3bI+GqVzZHTnty+d+70WDVA9ZYRWaW4wMHensv1Luh1FW83QDVqvPy3W2
Pjwl6xMkJkLwoAEGO6dvlLnnwe9B5kXHfq8mlapumExjsuVtAEaAtd6dH87AlNDj
lfskRGp0NSq0qalI6H+K/pa3pSoQX49nkRGy+KMYFg+8zYUBQvryKOLl0Ler9Vx/
AOcdxyHmvNawSgZ+JYP9j/DR+4hFnrK4CmnR1PnZQc/Jsd2HmrsbVo3CCBxGvpVr
Gy6fQQ+jv6IhcNCkKPNSmBFJ68D9uOcrUsX1Mq99eHq6HpYc0cMWa2S2lBpZ8wU3
8+znatrcqsgvNRcRWi6g9LLWvarWvTW1AVYvucMDNXUx1hmiSKEnHhn3FdAuerDL
J2qyAD8QtRoYVuvg9dCofiHzxhW8ueYc9Kw0S3UsvReFp/b1gH0YxLHIVCrOJMBC
eW9h7fJL5sFZ6XwDDElGhtJ6csgL9ddOw5jhEzghOKCMlEqLMKwb37Tua5QMKdRa
XK3WeiQ42Fo/EhoVy7Gijg7HTL9DslGRcObtZX2VHDhF8KkB/TYkgFno0mvdiWwX
UYZB11MYYwPZVZRmnZJsQZJzh44GxmCCWLFMtBoVk1OR36tfvAccD9qdG4iPkI7e
YVMV1OoSQb648wJTV+QpMPndF4hCgwfQjHQWFecgbVnX46g0x9BYNkRP6YtXGDUx
B9Dr0HnGJmyiDpI3E/hVFZqhAsHHN5FsAsiQyF8Lmq7kU7Bp1+YrJtgIwwgkbbrg
ASGm9wyyPbGSldb4ChwimrPj5jf4oAE3FI2XisApn74xce0gJsYd5Z77jlVnsWNZ
rOA89qb8oN8Xl9IyzDLapGkWjTtjCKQvYLjXtbNxYGcSQg0V/jdcjtHTHEVc3Ke2
PKGcIKNarIey7B6jkkBtFz6EbEXgNJt/NUAlyZbQc58eaZdPQsU5IiPEw6GzU9Qh
ribwuaAuL6GDlKUOT3JApewvBlGxsWfm8bLPxF9e+z13iCwCThaJlVNtvVhvgXtH
n0Fy1ViLMUNO4VN/TCB73WwAVN5jLx6KK0tlMhQ0r6ax/Skj3lV1iVqfzurEBlj8
TxQHwQuPm99ufHzZhWTwW5XT1skTEviHiRbUI6jy0faSHOOId9UtFM920cZ/pmic
QetEtKwtOu9mmv/aDS/PyhXAUN9mHVzud/KLWb01HuSS8ONIpRXmMK0qt53Aey2t
`protect END_PROTECTED
