`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aDKF6Oyx47Odj4R6V5Trk6rvV0BTqftlSQMD/4inYWJDRCpTR0paY/B9hYkx6REn
Cgk9wp4q4hzix8FLpnfTGdNo1+IxPL7s/gij9/6DhRqe5/X4m9U3uvwmMIPXI73C
M3ef8Bnx/SFwWR9kyzOGERtANtx6vHV7IV0xVw4L1CWeUmsxkVq4zJZzarTCnFPn
UnC8g1So7C/lAdedcFm8oppmrdf8+YRRDhiBn3e8BPgS8N6vDlVPNMpExGtfRBQh
ps5D3FtGzF0XtgyjLJJuPeEGdlKzG/8Eo2R5uJowllu0Jifnx1m5KO7IMNlvUisx
Yswwkd/abmot/fU90xksrdaYIR+FaPuE6X9aoCjLkmh3+MqYt+ffVOmjw0c7rZO4
YX6Zrn0k7OKWU1ECgpgT2saKe4M5T/VocpIYtOl/N/pahKk7qAqnuemDP8jfpiHu
/G6Ii1Jrg7fbyjr4FQ4Ylyosuu8jQzm3GdsV7p5sh+BJELCDqrk45O6k6Wfqd0Ur
Ej35D1b1utwsMw88HR/sS6DbK1/p/nS5gbKW+mdDSMT/FdyAjIXGEo+ZTj1M/Tu3
EqCZi5a/4TOHpISNGWojBuKMk8jRxlMYnqBm5/+bggEwIVD/G2QRqn/ZiI6flyM6
vRFNVLtJIJ8nzjUNpmJAWKqsCv2HmS7eXNL9LrLv6EJetz0bWkJhtJ4XPJwbmQ3O
pc9TlpqGCHIhEnFi6tfTNW0H1eZhUmMjN2gB2Nd08WZmD4vuuf8ONzR7Xw3RmQln
XCcw1jsr6mu3Cd337fUb+lQhthJGOmj5sBtlMbWqcBd/UBfVIslSWN0MWe7PqBlv
E/e1ltAWTFk+ABFC0jRCbg==
`protect END_PROTECTED
