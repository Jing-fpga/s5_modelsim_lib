`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jhp2EVX81Mp70tYPjyTt8r/vGyOQXCXxUgZXVPdyf56DBx6BwPPb4zJQVdUOylML
BVjKcdkRbWDgGASoRx/kEAtNwnTfyYaGnf0JCeJe3RpxAQyO+7QNoHD6AV9qiSJB
C2Abg5n43nvx4cckTXGhAaQ4pQEcmwjAB1XCZnWQYRx57ZCmaKOqlafJWfBYT505
QuWbUvG8wgIaZyX5qjWnpiyuz/iC/Kq5iWbju6JAhLf6LO+HBk817Zie77hNA+iw
jopB0cF4lB/IVr3RGOaIqsv3YFPlqwYdnv0+a9UqzmIObEeVHDimun8xW9OjWV1m
0QWv+NvGvmPE0lXiRQtC4CCT1MhzJ9h2ES0456e1fqb73JGpJwAbd97Rf9DQLlXn
oXaorTF5fxOb7BT/+J4FQ2dcrf89cuE5We0ehxkKnL9Q35rpZ9VN4fF2Z2NhtB67
62+A/lSCvVw7KYkY/RIjVvUbanMurtJDtWj1PRwuQANToQwM+DrcLBQlEBO1jsA7
dRemKLsCvKmdC8mCrM0pGI8DYylnd7wGTn/RX3p2fGvQR68U2YrnOI89fXgL90mf
TxjFCZ9qDmthjm3bk0x4jYtibZWg9h9n0tz1jEM4motL1eZLFrJjJuR1hFXABiyG
JJ2/uSc+sVr2FGpp+kc0V48F9TKlwofLzE1ENU0onzhPNgfEJ7ph3xfCYKvLqsku
Mn7azr6+1H4bj0oif+T0IvxsvUMM0WAKIRwYCCQKvgK5tKCy3fhFN1nEFpZhc9+n
SxyuGk4R4+yjHsTNCOSthZ4F4qNu9uHNAjkpc48GO9ui7xyolRdd9nJb5aZ/4YYb
br4oNNtJ4nkrcPgBULs856u5UfPBkWbXMmtOTKZFqxXSIPVgwHk0RGs6hrRXXPQd
Tlh67yI3+X6HknVnd0hoW5AQxBM5HjbdecYH0kukzUd+cDgXVffA8RV62sO90axM
NlAV3zgE9Cb6Y6c9Ics+Ek3Cgp5PTKPv6xSqNgB7uOFRIeQGEZ321eLNO297WGTE
TgdqI62L1YPu6PhCCGRvlqVwmcVPYEbVRhW5GWNclsJ5sf1AvECJylRySNxRvkY7
IodHC0GGi4Xz5Zun6qJaP5LYfbq5M9AxhJAxGpMVc7Xhv5O2dr3FJq65JVLbYIiw
8BMltUiAecoPOkfeUPXMxegP7GcB+vuAJ/Gpw1l9DONAPPjzDIKkhxi+R4cOLm8F
R2oz/HM0UT6z2Dgxi13iGMNMJ4QipqXubCrv7TQ1MQbvyzsKcTl64U6lWcduyaOh
yYhhNTQRpC59UH4/2K49fIceggqt4hRG0P0QFgKfcWpwsViIquVRpMGaCbJurMFE
GCC03u47HJEXwo4XlQXW7DBHc0vSwqBuX1+VplPupfv5EaiFTdZ4D+l09mH41Jbo
tz4/f/PTnmmx57lRN6gNuhCHjSZmUd+32eXa4nkZyzbnWq8XcCxoGCRtDIdHQKKI
rgmazRoLJoWhxWU+kSK2I5CGXQHYJVK2CInv3EJ5tC5fmythhKFmrmkmRAjteOWY
u9AeASihi+XYAcQB0VgvDpjVoPrQhvJ4w4sYl7izY3qNaDqxj5u//hiKWTSotUy6
+CZOlc/11b/7GjtoI4cK42/0JwxC2Qoa/McuMRLjLLerukZlPDUDzVRHxKd3RZte
MgVOdCI326uCuGIjpV38pTnk9Z+ofIQ4g+DZ3121xNUzDDkWRBFSuJryrzLWWwPr
XohEfaWSImkIl+2GET4XndgJ9phajdqVgKL/Ooxsm3cMtcA1oHTOjOMNju2n5UCk
2Cs7fjnih2XFRvTEJMzRxOsmuvXYlI7iEv+bDsiJVKFXqK6W4GPdwhR7zd6sGdli
W2hTIsqvHQe31MHfZRmHEJnORk/oUriVj5OckxJl9w/6DD/LGrXiMXYDoo1FYp4f
lO6PSCS9dpMZkkOhPJ8CYDQWOs/4CCZTrDun9Av8lq61AqCq50IfY5rIO5YU8dMB
H/k8Hk3Chv8r7MgSgZbzC/3A5UOgk6M15h4KqxdRxbKi/5Fve5CwYXqj34/fZ2bg
f8bfULYv7Qm2ri7tx8gWfthXHykW3DRuU/deXw2AxSn7dxoQlSdC6CRUgfh28swB
ao32PHCPBfSeX5cohjBafs5lSi52jbCm6NXFizWu9lT+AAj8C7kDyEpUq56ajAC4
pqzdnx8ToNIjmVycspl1D+3mVfLvBF9JE0Uc+2rzNsMpp0+zLAW7YcIa0kQtbYrz
tqBqqWZEuRspGKWg2hgJ2LZarDVRVSpuszlkCvw5Nlpiu1zvIILf3laQyY8EHt31
Bo0Oez+0B7FJHi+9XNgv0SEJOYh9ce5Uk1VfjsgGP/5E2NOQdxB3yHG5W7J4MZfN
qxcSU/46QX3B4TbkNOWXGEzT/nJsVKrQ/GCupP9V59GzLwBklBE/4QXPF/cBxti7
mSbm6q6TtO2b3J7rw6DISgRpJ55Mj1J0jwV881gqkyHFYLy3OPeRRHlzWAbG+JLc
2IsiakhT3AHktS30uspYHwq8FyHMTkvcIaRwae9qVuQIN4Dc/tXHilOAnVksgCpk
AfrelH35xR6uBExICDwNaeUD4X2xnkhBEnYeRWvE+LCvL3I8P4M9AUjtOrMHG/16
AWq5f073CYKNJ8cRFUIlz59pBNPaPMeUBuwy32ZWClPOcoQyEQ5Z+GAS905wy/mq
3a81IZDxgN1G4tUId/D+evC7GuW44/sI/SOdYaMPi5soMl+Fpp2xxo7Sj1NXzf1P
BPCheGu7IjjLSI5FFRC3Glsq4CjQWCK+wBizwhmCbInfVF1VDZqIP0oi/Nk1mmEO
Pam6oBzG44/8e2BROC04N1J0vE8O3rdlc6A1fzgriJvRQxOZZNWjIBVqs4r/Jmfb
jj/9eZosy7idM3uLYEU5Nez6mNh7Jk5mXY4qijUdjuLxSYLKtDYR2qsUOjZCJboN
5heGlX2JuQir/JLjD/AWGrzZWWqEb1sRqsqJ9Z7sCXjvK+fGnwXwxUwXMRj6nhYN
O4P4bi+PqZu3V+40G6LS7u3Lb8PDC+fvVAsa7gCeXhw2eg5deijFXbtU4E+XeBB5
QV5fZxB8hv6mir0Z9Ei/IKmGHtHEHa8VDPOgkDI8YXY2iF851lGRaazUJDF0fAbp
zQN4HyV4IT2XJ1g87DhiAn15t9/WDygCJd+uDto9TfqQxw17Do9cOd4DrZYDC7yh
LUM7iY2C60zrRGzZgLWoMgZZzRdfW1UHJAylyzvGKcVTKQU9kBW6fQEO/R2YFC2H
5zJ086S2us+0MO++baEvop7A3NeQT0+qCjlCVp+8msh1UF0U1RxvGE02wiSuzQIR
y3InLt29o+Y2LoBzIpA/jLHdxo5WOMANdnDqt0wZnSM4ORSjf7oc9AelaiNxTfCM
CHyUHZAlIeJ1JpKtfwrP7vuqpunLskKJwphVrncYRZWNnxhLQSQKNjkmaRY6KhGU
vHDe6Ci7T8W0DHFF1ohfl1J3kAcuHdYswhJ2ASpwYUpVLK+H1EMivc0+VSv3r6Wc
///HCOQGObe0ETTOeercKohbHTXdjJpC77Pxcz3KLOYpne44o0/KNh+GDJUh0ujF
Zx9dPT9wNoDOLXaR/Uj875FQ4BNUOXxbzmVpCshG53rEz7jiQjyGy8208dMsp1L9
vzfFetLiSoYApnxe5vM6nkdbU3nxxL5YCwAchLs+29fwjduBDlCSG1wkR19o6Bh1
x6OFtGrmtZMkNVQab20JIqpa35P6miN5x5e0ZVEYi2zmLDtTCNZor/KcHVqEzUim
XSOCLhAWmV/OHkQBcjJit4WatZkaQcUdXX5qU8VBrv4h8Hoy+zwEylKc0WAwa8O7
mcMZfMcanUWg82vec54L9IJrCLf4TAUB390BFkZA1d6GgFXt1+dhdtEiNiBdGJUE
lHsA1DuVdQCNp3hJmeLcSvNsTTgs5eqwsmVdXbKPysbUxA3DPICOGcpHwItegF6p
r5HKzI+rX9KFo0v3ljRLjoTaRfmtsxmMBflzW57L8BBVlwYBasfR56jXPXmsWDB7
45aXaWdcB2DQygNyeBCLCeTQ4/a8akoWqYRK/QYawtlydVtcSXOV1xzZ8RODmfnc
oM+SzVQhNiH88frE2J5uJD+0zLF/Qc8+6+uQmesIQbo/TaCKdhZXs4kftH+E2EAi
zRb1gndiTlPcBOc4WOjYEtTRkybJHTWqFfjybEOIEvlBxiJxC9LiFBH2tQ/SF1eA
1K18w1tBoHJZhyhRWcR1zqLkadVQWSy1tCbECdDHvLAInnkGbfMHjRuCswH1nHde
qdRRksIdDJEYhFsVcom+l8EFKpn1yPzVpQMu/JNmn8UCgF/W8B3RUVZrVt60X6u0
A9dFn+79mQXiKAP2oHw4U1VNc5c0CRBKLQHVPq0sGSizjV+h4G2+BptjuSnh8K/B
WLheBF+2UW9znLYIM02FZchYkd/Pbr5tNMeT7SUhvztbgHOmn/XqbZ02vmdEbHVx
2YSh8cCtLBb+iahYa5RocW7lq8pLAE6MHldKj8rx3J3qNegOktRgIruLZzgr2V0g
gZF49ysnT/4EV8YW9ST/KySvoMvdabVfbmVUPuls/FT5V6S9AHWrOXvtQKauLvyF
zckBDIy3dyw4a2GAKVM9oF0CJX5a06xNf5tbwmmUBpuipbIoNgyt1OYxkEndGqh+
Rdo3+CP19l2e9NAAi4z2omKhABFUR2/kD7OEo4BMP+m56L32cgsG/55ySJZH8M2E
p21m8CWjwW+riP4c4jI9T2xYyqGmLA8ERi4yy1aJTrNNOX8jr9jDTg+h82Vv2ljV
xa7EuoHisqA1LkdJZfYYk+TwzIpy78qdyJBCsiN8fNkuBZpY0BEKeM+8KQ8V9CYI
OJyaSZ0Toe7sJfnplMeNRO9q8eky5D+/1sE/SyOsJ+Uwbh1djMT8Tftj8guIN9Vr
alOTJF+QYM9ZHhZsTnZ3QmCV+aTckqSIU1JSpYCgeIRuuM0lI9zukzodrCn99MiV
pir5DfO/ezAtH5St5FQ/z53yEAcXKPwsUCmxmZL0s/2LxFZh5PmP7GuB0t9M1Unf
Ye8t5VEBCTAVyfP7wLLxIGoXAuCxXFr/z7b/NoZGBcQGR8QoAM9VmQhAMb/brM3P
Hg22rgj6t5K+Kut2Iwb9dkbF1Fq5M0yBUY/GvT9e6ukSB2rqcAX9qgF1JkJ1qiok
d0uOL9oLLeA4Yeoa3qMVqdYIyeG/X8Hu5JY+MlgvXhRMI6twjkJzvFg1+RaOho79
3LZS/WCN+yggWdb2QIEKf5oQzZdSdJQ5e8VIQDOa9XVhkvPQ67lHMe0nrkqx4Fct
+ENNhaAg0NCdS+BJfhspHo6+MS2C3hGGLCADoh2UOk+KGvqNGfMctE98vLAA4U0s
uu3t26UnyPrkmJ7lfnu6LWRodoefU/z/0CW22goYsl5g5kqspuU8KXpFaUz93JB/
voFiMHjOm8P0OTFwEHyZiHi5T+YbBNK/ZACMwkEsZ8Oym5gR8pH/XdIgA3/7Ef5/
knWm1zuqOMhsbJXja3mkJoxDDR+g28EbtNhytwfmobbmULlY7yg28JbSMFiTHHFT
agGVI7yhbA5PwOYjK0DAgrp5H52ero/bTDl4JLnykY8MRnpm/tYPZyv/iD/3E1qU
1JDZ4+UwMmfU2bVwdLUsL9FMf+cNuO/MVfVwhxK7BtToMU1PTQ+nfQr6WeiP7U9F
D94ck2+pC2RJo6CuKDOqEXL7rb9mZkrSqCZNO3zheGSnow2WmVEKfienVuSKRhBK
Tyj7wG6S77kGrltauT+0uaciiLOSajKOBmlXqe9TOCmQE9ciDcWX3DXmIsNeS8U6
dYm09eGMYCB6/w7OLgRMPs+/tGSuP2TIQ5NJbW8ihRiDNvqfto2w1e5WgGLyEEce
0yEPgA7OPLlc9WY/0uCjp2MeKhO0ksek2eWziY/V8UEH/p0AbmorCsW9QvzGJB8U
xRfhVr3oK2DRRRjjLeWTIAuiBpfo6KtYnDT7ll1OSTjfhI0HFfauot54Pos6luWU
e2EPVm6lD6DhIXZqi25FkXqSQZRp0bWEJ+AsHW1zovGf6Ui+PJAIbDPYTqlroPb2
T8Hyp+zH4B4Yr1Z5mY5zgC3TD91Glttm8TRU3KQT8Obqt9XoyPa55VhaMvnLnEiO
9/YmZiY55o8/PZpChGEMhM5sPzvgYnmdw/XRsS4yowvwMfWrITna48tzfF7tIUQA
A15JGr3K4TcPeXMX3yHbD+x5gGQHI7tUJHMJ14zV2BHvaNz86V1zv8v1KQbLULTf
GyldIeL6FKBJX4rzstK8/aXY/EpXUml/HcwT2p3JBszTk2PLk0Xz6hC9Y3Q60cpg
t9NOglNK8B0eUOTRxIx3jVnyl1EhBg8WnpWH/8jqj4H7I7zASYY1mLHExbnnz4JB
QWr7aQO5d5tWuFz62Pg4Rd9O3Iz4ROL2FMU1sqYJQljvcwBD7nXVl2QPe9Ks51eM
fd7WiaiWs4Kp+LmxsYjxyFT5dZf1g+ep1bgix7TVQnJQaLdKDnljWRbV6EL6ZJ9s
FwvSFhREgNPE8Ppoc0TqlGcPrsPn15z3OukMzLH4/VKYM8+JrgzpataRphRURnxr
1iY1/CH0FoUnxEm6eF6ivRSTPwFdqVn6BXddov+rhk8borv2RUJK9ljPQW0V/5JU
BI9c5oLeFgG2UFkjlJMI2E1al4AZRNkcJo20bCRvx2OkzNAk3THzVlz7gAMF6r6f
a/WYKVTWGFcm5MlPbETzOHU+HgxxYcH6akqj/WE72N0ktbnN6jlwaBCMCEdC/rgT
odZR4P4Lnlg9RtmFxInrATClo8RXaRObSgEaTUzj7bfKyTpvPS+M3UFkxocN0F/p
+YD/aCfVLB+h+q3iA8gUcFxVoQCNF35QPDJMVFkcsq1yYnS1qCgNHSvAl2iww0bH
iJKBVzatZZ93o6NqkfFWvpQ4G3+AoB1mmMseRve5HWzNHrPl8jVGXgaFHcC51tGL
F47CxeCYK4M9G47Wo4fxLEtxpXs/ODx1HPyP/v0y457Wj0HM8BSHjqgVeRsHgSHh
Deva2K5nd6NXOJniXH6NVgxszake1yRZU3fBwvSzSJsZTtny+Oh/t8B+lVN9RTNa
Yrr/CP1BdjOFUKCbGP8gRDmDQOu4AAEhLivrRqn/z7seUACGA0II7A50tQZ5borx
pMitcPDciGkwQwRdwMY9jf2m/0PKDzGb7NpqyPPVg+6KpaROv635/qLFrlcJ44rt
mrC8xwOU3wY+WAOugVj77lkYFdR3ul+pjrwdxljKd8qjvN75mOzR5SVRKYWZzH1I
bk6LSJ+usTAxYq5wELh6PlTMk+3RtHstrHyoJb/jtZG+LHpHU9bSeb0dgOWaILYA
X/bDUU1uDwNXN6yGCG1EJhBt7xxTVkKD3zdDd74WrF3SZ0XwIW/qiAd+giO73Roz
DhsR5tFMg77Wyp7+C4rXw300sAsQZrHtQ6W259TUnOE9/va8oUA1qfjPATDJCc+w
DYjfM2G26H0m/Wiqp2rVzon+40A3fJXYt++eL8XJMnqeM6yZbAliRHhPVI8jM0XN
hr5eQLFVXr/+Rig75hTAkKnjjFzvl7E5woRSAQHkYCqxqojNnebpEINNypuddrQ0
IIu2wLEg4Zu1nyZdwbXBmukiqkLuQ+W7NoQfitFPGyRN7p6Qm89f1QAzkIrTCowt
uhtLJoZRRDJ93qL7jCl9HPtc1IXXKTGjGBap/20u2erZ9rH74lh+7rP0GE21UMrA
NxSxU93iPG5C34qutvlAZghGkhy0AmT9cnPYWALT8EwLa0MR/SFvCAMWCtmvd2ni
xhg+g2YUr+XBMBLETdfnV9OQW9LXBN1KHZ+KKx5zrkWbKm+eJOH42Tvv9k6ufDdl
QGWu3f4ojTBS8x0fqOyCPcKjRa3TkbHcT0JVgF/xQfcaXId79YYfJH/BLsIqad60
rgX8/TTYagbkbMj9Vv29RguNuebcKz1YXCQM8PqUUOVt9AD80VgYQGEdZHzTSIwy
SWQdIZqT3noKdPRxDuw3/tLoiItxuA0fEq7D0Coa0h9zjPQPT7y5Ac0V97twcx3W
4M77m/pcb0JrjeZc8/j6yhJZ3IbWu+x0YtHajb2RX3GuLD1fos7wKq3aTeRNkSja
6S1DdeD6fdSm/FHKpHpAq/UmXA37M5i0jW32JdBiAA/5gYj8TbuHh2+1u5FHgbq2
1+pQ1SgX7gSYH7n5yko2QNRciENWeqQ0NBwnkQ8WyMImLDgXJCSkYvoiG34SkZUh
FEfuo84IOApb8iyiScePv3WyL6iIRF/wfV07u0T8t20194WVKrfONwIzvBeNPx08
kVmEyYig+hE/Y8+kWsecZaNsvlcVrtNVP89f67UlmDucOktO3L3bX8IpU0QesEzi
U+6G+C8TRPpVMm2QnGWcryd/EkO3fDurX/EYjt7XDbuvhh1ZEq7n1dwzVCjNPdLX
PRHsgu0K4mL6NFcIsmSkWgmPygpJQZfx6zfEovyKDB1jT435d60QjUTZFRat0Z3E
lcdGENsrLbDSMJZnys7ZTweviPZD3xy7iFDd/r0s+oMmXK+kHID4Xh95vRq4hrjj
Zgkz74kkAKjNr/rJiIQoszbjOyCGYILNwWjkgvDj1L4v4iZ6trd0dQogOfAxqETV
ZOHekJkq22EfszqGyMY0Vj3BXIt9es5NFVjOD6lm/L9RjOvb1hgISqrX7LscPawK
k+0fbmf/WYg9MUPNI3aU7FcjTFEbKqT3AXH/yObcQ/hsDA6fyDs42NiPekzTl8fo
cyBoQI2eK+IRJDm+rM/WYZR7KWAhlvmlJWSVLO+eJYyIdr2J9btuJ2Eipsb3epyr
X/03+gUcjqf+2Pd8iU9CZLkq7N9Go5POsyc3M1WozDcIxEEKs4ecEvSsdw+t7adw
NvjRHWk9X8vYHYfxDjWtPUcKk2f2dhqexTq9+kf63Lg8eQCie+hxOsQmcZ5jnsjE
LOK8TFb2xDOkIiAb3GcdPSGzq65MGThMBBjZF8wM/VL4ZPDLPK7n1POmFNZcUy3E
hPjA7gfBrp9/nUl7WrN0fkaDI+ifbDfqP8hQh1EGHnFQk5stK/s9yK+k/soZjb+b
hNSdefMCACm6yiyvMahR6M4cIQ073injpL7PM3dL7RPUEegd+RwvyShzdCq51oUz
tKub0cwdd1fqgul10MOaCyqf3Q0hRzC3fAYN5ajwuhoVFhJ7yL0SMguUUrkg2VJm
xXnn08DYX4C5OJrQaJkyceTshq7kjvYq7lYwvuuVAW7HVL9KeWzL3lzln1QyImPN
z/DViN1XC1VVutLEVKylaw1jOMQ3wBVB5AtN9LQn+NR1wfbKg3Moy3t0yUx0MRTd
jmGNxJ/wFWy9kbQggNLBM8XF9CWi86AEBYtPiB/tmq+lOZWdIusTAXXdLVV0ulOp
CnsbikSlqt9IMX1TNPpCy8IRVB+mved6s5CnpfxMOtjx+a9ElnkZYCSgGw0SE7dK
tK4691Aq4DiIat9+1HNyp3dmqy2OPvHz5or+nvkoPCbIjHNemav03izpE33JHVNQ
nl9cjRg9pXoMX37FzrS1lZsZdNC1Hh98v2WDV0nZSs15JP0rSwrPulCFQsTfZjLg
7JTysnYFx6blFJm65nfhE2j1GcnAal9ZSLMoovqtDohseRGIJTLwRO3FOabCLjTg
Jz3pUV9oPI2n1OAYHp2r0lP8foPFYJGHPjyys/gAuP8mpE71/cA58PynSKq5uzFe
1kC4F3uOeLdRW/sCziRlcuHrZJlXzQnx7a7+OaLjMGIRXXF21lEBFvJ1/UbOBda8
NMqSivZHDzpYdeZU/Y4KzIwH/xTaJMurYm2lBysEW8bJ8xzF1Gdr9guawzqETUT5
R5m8WE8HsUNtJ6ZxhgUHaLqtZzwt4LjLWhYXSZKuEzozS3pjkY4kiIxB7jQ7MNu0
Aglud+wsE+rTaAWPlXcW1xi87sn4V0wjCmnmcSq9gfC4F59MtwQBZGVlFCwd8x7g
sJqmOKLBLo5g1MdQ1QocGyKBvP6OEozwmPO9Se72gJyq75ctlnqzAmAQ+jO2C6UP
zG21baRPWFRW1vMXVTvH29+oMpFQ+Hx/8sBgl6qmRbxilk9uON9puzfqriuIjfWx
SpuQ3wSEJkH6yyNtJUKaqXF5oD6SUfgsU5QEgkndWVm/fVjZ8jod4khjyNZnU+mn
ZQMk0yWb8cnFYe7IQZblsfYdfPpO8rctvojbssWHb9viC2YVTtPPpkVfWrSb7V0h
cc/izzBI69tFf4B76ET8NjxJI2e5qSYQKRSBHANJqx65BDXaLbkKGBMhad2v7BW/
DZkJVuzDSVlqe2dG4bf8YT7gvoQrn0940wvyyXxyXVJxa07Eysakul+HI3guBcD4
u+FFN2SfsHSFxbwdxHVxAiVnnq62KPGYTLWzxAfOkfn89WI7CntBqSkPcy4pxs2l
SetQEfxCTYmWouKuJ4sEFw3GaICyKfoy7E7kfvfDMI0Lhm5xvJyRhc96R4HYxEGq
UZnG4+KRwY1fiQWsqRngl9cg4h/zHjijiWZGvKYuieA5RZCW2cni/TCu2qoJK6v0
x1HG9gcwntTOOhkNKQm5rNyKD72h2M+f721uJgHNgRH3A7UAdvFl1gzcp4pFuwzB
6Ku1JdMq/2VDOlyzFr5SkdFo6ZYrjsh9LkMhj+eaiq0w3Cn+sg9H7yPYPMJCeG0w
3WkaMChr1I7ZvadY/Q2lg+Z4ij6QThpiYsgmd55RVgPewd9aJPHH3pajZHPATkNS
WDXop/ZLM9p9OcL/ax7QwZ9KMNucl4BqWOp8RdKnTyNmKeTdAQTtkaT7HYjurvs0
duVS/8Rt9TU6svn3ju5H4cro3EZ/tvCwwPSXWTPk3+CoOFVC0M+EfI8NlJeGnkFx
99AF9Aw50tvekyHR/yI09HPC7mFqnOXbfpV1AS+oR/MPqIpK1erXhS+jIMWLFKQT
y63Ti6ry5SLiS1pMUkEYdWV4vGJc2bjvFhwTxjj981kOvBIZj4WVS4tToq/+TIv/
DU3bYlacXjfpr8bCwFlAMU5jYWyxgI2BFQVn4cRcZemW0adBfH06F9XBBST/kjcY
LgOPCIETUpR2jQ59rrIYHid/ayTh93Ov2bGWrqb7qhpqSdGhYDroLrlN1/omUZmd
28rpsMq/CcHtwtVPHwX1uqjE3vt9PlZgp85AY6V2+YDyeAOxXmyWMGoDZXuDzeXu
imDjGhybiItg6hCIzRVmN3OlyArbf4jQZfSjK0mNpg5Jek+9GDwnhRg0UUML7h6+
1NFpnzsb/1u75VV8WfcsXfpjEHIoGlZpSRfkx8IfToF1RtlI7G8cBmXWOM80ROut
2SWijwU3AJRyMh8f8GICHZ6L0aUfH2OGQmsaC7qMV80kZ0bdJOMG9M4hDVqJuG+E
gvoD0ipU0lMjQ4XbVIL1oJJovAVlzZjJ0ODfpLQm1h6l+9APFf4ApEyFNYNGg+IT
9jDFWwLfgaZKisfmDrfw00gK1/PhhkQc8C0k0jcrdzMrR/MfnLO3Y4nywNDo3O6V
wyR++HOzO9GkkwJ/OkvT0qacKMeNvjOrDLE710Kbwr5DRZak6hfwA+/EpNpqWNe/
Xoy5gWn7uJa4DwmkeEhC7+R8kqZFOofz2ZBBGLFLrNWBxqTzsjtYcVJYKRy3SgZh
oy+deAUJhXt6j2f0O0QwrLdsTkv2sKmc5x0uOn7Uo96Ws5oRxOOOCRDStrbNpW/i
D8WbP2Q2Ekf8kNB9kZcrXGkPwCQL/PZzYdUXbkg1t5y8cZrSwfPqu4Hy0tnSRqDM
DlLXRfYLFGIgdyB53hLn+paJmZE5o2H1B2PyIag68hqt6YpEOfCvgEYg5AJBxd2X
Z6/kBI3EJBZLUe90Sa/IgH4h9NZHe01xcBw3+C5XbxQ1aGz3xWbAKSzeTzZMG/xF
6KfJ+TED2ZNKG/2Th5jgzqklMT70fEydObSCTWGb7LfPKCKYU0ketlYH+x1QXWKJ
rQJLqnupRCRE6P+6jRmQnbXUbA2B7TDcF1VwI4CAn2qoRLo2VZgzJsVLDyjwh+SO
QGvFHK8t/2UO7fiKi+E9f/qf1cl1Q2Bz07fjTk1lyJXWWFMc57KqAxrcor8f1q1Q
xVX4c17mFjqXwF/Awh0LOC61T7r5zEjHVm6+mwzA0z94KkNB1xlI3Qs2JwKFVS5F
PTWyxTuhRtF/dwL7Rsw+oP5BbHiIPQjWDau/SXRyT7KZIkEqLXxayImOwOtIdNIS
w/O1TjBYm/riw13qvH07En7MX3BjpbPstur07Ccfz+fQXDin0AmO324vNqBb/5c+
gT+5X2aQ7n7+ipUZ+CmJg787qy4m4ruxRsMr3oIv8FawdDYT/iO8s+b7PM1YyWeQ
1XwapnzM0ZLsZSXzYJeBg9wP48cTi4zlTsbDvT8sE5h9ZGkYgxDEqlIxIagbq8UL
potBrDFmeQGZn8NpXKIouIM+ZZao/2LM9M48WoyqfHvxlT9tNkSgL+BSCDE9Z2cZ
GLjZMmuqkcSd2yBbH0FhqCzoN/gKgmx+tCK5a3prhnQybcDvhs1yHAMiLis6FSrb
VRcVbdAJrH5Z7GEB764HG015nbT0wUXUsN/nkUz02xw+wPkCCPnom5txp47Y1gA5
SG7mE0Mh/jhWYENmPrpXWgXue9eXJOPHY/04k8t0H97bqljND6qL6eD8UN3pOsbp
tUPNArI3eskhTeURcPvLT93HWHWqaXd18V5vHtM0HxMoXuTpjJ0O/gyEMmifKNXV
CCS0UI9zZQZMOJfHdmqLFmv9HY4vDDvVa5dNvtWEAp/2RUTAUYQEM4fAinFmW4Yk
j+Ml0cSb4exMAGNAtfo0JOvNvrXhaFQ0OlnShWPR6/UDlhmxexab8ejrLZcrS8If
piFFPc7wv1nXM1kav2n03vZP8SiDrcXkq6TlnWyYKbp67lCQDAdgMqerkL0nysPB
kiVf/GTV/PS3P46ywSiF4GmyefqW66mjqolO6cogHp1na+onmaQ+xvImoIxdpIr9
OQ0IWeOT6C81EEch9IV+X3OtD7X8zVjZg0/qQllGStCgdqKPehLMWh/hUnGBF+QC
VHnZLJJrqZMXu+knTtWhiXxonPcp5kk9qheokOV5P09gYjK/NhV8Q6qoR2poQ7Ot
LkkrXpOUvv9vstojPh9eE2I/QY1W1YGqbVfoehj8qOZQpaDFNkIAul57FJbUj2PW
ldXrkQDRIoiN5cFedc9UOD2AIU1tQgRlbpDQ1FK3ND3aCl76FkufTjrxn6rhSN8r
vcJy2iosSWvge6j1bWfk7JhuZPatMxO0j42hWP3KoHLjtRMK4hqISOKuLpxEuqv1
AASxxxicpqsyR8mdumie6Vn5tN6LQkQsHHQEOjIMtPoonsSie9HsomhMXXxoSgBR
fvMWedr9MFhzd2A6hf/2+nakDQilBlHI3ZBXu7gMloriNH9LA0V2NDpoj+VoOLIq
NqKNRRKUqf0oNS7E6iJ7ue7let5f77ExUDBqP989kD9+dqrrWZt7KJvNyvxp7muF
gmuvhZgp81GnFXoKDtABzjqvCyZzJqClyGFXhO8CSEUsanP5tIVOvlB4kErS274q
OL5AFLO3awUk8fqoPsebRdEvRL8U4TL70EUOSw6ymG70NN5ezgu/5h6n7IWxd1ee
M4l6S9B51ZOzcyfqvMZXyTZIYrZM0p3uBUV5Ogv1iP7R76Ch2ynbJT/VHPoHCUUa
YGiL/4u36bqaNy+BdJ5QnKAC83qbmxWpANlZK8pRdYyoT89x4VRkB4D0bCBhUrOH
r9VHvN9RMr2WnzZohu3PPOUvrVPDOqFYN35Na2cMC78xakZQIjywnE0qEdKv7FfN
YnfrRq0fi9KKj6214zhaHJiDblLayRtz79j5tfJS5lSQeMXMDgi9r5WyDbXt7iRV
Ie4eGkUaCpZL50OKaZ+BammcjX7BBuzJTEfva20U50rfStm2A696J0dcBy3eY/xC
dP37vzBcHEwGfP+N2FkSnm7wY/A3Vh1Mrta6hHxd+1u4cbOAU401Fa2A1stY7aAe
JmFiq8LOud/SPClVKYIr6PLp2xxBLBWtZwsttW7Y27oibbM/KCaX1P45ACZHt0iG
CggQe8dkkMnaC6foO5ETB0wmAobGlMMF1hvo6mnTToxSTcHhPirZxFk9Xc0AIc0P
+hXta7q/myjALZRnwwa5tLZZm5wNWjaV21sVO170R5XXYh4XENl9qkpQSIYkIDcv
BxZ540CZVs93o/nSnCoqRSFPqaoVQoCyzaWw8dcKQpxAq6ZtrJ/h4vyReu0EqPgW
P5zMRAwHyzvk+uZIsmgjSXkIULgLIUPeLqQ6+1jJJe2HM3gdaod6Llvt+u0USC3H
5k93ubVim0GhbSQhRQNKxRom7vISqAg8J/jZv6RBrm3NvGKOIssMVa757vYfiN25
ruCjAuVtmAY4xCL/soTlNenbmmnwZ9GGRdkWngGxjrH3DI/kkkGZ8q4SUVJkJcGe
PbK4Hd9/7OoKde9lptcZeB0g1bLFI8+u/8nsRPjrnlASask6p7XPGXDOjAhbGk5B
/DA2t/zkoPZCwQs1FC9xCX3xlBLM2ntvrjoMHbj83YHumxSQb89EG2gL/d+MIHm9
gZu89R1wSQNSFPxcV6cmdzKMuDooHBPi39QOWB00K8cw1OV8q2JuTqMwGpDTI2Tl
aOsqChwlE7ebMRcMhX+B/DjC1gZeZ0P2dRCVurAB3lPdLzfNXnTjPtHJ+D4QcGqu
hzj6qzMgp7FkkdG8RdlhYDEBTNtNOUIcsfu2rvTRLt2KVZkt6M4OiloiChRvpGml
wXhsmdLjj9givy8hN5XRvMcLHY8opmmJwXJvZ5QvtMyrJnWSO1VO4aI2XR8TDJTP
LR3GxAPgtAzE4BBfPdgJJV+TwdZup61j+ollvIPrARMKOpFFxua37OHSoUMxsCBX
WFeE8ReA/atyRxBwJ69o+zUso08gM372kFB4mL+njqNgH0YlpyUN1K9NQL5UYkKd
eQCDl+KZ48AyE1aBXBI0tsE/rOhQZsW/1vcrFy4RYXlfniy4S3pxM1ujjyBiGR9y
Rb4AgYCqRVSNLtLMnJYDipwo8C2DJDLxSr/jvus9ayIS7oAeUw3TH9raPbAnQojr
uwk5359kQ9RlJ9D5+v5FiKdqQwY5y2jbwRl8vPrp1Y4VGkuMDEPocl/WQg6r/lxO
wiBJ55TrhmPXBi0SbLusGWRZNuEUyxCtUEUAqDRrnKFKxi1jrk0Q9z84JRo+8+CT
sfofeHtUBka8hEdRA0yoA16PWGUhi9NR/urUVwqmiCNpOkI+ya2pbAuI20O6Jnxa
3Au3KAgEdnitsh7JqOrKkyfywVWrbOr2Sa9tkpn58CfCv8wvWVZEil1fzLeqQ2w2
grjgt28+1UuM6FhFHGyis9kXXXLA+IVCm74BwpbjoT1VTzlN00TLDMc8nBpnGbxt
oGyaPG5qUzJrdB+4Ajzwc/yeb1AzDWWiEQ15p51qiYpNaOsaJ33wRCGsUsRN1/3x
EtRaSxxpEWJZ+TQ/qGQMsrxTbtIUuwSAc6MivH1Z/dHE8CHyDH42dctwrcA2gO0z
SCJr3N8DXEwEhNbUNlbVGdTUlolatXdx2Ut7wDGH9ujyS/XjoBxJc3oe7FV5BQ5H
Bw7a6gigS0Ni25epsXZ2ZAspqyrMagPKPgLJ6zYZBsfUh2vCcwGVqpFEoq6XuZHX
ysVzxeGVy4kMRv6Y/w3CpWAGAXCw4jD5QWswB9U3gGc7Nx+qynpqncbd7Dbi09Pz
h62SpP50jl8Os7p+VdeKhI5yfoilJ063PHjtJV1ZB5viYZP/IGjmywcnsj2PfmBw
u8SGctv+pqnx/IAS/h2iq5DBxOanLm83o6/9IptQS9/rL8qJE2IBzXKraVLls4qa
V7AQH51P5AwKeuBckjxqwFqRUB3PJ5jyFEXO6sGXKsIjylfJuUJZvLurpNHygMB0
isD/oGkzgaFPrcRPjzqTX46UZFEfRKRi/BjuxIj7pRbTibVAmpHOUIVB50y3Nqom
G4vZx9qDi+jH5QISslEzycOoKfM8V7Txj1cwb5qaN47kByb46Rq4b+bfaSjMrhYW
rDNz7YTKPlcUVYzfmLwG9LjTCqBWJVIJlEc3T1Ge0q+KUUzw9oeVfgUsivobkn53
+88Zhn4mYMImP0ZMQVaFX1ceARvlFK7S/3FCGf5CsXoZJ/v2CRjFL2N0WwVczJnu
tiTddzEk3kzjUgsBSwrZ4hAhCHpkczWfi2Shg77cDKq6tadsttN8ussM4RBP6gZX
GmHmnuYCWcvsTpC+vGg0AsEvEJ4VWV+f32VpRbFiYCiPXpv6fIDp947l/stzTe7g
fEG4doeCsCpD7J4hRCBdJ+BkznH0vepVBMK8NX8ThPqylJfQpIbVzVspK5hUrY+B
Ilt0b5fnM72N1bVQbm4GPk8A/v2dZJMQyIRyYdYLvXUj6qc4kluCYqGx3CeInNVb
dVEZxXy08bXAqGUvbYz02Ipy9oRYM0gNePzk1QRm1ruqHmYjrO5h9ieVEEezlGeQ
x6VGNJuwHYB2SIPw7vu9XOljE6+BdoqWUxklOJNx35zn1OfTK+CJ1C0m5Kf7s+7i
kQxVJxC2WB67zOX1xbOtaxCNhzXuqb1QMllaStu65YVgl5yZaF4WvYd5tlDVQyZW
8LKbDhCPxw/g7/+7sGK4P/5JNZSgTJPOegRdT97Q6BMw1SNhmgJ5Fruu4fr+Jjxw
mua5XeVG1rTFzyuJP0xD5a3vorkYrwTixMWORrOMYv+ChlEgjRisXqwydtFWLmbs
uZ5w/PhfilmN/PXA0G2sGadbavho0SYhsZVFGplFPkw5QH/CGhf0olhSjao/JdcY
U62tAQMn2AgnXXwGlYKxP0uVq/9JX7C5HwIOnlp7CEmSnTOqKosIyXbgkVM8JsGk
Uw31TD9da7dtnF19Mwa8vhHnJ3rXjopDhv/Xr5trxj4M+W+8/66p890KT975brhz
vn/n62b05HsDrt2EBGsu2GgsBFCxKueWzKmDjFd5Pu1Mud31sqcR5M2m8aPbT023
uy6RMB+UuAaz89bhpvufz4etwymx45lSQWXnbGhBZd+LPUJlppYjD1CM1cKPQenW
cEFIKHgwL6kua+FzBIvfNg==
`protect END_PROTECTED
