`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/5h9ay9PTO9EHuMsUKnWcyDYXVH6hLXfYJxaE9P6u4PkHhsa99PrrTLVItH89J9O
FBlr26we7k9pOVj5N4DsvqQNxa6FmhQBd5bN2jl09uIog79AGZjCRqasd5tkxvxp
v6XbxUGBrmn1ukrAWljGGpcSqSLULJsc/DaasoGoqT4+JIW2fpp7wqdrloHXsFLy
YDdw2uDzx7IfzVLy3HZrXDlG6RztAUO2+2KE8xomEgOQrJe875qNw58ufY3mCXOM
06/OUaVMiUdUjYcYGI00FNWWPu+vW0adJI+v4PJD57gM9X+NYqNZMnJFmhppXuNI
tvadEfEa7/B9EZLuCZynoX6/yhAkucVWNACTumCPh5+wHvpW3P2/rwNgvHFMiubm
t4Wy3ddx2esL0NJeyAjRKFl7qezeba5cW7+PrDqAkb5R4Xtm7OvpKtZOyA5OJu/z
ZYv6gd94EP/3uOCf+YeXh42zIAQ/6bLKI8PYpBTxwXFsB9byJHLkrmpPkFV3PqWP
lxyM1l/om05cDfj50T21bz3cH73mj33oWcy84T30fJJl9/C8vl67cv1BuR4dr3E5
jQsX8yhOPLmzi30B6dqpUr211EZ7X/XE2K/6Qi7Y0IUXk2DTQE+kkIgjLWMPmnZk
RSYp/pk8H3msLZscpM7Wfooz1T35j5nDFnbzuwpiP8Pr/E7fzciKDx7oZIQymp05
pnE0ZXkAcQPl6fLCnBXf85k+YT/b4vmMf8DLMe2vm8Y=
`protect END_PROTECTED
