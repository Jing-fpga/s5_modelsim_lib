`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MzMu5Xn2qAjiawmB4iw1C/GibBP0TuXTRQCrsu4n9X45g8wLaria/fWRRnrMfT/C
vUX3lrDNkGRdZdjchnyGs8Wuk2cImJRW4kVhpExuAAaIq+blixEG18SjoE4xqhC5
9WJFan9tr6ZG+i6rAAEOPXCWwAEc6rhrNxUy9xfZ+Qkdz5KfocbOz1ul82lkZOgD
7ttEXpxZdsIvntFs07aL0vPKCmE9lzyJY1J3CxY+ckuEX+0ZsvRoxkLEPXo+SYZW
egLP2LThbwlmlrkU3rm3m2P+mdL0UQPK9oO7UyScMwNbSV6aSj/ke12H+8Gu4Cal
QiBadfRYj51BKVqCBNupM2UvVp0PVqRt8PSWQFZcLvcHjpue6h6Pef4qGZsPvQWf
dhwa1ksI8DAYx7Yx7eTcm+K9F6bOOiY243DxmixkAZk0q9m63PN6wgKuwoaOSPTz
k8OjWGPr+w1yF8PX8jrqldexvfyKwHcu84MbwwIluf6Wj3MgFMv2rnHduB0pAPM4
/1vBo4YsZ7vgZvRWX8U1Fgq0pTZhwBl+t03Wxktka0SeAQMjjf8VSUprauMryfn9
gIsUZrMKLzIgUMv9jslgQpIr533/zUQRj/6yrItk+ylKeYBc74+MiQYUJwzR0Otd
jsJ03PqbZIesi+/cwJylTl1ZgDO4W5QOxIwyO3IsVaO1AFpw8wKvksLXf+khQswy
LstZwHP+bTifHxDKluTHvzqNjXQ8wynghdhJLdyxZDcjX4o3GMHzzEKIH73b3D4P
NFcH9FFdgD/3egBIACG+3o8/GkRlGhVSlIV40NyO2DQ5fVUBWPv9Hunt2TEFsLSA
OUlw7A58WOdz4BY0Uhf0QFIta99oV1Z9i41WquRxgswmIWwuoROPksQAJKQ5cpKB
kfcMVtsf1xT+XdlUDandLVOdyzRgyuC146ydXDJ4FlI/eiztk1rlQkZ5VjbhYNY8
s/egkwK8RUlGj7AsWklgkvCNtFUiXw2GgdP4DF10tsBYbhH/UyzlSKwNVKHmF7yQ
fWtO1sZhjZPDjVqWPaGReDxYz13+ppMkaOxqZ8J4RJU5M5aoG3yQyj+Vz5uqIo44
6EmTuD5tn72ZG1Jd2QiC4ZT5IWSVP2Rbs5up27rvgwMxY9mznuGbPDjFSLLzz2Rv
BuFrHUjkpxNKtJ4rb9xgZUw23+AQh6u/xVbbhNPCaEKN19KCHCqk83NNOKhopjaA
gayzTDZ43pb1dISJWTjzaQK7y1g8NFmLe9BJRJV0qMEyOI1ckn+mAU6qVw6W1Tza
TeAdc+k57tbPxcd+mFsNDyfJ+vBkdXgfrbI0337eUUfxLfBNbZuIbz/QW2uVQ5QP
JUnVQvdI9K3iyjxHNNAuq9WlWeA6NKbT8Sgze19T9NuISdUDx/hnAs1mLQnz0Dm3
CmC054qI7a9//vLS3uX4bWFs5DW4/aJhBOiUHvmKaSRKv9aW/FqgQPi5pShXVPp4
gezsdj47sHgv2b4dIID9QX3/FaTxQzEJB4hOeGa3dly8YInn1Cqies+eVr3kBtyD
0vD2GAbt11Qrd/BPRkn4ol1P68USvQIEq05Te59iXx8++3Q6VTfr+bQAwDKyFGEv
QSi2gwTHA41MM8IgkvG3QOG2T+RAr4ZoTF4LJY4LQe2PxPUJwBL8MYdkZ3TAf1jo
od+oWuaRI48K6dwzb7tkrt/BvEHSCPf/r98YKoHTJAdJsIlFiESOfEIyF4AV53fO
RAwx54pN2bKIEpGE+FrlOZq/hB6cpdCpp2ivo1Bobq8VureSIHYFJGgrG8J4T9dq
A3kgir/Ov5VCg0Sk9//QT858hVPGoLuzv8Tb781vsxVrp/PwPWkWDa7bUfvegrlu
CU4dn3SU2rmbbtonlt9Jb3mdxrAnYmCy0rhjgPNmx8dsjdXpfCwYZw9Zfx5ztkAI
Cia0cqvkrUCpzWb/a18qMI6gKe3TxAT4/StXHHGWwBe7BeMaE+VzW+5ZvZiWZFBY
zCFnkRkxQ6hlgbGo2KvKyg==
`protect END_PROTECTED
