`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HBuE0XrwTETFbwRl+qicPXHXNBMvRwvEIRWCEhgaZXBP3dJUowndzjzJXKAHLfOL
LaLREqTpMFo9NSlAN08L6qieeQ6rtpVe8/VELVdtCK2pXFSfNi6P4asnmF3Og8CZ
FNGYAuQWp871ntRGb1/dd9WLIlKZ8vYYoION2vVwZbKmyNbs1YBWBqmwycFOEESr
vV+OrlxiNZJIeEWy1MQIAUm5ClBQdHTHNvhTK9T1ZqZ+k8QRemZDp/IJdDjr01Ne
aLBzYUaQRpbMlQrjXfCIHGU1p+f19fu9GtFN8A25Kuf7MsRiAxLWUnoERrSyjWz8
HYiAauQgWm4PXarYlWlVG3aWdPkgSHBlE5zLS+2PwvDzjRFJeRu39iRboKxkAqqk
Cg9GjlCYbaWrrMAbDX/d3FYVf97KULLyw2ickKIOFY5ZzUVb91h+4svxYGZkbcrJ
aX5ifPrpLSmK17R94glWA9BOW7up0mgf2TSwbYktJvugf7gImyi6ImqTkd5mc2xD
WjJJpWwNMmsS6La5M/QDsCJRGGUM66D6OI6RE1IzfpzK9Cr1QqX9QmS5bHAAM44o
QH+i9BEVI7NG8SNnZJxD+c9hB3ibQb95bOOJg4H7CuWkZviieXKbbNIsLJKFsWOl
W1CFZIP2P5UHQX5gkqhgOrh9m4IWxI2CyEhGEi30DDP3vpqu3tVx0HzqYcXV5pj8
ccetOg3zSfFRxUbYhrL1omjkAQXAvJ88v0fYiGd5K2EkzTNkqzrcOrjDXU+mT5jQ
g2TeEHhk+ehhxmPXoX8Cu2MczpT5wR1SuxGNjAU6aNVgi1LYJSW8ZaUevoGYEezw
HoXu/BsyegVHxpDJAAJNCt7S6+Del9bGrfm5cffRLAM7t83/6uya0nI41rMQXOfs
ahAaYCW9jfreAbKQzxG8bKS2fRYRW5FcwtNyVHzW23MRQcV6F3rhsmwYM3BQuYV5
ZgyjbgVmLCuKDb1ZNLVzqQ3N0V/QGo3BCkNQpmAbGp3yzZo3ZXHUmB7uTxYx+4fl
3VI2+ktgsLs2/6oNyVckJjdBMs8cA4zn05NCnYZxvNXw+aZZv+ip7RUfqAxf+0ly
GBLICiWcNRn/thfV4klMONZeXbYRMq8fDiqtRq1I2+SuCG1yza7f1Wbb0gTBiV9V
L7VS+gcLIS+/LcAKxdhL1lKpfA4KSQDxQitPAWFhC70GT6Drpt84089ekUOgYM/o
UCJKDIJiZkG6qDY+sxnj5ymfoDC3eoSBy3mdEG1GneXuc/nFkUpmWO6OLzOUMAfr
zkU+6RfPax+vefcBwCNFcqwM0IU83xvpcvkCw7tyd0m23AVxVZSEA52c/v0LTZQY
bTt2A4PxBQfLDLdUePCN1+Pa7ImmtTaiVNQl615e8T5sYbg7EEsRRE7u+9osBRGg
Yf9bIgL233bylG16M8n4tOfhkn0ge+/fAH7leWbu5XGjUFDJzvnl6rsSe3MZEYF6
arEAxp7MpCdsUV9hyeB4TiXfqEIK5t+Yuse6KP+msIFPXzAM7fOCFAHQdPKoaEZx
9vtdm/1fZfRrcd3x0fYluJ4ELhIZw2Sd1pFPooAQ30nOlIJq6KJTdC+xUXRf9lHg
wIEj3Xfc9LRQpUL76yazesO+Q3u391ezXaW33/PBfycyDGzs+1q1njTTEhlkl9zj
9w+mGZ1dxG2xQdGj4Cvg5O560V/b5+rCExs8atNLpPd5zv5Ty2LEevRf7JjcMPx1
Z1NNYWM9bYcqXPK0EFBMYUzJmyicVUdecwVKJboTZYkMhW1VaO4ed4hboMfqcrMH
yNbANf3Z3IKehWEEECVfYLcTGPGXRfAzIUvdT8R/nixgLhzbapyi16N73yi/v+vC
MXPPF62ws3H8gs3HtGHQjF2RPUTWv41UIHVKmVKBW424RyNt4gmlo0bJtoyf9LOZ
duQzAqnh9Lq7iT3xB3uaAemIG5Kj+dVxfN9FyUf6qJjMI4Z7jJoIR9da/zSuQifs
mwMnGbLmJwtZfO/+8nXoMiIOrQP0yxr4xxDCmcsicYfRDkG2SJNsTqGZUlshvWVm
1iBRFkP/Gk3Yn79+AAxXXsWtNyUl8/9pSQGINy8xL969ezhTI7tan04iXGm/56uw
8MCRtsOIkG8U4O2KlIQIeiujyRsblwcN+OoknmqIw435/NIvK2x5KOmkQ8DuY9k0
WtEEu3iQW2rSLxnW0Dg0KIZLtXpt77SFQO7TZXQmf8pZDosEfDmUwVSgvbdRzrwU
OGLmMJeYgfsshutvE8CN54zCQWX4PJsgQslwvUlw+WvA5ljHYD+rg/6PsVxhEv6c
8jObLlAl/Zq5LD70aU2fBcYKBs4GWEfsd2TKrjRLMEgxwv39mulBHMCjweSdo4Vt
ZjRtHxJ6URutbGvRiVOtGrzDB8Su46hWHd6sqj/4pmMEPq7pD2fS7XAVepHJ+jb1
sOyYZc3lRwFH7EVJFFeejesqUcSD8QG7qGwkbB3PxJddmXdbDoZtvLpGqvfFHSbm
2NobWmVuk5ueS3lq1bp+xrpyjYN61L517Vfqrq1ZDSCNpcg7gbpwr3j1sa9f4HPG
kuiK1t5lOwXzo9TzpZkf+v7qickqXA4gy/HoEAj/NTFa6MbxAk7lBYVcGrp3R9LV
zJv+iXNjnIafwM5EKfE4/QIssSx3MdBw0YoS0C6YlrEZbRoEKdnyygrhECCTV39R
vTjgkEqDAo+AlL+NmmHk1HHE7+I8BkMfc6I5TTFBPpOt9qaCr8lZHubAgpgFAjtP
Dy4P4InRE8YjnnZEbKTIk5Mjb5Qb5F9i+LY1FUgvi6FePNWT1xyssN32nvoZo5Kz
5ILCOgywCyw6GEUDI0A68j+b6aQU6tupz4zqq1+019PbE1h7koNSkPNBJPEoc8fl
jRv3qJMHrh38/yZjRxphfQYnymYnG+90ziQ1NnE10FLMyo+47AU5ceKSCWa+TYWM
r1RSpvHSBDZW5Dd68W+arIVjO9vOc9b0BiPGNgUWtq+Pdw3uosxuXbGwodHIbxcx
7qahOF0SotntyV3d/oq2+VYdptfU/tThlJC08LMIuUfPcpFsyvNzLN3Kemd8slgy
YZZM4Jq5OTzl7IRjO8ROsifgdzR77FPeUsBk6jw+temNbVJJjkcMu0e4Ip4PaQsY
U4Z/836tbNs+Qe48hWSkgyTbH0/FCrwvSLaFapT8OCdnEKId6dlW9Ej1FUVi326/
RkAIdCxx5UXc47XyjkoDj67vJ1ZeDfUIIBgii79GFA5vog8SoUfsg6xQaL2I1Qmx
phmhbWaBtMcb63LA+L3yFbggrI6TgAnQvzc7pt/VlUWqYjFplKKlABYJrDCkvx9P
X7JU7Olu4rBkCJMgs0uI0WfdKc1PGK1QAyMgNA+x7X+uYTchPVjOPShGJEADuwsB
VIZxBvPR1uJbD5xOZ/TL6moGmDLbQ2TSHIBnV5oyUib67Ap2/y0ruLI+9RheID2p
oMGDwBD+bIVhi/4cWNYbAysXdXVvFiDXO4HPWFlq+O69WbZr5+SNXPSzvNNkwPcd
iRZWt5WCToRlpQqsd36Bcg+BGuicVsgy1TJSi8eRVgMpbrz0ir+PQb2AluTCKK8E
1xen5ycnfGUJTNtjCpKoqVaNcpRj/+UGFmFw8yKS0h00gkpGYxcfkVblRaRp6Qwi
FI/i4fU42moAN1yYqa6RxUWPui04Yc4ZPU8AS4eqSLz48CMO0XugHHfsyhO8GJf7
nrDRSZ1TvfCrxxidcM8rOp7+xSY3TDNlRUiUFFBm97ozJ2QJMwNjPdvIYoGYt0E9
P7Q9jRIsFYn+PT2wGNPXQQkM3zM0h6pEUBKpnEKOUXK5srRYdND5CkCQkWZUPIpX
JOz/x8X8/kmq8O8UVRXIYBlwJd+TGg+jonfN3bIbCs5RgQlOfN7V9zkn+Hkjodpv
gI5ypXOTpEaWMXCcM+OE5dPMcmzd0CUdbHe9GLroddUEvFup9jPnwS9PULwD83KI
bT1OkUZB9DkXxQTQNDBvu7FOTUaecDnmma9S9ppxOat+mYsYGEXinvA7r7Sz5DZe
p/kLidM1UHF4R1MN7kp1jVsieSA1gQj+RBmD+u7EgTXx1bv2mBmU5x+xUmn9CN93
SAubNnt0IwcYPsBLJfGDYSpgQia05P2NKrPUQ59FWAehQaQ0p+s4IeZVw6GehYlZ
fmFbSSnjF3lP7S+cD1hmxRYdOYuu4iQnVdYSEpiigXzg1VTxAU+MGMplPbaOqcOn
wdD1Gh1gFKaqFt2Sr6fSIh1eSG+lSmlJQKsQiioy9RBlUW4+12roLl5Tk8shwu/C
cEqWdeRs7I+MRo2upjSoqfL4mPocgECrfQkLZLU+IknJs4pgULGL9eLb7/q2vHcI
zkG6cxudlgUKwu93PKEc2B7yonNL3FA5CV2eDWi1k/omWnNh3vYOq//ozJd/O1wB
8hQQzuD9JFBW1vc8Bezy/0PC0HRIr9MG9TeAr7DLeh+ifa3GJaGB3Rx5II4RwkBC
9J1+6ksrSBTeIlrwByLwYhSt0dARvemkb1a7RnKS+0SDjA7ndH1Oeif44a6agYzB
CNZkVatIi7/GeE4FW8Ld8w1G4CQsjlOD4nUri6USXa1NWMcR4gSGIPhsFXH9ur3Q
z+wuj7LwB2g54IX8jlf+r0mhw0TzJAOOFHKX/Fnh39+xZD7FX4RgAoc4ME97hTly
WEBf6RDxvSpw72sA9uBspHhFxKCuha+1piqlm/c0e430zmYwM+4Quilxk0EXQhLq
NkQa4Yd40/oA+bEiO6biel+1tLeUz84YY4kpmi770EmxWmCi8wHJxAyuBMcsIMzr
JORBa4DhA/75pdQKbi3i3MlrGvxS0DT0JEEzDE4TZRI6Bi8qdciEp9L4myu+fHYg
wIHpxn1kf0/HPG2HjmhK8JtPHk+l3MUhGUUtcy+6NpdsnGr76ttNPWjD6b2Xaew+
2nsWlSu6pV/gNQSu1a0g+REzlC0tdzxkINedubORcz/NCp72sbxfBdeQjd9CaFwC
10p+Dg6U668O42gRfPRSh6fZLEH75teof8XM8oiKnpB0lehFBea6Y1UqDnDP9T1K
6SjwEUHryDU2vzUosF/NtqpBsKaPVkkWug8uuCQ2akTx92pza1tXi3/22uiJGUhb
gT9R8NDrCkmhE+nd9RLh1/Thf07S6KxExdInDFO2Totlz66Fpxo6n/FhgOiFerWM
L0CrCC1h7Wii3KOdLAj9rm8DS7w7ABg6+Elv4nA7tqCoubDYH/BzkXFVVeExJJfC
rvPFIoR9yVajeOubFCLj4zGuNTECtfhunQS+1VeUIPHBFajFaPM/TncUVuiCGF2I
ktj47RcIx/LliJaAXf5/b1pVlaBlKgCxiGwYYWWn2Fzp2SA0llNZk5Puyk6LXFwT
YsZShUGHyaM7yHGI4KaYFhHyA2Ab4GQdxCPP7xCtYPWP8Wr55Bei3oZ99WtzivsR
5xw1i5VlQ4m2AWRHbgLNqmOIgb9SaKwuithzEaYQz8+D1bV5oupw+eXalqWFHbXi
++f6vLGyuWr+6eAC1T883oP4od9Kihaw/kZ0g2JoD+mnIpbPyjdDrfRdJVmR03pe
fp11fwXwl5xCMi/Be1knqmv/uNERQA2l1PR7bJu3pPXcruXRfuQH8xmQWBgVJcvA
aIJ6Ej9DbIxWaM5wiPZ6un1zZ14H4ekg8TZODMXtV++Dr6x+Lr0uS6j2xg4isfEj
CGazQGCfwwvhkHaGMSlKCGM15Jc85+8y1HDW+aCp+VYyyp7QXmYmRrbqAmsRpwq7
eSXzUvE8Aao/zSM2vOQTZO7MjmGFkIYHbdTaGJE2pVZNVDXjbqyFvkrddRDn8v/7
grgsOopRcawBt+H+n/geSdHycMIrsDJeIkdrYVPPDgA8Vpb/mnvV2UQQ5sa6gfiJ
Nyy+0FPbdoUEoV+KYJou6zR+I2OaOA6WhpoV4w3jsFYOcbca4IcT/YnF5uF4wb6S
vnRtDvjRZJ6roeGwqtCLbpEbu2FE//ZJMaU4kVclfHsLY045U3KN3zMuLlOaG9v/
NWVmR7zCoWmrVL4EHHH1AXd7+zsnNipA1hBvcD6KD4RO1qnIHVqvXsYL/uByCCPa
fjmu6+GlqPiXKieeThkBAtrYncN0x5ud0JLsPWU812kpE5SruVKAC1N/XL1hzKZ/
Az0hn9RgrL8TDmj2QogcbgmgMOEDhOWGQCK8SvjQVx5b74qWy6PtkMSotumBOZEC
H253DMwBlDauoCYvmoMdUZDJVuyIgbIDVRPq6qlz6Tou6d/xk3GEBGvphCoOqmvM
aEm5uRyWcdWAwIdc+agOmmymRabB0Qr0ZfpoE9nmEmEAlGJf6julkUUGL+0rQY2s
HAGv09hM/f/PFVIU5b7Esw==
`protect END_PROTECTED
