`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zAtpyZvebIiFFyp9zAQRGtXU2lKH1OC847S1dPK8okwl343FHe4+b77K7HT0DQn5
PG8/lyYeCsxxG5onngaY7SsSCo7HLDUdj2G1sJZ+CIOEQ5H6loSBBkIEeprpQ1+3
Vz/RVBq/c/O3scaHYxorE4uyqEicENxhvCGZ2Cmv/MMuX7b2d6ee/P5jpMmLPJnY
8eBbU5/z4CXEPo9zhQP3KD0wJL9fk3bdgNCQ3GTVDTuA1RgAiEcwWUsRCeBy33RI
NNcVwVm8oDdNDlwlrm9M99zd1Cke3sLFFlS1AtoeXh9pTD0sWoziGx0vWhEGOH+4
eG91Aoz9PPlUyImk6bUGo4xUpFDkHWOK+xGwsZcts+ForFnlPt/AqmrCJ7zJLyJj
KPSuBD4ubUyLDJZDU5Wg3hXB1Wz2HSvcQn0bK5aLASqlbrIPaAJhrUSWNvXnHWMa
0Wfwz0l0LlQLJvNhrNU82XUbDXLujO/KJGYmPtLUO70fY2X2OzmbfeQwFuqSzUar
rGtFoi/uiUv5St+yDXTZacD8zNHdP2ytOeWjdvKPv9HE7u18WRLbNTXHcUylewKv
BhMjKWk2KyTp/5mWEouTXRIe4x8+FlgaGuhgiX60PUQ7z5mSl2NGkG5atOjdUifA
NROKDKQZfVXpVGQKAgTatmsb7L3hUTt5TKGRlfE/nSOFkfifotBAdVMSNW2tdOFW
zQI25u/ueSlTqIKDGAmT1vk/TR0bYZ1prAtUYOgngy6kuW+z0i6EOFy9RRIumN1C
9AyFbUizutQ8tLCVHPug6T5by0iyprNFXkKT+hShYmOXjJGNcwyo52mqrKHKDwUv
c63cRZ9LlNpZHV8FSHMuKeK/KLIj1dLCPucwR8yuEfXuqSI7KqGb0VE6Gky3OeFr
EKuOqi3uvnjz7oxJ5NSWDXAG8jP12uKdOSWrN1E38M0slXU/27cWPdP7FBONXJPv
c7C9nYXtu+8m4HupL3lGtrnW0vwoGRi5kJNkUapx3jzn6sWNyQFvYUz3C/LGgmH9
iDcnL5mdejPgND2Z2zkXnr4eiSSaZ4UWDMqUOLQpWdOu5n9QGY47d59o+/oelF2U
EI/21Cx3l0vy7eyfL98xMAbGfCbVRaVVZhKoqQ7TxNtxVRqTZobaH2YgwdTw2Cn4
r/4fqAfwm7PBz8M3OWGS6NnlI2FVYiP4uT0lD3G3clzHFOh23tmQGzxqjEY0pIVD
P2sZB+O/zxrcLmyZNwXFeDDw8cd5KYSSwfktEJBIHxnXCGLFQd1HKNxv00AvueMT
99lzznIZQfxWEDYDNg3HNLdQqKDjWcOfmT0YE1IyRZe30PdF2oEBtc5gHHjHhMV7
tufmNvsTYsq/q2baAu7wYoiJ0nFE3EYuNzO6Vr/qI0RvJDgEqGVP+L70wmuBMbbl
wMIr1aInvnGTb6xP2QQPZg2DNeMoJkK4scHnzTxegQegVJeMKJeF7AtllO31MoWi
ZBRIoX7gDSegWMSfaA4mtM/8gLasKgh3ra1LXSXiXKBzZYRgZh85QH12Q0PimHiq
nqmO1rhTXcz+6G+uQ6lk1oo64IsKCnJ/RwCdqAFp4uvPrrHYu7mQo+hS7UWbm9zW
OWTIeVylrf3Cd2fQMA/LDyn2NM2AmwL2ruVKoq98wQCdESPxPQrfbs2oImBltIXG
idnGdaDopCYsvt+g8qjUVDNvjeuFRI0bj+rJNZaHmaqfeanKmnD2uYIYv7YXey0X
iZKJckPi3AzIjEHI77oJUAu54ZRm/kD/3QLYr66xhDNgAJwIFOGKUoEX5uzv6Y4A
2M3IsfZyZ9XrPURKqpMRhcOWbEPOaVLV2rMjkYtoFk0TuE4HHoqNvtsxAs7ogwtR
cf3JJXYuXPZ7ol0A/FaOiL448+7vKB/vZONjJ4aFq/M5gqcObJO9VISn11/+fVnc
3C7FsoNUFp8CAne6oj6uQvvUyE3acLvKOW1N7vKbbTyi+ZMw1PreV+h9q5bNRefF
uUyAswr2YZToqM/5KoNJy9CyRxnpHRZ/mVpSxrVkm9PmQcThD2IOmkgVQLcvP76h
YsHz0UA9Jl3C+0REpZCCntFgE4en66oP2Gh7F3kVG+qtGU6cFemj3ARL9NnU6yrY
Um2LTeiWIQAAbyB1fCI9CjeHrqLiWrlbFOSxsVVoNIznBwtSq4F10T29Mua42YdM
mI+BH7pCMNzDs04QmtiiPNfNZPDNKT9WcIHh1YaVatTcHsU75FS/HH3eCIAUAUJ/
CA/EltURI4C9we/Npa5ZriHZRzXe4HM1jkScLo586bOTAqY0iOX95WgtZiI7lTQq
t3Y7NzVzITncQudmR5VTLGVb7Rwgh5h9TX6HOEyvV07Q5PJWBysdPXzAXpSBv2XI
b8Qbdg9cJ2IZre4iteGpYNNrfxxkfe46+kblyCpyBRegMhImmSHo9geJMVgN2VHy
6A7mmvEbchARUUhQSGic+t7yIfmMlyNZGey8XnU1mz0DVMtaUc5xR0tFHuUuGhmY
H/SeVRqNI05BwP0Sdadv/A==
`protect END_PROTECTED
