`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/+VKqKiGgC61qBeL+Pz/iV/YJaQlKne8pVQeeT7304b9zpPfqes3IcGET0uJ7Gzb
WSbo1oxvXtcJZgPz0yg+snx1YvemYZfI2fORx3fShJpWo47dstuTSFsjVQW4qRSw
e/ir1ec7yH26LWbBAJKyxj/sDZqRPEoiusNZ+/3V6Nx6LVMQyfBASSwacEm3iujl
OpeWzSGwOWVbD+DsFofDeHauNwfKt3p3xNlECk3CLfcmjCeAu/Z+JlJFTjyLK8aa
JNUNJzwi0Mdh+K57tOK8FHVyrnrjWWDERqA4dtgX/gi0waTYreSlJMI98lVWuezB
3d47nZiXSJ2W0/9Ls2HQzxrsiHqklxbLvy7e8WcyPhvJEP0G6Etzh2uZw3qcN8Zt
cW/K8NUQyHgeuPQgRS5DIaOKroIImmsGC4FjM/mbroZNqpp5xSxi2icRzOt6h6Z4
siL4sJSuAlwO89v8pvSYP9xfaqecfHTXLcDcrIIIEh4CRRQoPv6fYvtxFiD0t5iF
xbG9h94IGH96e3PeViqL6gDPkaVz7H0m94Yys30FPn2uvQB9UhQBiP4VI+FcSqni
47KIHV3fPfxV5Bo6Eiij8qW/Hq8kkSBLJG0gj2Y+jDantV+/unVnx9A0FbxYw7Oj
4e8rJ1gwOsWvmjhR8+m4fyAD3J1hGKFRjOPq+4rR93s29zqu71cdiJRJLM3C1NXS
cC6qH3lTem7jI3M7q3r1UxKHrZCHUFqfcmBgOzl3X4bSt4UsZ1j9Sq9nFMm2WVCC
cvwln1QqhgFBZCBne1wvr6NrKNut3xj5rC2vQkOTvD/v9OAwi5I6YkqgxxU45H4q
4cy0aS6jkXXnExbN7C8/oGhY5Geb3a9D2q42lBU/NLJCXbfw/JBHe5bO6HpEIRzV
8lSFQ/M3bqaZMiDqc/yFQL0uWVjyYMSvELOWp2FC3p0HKlojhtKLWhaQWyKBysO7
2f3mh/Bm4Jrp0CJKac6YfXr9W/YUbOQ0l107633yklyfoz1dF0cFe9wMFbIbAfB+
ZO9BIAArGD4vtUgJXeoFMPcPO5kruroXLGStWPGhKNm5yz4Q4WDk4thX7Vd7eVkd
DyqLBJQLHulncq7gxNWqFy6Noj90KYokjQd+8HaIstZhCxk4CvVJ82h9Qbf3LES5
AT0kEevDLp01LvYEtyQzEECHz7U0uEgR3qTLa8ZHn1qrtKM1lC0eleeb9rKRhG2r
Z/rGdwJX/BbaA3hlfdh3UPk1nLm9/8e6Pj9CwUzb9ltK/2KbCpH9TMOMhQH7DB+b
tuXj5VxPB4H4gB0+QuQq3XDSq9E1g7Pht+Dj4NltSbLG+R/L4BIzM9y7NWEP3OJl
pRvglRPXLVFROa+UXnhkKx8AHFlbkEv+I8rWQIS7ICI62All02lc0RyovZgeK2ur
Cm6FtLucWexwdLDiCiaqHAhZJX3WkfbsuPEwgYfKkGzsB1QmrfCJOcERlMsFX5fH
c+Q5B1cyTwL6Twki3NP4WrUvevYb7Q/VXeVpxGS41vqMbIh3tiUl0P4I9ex4yB0x
6FQ4na3Tpw6sIMUbOX/D6GdeyUJeJubQL32zK8pm0vM+3qt+4qYAkc/U4dEdyBWd
ukH8jjEvHy5o8K9qBQNnTf121erVyhjtsa4S28HtfQNH8+NQPYXR1UA8MxY0W2L3
DRKu60SDUffMhl+b5e6lGyl/cDU/N50uffKGkiZqtUTVPzgXVGssXvyJBh7o2q8b
SLaWktI4LmTYdLTzcmctHXqqV1hXrs8XPRdgPiKMH1jiQVfrhjuZky7S8a1tjiNc
KikN+GV9rj00/TZw5K6oUKaH+wA+0nnMOjW+AokuK3tl7FYNfoeBIHqw+fWdjn78
tTMZeyJBJmuo1iUZ2DEMZp/I9cX12CWerjqXM6XtDkQqT6OeDNpscF7ATbQ2se+S
lnUZhkqpNhrUkKU5YI2595pdIeDeDIl1/LjUlIt7Ww0q93maBZUK0zsdnk+2vr6F
H2EIThCMcKFgy1j/0aMmyxMWJiFHtkpNKI2Ss0PIJQn9SV8e6L/4cbdNgVLoHp8u
zfAAGmxH+zrGcDauT60f7L7+tawvpgjsXLiAJsu+CmmgjGvoaguC3Bx9lGWlbRX9
oCg/GaGkeOkqlj5kCsXHaWRCgaiFv3jO7fxuFTcArmR0RVMfLHFXlbWzvhAoqzZa
2ftT7StPq8qrn74+F/1Tf1uo7Jh9chqQAYKBo2CIPOa1jlMSOyg6AR45DO6kz+ip
jrPvBWX5WvAMyVVX0D43ivTFEEc5wIvFqel8gh8i96my42cH7RUITstkPPiZyyTM
lV0ZK1jwOxIlCUrQoTpvUTyBSmiGR2UHTBjhRaK2ZleCPrB16HRPrwEFzZCillpW
77YtOpEBccXxyUV8oCXX2dvW2sf4RTVRBsWSaDOplmvLaIWPez92XcJrtjARwax/
wlDbmRUoBx0m+XderIwq7suiutBcrnWoJHgn/ghIAFrrQNAlPXhWcr6LQVIgaxFX
2apxTSlJ2H+CNekzrUz7NnmQC9tkN2fRlr0xFDwqGX1iXejCDfxr2xmsnSQPaVGd
S3ocbTT+BYGmhf9yP8MFT3GmlKiOWhgGjqy4+v2TOaS389K0eR3a3akq23fTnyaB
7yMfyKmE9P/s29OCViSN9BbHNBIoFxRd52tkOWnbZxNKWAIuidqssK43zUVmqD3O
oxnwsbsANbh+JYRkW3e/+h69TEO2kuqidtamitdHc/ldgINJr5JxtdG/1JBzlq7n
jyzxH3cwFGxqovjnWKYik8+wUlOhJyjvITC/2Jus/pr4OHfp+mQXcMX5EZXT/VJX
69oAo70hKqz3LaqthlKzz90FhGdClI+AN7n5FuM7OcHrjepBllDEs/6x+3EF88//
TdkhTg7Pmzox+vT5CyzEOgIJ4XuVAPeBYHMh1ZbXPRTPWl5pOCH2cY9yTJd2UQZP
KL+hmgFkUgiot/0Lb28Y8mzbHTsodifQm5ZRB6Jo535+ElX1KUkqD/It8VKJ26dz
KYUa04xZ6xXCTVytsSRxRhmbGHJG+LMl+LsQjVl1H+b8Z3WDWs6+Bi42y52lRFT5
+l2NXmCxN6h30qil+Vb8TKqLbrXoXERlwZYzNTeuM8ALK3SaYBW+sA7DmdT+BS7a
DtzUISzIC6rEITzWeD21M3SrhUGWV/mWCOAWVFjuLJ+N6v2H/A0Q8n/djDDjAo+0
caY9/RSmyP+mE+alV0dhjtMATmzzZL6DUzhgtfWUAlfSNMWbPapdmshoivm0lgOV
li4XJZheKOVmLIDn0+Wv2OT6CwMR/sYfHucgn+p4/cNnCDxn/v4aElXnGtMSfcO6
Wt8Z2WzTaqrpZ2g0vwZCG7RArNJojU+kAUlEeEC8ildUs/HOyGe/Fz68Pumh1Rzd
AtEuZg//a2tSXmzoH81zvwqAK1OFzif/cTn+5bsElB5K7SucJ3P7GLzp52LCRmZQ
Yf253uOEiaA2+nRZMgY0uEzJgRGIaX1rCNIlWJCZM1Nm1Db/nnBVHKNJrTAdawZy
bRD3NpWn4VvAUcC9q8rNmqDxvIevmCABFH/r3lLnQwyLpxHe0EaxQrBBPPzfSulZ
AoVptcBbCljX1qOCqxgAfQ9oovAygrP2OnmYEaWf+nTYUlKkGfOemwbJ+vb+jrUz
mVbgQPephTpYw8OYrsVXwHQV/CBLS7p+YoDBqB6zSazYFQeD8p+b38kgy4+A4UZp
euDvpLuJTnmL9Uf+o/MdHpxhJJksWdvoUHpywPFGEL/57QQLOMcqd+feNHJUUzra
LxKmRcDBU3bd4kQP169i0yBp3yBuz3yilXTkkoUBNaeU++EZiKBdm6Oq5o0d/2i/
iK2Lu7sOaadmWCa4QGnxGq1ijFL4NRazXYaQTkao+rbiNNFR499r8ibT1Beg534n
nHcAcr5Fu0x4NfNjFwiKZDcozN+PaXDnpuSuvmp+T6RsZovhGpdVwnQGjVwvPyQ3
ByseDQ30gy6vi/vo39N3pe6HzO3BXD6laGKwoVU/RfdBXb3P8aoXDCXtTcqsxz+d
NU/Msxp3/1fqm2vhzp6y46KhR+TYInUM8kCUNaq+AWHiMruq9+zvvqVzwa4JX6NH
tn6wQr/u4Ju3vTwBI2Ve+r3381gMTr6qNrKl9mgwRahkfwvz455t+tVnI4I9NNZm
Cf97xSeVdEv9WXtVKW0B1ev/1sTe+fecvvh7AydlTNaa+jpL9WpL/FXDepC3at9z
rm1wBaEDpQ5RhcSFRlTvPAXClDgqXTvbUqXcVQbf54ZdIVX29I6g16VmOI9BdsTa
Fm0U3JdvOIDWr5S/5pu7mQS8Wdhy6PrNOk2Og5hcuornuWDqxufzXbO/EIg9yriT
gGtPnyLHYklCbeW76I/LPk/2883DauYaOtyYX4z+qmdqseGcFExWvHEcGVDE0enk
RR5D9/Dj8gk6nX9JFq3G0SWLqyuVFDkfOR64H2vrF0cIHgI4kHBIC5SmpLboOyrI
2sk9DYGIyaqJQcHgk4Ybnk1xyze6DEfxobSRWYk5RHh3GKk8g1Hlvv9R83UuvgLy
xq0K5XApXfDXoWWUIsV+Z66edU6I+4Ar2rxRbXVjHLIQvDBFB4HFNd78sAXFrQ+M
n2vDDhMlkQzuE+i09tL4eZZboI35Enp/qSutE3LZz7e4vzoZj/pDuezYNBZgxHkH
nX2d08iJAf7MLb/40e0Uubnm/Xf4R1Li5B6VJ2NOtlVqt1qgu7aRSg+3JDvxvDfu
p6eoJdDJZASxf8wHnl/yFIF58CEx+EuxoUSM2Q6LsW36bAT9qay+eYa2LBvyEN2j
Jcw4l87kAR3VdvKbUmMDodO5Lqb6R+9xWFu4wL55UsyPANJcOBjop4GkMHbnQLcZ
CDT6Sd6wtis9fNL3JkezomlmS7WSTv0LSpv31FAHPNmt0NEcWdm2/Fyq6i3hGtNj
coUWcPFH/YXuIn1JQZIE10Vu0oOAoQBbQxWm5ZZw2AMpyquLt0K6kkfXVB+n45/M
NaS23Chh1JtITFMoKrjb/jbUI1csxN4s5ko6ZilaFHneSO//74kI3HZV3crQrhaF
lVdSWHJQ9O6HLbyxFjhqaksJvhbxeCsrd+JKMXscm3qO+yOcbcK5e1l6/gF9p3y2
UN+kmYmWUN1MkNGM+bqIAhcFEGXq3Ymv2HciLyJwalSZ4Z0w4udE+cRHG1WKJUNs
72mJqcNKtEvm2fgF8TqCVoH+y13SVQL6CcdI9vnMtzO+XbAY8tgedSeqSdpPBTgW
AfqVwQ+SuP4OLnewtxEg/aL/EKFKvyZTmGtDSYqvMGO12nbngSBLFwOSdqwZlZou
riCq1R3l+7AWKrbTOxQcy2B8kTCkl5Xx4rMT7cUiCPjmBeYJcNu3BNMWreq8SxkV
XmoFj67au+4AJbKeqd4+uTnoVDysAcyIG5jrC/pjhaXLAuFjt7KrZWwQrre9j07v
iLrPtMVxNAsqj4iTdiowPyIe2QKTC5VWClkOSeSmlmYsNXh0VQwebHgeOSLii+41
97E97IRTP+lYheLdyTVEktcYCQIqXAFzfCvtSiXJ40AleYXeVJy/ehu6POwjSKtW
GZMHdgkgXG+/fW7QSxbhE33F4xb2oJGiRHecEdlkzZK7o/KCpHs6Wgw9Km6yCa+B
t0J/uKrIVJFw11qsCooQt6CglIFavrXl78Kg/LTKCJ6obuGevcZgB9sbWpQ1K799
g01zRL6fXJjvsRoMaXPl6tDyqOeElaWJUhpb7Y6D1qUH938P+p3dN5HORxO/xfP7
dtf9wFMTTkIHspTAnRAgFj6cxP/SP2hJYQejv4+dBwIEPpQWkziMAaeF236oVNsB
e2QMVZ5Mi9q8hr8aY3Fu+imjDS7yy5Zetl9lfiGtAGVnfME/UPQyq67XEw+lglyV
WON9I2dBd0vwzk595Ek2NDRUTygefwjBSfK9odwLEtfourI8exs7u9CqUCayPdyA
S49+QoUkHIMPIZVcKcqKhTYu166eeqdSwEUuSGgb9JnMQRo8CwKMYpqkNVRzkl4d
4JNVeDY7fTnjWUKL1+ieuBnVGc+hoHsMjgs1X2kpuWEnLxYZ344Aum5QAeaVqINN
jhMJSpWikuk3Airo6q9RFAqs0gPFkmrikW7z8/cVhmyGb8eVZ7GFnTgVm5qAAxhl
W56R7pLvmANjEsTn34uYTilaysDyUUkG560kDgAIDSa0RlvkQrtelpDEANTcifWi
84Dlt6MWsCvc0J8Z3bUZl8ZbeKi2P19Fk2OudN0Ah1XJbj5SHyuevCUG//IpI1eV
zyIGZzgGWTpQrGt92TPtRO633yZDXSJb1ZJyRUZWIF5dEr2L84CVwCg/fFHbpgdF
B20GW+J9PzDu9Hc8EI9HiW0ehfcaxL5Bt3v7gA4nyc5prudakCgSKjBP3J33jmGx
YnCQpMnIHqd7mbavCBAZhVSknArZHnDjmgpdMBo20po1Tol4zovWzbjtr73owBhy
OZjrLDTnKzgMJ41NaZ/zn7LWn5qedg2+Ptt/+7zmJToKx5SkvJFHv7NqkCQ9Pxsx
cpUPLCKefUAJzsb//pjYaLXbxrymlaSgJleeBVYMU8wcaL9uZ+JNLGvrGFnDesyF
QMrTWuGNu36jhAO1X+vcxyHHIzrCetqloMSVUHfPa/fvG2SILrtzHReLKWRAjwbg
bwNJyLH5nbBZXyr9jUmDaSCYu/qFWyUL4fGmN3fOYfJpxmA+QzD//aOQXLgMsHbq
DbMvSNId3NJQ837hXrOA9W8Yed/hz8h4J+4XhfitA8aBdRApX3l24ZrB7DzbRYjV
6DRgNYPGWRfULOwDaM7Zyuh9Uog8rxHnQQOciaP0a4c2rIuqo1lUn4dbCwWDD/Ke
a1MHD0dbG2AAf0+B2DiyoPMsmxATgJesI0DWM2876XabUvJazhryXmm1GrZFaAHK
OmUIhtLgtL6xq1FTIZV786KA2sfC4iYHN+2ZHehFVRotPqj0qU5PtZBUss/do/eQ
isjpjQtdN36seRLZbVvmI3hh2FSbWW73QvtfBeIYoFnwdzl+GFUh9UGdI8kDVEGF
ViELrdENAjFnsIu0r/Cz/yqLY2Mvbu9UFWcc21chMjgglxLIaH5TdYGeCka9dZqz
O2C+fC09gNertiNEdbH4ePG9waPlCnq9MJPyQHWrKNSl1TqZHXntPQO4sZFV0bqr
Lq6gDpWFgisLJZi9E+0DkW1RaBXFHZ6BwIj+8izWIDd/t3JTWP4+meWLN3tYZaIW
nBYAR35AllLJw894b5dzB8chRlPE3Fmol990ox76MudrRHiSrJINa2bWvhZY6Lnc
RcXCw1RHlJRUj/EL4gxBibK57YKYa15yYslL12A7NYN/yGHVnAJ6OPEkvtYUiVAZ
BxNVeCvVHPWHXiSltCgRSWUfK3MDg0HqwTlGGJdDNj0Q7eAA4o0r6VSzbOoyPjBc
DBn0DmyMv1Znb5kVbxg4Xv1kAdWR2l8xdZs2gJ+ONhUdH9+Xlep4ezI2YJLqK2Mi
4nWv2VzCKHykcr792y3/YIRM8qjOkxeWKudL/IrzDXquTi2R76wqNbCqCqbBSXeh
QnKqeCaSPmTzpogF0qQ3fDX1oEcr3J2PiK8Hd0fXf/6pNiDd0ZF8vzgQlD4SuU1P
oSNpnLHboZWjiuwVgMVBFL2Ulpql9pEPfzv4mMmTZ+DYLBMGfOjvqND6XOax/Df3
rwMkRHeTaAKEUUjWB0VnCeKvbRlm3i2kgBojZXhIcEQKhiDx2dGQpoMY/8baj5aU
y/TB1wLnA8w86x9juO9MY0Ae6j0t2097dFT8wBMi9wsp35MVEYrS+Z5esxte2syS
piQNxcUVVOaQMxyREw4eCsSJiUTg3VBRFV35WYr1HOTTziGrzK8pHtlvtAmZ4Ta0
POhR+R2fdYsha4aD0pXMFXLAx1VcWB8x99M0v7wLIfKd3YeFOLMwPSi0rA0hxqvN
vtNlp03BJcaQNJ0z2cmRDdafWVAtvdHFYx6qmpfD/IjketHBVC6JltxJwJyssflh
vTbC8LjEYfUWxLhIDjTbnNZnkjVRZsnVYsNBFkkKCQ1WAquQDw8G6s0ehYo5xCeM
wU0Uqn5cD84ftyuNPXXe9KnBKVqSUC4pnYkEvLUaLtcLiU+YLjpp1/e4Xh2ystPj
pCJtdVGcjqh33z9fpBRMloVsn7zfi7J0idcqeew2ooU1JfYjAge4CaJ5gIT30Yyx
e9QZGKdfO7axQhP9iYAKa+EWKCX6G0haACy/oGQ/EJE5sHCK89/YNhlWIUQc9QKp
jA0wTp6aP2hb2FDv3yBDU/ZNFKBwjPiiKcE/UM6mCoGDKQ71dCWzybrzX6k6Y31o
TXFrzfIpNvRPCwKySbUSghqzJKKtm3995GwW1WzMfzVB0rj3UThwU9qPOTzs0pql
ciL4HOe0YPBArafbrkgTqKNfQmxVHZuiO/0ZdajPUger330spgSB/4sp0NnDaiL3
73tru/DaTnuvEgjwJ4lWUli5chVFdnl2g9jBNAOCxsYXs3IQe2PoUHXLKueYhaga
nc1egLFDL4cwfz4yPPpYAzZIhUSHWbQL6CG+MMeHNhU0aq2RELqksR6bfSrEU0ie
/FM87/izq8fr4OaIJ/2wbV8Tq9x52xJZ1rmEUM2J1U0sXvHdljmd5tMR/bE3ZXsA
5YMO4ozLOziDbNAAj0rZfetCA5tvdgP2AN2nwSWwWQOzJtjgz0MinLOE3VTBbXOV
k2cxvv3ERL2kMKB3Fr4ODqOiwPPZO8dtZHOJf0ToCcsyo3TIbrRMoFxZQH6SlkAt
ZcCOHcHvke1Sk/c5/nRnhbph/V475c4Tk4ilW6OIlfkBGGlaPF1BGwUeclLpQM0k
7QorqEcnToswsfKNoiB+E6GBj+BKnyf/3menpt6N7vSdYtWrRG7r6y3zfi3PZoZY
uihtnPAJgGWqEQ/vqM+TxWHwedZkxeY2rA0yaOOsaQ3e9mmN7+xcwKJzPeu5HpvE
F774lR9ZbjR4TXFFIMpljObztCStcdpkPdCgUS8GDxXVSrxn/1dwJoJjEy+JODyt
M3SaS62YSoZFdrPeTiCIV62VQcSfbV3wx1Jmwyto5Edvh6pAZLrczTAoilCgJ7lc
Ua2zTDKQrktSxJcvVyeKCVNEuJCdRdJ2DSBqST/8plrdOJJFs0IduHuIoNtKKEAP
Y+4l8s4Hs4IUSti2l0QfejTXBGoMJPsPOiTUmkSfcalOUq3lW0OsLNBY0Za/kmJx
te/FoF1PBaK290M4bQVBBpCgTzzlaqWFZfieT/4rib5gcOfmed7PM87ZjQt3ZYUj
iErg9mH+WdlLY/++v4zzaAgDI1S6KIGTQ6RwMerriqE3Rg0U6fMlpWWNTHqpAkIh
FtJoHxelSLx4vyJddFSy/Md9RBwYifN/MYDyMgnV55WgFfJvLh1UK8JDiQc10Epj
w7KEuYd36cEsOr1gT1XlDZ9SquOw8f07cWksdTM2/0dcFOZZYL7uC6XWZA3ST7yA
lp12Woi6wfKjMztUOV8Yr7+0QkIVeErHmwji6fUxIbYX8yTgRtN/CylWKt3Ob19z
s8gYeR1d4aiew9g3FG07pHGGdY8DE76+Dm+TXTH5GEoWw/14ybrHUHouWeXsApM0
dNvRnIQnedv2lHHw7MCvzRlfweAK3/+lDQM2uz/8JvEzWPQ7Zd8cOG8OF7McgR+/
x6tWaGvGpaMrfLrkfhunuUUs4ZAn3hvPorkl20TW8v5Drib8tWZhP6/jPdpvnnsY
wYtSRBLobXGQc7xP9pt56YmZUnsj2/ttAG2GTwi3pGcPee/si/8njp8PTOBrvw2O
5hBnEHACRVJ/Qs4D0PzPSX3hh0R3bpfMm3sC9QMy/e7UwHJee0fUh7FtlIbKEWHc
Xf2RKKcRnHvfqXx3GsXWbLU7uHgjJ3bLi4YzVO9qsdI2TqXvyeCZ5KYZz3h8buOo
9xWcDRC5i1DJp40gK7ii5k0cZk0QmfLjBJ2Cx3NGHjpTjRoWxHuCtIIMk8GFHCuD
IKG1Ygca6ylA+5bKPL3dCnXI6xsyIf842KpkZWRdM5AvMezaCvsHST4GD1JN0Inb
tTrssZ+A6TeRewhxoFmfgJtS6AaV/P1LigGrmkGQ5MD7Dj2sQnDcgSYPEF1/WNA8
b205TlM/lWAmdqCjYTRVfe0qZpYEjp6rpTPbsnJymeGsX8e+WCPTwit6fJDE/vXi
scVeaRnNJhkq1mWGCURMf4qk8ejeBzOAYJEQdE804IJpY8X+HgZ5CW1MVNdRO5vM
wPFIdgSNStwRLmPQ5FgJpbYCAA9ggISN6u3+mVuHpH1re6X0hsvP2N7KiS0oHv1o
dTtREt615ATWGk76y4686ojsAd3kO1gfbKYU+z0CQqsm9eYHlClK93GFlmaY0kvi
WWSkgIMiCJE8a2psX94DVWe/ZBJ7ccCNi5rjdkIuMsN271TAhu9gkGE1WIak7r9x
VQL4geGkbo+YdG2lhqNhWWQQxDUaeh3/tUrLrdSICht0RYqzXOzhVbfSff7W23hw
1ItA1h7niafyx2UmoaQRTLSlpAJ3AAnMQ2ips5GR2+K0RbAdDAFt4qaIUi6jbobK
7lNqL2F7ZNAbKQSq+DQnz8yaFJ8SIRr2WIECY9ahbXEIzAGx5WVMMlT5QGa5rHDQ
EdWz+xVJhAbXGh+1JaicR6fRa4t1lczSZ6aCHIdZjGyIimrWiumZMwR4axlM9Gcl
uoRqO+MpFlmwHaUReyj8De21nydqHF6lTg0hdZ8o0LU8O9iKkbLQsHQjyFyLSq1B
05cTW+tI71JapE7xmJxyE0u8oHHiObxKZ4SoglXwR8BlbNCp6677ovbDrfb0jK1p
Iv2TOCCJcQNW1Oe6bSqV+6yo5d3TYoyl+OLtbdAw9m1ao3IrUmxW2UaAdH+F9+0l
BdtdXrG1b5p64MciGo9U2dvCGhqDbEzlI2ouYw/RUJ4J0XkdNGyb81DyP499XHu1
5tQg0nEHHisMMEh8rwfnUapSdgb1PAUjZJwUC+3nesjff+EPqCd9kF5AJvN+6eoR
cI0Ia2S0ZdEa3RarsCq6NpfO7vYLg755gd9Hfc7c8sdFqgaI11XVuenI6RSY2HPR
AZWQ68sW7vkOwMv0csl9nU0D57m1mgz9m9j00YMdE/OtB10xcC/Of6LG6yDGG+VZ
Jc1X0rLZTxcNQBZ7VScMk46btjTTQgQpX5aiJ0eGAcWMn3ZI7OMUSxAfyF7yFWT2
fsEefZ5WNRwtmWjK4RMadhQ9P4JJh84+23HJvTLW7SjASodbS1eRcnBt+tXneuKq
2n7q2ziF7tieFBTzfRoVZv8hsOI7Is7qjXhe6th0pkHfDGry5VbHveMdw1HE1T5b
sfSq1PQWeHdYa3Ehxa0rqzHGJDW8sjd/b2Im7Wfyu2htdRU0UZoCHoUN+zKyUyAA
SI+EFBI0oEBQ829OTahJxzYkNluxOHKqhWgVTC3HmkovAF+rupe5g3iL93zfrfJu
eGqZFP3OPqmG419VOF7MzBqMfW5j1V8lkCME9sCBf6BVupX/FgQVnlMaBfrvg4FV
G0bSyXkwhsJXfFqA0DI9l6ck1K5izjXLziEG0HMByqvqsAVYAFQ4s7a7RnGWHmtC
JJ4L0yECTqDhJKwsH+/GnFBgRmtEZe3aMwnNt/WUyF36YS5Z//vEp2rJJ27lqN8B
KypWv+DSsHqU3Uy7e+KS4q59R8cIYT2rFLjM3dhe9Kr6YLf8LoJ7VD1NYdihMvfG
T+NfmRKTuRImN9nUucaLBlX85iXKhrYsylKJzzRHCwyAb5my8ISu38n8CVQZtPdi
nozqSIi/6859YDoiUR/xwv21hmiAtDb/VLoYHTxT8k9I1AVMCQLXLN+KPlUp8bFr
Bf7SyqKblChsOcSX+hvZz7V8R2/DqhvvatkV0alX0W0w3zQxCcL7LiEazueirCVv
RpIahrSsCpyGIRi5LAdNWOdDglVLZzj/vC40oO5wqoVDIZKv0a35Rsa3ldkngcpp
eoSq0VOTGbVXWjoPQ1POYW9y1BBO+KX7PaPikiho+OzRSjo/fJG459xgGnfrRhaE
VoTNaTmmFp1+JX40gOxuDo/1kOER5HWO7Y3KswIsqzaFqbvzQlUyC10WVTlAxqx5
KUpsEkzAqc24TWXWSt/00esNbCDc1z2YBXK8bZ4aOfHjWO9mYu0mlnoS/vGgcbnG
Xk0gnpDQa3/ABnKzyHAkDGpzY9YcGnVX6JU6qkICoRfnLMiF3Jz4arZu3qYFojRW
oJxkKIpPhGncUhnwWITYu/O1u+syQnuEnciLrmuvoMcs1Z9Ez621ErkHPv2evIM5
VdQhrHVkbakJrUY6u3ty2MQviy1mtPhQbGgZ4QS40T01jxWSCJQDKKzYXZAt9ANE
WER+tQ7NOp9l6jpQ1pR9IJJI2DYA89eHJXpHLYWBDCZTmpz7dPny197xm7TJkkZI
ByoSDbTxwvQnjj8MfazOkpNRXTCLZN4Lp5X3RrZRKAuGV5Anv/F2wdUbckHI8UJD
/KGRPShBGSnR8l1xQDmxZh3Ej8E6O2g3L2DkK710i1RDb8Yy/pU2khVlQ6TZP+Q8
SYDrcNNG6wIbUgkrYLCDWjPxTxopyeOgeVGr+rqtc0Mz5hqBkARV74SEAtqo2wBN
sfsF64/MR+p+50YYl49rOl6cBTgVgfR0tReqyGfLdrfJ74gp7cYXBKu3qgycWoQE
2+8LYC2lQqBkfvox3wQsGBQcR5WZnIlXglp8caLTGykYNe2arToY034MD85/edT3
w1k6US/WwsPBv5ZdJZn53uy9O+Sgkq/w8HNt3HEie2W1mnXIKF8601V0mxnu6PyP
w4lZw73tlaK3P8gaWOM80UvfInA6emqlWH4V8M5jNZ6ZAfgsTqToTX5TNwBDk1zF
bNzxYVuQ79nC96UyJs2R0G9Nai7WfOC63ldNH/7dhIgBUwJcHCYrI7G665i0cxl4
meSmgrBF36Stvd03HCQCk1Rv7VMC6ONX+P7rGwPbBEjd4dgvNUP7EVDG/LyWawS+
Aui2ns+y3CO9IZUf9TY1GwbOwTWPVccyKq9ueUPIR4kG2lccEZelYllJM62VqEIV
3qBHLf6KuirdPI/E2AIq3tDFxoFODb+u/5pZymH6jsTnCFxv0XeVgmfurDDGCVRI
6RlBppHFUPYVWmHD1X7rKhSpga9a6knDcGP9y0oq+IzLRUAdregM9DLTX/jwqnsb
StVvkXhDh0sgq9oO9Cqt4WLccYl1ME36gjm5n26r9twmEB/Vm0pRIaPYJiJIrzzt
zOmQ83cPfhP472hxMfoVce7WEiuSOPzQeYN+9YeZyUAgaielnSIePKcGbxW9mckx
XCqaGQy6GrjXytoAjlkotYF8VhRQz+8bmRf2x0HRDcrubFzjMXDJurWkNDHlX6xj
rBPFHde3jiZlgiZAX+pS693nJPoGvnk7WvqsiSnFmLtcByTy+W3chRweuZaT7h5k
ddtj8jR2vPp2yiE9IDzPHTR+h8LWaW9NN4vz4abFC/Vex+t2DQm5csdFHALr8Nvz
8byiYG2HlOdO81K9vh803CVN8MitkoQSSPs7nGJGFkJdYDkqTUiCaaRgqo9nIFcL
ImYxqqkhm1t4J8AUP9ufiB6AyXJHBpofodU8h8rUZQ89E7P7VTgRn4WEANWOF4Z+
t9z4nhFwBOHFKw7oK4n+gkwlK0xTO9+xK80KHqRwuA+eZ62i9Zl7hsQgK5r36pew
5D5ZpfVlGCG+LlqQh6YREURefwPwPx/bie46XrjfuoBPJJKp7DAv26gHN0U8ZfRT
5/6OtnONKAhHpUxZeuVtoGQRyvm4ifXC1oPz2hMdZn5IhjdsxPtBAE7/ZXePg2h2
GEUjfhYF8o6cfMJJG9yu8LxB+9uiSwXB5rj4DK6lUCpVaPS3v3EFdKN32+iQH82u
OAce3zGzO9Wq0rshy9akAaCqZu/PPINa6br3WugBf59Wick3DgUA3gV30JPdtKkm
Un/6tTK1wPAnOjwkFXC3nJDHU+AyzUpgBqd004CBBr1EMlfcsUMAttTO1z1rcL9l
bT6PcRxFaG5EVpRtSya/Hk0/Ick2mf59lveAhSCmzkkkPMjX4jx09Z2UB/oTjGbY
m391o4tpUwCEue+K5Mm4Cf9xMAxP9Imt8qjSgH/1edUICuIQrUOf43ChOJP2sNqk
5T+Pq2bEcaOazSTVcrKDpxndrGT0DvpIxSjxIEvSwl6vCO4dtL2tEhqqor69QfBp
9/46uprvXQhgJv9qmx16qH/CqASbmdhuHlrWFxRm/PE7XUSyYYCpF7/bjjYuzt0i
FPgMsDCaIkun3ESHl8yxX/i/TaKLwohLFumBKNrgTjKJkYjGFPoG9QIsYMlnqs+p
5HA2Vt9QwhW+LGDtRQ2hAskjeiVEZXl5t/iNoOt0eo3zMTUQ2XVDJoXfB6tYku4u
dS7hDXK5vgaJmERTk2TDPVAvQrrv2eo7eq5utOg5JbigJ8BbHmfxtjTHypEG3WK2
LwPqnpLJMWcsmwY8p0RBOl7obnY7GoB8anVu+jyoaItYvTYJQf4hs/MJIUjVtWYE
0qqs+e1AvG1QoKnVDjk3EWwyolXSLOYw6BkpkgqdXZAiW/hoPpaVvKs1c7xrAaFz
aEqfl5E+n6tvLn6bszmowphJLIdEj+xH+n0Bl0X3Tg2CvGxHzuZdmfCbeAakJ9Tv
uhwpP9CP7irbG36W+cqjAo9mFfYSRN4ZVEgM/0UYEduK5UHLh3Ix9oXvvu5Qv7Sd
kCWn3dVq7AWxRH/cHWITMsAwVepXm1v3zDs9M6IvuLEG1QVYtJ2N6NdXyuO7MoCw
iKx3/AUn5Z6gbkwbLfzjXxOd4uAMO9pHL74qAJwhMTRQMjUofgts9Ma7HJL1ZmAK
2kp9zV4KdFcApSUHwG0Aje6i0+c4mA5uz2RxVhicM+ZMEAifK7/K9irri9z2MVs3
0Aad5CHIDdOKc0b3zwu42znLkzmIeNQQRaChONMm30sASlCsgHeUyKs25J5B8cBi
3H2OgOGaQ4DBRm2hoMT6qjQyeNVUXzBrv9idxbZNG84FFbhPeipZyYDOQcLPiS6F
Q4aVcnX4WfmHxdeAOtgbo0Xgo/9B7/Bx5Cga3tGRVNIapyOWwlPeSqqSzMTEqjPQ
VIT1s/oW7PVlmBU3x64PqtxvUDvt0d7yUwPeNfOELrYdIU2XlZNqMznFjTfgxIX+
FN2yNr26UrW6MeNPYJPVPbhSGdInbnjUdqySN3GGa+Z2UHWOHatBf2wXdnNoltyc
XVwFroJyrjniLsQjuaubUGH8ljShnWKFQoTH104XHPB6Ng/HueNZiUnb9UlIh5i2
1rhmaziU5ZfCQSSLSYf+QCTP7mmbpe7p6mCKbON5Hvk+7K4pE3Wp+PmSuD5i5glT
PHxmzpfUzSumYNQ1dR6Q2i01DxreuOdUgZaOc3tHELZlVlpv9eE73nfhu/Uy22+O
jDXO1SE4GR0DKpJozq4rKI6MCjwDmENxJmwCnTc+iqfUz9xaNVhaX6e7IFd44ktJ
NRF2jCF8uPCwvIlq9pMq6DmKQ/USPb9pV2tKZ+rMN9lyHCFKdz4HTEaMIm8MAQjo
s5NXyneZWrq18J4Td4SHaz7DsgZkIKMkcWNyCkm5Dy/3XgboWfiviBy+wJkxzsJU
kbNxRoTmYX32F0Svze2y6QFy6tEjFHJOEU6jcHSWzhyCuePHYLRhdJY02rr27RAw
MqHdVVkh2bOPdL0XE4fK4stqwXwQNs2iNGfaBFWYvm/xlNZmSmH3jH1phaHOxF5F
qLBwZJhRq5uXPc06f1iELDzNhrFWW0YzJqwpuckNan9nmppnoxQVZzp15q23r2IV
4rcSenUqTA7NJ6G0+Gpz+b7vMX/JGqmoZWH9AyAbOf9/RTU+91ivQRU2Y1bV2nzd
EudLn+g8smAbWCPunrGTiw3nKy+S2dCW8KsF5HqoyEL0+0wGmJFdDqkdJdKicrjs
QIAac1KlIHXU7Ltjfl+YRa+lgNz+BabfeJDON5J84nVC6gI3h+fyX8TdouL/T/l0
8aq2iXjiHuuaIWH0x2nJFE2YKXlkiWW892Tk9idroyS6YgMjrmE59XRYrB/O46Id
W1GVgS4+ShnODjWlXSme8EyuKqbDntCnbSFLq1cHLFYuYdQMYTzwt1UX1A1K1OfO
ScLhtfzZOF/4NBCuUIVcw7kzKYFNFjQ6eGXZKOae3Z4GGpW1JFc0VoGZBlP8XtrR
KGNEYBUewGjobQOkbGroBZY178rXcuBlNPExp4t/iGcmwRQovfz4v7MbMIKJFlkx
VdD8YBQBEI73vEBHwgtzuqIuReGqyzLqxbWJQYoZU18tR9oJuEIEGAK7fXxF2rtD
IKHqaZRX73odk6hJw7X323BBdmtqt3JC7jHbaZ4QwPLsDJir57kDSO0m+5ARYmrS
QolIjmPma3el6Syls86XvrmWn2dni83TNzIT9sj/i2XxVH7/k4REnR5SXAoUDrF6
r1wP1J0gAkr02pWu7NzhElM1WK9H1dRYS+w/WyPSpwcJizGIGYxr01rmdkz+sqZk
VX3ATeXnFcMmkpNrcIMkMvURB6NGFvVK4u73u1C+CbopbKXnRMYJV+zJ5tQ7DGDT
8fyCNqUefYvWWcSkJf1dMKSeCYcYhQCJE2H99WUbMQwNXUe1Sb+llmwey1lDyUQd
uqFHXV4dGbFAyp3Dg/dDUm/DaTOLRhxQB/e5GEoCn0bNPF/By7ueeLblqWb9CQB8
qBT7qkUU0ZArFN6uduTFSEbfFgRAMgd6XwD4CNrxlx0ALACXWTgvxXwmY7QvVhuh
EQQrwt55T7qXbPb4QwKTal5vLHzC1G9Vkzq+XYy6ZnvQxD8wLgxtleFS89IZ2t+R
bzFmFKm1+Z7OSlkkEvQr3aejfb96UxCw857BLgzy6pCeH8xpyCiyl+BlFUBgT/ZV
PHq8BVc8mNY0BnwLKYOrB0i+kJWywdu/hmGMGBzTmIseC0YMPZgSKDGxvMvML53Q
Saz87pXF53s87ba++9P8SYt5oHYgvgod1Y175eTtOGBG4fZimv3WSHwn7sDF/EJS
IlrIiU+Gf9PXlPAZGAEe1VXau3VlqDgGnVi9FcPtxmACQRoJd5zYPtVePyAqgov9
6uHQ1r2SvdgaL93jTLvJwvzpAwOXK1zA2AJ+Zd0uuC/yDi29hvBd8r+xGy9Qgl79
uKjOP6Y0SN5UhMdbit9HvF2HbqK1SMvSKiCIL8lHiOTHI98IBOlKt6zR0GR4zkL/
ea+DQW2mcedejt2yA+/caj0v5K2i84WCPyN58nbVENM/V9xOfIr7fqKg/w2akSJP
vSjF0/xEgPhTuQH2d6c50KKjuOco5O/mLkW8LZdgT3oZn9NycdIDGg7M+EmNQ+wH
A4bkusZpI3L/8r92nYo9D+kM8Y9rAJdK5IUZ/FHgFBCpFbCWI5XbSnqdaqPJbr84
ecSFt/mRR0tHEl8eDovauqHiqhL5lsJqq2rKxJQzXFNyibdu+TfTkL/5NktfxIVo
pI46LoAV8zS06ZKlABbvs6iTCyoD+6btnJeBDxG8hMk33Y6V/Po1XrhMnuSxqYCV
W/5UnRkCShvlQCZEEkWEExNWhF6f0DZEINyQEiEmpSvmnlukO570HxWGTN38ldRP
EJrG1hub8FR3C7lsQlTGG18G8VfqcZuPzCVBI7nDAYzxRSCQzZXrOpRMGb/FtzFm
xgZI7jgotYyzE1zxKyx6/IljPJCN7t8r3S4pFrT+Qyhx8toSudSz8w+ZA8MLkVtN
z4BkUQ5TW4uZCObHqLcdnc2HwPOq/kvuByPUZlT91s+mk3Y/fsblsVr1i1oUOTIt
AZUo7+mYBncsquwGnqKgQQ7tMhG47wY5jJJvHbb7xJ6mkLBxnag6vUU99bThjtax
9EtFDWmOf7XEiaQjZjoao2BBGz4h+ostpETaovpEkpDNXiqTHo4owjVEy9YiyV9P
paA1ZtAXB/cif6afaHGEexwJNXzKOchq6iK57Ayn8jz4bLF/DpCKIn6+B6Acm6m3
xVEtSP1M6KVQZcaOxVzbTKx8Tzp9nw6HK2SPTiHZwR+Q9tfIOzsquE8kQ2ETLD5Q
qzZFXCC4uHrTMh/XVa74Dk1tnO8Cz2cwkG3VjglCZgqXavaHGSiDciwStahvMtoO
gDZmIUxgyWcfjMfxzb6KBVqFPYOGK+2AC5JzZcyCxAmFhB7YwloHI305KQ6v+Ico
xvb8TO31vEPvsu0+VxPSqLBy/P7z4mn7ZGM1oudtcyp996TlcXuaKLi4jHDBDOiC
VGyf7mLVujq9Iwict4MLSKWK+Tbi60jF5tlQgMNhsPbUMpSGQhZ/Fbs73iKod72c
3TJSe1Sg3L4SW6xjVfLZ2J+/6E5Z1/hFxSVIsLcrR7+n5AmgcHavFD8eSwzU/JfC
2FGanc1bNWyEx1wDlysKepJRammpxIpg0U2Z+55vOBQgXtRkqurtUjxKFWszfw22
wZNC2MoEeoXtHeqydUrWLLGC4vZC2SFTgsfm1ulZ2l3tSMfkvvjKxvbrhcXy1LKj
3cG/fbMIjJK522VH7HLhthE6XVLS+EvtPyV8ixozUr5vsq6dg53p02HFClSD+pac
uOKc3UUVQP5/DKo/yHBImXKcqJCvfk7KKNyAPcFuU45eMoSimOiFE64cmYIeoR6+
RucAwDvyZD4GWG/46LFxCHXQ/33kD3PJLb3dkJyPWM0jGW+hDhUaXwaG1ijVbPvH
A7U7aPjtC1d1+tsF/2Scyy+eK+CBDOdS+azM6rpsGKy/bgwRIzbPE3+FVsOgJF65
aupR/YPuElHsG/IjSMvbOYYASUtFnOa5Grxm2mM5p/LepZLrviccSLqGgsYsqFml
LY4MSElhMaiMWpLVDsdrUDo6YQ6Ts4LmYaFSrsaISWlxFrWHJHNyo9OBaEBe+qYh
ax8wyCOHekvq+RVdCCHWzlVpVrzntzCc6kx2l3dwcalha+tRDz2jbtMvzwUccMpg
Wzp+aVRsvDqm+O0qcuNOLYSc7FgIlmo0nlvt6qTThYsVxefhpP4zVfFVZ4alYVfv
6TNBZKQHf2iTsdz4AX5ioqDQ86/GJ/nGNcwxUdbrWI3o5thoRV6CMZPUSaQ3JJS2
ASuvfb5R94iabCKsWEFwr/3JWRdmqQsQ9yZt9VLiMQNN5QvUWCUvILhB1h3oL5m9
HlnA7TmNtgU0TVF7T27lpicdixnDkw/2AytXWFB2aVIDkH2d4dv4Fs/vfKSkTK8Q
Nc+SpgaxssAApx8MtKwSihQZEaQAivIyDZQoEViSJH9dD42Zvjl/InaYYMpl8NPL
vXyxcQl3DUW9E6ZoT8ijc319g4EOb/oU/PJmNcYT117iNW4DSXRSyghb2l2DkxCb
V6x8Vfj1cBKmWYryx4ORO6JpsXdalXgEl/FmtsPOxckYKV48RQl0pYchK0gzCAJ/
leLnv6+wQbDusBDiF90VmDmMphMSmOVdo7S2MZRfmdIBa0laMvOnxF4YEX4VJ+An
tnrA0EX+9XLUbXn03yKAe1KTiWREDnhTyvanuyhNQyRvWuDchvkEjSeOOddzsJ3g
1/wDzOTlqNCn85FeQErHMzr/4nVU3UsB8bd8UVtZupguOhebaEGthH7R0UBluxUs
o4ileQff4+mZS39Jm2t3T1X7i823FQvFJ6xIGdwN/OIyLtgGfj3a+S+7P1yC8gek
Yuo1gvz5cXfggu7TmXnU4IWjeFSnMVUhKPMgZE9cH8T56/aQCJb82g+iD8gBWprG
vZOhV1uwLYD1XW5U1ude2lJfbJtxwNLl9O0o7g8KPyT7+tMFz9LS32o+V7wiHSj+
+rnvi6yPfydJAAC4PSCBEBjB4p08I+woHYSNUbdeCzrafKxEuPypaNFwIVppcv8F
crWMk7uG2zWjs1VSf0DUDjhqte7p4DLVG7TNL+cViVUWKmRh5hR3RLF722dV+r3P
0rPEYt/ydEVOmjsjwlC02uvR/S2XAqvEv7BxLRnZKNHiNCFQyQOITI0HjSXzZV7W
vFh6mXFSvhLY4+w2FcVPmVB2wzyf2ZnKRYMz2gG2XsXk5OcXfb7XIAcRpuSfmPp1
EmBHoBTouR44UfOJ+5qvimRGVvUzKX7WL/IvW4ZOrlRjJClqYC20jKdOMxghGNbu
erMRAJI1oWYjKsU2UjjzmluPyIH4m5AAntGdv3Do54Cq1RzYnJjYl4cgxV6QOroA
lspyXFMxqiZZyAF0Q6GYmakmIUO1AeBFip7LaHdb4sAiS+AgO2ofcIxitqR+CLas
dtD7h1B6D21OCVnJdHWTOlylxnyixFr+yr4/e8EZcfis8lPlLKDne0Kzk1/AhMB1
tgQy9Zar9XDV/ZVD3qhIRJat2nUE4soi+zcRusxWoMBStTgrRSps9fVP3IXaN8+H
x8QjNE58m+c1ZkBZTUEbMDYWMTyXMfnVqimVA/WB7qDIfkjfuM9EFXMaY5MkO97v
GsK2mgPc1bvsmKdN6qF7dB6m4hXxjqIStEQWHtAopa/q+6w4IS02aIEOmXTpiCit
NGysFqH74QvxPei0FyDx+6VIQsV5vyBxW6bg3zboq3qf6Mbr+7Gu50eEXWptLasH
m54hm4g+ZIFmKSe9Yhtf7AaYKvSujIYCLqFnLtBaa7DzUM8X4nx4jT2yX+HLl9D+
E9xYNKQEY2qACvjDTrCvJIGWXl0qwB92KFEhipyDFLahc66Fzo5Jts6y8rwWaGIb
ksxTGWwkxI2zEEypgrx+yqR6nXmoczXCWmCz4/V5SU/i5mS8eI/VYCMv/iBpI9y0
giVFtfcdF0flaeHbr8+jn14nct2YWl/p19q2/xcB7lRQITrbrHz8dJkcghBg79FV
P7qyxFt70MiabTtgRdn6PrFC6IbyE/q4KB/Bm7J+OGHlMCaVjQU+5mgcN8je3/ix
276KHurwrZ7BU8HhcyOi/JxHD4SEalk73/MRiA3dBoJIlmbYRO6pPm1PSxYAtD05
xrpK285CqPi/TIU0BG4c0dvCiRiucovxS8U3Y/P8XXOufmQhdQfQGnIOnV4ydWFX
vUqanTQqq1NZewpNbWngd5qRdAZg5Gk0bUsLhImUYRGeWaTS2FOAhBToNUo0cnoz
aJetPPRGWhDsr1tRnnYexJ5v/4Hspk87/H7sEuIlftME9BzkFcnQQ8uYTnNadMU9
ShMDk/atO5uJ4/vrguQEh3oOyLKg/GtmhJnoJPk5S7w=
`protect END_PROTECTED
