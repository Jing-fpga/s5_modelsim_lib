`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9qs/2cKlxG0DWBaTba+FcBsskcHsY12SDtGrw38d3XBaiC1U2036QOGa4F6KxkGj
A+nk6639biMAyJjAXvQxxSnP5V+UZIl/Ysss15UdWlBHxOXLZCsaVUwEPMhS+SE9
ZWuOs7sgYlSAxkIE4cEjE+l+wr+jGiVkvM85cPKKEXtOEgr6AhjE1Vc0cVk/XSuV
ydyRHI2eqxVKlh4oDk437YFyMHPM+V/ODjzT1/7IqmVnro/F194+hHpt4qMhQ80C
wW2yghp46eG8B7BFxpwqIFGVkdTB1LAdsoZ1VFCWqcFfd73ypw8iNVEw1EM+jk6/
vowjDclp0XKcATdh1Yl/JhkNBW9nfgczWwqrlJNAy6cQB5k9Z1T01pbxtVkNE86u
mNA3CVEmPURbyrdd9QY67tu+oPLlAiD6aZRXNubNhtMArZ60uNLkLExRtmuisVep
pASiBMzbMabM/KHuHZFSxB/4OAkt5Ks6zVdNEX0pXbB02HxWbvxY0wppwBNAO1sQ
KmulDfX58AWZyymyyWw4j7Zmc/xa3Em9ta6ztrq7n/F9UuoEP/szrPcv35dIPIZn
DgYRT2vQXE0JafnkA/rNY+nv5atvnlI4iNioIPChqrpzixSF9w/Wryl9BkIO5ta5
P57b2ZlBOBA96coXJOCVWnbFsPcGi6LWwC02igrl09FzpFPWzyRKhmHiWWBfkJYq
WRa4NYXae+zw7lKQyPqVpf+N21Cv1fx42MCzYD33U6/wX3SJwUqUcBoM4NF7lxJi
VO9HRKBGnRmOKZDDOno5r1RpT1D5+6pikG8HJ+a3wGuS9/Caxj0EX2a+6gjT/h52
QrinEBJJfmdcxE1BzVaLwfHSE66OxyrSx9mcvnsw6u3NXIoIY7TpHToDNWxyn4w1
nhsEL4d76FHdFwu1oi5/yeJjBqNSFd7L4gVXDUrFaw/Nbb8MaSBF+4qe8qku09q7
7Og9GnCr3TNyPZbjokXr/TXe4jUnSRXrDgWs4CxswcdRLjydUDLvUyatVi16B5Wk
dhmQOixOfvswpNvAdan7zl9v43vsZ67pAW/+knPh6lcGjsDzd+jJ3JrrP8Yiu471
4QXTvEoDsp1lnPXoMls0I2mQ/6SZleJIJERtT/BLdM78F+n8BpMLih5sJkhKGJIU
l9H6tjqr8Ejsa498fe+jSAfwCfIWMOn+Uv4DajYpuPHO8MxbMB4PRnJD8+pzPFBb
oB85l4/ittzYCJB2y1jDoB9EdEDnhOeqHnMYxlyMWAx0JgZ3JEPcMPh0tCf0HtY0
+xE73CDjDGXAso6pRV9BEwM1Ff8xZKAVRVl6/XrqbgGJJCsBKuqr8mKM7kom9KbX
bncORF65modipdkHRBWlHPro8GRJ5aSLp8NrN95h89Fp3RtcOQnGkNxcrQN6ZYB3
31n+KEYIMeKni2j8C2bz/IUsvErwB6EsJdtsLCrPZI/tWO/cFztTseAMv2K9aWDC
2XKPsI+Y/5MUA8NsWdYfKGkJv/gWrahYba0jIUULBnMGxAAE/4bIpQeDBBbW3VuA
hx+JC0P2d3J3+Cx0ekr5pylx8bLE+WdDkIjF7VC/i3vudebdKEGDjSuDdUx8tosY
TQ+fYzZAdwkNKoFaea49psTgjm/TmJ9D5ayNQDuCFMukFXeIhDU37dm1mbwdDemA
9kRvAaVIlArO3Ic+RMOqQfgDTzTI5+PSFHuHhwtL0zzuZ0nI/jUYANDBY7xfUpJv
nnkU+oI+toBfsR8WfIJtViF1qyOIpmmKX15ONn1kzkk=
`protect END_PROTECTED
