`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8q6Umjq4GEpQXoUsg4D6K3cU5Uu0Yn11gOq7CEPQjN0lIbzEFf2kwx2yHKtJrEdx
nYKyFwWk5eXrOYKuB8uFsxKuH7FKgYQMnp+oSvobOv7TIuHTyxYyyTPcgNVDY8TN
urlQsbyCo0u0XH4LPIPrRynMaCtiIvVGHuSzE4ST1bfhFLb+Ycd3WMWyF9IoXc/I
hAlWc/BmuKf8gOqPtVz1ayLOfjGswjQO5X0fSuM5Bi2oBFY9vMxsBJAyNAA+eKrl
HLUFVkRxVdC/BPq08uIFJ0tOH2c32V5GjarZTZ0NBx9lsz4EpUkpZY+DERTVMOIk
+PB+7JU+mOBz9rXrk7DKERTJveI6f1YCnIYaC+lvPzhUJUG2jrekVK7vCpzE9hI8
/2jUm59UwpzxEeFivswX/SHbdfTFZd4wsTIs489KfnSofZMVlPXDcc6aaB+jvQ6r
XYon/W7Qn4Fr8oZ/obd4pMTy4vQzD+vGRFanoVzyD+U=
`protect END_PROTECTED
