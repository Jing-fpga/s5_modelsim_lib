`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xcaJ5x5lnkvJxuijbGhFj4cxRiaOL5IE/0ETC3Fg9l3rfc0crTEGLXNOXbdg1MMU
FFZEK4bAJIW/K9pV4e+jvTQqfKG6/h35XvxJ1LJOEcUJEHq/5F/eCIGRZU3sMgUD
uFTuRV2auAQViJjaiMg0T1Rnw3ZyWHTvsWa+jmRoUqK1w2HfAP52gGIMh8k+uaDl
tWLUNWAT38pjWqhM57aa94Kq4YEq3aklbmruOsu0MpburMnwLXNB8nZAXlLRl2QJ
YuP3wQc0WxC/0SHwc9ppPqAuuEoiiC2DoTZUG83JK76VQcBL4pG2dM+LVwMKqCSU
QggRYN46Ut7G1ZSVP3c3fkz3X4IsTsrG9rg27CRt5Gr9/9fTOEJyUYKdzXVmkUQ4
Q9AghaIGpuN/KHF8Ca5mwuMdXkTre6D0sQiXe2iBrt5y7dfXhV+k6QKscJyMgjs3
kh8GguE1Q08vOt58HI023ikmOFzHQ+2VDlj9nc/Xf1P9Uw6BdH3PpjS4iMELPQSb
Sy+UB6oOL9KCO7jRMI13g+zA5NeVd9cwg5twJiQo2iSej6VtQVucWwMqc0b4RCl/
YIq66O/7weRgSEnTsGeOsG40BfoMheVEY++HQr0HXO+/IdVaEwWJpI1ZdhoySyG1
XGx1020hQvQbXoNROzC/zh9Vky1Hjmkq8X1e/jMOIDg=
`protect END_PROTECTED
