`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZbyTbfljBjm5kEOclWJWx6vLfJUXPO5MoQQd+EpZb0V9eZj7LgWW08FEUi1b+EW
hg99Fmc9uvBcc4G7HAbbjJSRya2hq4HHFctoTRQBXycrnWW8dgzJWXB/Of7bKk4p
MPJnmENpVehIeeUpCyZb03aP2WK/sUEg1Bvxyil3AHS5WB5kJh9pToSEHgeH8O5t
ASfRNpv5p+yZu1PtvJ3aH+BBIzXYI20PpfXz2XhXlAhNlTLkMPFzsZELwPMhUjms
DOFDulKE6ByGQgmbl2Jie1spNIayLuAIqqXMDCJb6DDVI0rKUX8mjkC/1qndKQ0R
ikrIsjeyiAxyZ2sV1Bb0Xbk2+SpjoL3CWUa7GCJSWDmkFsZGryzncTMVred2vybM
3DG7cNAM0CTGPaqPP9r0DUGKfZLzLnxH316OiWe+tKClg65jbIQBBWXRMJoF0qca
NziiDZbOAxUtBGlDasHIuuB51x1VeiEfJp3iFkFDGZ4qhPIMJKi28BLo1xnTxM/C
CVkx4fx4OMcacYJiGMOtJZfvW76rc988S+/iDhqXCGmHen9EqpQfto2LQLBK2POX
p/+jwoYxtDe0LMRyRi0daCK17nS4+Y/2jbc8DSj2tPKdeDMwBEsvRqrl5yv3IC1D
bsAmiK6i0mj/5KRpFTzUumkxnOkuj9GKQGts1INfMCT3nl1hT7/aYOabPQx8knec
YNxqYJoi6ICefbPvyUS6IeQg3IqCZxX9xIK3F7HselM9BSQGYelMhws8OxABcPfH
9pFaj6KcLFIvbRwGzjKsn+Kjbq26XHBuQFP6hOa1MtKRu7kkdEOq8QTRL6zGlXQQ
ETh2eYvmEL6gtlpgfEA8plyOe912LiK2ulbLcz/C/jvM2p0z8IUp+AcYPD3q2V14
9Gr5U3dQlnLAvqGMDd8u38j1ClZnZe3CT9VS4RF8vrVkXHlH7uzqdXZvn+ckrJpO
/HgI+QKe39dKOXed6KqxtmxuQUpuyF63O8oq4gZ7lB1TfX0XEAumDBXIGSGDe4kx
ygmWkouX7zVi08EKgisRDiWdkUcBiU6zP+KPNtLi86v884jYr7q19vP8b0EfknDw
XFMwNEzaY5bK5EPfz9+ahGDZr4VhDKTbuumhuFOgbD721gWfwpGu9NjbRc0/rYX7
EWTpcnZZmTAggfs3zaq4Ysj+ouHGnnE4vECmpY5CE8f6Qg5j4E8Tad5u7WQz/GGA
Jivadj5M03+jQ4XEP5xHDcg5ENng2AXRakt4Juy7GgYFtlMaS+QdJubaQtwVv6zU
oCn9Ivxyz+Do+W2HoPguB+YN+REtGUbXKKpR1M+SbHuPu+C23xZ96QDXnDfXgB+4
J/xWFlEifrnoF6g2pov549+4bb5/PN8IA1SiAQ2UIxJd91VonQ6Ln3xTS3tJ5KDQ
RqPCVpHxg1ZuqVcvhlFfNBXFmQQx0fEKb163T0iHGMaQcwf0Xrkik6Houov4NTcJ
8U5+b98JmpO0xsVtJn2hrhODZvrJgv9sVQ73JkArmL/aIe3ladT3Hf4XkYrHeJ4m
k0GtQVbpy78Gzfy/YE11dA5sUbCVIYCf+q0IKpJfEa6C2+ckP+1MAKpvoVhul0w1
yfQ6TU1QULfEwroVSpXSyE0kHb7Fxh/wLlLhMDJTrI9mmANvUFVimfzDQx5RTMlc
y8kTaFuwAySO424JpdJ+Wp5oCcc7Q1qaAB3L9ejiNJJSSzsMh3EaNhp6THp9ry5g
wAaO3MdAZsYPmfKOccZ+dw==
`protect END_PROTECTED
