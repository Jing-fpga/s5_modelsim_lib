`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OCXvbS3Ix5ak3z3QJqeDzsvon/6ada7UZuFLY/rp/p/mMHFp1BfLqLEg9SR2yn/r
ekL9jzeG07/XYxpF4eanld+oEti1ZjjNyZ/5vYZqp/QgFW4lQnmagZWMEILNdqzk
0/0vrLveLK0fdZ6S0i6HyfzQD2nziFd8YyEXFq1PbIaxXy9o55zLLvjN7C4LyXOg
mVjS6DBmi9/LqxiiksDNoA+sqVcWp+TT47l+rr4tkP+IyZzThKucFYj+rwBoodd0
TrklX7leFSU+Hq1GeJmhEvE7ijLDlXR6OmI7IDrTL2pucGORX5UYJDO9ECnFb5a/
MMjLb1DerT/3ZquRKCYcXiF29dzYXzfMyhUWjL9DkLrX7+SS30sU24HxmDOwLaI0
4RUsAvyOYqgnpQ/5oQOmodajh7QeIcxSZ/cBnTGHvjbR35/ysnUlJjgiXDqKTU9Q
LezJEiBfGjDwLXqQH4t5KJchfuw5KYo4gwNXxDC5fHDgyhAJjPts7k3byxgfhSVn
gvvqqpOGzPAuP8smWeWUAL+bIei3zqDQDhd+DvwlZCGpDSuabNksL021yTJxUapD
ZSHo3WgB8/55KRThgkYnNmR1lE35YBFsrXCG7QqnCqPiyCOVrYpRivydZF511IvX
yB7mNYJNGffmBwVG9nYhzuavHuc3elhit5fMXrs01PCm2rvgwyia4eHaNPpLKeMT
TcBDAzWH+8paoJcYgrj651nESAaa1NRDuvfDWbPEuCEHF0eG/Rt7/ZloPwdP0Yxi
WEsKL3/+0qIG5Uon8GmLGf9m6Kd/OK7O4nepD80PFVeJ0vh2j9gFQig3Xfhi7ni6
P3R+1Kvc+gvquhxOQ3Ijrw==
`protect END_PROTECTED
