`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ii6X8CqUE9yEpXjKAHStXlTZHP4ecXxp6IUlA1Jt109rkCnSJBjeRJGjkTAJG4vq
4yF1YlgU1Vq0j0vboqfCB3lBsjNbB7j+mxA2r0PnAZ75qjYFbRx59dQFhiSuCUQL
pqPd1REdMMb5hORJ6g2FBKMeLodZC4m5GVPRdACKgH6sVDHnfjMgnadgvQjId7lD
GNHaX011i0c4giZjDGiqZ8+O6ELvIIIHFiLTNCznLv1K/BK04BMqov+OXHHMMY1l
76/C9CS+biQWPmy0zFEyrTz/q8MvpxRBrgBE5SD+oG+GQM2XVNv57EhXdTiNcOk+
C3CcwXsRUDzKqP9Xl6CY/LfsS3lD1vJ80PjaHvQXce7H7bSlp5HHLUdsC1y+9+Cu
5toy8pXebBm/mLRmUDQVOvgmYUEuPAafnr64+vrYDOzdyFSpkuppbpQZs4HmyEZk
YbDhF+1bPpiifrgB8tV7L95yIP970d5SjvvUa6vJm7VTt66f9MnJTDSkN0Vejzht
4jZfudL2yRQN81hwkEZrWc+Zkt13qV6jVrJskeW0uVsOxsYtR1Q9Ig51VL1FGgok
QfU3K3z9FqckqBoHjrK9q47i4ClK01gm8QSnEl2UxfvQR0XcmFJJx+y3gifnldWx
f/wOy+4HKjujTERE3YfPTX9phRPTDhn6jDdqx/0U1lXfMGLJtj+nwCwYqmX7wFk9
4MPcb1YxWhFZJCUHYHLaA0/BU0DXxW2xnN061B8AVStq5y/VuyeWlmJcsGZugqto
PPrz4iEZ0rD52FDxHim/Lu4fTx2Lwsnr6pCDJ6gOZ/TdVpK0kPtaeEKS494rBU9U
SSOhYPES+1NRDsjxwRFf213qn4vdoN9650/FDWxzaAN9QqWbB4fj4C4wTApyAGVJ
XtJG7amzeGzuiCoZadzFEOkaNkh/C0Yd6Y+7Xsp7ROJi8M638oOsu6bRjt3d1etA
ChyDYBF56GFHGBsA1T/bTjcFkxUchBSMKjslGhfANbICdceibR3G/vqAiMuqzbLi
82P+uYxH6Q5IXV2/XQ6A9uUHeOgQJ/alZU4hufdH1owFIbx04hxnfxCxHjjJ2y4j
sBwre3/R18cwXbRqC5DesqdRcPFBPUDvlDLjQThUPZUQUiM0PXxEbH8EuYX3XL9m
6tIGgEmyYICP2gLl/zzi4FrAVkY3D8VSjD5vqnhILIo1Nie8zg2XEhpbRLyqwVfl
GiAYLyr5mFdc+6kB7bFja+mGsO1WruSNzvsd587Iw4tfI0tgVyowkFVReq33NtzO
1F9m6T88JOWLavV5RV4rZRZz+/xSvJfnvnOHwopQhTbaF4auZ6JB6bWF/Jfq3usD
Dq+bvdKHJ3UFEMkNF9cbgqHn104yHSvD9P/9zIWSC0zcVPrPffiWxpX/s5vR7F7Q
eXni8HS5f1nXQ/Kj8MzAluLr4HO3Kezg0yGNlmxkdWs5/jOFP0dTj5NtBIyAJwuy
dGCt2RsTIdqzwavUDbIUX5M4O8Rghu5qMGCXxiRm2nFv78XRNJbCmip2WNubdwcR
9BN+M+VhGITY4025k8oz1v2B12dkI4xF1hohjwpPq9G7q9oCQWPIbGaKyVV0lg+e
97nSit/FNo8j8iBY+zXv1uxH1uMfATp5O1OivGGipl8pmpwwee6UpFXqnmNSLVut
lET6EA4nwcJE+lPD/D2bheME0SGxudytzuBvQiZRPoihB286b8VeDyXmqu9f6L+G
MQqQ+xGz5qkFDS7gFQhmK4J89qSvavJMNe1PiznxYqDtk+YF53MmpxCyQYwFihDK
eXs46NQUpkvAZbdYuwaeTz3gppOVM0Yoaf0HwNHsIvwN8Xu2pF0yP+zBb9HHuitf
DjP7QMmB58zvRWCeUuUfWq+Xr5kHZiRoDWk+5U6uo1ZuWToD3X6BtLrkNnSmExYg
AFdzt18nNyEahZtMzcbeCVqIss1gPoGYMHDO1wYcnuzmpNK/orM9mKdP8jex+aXD
e9OdBORm01v5dKiiO0R8ko9BblMozFT5og7RG6PdnS3vCqkZU6szzpT5nRl6zsbC
oUR9bsdYv9rWh0IxLwi6AtpRDH0yrdPIKQTvm0tbkTqkbx2iSR+qFIBe/pqEo2fz
wAJY7ctsObjD5ENOutz+T4Xk5zgbq1hhWbTYPYjFXM9psulY81yFK03gz5AKEQ0M
282NjQh6RICRZ8B+uNR60TEuUEeq7KUG7HKwH9J4q1Z4IfIOMUm1UZqRpuMxGiqK
EieuMxrz1VYCmHcmJ9WNnqm/UQKno2Xc53wh4c/Pp4u0cyM2MLhdvy+motRbI4wy
gpbS/Z0y4kCl/JKnuP3kQLortbKzmHfEI4zompBK0nBSOebXpEMs4uClOhARuFcU
SgP5X+ytQ70ms8jNY88wovEtNAn1+BBoSm4uMdemJi51ZXsyoOI/lzVmUJ0GD9tw
YdkGASGcfqsou7ddDo99XV2sSca5l29+uAn3cq16/DCTl9FMkOlQz2GDujUwRIP3
1nqi3t3a+AVKjkRjRf1Ed2SO53fHE9Sitl5A2pOY+hZ3+96bmihgJ2Te7FISZ/nU
70hoGhnYFwdP0c3uqWjunSxyf8jSNJtFJ+q1QjyaD9TnnKoaIPxxtXj2c6XiGtgq
cxABwO7zICSybzCMMZizmbVxUcAHymuUABo2sIn4d4IYFDfM5VnM1cyd+O8jm9qw
RP61K8hJ/BrRqjluzxsIyeLphp52mxjdoUva+fWaHqIdLvsO0uYR/ePIxT8+k0z5
0TvKiyU5b+Va7aR+6TIU02VlqS03++wmIfES2J/Dqx3gBDvGh9Ut66SKZP0DtTYM
FQkfKlt6vgTHFI6GgZY9poE7eSnbY21IyoFL4AwE9vJAKgP/cctfmW5tsHB4Xklk
me9YScxmY22FhKtJ/jWrN4S7xUQivMAc8uEmzEoksDt4PwyZwh+7ChvyetOqBBP2
WaDHsC6TBo1BbG1nb1RrajBiG0hLniLy57lcgJbwkG2aE2LWlKI0yTbw3EYi+2ni
KmD+CSjKKSuRRrxKmzQuql8xamI7L0XMiqA8HG8zL8Waeq3TQns/TB3cEIj181LP
dJiu6//OIiYUnIv4XCT8QGjZusn4vdTV2pg1qwoIqIpvNm0YER+6XXQAafroY9Zx
CiGzW2LE9ogOi2ZOALhZShT6IafVim+3UlN0lzT3fMpzEiP0LGIvxcQ7jdd4HwO4
7P7c7XU2VSzjHiXjqwAIXD15te8S24ArJaKUl4fcX/oELrwPNTMCXSPY8t1ipzT1
pdR4fxPyRs6hSpsOx6wDjK5R4X9r8zimElve7v4v7dJ45D8zXj8LrHkzm8NLu1Aw
j2zyZAGtPg925oiPsLaMP7MabpNDGxUbkFYGn8tvzZ8RiBC/77kqJ4FWu1vjtADu
MnNoZwdJOyn6fOW1c6qjPQz2tIUJG3gQl214+MHki1OtNVt9XE/yHgsk2tyfG6Tb
PWnTS9mUtnKcBKkwso0l5z5oQYmhPTu7nm8+T8J4rGQ16y/s+e0p+qvWx3OFHa/x
ldw1s4mcuRQx6k/S9fnR3lIRVIHs482e4FvnbC1rxgYk+N3HBPBWF7iQcq30PDZb
5cOlJLWuWt2kvE0A+0vqXUUjXN77+qBeSneJfSPjOHFRXd0aFFPoU8aKwKkrPt8l
aq+6VPI95bQZhZJS+9aLqYRmjEfyxVdpN5LpqlOZA+FjOJ/P80JeKucudKKhcxU2
UZFAo7/ByjubmGlHLTJlExltGv5kllZoKhG50bW/5Nl9mzCC/9eKDmcAXj5++wgm
ZH98Xee1OP85XKBM7BYyB5ouTXQFGfG2QN/LfxBPbQL0BwTXoA4HYU6Plh0eVMXX
XyW7q95OKjt/UEO8wB7k4t0XUNlw38rw33HcISNFdJpw20d2xhIAEBRx4GnwQHok
ROPa/IaP3MEKj9icQwuhOpjfC40RlzKTii+KJsD/R63G5YO0QBtEL8QW9gp+1PmJ
eHPZ0xHQxRDnqvWk/E3296OnjcTfndDDO9upjDo9vraaBkg3+KjVyRP8pbI2pmS0
QU6IlqRDwFHS218TUC6It0XeS5zY4fZA7kIsgDhyJg/s5wLMXEhfXVlzsljGT3xF
Q61N+FJfE2nHp2mOP35AydcS3zPoG7qEuTBNgTOfGbiNeNELw3CYY2JCIyQLr9PM
aM2X+l0vcece45P4aXGIxm6hczWgOcC3ewZINj/mUma3dOffPylXPDU4Ls8lRLGQ
P5ebdheX59ey/B/CTNW41/Y6WgX425iuKgBUrCGsL1Ok7zUvGcgllSvmpW8dcy91
x25n0l8VYITey0rrL5vk/O+riRoY/kElr0Ktv49LrV6pK08mNPfUXxm9gqUUqyOe
XIe+vD8Pbs+HeA5GgW/7XSLriY4J0+WX/LGyBfL+aMI8xO8PANGo4c/YAfbjqjWH
N0I+z+jaerpc7gwkdD2w3Qmd0Q8Vnos+E7tp7BvXyymFLeoK+za7NCU2gnevm/ZX
HwN8mnCdja3puzgUhw/cyPJRrmApGYLti4mwTtU1NpqReKYja5iVNC8AL8TUW6/u
hPy4kZvkix2sigZSQJdZkbeAe8sOkxMuowoXz2vH4bOeVdYMTbFoK6odRrZn7y4I
bHJcb905aOkoqz8ccCG50ewUg/+a6AH8bt/MpusG8BIIyTYVKfCxtgVQ2YgAHFw5
bmjIGSqsitlN6JSFCufrqNh++L6CmgjI2TLneNghtMmE904udWYY952cYGxP4Eez
MEAuTN2LZBBtuqtEY86EMoNhh5CYH5QQFwP6xQpSDQbG4NKu2IvQbumNHR7+9dcA
pvlrKlajArop41U3ycp3/XfzUMxIRJs5WK1OmwE2FTFuaJuh//h950m6i1E84907
oCnd++8Ej6sSKTY1qypL+iU/zqPKFCft5PcyWMlntRcA8u0/fGvVV1eRCpLi7mDQ
I/OacF1oGjO7c5G2Dry30+VRdmlrssudEX4Mw8ZixP0i7OnbzPaLE/vY+1wtQoXP
TgEcVBKLkfRInup8gDfXbvHb8MlbtTLmLFOLet4Lq8W6f3k3uOWeDowKBQX4WnyN
sJ5g4+kERkcH4dem6q/dHpLRAsqfd3+wOKX4MZgrJi+u2PZq8+86aDlh8PdRCy0N
V2tP6CfR1bbYT9uRfjqLF92g45PYXvnypmHB5rHUU0Ecz1PRGdTDC5oiCMYNTfEJ
xNi+tjJrOvxuvA11cfkd6U43mA7+4Mzhr+lw2TkuYIawjvLAOzp+yRUf16PsrsYA
PnfXeGuha2LvWKyqGb5MAAncArJTAiCNxWGpyOOHQT1D9ISt+CIlgqJ3SS5jaT3E
aQ21o1P9oLV5GpkScyBYlw==
`protect END_PROTECTED
