`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GwH3/Tfq4WAVPVPwqhJPT7881/OUMBQLj5WLXKnxcyzhpZdmNMbyQj9Lam4pvMAW
hneV5Co+gxJHkR8oTTJiJLy5T1tPBZSsV+0nuQ7ko+C8+QT6sZO7CxBd3YW94oVK
Nmd46mcxFehLvjoCMoea7k1Jy9Lmhn2x3d2Q40tQ9uAlN+riOs7U+ttiIqNgz3r4
nOU/7wIi8YkFqoJ49bRNYQFURNL1/am7FbGbnjoWpUPZH75tzzAimovEKwqsd6Cz
JXNMiGbeKScuiv3bhMXl9f6e7bala6SaNm4wZ1WgKNFMPbjTxC1tPFTqDIONo81t
A+OMVv7X+5uUbT/K9TMvn6Gp0x7HAWhhVcGpBznatpGCK96d0vabHHY1Ia7iPqIo
Pd455zdc9j/w2XvK57jmNJnipZweeil2M0LiC1sjOQhr+b2zF+VqCd07u6Idd855
sk2ALM8x8CDP8xQ2LaCKaQXBTW+MtUqrYSNMSmFmN9O9OfkSk3tp3+F3X4FtTfIq
c1azaB8k0aXGwoozV5xhFNSa916MZGzDe0geQxURovHkl15DiqACrK0X+9NsLgIS
qLYQNX1KnTobrhXGRJk49GGR7O+Of7xm9KmpuW6VkO675PQKVREOXp6vA9wvD0PJ
buTD3E/3gV3hiBDfwsp5lVAwDJB9MUrL9aOD/4Ykn6dskO2hXMrWLOF7CXgSbqEI
wqYDC0iLzts1thXhb/4IDTs9i/MMq2g4x+rNI7Pl7N86Vgjp61/WOWSM3X4P2a0W
CCrqtiSZgrmbt8Gizld7kMF1g/F2xwIeIV2VkjSQk8L0bB0mOte+kLKDnrQYz77y
eY0c6cm3fptZx42CdL3XaeAM1px453+vgy3T/fr3l0S8tu34T5gGrO7CUGINoAsD
/VoImAfk/DJDc14TR2XtNFxphqm1t+dzzNNS/KEeuxFiLakbxG2B7EljAprJgo2u
rcaKMFhfkJoE6ApXOfaQMDPZzQ+kGJi2K2KLkHUIsN2gQ2mcSHN5ed+sWDzb8uSw
9C0NOhamaEhxmqTL8FiQC6DBDxuUA0BdETn/Q451YQCPll8s8wzJgy3wh/Ym12KR
/AAjMz45TKifiFVUxmKWzoVDJFr8HNnkgVVo5uoPOQkQhQGXce49Eg9KHW/BOn8t
m93ALCEt2XMNEyF3yg+60BGH05IZ3mjMVAeLy6UCVJvjeZGXqUy6vknOGMUMP9MD
qPG4quB0cyoRXPWVDPs64JEZq7hI7KJ9nCTQx091jGqsiC6DMfzAfkzxZONcsTJY
qWfS0XeH871RqAHlFdc6WZe4TFs1ZDKZcr3r1hNXflzCYptyUHVZutUkOXL1hUaL
sItk8ffH7F3lgeKab7OM2r0tlzGNltXWuKIQ39+hGwcthgCzad/Y7AwlpJhBdv/A
G09+5FvRUcu1fPNVrwIS2ibw7jJJoC0IYWR0JxnFRdH1LNhjJHQICbXYuxLBM7Z6
kucAItW1uYOmYkkbTKhXLtlB1hzJ5tDjA7GGcnU1MIkzy3BgmZsgxPhjAeNrQDNX
DvICzEGpXiFWt5wePeg7ogele02I1K9GY4LJn0vTynDpikbo3P1h10GaYlDXqIU2
SrK7cLOE2NHcaviGnZeUN72BpiLuwlOr0bsbWVAQ6UuKVOaaoAXDPbx1utqnpkku
XP0KIA1dDk5Zh4trdUlnNn9DkeiP6fEKHJZ1hxS4u/m65/3wN+023Dqg2K1Lge2F
3INaG3rfqiOAjfokS0FAKmmcvsmrAua/a73gBJYKzzMFh7NxpeBKq8sh6iLPWI3p
P2Hvl83kjHsFybgCIo/YJzM9jTotUCgi/5W+bMSMe2npWWaw6NUP+n7RNYBhbVCd
1EMLh8zctM0inltszhhd21D2aUqnzDlMIDEI+4IrNkHGHKsIeRPqme7xcBxiH1UK
nAB0aN3zUhAw9HIi9G63PSpg00pJvKd3FgZX8HlmXbzgz8JaUlHKSSvPBsd3adTv
ZEEK8eUrOHQWN3bv0ePuwSmQZkuUPQWv6Qxx20PYbLxPjzFlNRws9was2xWDMI1d
qeebj/fth7VwU/CvLMr1YQeG9dqwGBMZh+5Aw+F7L86tl91r5wm3uVhBn6KNKIMI
RvEZ4ireNz3ldZ1MAtyF97SVyJjPA+I4TsnX5taB+3JjNhh/s6xPV1pGz8UqQS8P
lxmNMOaSSz8SbaEG54IewdFp4sUzwdKsBH3nsn05mJz3PWwGwiciYQBxHyhqCcmB
zXTBnkluoKFYd4G6tXsCscdHyDVQSpcPfKyenfrc+04rHJKeBVd/TYNEcOvGZ/dy
JgEEmhs2VrHr3dnZpAkKzutOL6lcD/uCO1AcTgm/RmE9gP/w9XxDatwcbnbI3buX
YWYafhdv9eHZ8bcy9Yx663q43wYx6rvjPXXHcIpEU/JYUs6ZBTnOSJ4SBaKZBisT
G84J28J0dHa3673BD/u6STDvsksVGP+ZfoIiVKdjmJAALzaBV0SBXEHwzIj4CIHO
TaGmO0h8HzTj9sO214rYbGsebBcweYQ0SG3s3AtPGyZk8mKwhczU5rYjwGik8AkR
gT9scNCHuDNnujOQgoDnIod9uglFn1iWp9SN38vt6AZTSqbhkHZC7yJWY9fsoJyX
7DyNasZMAx4AvLw31f9KD782cVMH2YcPrBOCYCBAs9M2SwufumSSnnfuLhU/o9Om
97zsqO5iYbuCELoggzHBNz2Ck6G1BeOchm2bvcex8ofVEtOsQXfJ3qfE0Z7Pd87j
ctZqmysbM0yd8kUb4w8eTHIaQHG2KDHqWVdmzBA769X9dkCEznSh9GSlTzT8Dx88
9rJnCumPPQc11y2ZNQrXC0rW5WfY4pOqhnsTR85zUTTKkNhIUBdVN1b5a4ELLtsN
DInOzkEtFbLu0a9clfsyajUjqoOjlX9ES9QIupP6J+IsLVXpToOB+Wf8MN7oqwMf
89UfvRP2XJmKVIu+vzEaf5m+imNV0uNGOOnCoOKKrvG9vp2kHEOFTwHvABYhJQg1
TwOEqBNuOZmx3JgARokm7aHRXBby9BBHvzFZ4oA1DmivqSnLpdQIUZg20duSC5l6
HfDTV4dAtN1jn4I7b1F1GsIty0ldS+g/inCX6RaqN2Jn2/tE4PFgxEmHMdvYeskN
jvB9xllpHatuQ5M0Y3UsQHONb5B8W2/b47hTDxCY9Ji7pN8QbLbLVWdEr+GA/19X
BDc9IzqVyM+rgQjk2NyG1UlO/w/m/z+uhvlVFBPpUieOqVINdvIzgmj+LJe6yFwG
cDfJP9E6ITazTdwaJ0R2LEwGA8OwHB/9/vvwNzD+XLMakQonTw+t5LdpR5viDIVn
8QrmhREi14focin+qyvQjQORRTMuvzwSYUQ/0yKl/CW6JTPBeCGOw843A3hYVIBu
o+IdUp9DB32J2aS91ptplUFsLxMNV8YXytt3W4uNsG8Wi1FiecJTKeC/bmwj8J9h
48KfnkMUTqzs10b/Pwzk/ZYtrMjIpeDSoL0ZW/7x3SYc3YNYu4SNHEBcnf03vjt8
pA2O8qiprmMEi2uiDSXdmDHkh7spRbrO4QxavtodpT9hyJOsunVP6gqJokMnQCjg
i7JYEa8hLW5aIdAPgPZZDC10jKxa0Ek0oIaOIxw+8BDGwC52GzUDj+Vf8IS3eS9N
0o9dcb0VlEBdbijpT27Yg+I1LOiAeD5J+UxBzfeR+somQU5/7x7r2P9FJpSxhH6n
T9Ye+udiWxsT6qH8lV5OhUBIUgPbksf9I0fAE08lix4uZTCyIKvuM6rVkA6wehzg
SaRoOPErGoicJBeeKtRKFLfMWsuLgfZ+DZqs9V/73zfMSdOGcmm/MUkgQMUQ4nFL
m0kLWK+RDQ/iI2Io900USgD3QR5hzkaIhYlLmYunZEjQH88jN7o893ehC5h+546P
8BemV9u3FKS2tgF+ODj8D0VFHA+drYcHuPLyOuwuvugMIQzu342fkhjW4h1Y1O7J
h10/btQTC+J6jd3P5Sdvug==
`protect END_PROTECTED
