`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
btXd3x3jJ0zG6hpwXXOAIYNbriw34FTNz30SKnpBwrKH6aTbA/PfbX3Dxqyu/URj
sP4WUzJlh1gKfghx4n8KB35Wo2dooL+YUt6ILe2mIcbsRaOod4cMdmvGWo8R4Caa
wzfnuJDI1UrlGgxcpbP6RML7YgcyvgiQX78R5LZ0ode4IWBltcEaY6oHRLAEtpWG
PeRcbl397ipK707W4bi79+6YLeZW9FhhvKTGAOwq2fWbaBxFtiRi0w5pgK3mi3NG
1EH5IuEC2WtzVL95oSkxVDhnF2Xa77BONvvZFBTlkG0w7uIs3yo2wvhg60XeWibx
7JJADGyeltdKhZDc9UOSsteNlLsWyjAu2uZam1pQj0qJ6crAWD6gBuvHzF0wcEwB
en11pSocMXmPm1bZwLlz2QfFVNiagDI79Y5df/8GVgE8TGhdezM9iLEfrHMbXvww
Sqcag3C2SpYjwqmIxJ2MSFyJQ4Yf2Sa3e7Sah5Atc3WwocvdlHhWNu45Hc7XibZe
XzixbjmIL4comzMvkGUCCjqU5fbOsS96KJ5ghDVOPaZ5H+S3OuAxXMxOLSelIFba
WXWF2FiSkzOrnD7cibBkJnm2apcwowr1mh7QEX/2jTlRoi7OQeW1+RG5JgKkPZru
5KuY3K6Tg+MhzHKwRpJY3jtF5oEy+N5Z4dMu/gDKlykwrJLRFERdEM5eEG2ibKgP
Xl6HbOz7nNMOkHHVcTQ+EyUTDbruv+Zj51fgjwndmheySiz5LCoZDGiGWMhfmdRN
D4I3dNgJF+wf4Rli0cinl15vENsN6ToT8YI9rzTISShM6rqFtjJ9xx/QvOtoe2Y+
ug9448Xi+uziiWf+w4xiM0k92S7mJrTs7BGuuN0ixIH9dzeUAwaQW896orspZkYx
gXcohS/J1KFXCtXhmI1nCuPv4dS4j56ZmUfPuvRrsoMfSEOjB6vJ7KovruAuO/s7
`protect END_PROTECTED
