`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LhX4N6aSJkMw+GVVB3Xz2flW6sKTM5zLxSg6c4C3v1weJ43ntybJTz+vxuTWhBk1
hTvf9BilcqwGEmLCnXCDUzINKBRIjzcKoY6tfhaedF291W/IICkUaNAZinsVXxi+
n8L87+HOG+ToeFsLX6s+q1CGzTePC3Cs1evNdH+fpM/ziR1qfo5ysfHWPhUUqsoO
HNTb1vkPEMu6o9QjNtajTrInKQ4XvXCZKHcFikQvOD6Dvm9QE34FF4TmFYenkImr
WfJ2a7/zllujsuquN7gWQDXtbbd4Dd35tfyN+CMR/QtbZcXP3ewYNYb7dBNTyylc
26kV5XQuC4lPMJomG1LJk/Q18m00jh2lsL2kkVEPCMHqmOzaYia+q0zc12vMjS/u
UDjYGpxXMNvb0nqfCq65ab2nBC2d4uW6G841l/Hk3KyyrwnAqyMyvjDWg/bdedCT
+g1jmYmu/4EpWnZ8vp6gT3nrsi2X97rz+G4V29bGzD41dRWVFsYWstQX3sGdVZ0P
9z8pirfayYFPn/ApaerH/pLJ7vcJrOIMHJGZB9sVtz7UsybdsQKdB+ITNv4cyaqT
MyuDWlOabtck+oA6/NZw9dBwMKogxGDkvdVIZyWEmm0vG0svcaInpEy4xavqj83U
sOHacpuPbTLIiS7feQYiYxUnLsxVrcXqlnsWnDExJkM0hZIZtzQ0xJZ13mWa0JTd
NVmRoZCWAVH7BYwACi2NWeOGquT8KQ2TIHUnE93NGw7nySi2Z+LYKRJY8YmY0eWP
bcYbGdh/RnbBGE4zzZiUIgVOWZg5V5iTid1DhahBjHAEMAu8gEslKkWht4mqeRzS
RSvsiUMq9929e7sIjznHitf5InRh3/kvkx0gO7w6bXtVmAV+yu+iBIyK0bDyVL/y
H2cOn9fUUf6cbSuUz4vOsKWcghf00oqlSG361yOIl+pzjKjkE3PzMVcVs7G3J9Cn
tQVEv0Y2cp4ahuKPCJO7QhOhpMl4TWMchZ8d18ruSOMplh4UqSt21ubnI+l/7397
6uxXbZxX0td4KBZ1UpYIOaHYMJHtUiWzHPR+YMF5qvlq/anyeY4ODjc8YdtJN55B
6wk4cCkXhRdACom7nu6Lt5fihTAhVts6hNgNa+KRfWtliB/75W5DjCivNCCTWfdu
htV6VB4kVsZl3e3hcvD9PGN9hvux/EJP6S7D3bUqIp5XtttxDrO0207IaUTTsML+
K324QEF1td51Yqh8zEtWyQ+6TSxYCsfpwkcFu4RgZ5+WGoFxI+L+5GszkAjciB8B
MzcL7GER2AeA+9/gTD9gwFkvol0fTMek72Oa5AtVDkv9XfuHZ+m8+971wXcsc98y
/3BgZ1yzlAySzVIb4eSDcvg/RgnRHD1GWNwHIdbnxWL6RwUEYdVKz9Nh7m6PaC8M
ed8YGgn3kJmSt90yAdbVmwhqhY1LB4R8qc4RBq3XlvXfthiuO4TquH/+ms1VsReL
J+QfyLsJ29DUB66cRKGXO5v9kYf0ZOiYPIL/KFx0Sp+her3h1BYRt2YWNKONHu70
JP84CpgEE6RjrKOPBXtXOvbMJVUwA71ruNzXLjEQCwxxuNcpK97QN1r3Nr1oaFue
NflSSy96hVzFOurf7aLnJQtWYZP6crau5UOrEjRQCeIZCPzpD+6YLLm0AxZd2epF
f+LZ/OHOJXxuZQnKGhUriBa58+WM+bsAIC1/B+Nbb8sQ3q8IXHhyQcUnZVs9DVJd
oEBDWSQ8EwYB3t3/sZMYBkjduNz7oXwdZdMX3gtzG/hwgIpFJlkpYzMaySPGS+uD
DEkunPaOAj36hNhVqEZYghdl0+zFj0JKW1OoJfjPtGAvx/ux/BYYqAau2a7PAcdX
N99k00L2clx5VmLpwxyH2U/Qz60mEXkcA0+2UdfCe/funeAfqhkbkX2YXj5BJEyM
W4bXSCdPReOp/ElVvFIfFcfPDOUyghf26jL7sgPtiVw3UX5waD/whppw4T81GB3O
84lh1RSL+34Y5HmSuu9gbHTNAd55Q94VOCgoNPLVM0GlFwqPub1l+21bQqh6PjQO
8mkzzUNm3a+snyagtRoX7/jXmancTSZ2488oqBFQDUCRH1MU13WhS9c4gfU95BHH
qBMBcvQtcHIchAGe5fR/Wp313T5jrl36zaf+kBrpgdfPDDzv9mtsL0RLDQq0slwl
B7RodQDyVeRTzOK2NAHa0xvlXGy++qqZtMzKz1xlcJi2uM124A2JIqO54ccBdFH7
NyM9+Axx3zr1fRUJrbq2LdDI7Wv1TNLBHozquLElQ3xARi3LEWokLxE579CHizoO
hzQimbAR9qtHUxYs742h0uQ9KNAAD0pT5Mqr2NqGOaUgkS/ZciLMdN58MFEMDfyo
dCLMS9Qw4MwZA8pvbJlLBAdMvxA+GDfgpwzl3CGa7HH59C16jaiu/MmzFJ9kab76
K/QUSNWjtjlEtW6noDLplUt0MWNZtp3i0R0hIgOM8rVJJ3wh2VC3p5+yvfCnDvhs
5sLEC0loL1xQogCCVaEerU3o9IgJYsuZC8eOkiZgJVXc+stnlcgtZ9he71aNR9uz
eUu7vU51nnY1TZM3fdKGqgF5KqRq6lmZSBk8giES1kq3ib7xegL3BE8vndjxjcj2
xPfu7N5/iQDp7oHmvsw/m4x00IcxmPyry4fLE7MVWtqvTtkjn/HuC1jeVqZ3yajs
pdia5ZsP/pcKpAcCuSUcMr83JmASfJImfA/zmPdIky0R7pmNGZZ9eJScJPRjkPte
jedOFqeRZ3mSeLDlltKUo6eBeoi1LX0kAtLcF9OliwCzs2jDvzhXkg+654uEWhAX
yLeWBI5MHYjjQ/PSpLZAfHc9lPhnWoiVfhWMfO3BAQWHozX58nmefxiDC8vv8Nis
eD7BEsa9rs4H5yRs9ux1z56LJ479wQ/Au/E21yFN6sUdyYYv8ggDah0g3KSCF5td
vK8rkIS5qeL3O1Myxqus5w+CbuDpbBTXvPG8ujtqEPshQwGl6M5+A+Y3CBH4UNow
QcLFBJPDu5YNVkJTp0WVN3PMe1+TsNQ1uEgF1ID5LA4htzCxIGqXynsQ8XXJ+yAY
twZHQFJn5nJYFOHI8KfVIYZFPDnVl4SHEJNLrTYouB9EHcZB88W7CfULU/M4HULv
gHTtJaYKdxZUqcEW3Eiq9D3chCo0ag+xpM6UN3Zty6gjYuPXELgHOIh7jTtfovWS
bs1fuQoqflMJ1g/5hPpUOpE4eUrP1wfXTJVJhFfGlAvAEJN0UQeaN/JWBizZeeda
fbPvQ+UJOPVYiQ9w+eI5SybwtekmyOsOrkDLyEE6I+OoUsw1jFx85mX9Z/RmYt4k
xIG6VKNvIxfbQD4Yku93d2gQL4zBHRgz7PcxPXJ7iaP1x0/RzFv9KiEM+eU5NgEC
axuT0AuACpYw8SbtJdWRS6DRNeNNtLGIgGYfdaf/gXCPs2FY6Q8DdSiMAVhyeO7C
Wfmf//PtU8FxGqMmYLizwPygAxewvldWfoni3r0C1Phi8+MSBepk8GV5YUoTEY+0
tW3L06cp15AYjKjoSbQV3XOB9ivwSujGZfWnHGMDptVy9i1qxleeErOr5kVnq1rz
cgvQfXw1fJrqmvhvDiLEytDLFPsRNA6O7uQF3EePLmuL/ztko/MQCCx+K0J1eeHF
X5OsVTx+nVaQGEgQK8hLNGMz3CF6ND4sp75uTsljhMTCN2VznpEp9H+ml4BQRfiG
OIgAuLb15Y+FA4gzG9LDBfYYoO+ybQCgQ9itgYIMvYgmUmSkg70J8aMPIV/Xc3ZF
vP+V5gSG+FcWye0tSKujPDUuOUdFXP6TrwS1NFoGSNa76A3qwSznGGklVYOno8zz
`protect END_PROTECTED
