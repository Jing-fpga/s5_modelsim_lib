`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8noHhCrP1DA8RD8mS127AfAZQxr8DVukFk21KX0+gp5tAkvzdMRMq60HoQVjRH+E
4qisFPPAnlIwL6yc6ji3i402sMdoj+aub1nRBGXORBRtr9pHUM0FHDAiMEhndqyF
YZnL6o2v41VeyuKuuIl2tSm/XZzTlmumBXjZgRgBmysjdYHOCnKyhfA/ZOQo+CEL
Wjo32mEayQZdyh/Jk4R5GSRwwNIcQaNxGVWaPxbXgAh8SeSFa09MHS2NhPGPkjbI
5EDup1gr4F/MYxaK/gItiFtVAUFVfxQbhn6vrq6EWB4yvKCUVMyKPNjfV94b/jfp
SpkTRLgHE6hepvPDo7s5EqmhfMoBWz7OaHj3ZxH2KTVraqI+r1+1arjqWI7PTbc8
3WLjED1DQ+i4K7vQiOU9ATvdMF+FCx/b2FaceNInpwhmxQ7IJXQ2YFt9FXs6LD4H
Blo3hyxvJYEb5x747jAWl1FKs5nvasow3WCT5ToKF0D5KdisX8lvIO7UD2rWxwgF
DBzeaX3XiwR4G2lRaSSs9yISCTvPnEbIosiExGv9qu9s502QJMuCnXXkKYoxMI+1
qyKgl1oKFbIiUxIwh2EZo9VBYCl2CXKi+1OrYizQIeKyea9LAnOL2GhVoTCefFis
aX/MbaH8ZPUvGpSupz9wvjhgqr7jMADgtclxhbN0u1uTDJT0b4gay0iN+m/8zpTA
EyTi9EcPA5qd12moFv3pTVLLSliFIWFLEmiqq5zjCfkBssMTIZRySA1vzf7iGG/f
xYW/Mm7UhhIzQWy7evTHEH4+tZ3V3L8FL7yybqOcuBWk24a1GLtkm8HTTFOhMzu3
JTYTLEEQu6o1hGu6Tcrqpw18npFEpXG9A4Fm0Kjc0xlAWQ0TpcIz7tPgn8g7Pl2G
M8vXIeOcgpUIPuBDlNDJcdmFEzwm/zQ+4OXLoV/a/EDtcjmxO4Lu2FO7qAQk/M0R
Vbinp4XpPztnYF0zz26lHaMOk62IRAjP9AAVEgAXgfxXRHwZ/P57HWT+EoNPfqwu
2T+ZCvbBzmfzYMTXhnnuAoK33SLtJHHM6XQr/YeIe/LE0aMBk6KeClHD4NKu4Dmu
3GSLjAmQAfnq8BhFizqr97zRfkhAcenSukcDija14uOGTcmN/czWEevODwrWtczT
geH6ZGG6iBihJqbET4J4ZQ+WV1CYSm+Pgh5YHeuT/kiQ1EZNSOYndTU/fEDQIeFv
f8eO0HnuuF06aP7avMCDP909dZS1JNhNhej8ngNXIPNZet5k9EL82gjXJU8etNy1
Ghuc/O15xpyzdzMJvtWm67u77OosGk4wBrNxCQErLLCp7Ji/KbRqkejVlpBG0W9Q
nGnk+aAPauuz/PGPOSnZ1T8E3FAQzMq0G2dmc2Trf72fKwgGJ87hs34E0SO5R/qV
PCqs9ryvlsDyW5V3z+fHzAf8vnE1e9xjGj7UlaliSS8UxylfP7SGC46Bo3/ZwX5u
Uy2/Ob4IjdM3NcVviaJmwduXBrdv0z+UWNJgoDlvd7N37eXkpdWv10ux+OE+MBkf
TfaixOHMDmlc+Ot1frkWriKykiQ8WuIP5sIwdmiFSBpKLIcJOuJO4wtuAaBFcnxb
dZY/FmCMTQPZHz76axyuqDtPK+i1hoC7BGrdXa0qyyNXwIYnm4Case5LMYTyM95E
5zTPMFCehFGcNp+0c1gBbXWUYLG3PwIhm5s3JtTlOf8GhZTjMMyNYZ++yWn4CtOP
oqCEA33blqw0pPtullfrq1rY0zRpFVfzg+FjGQwNm9vYq+napGA7Sa7SeNWlAkzx
eh6yBFmfP39hZkGdl8+vrD9hix/4ieKBtptGpCFHXtYpytFNAKjJczMZjsjTddDe
oXnhEQYuhB8m3cy3L7SVn5DwDV0XkwTVSHkrGUWUplNYOBGSB2pXPorX1YPyzyJ0
o2mqpbrmxgOtjxDAdM2iBPtpTEZioVhJkTJEkFwWFMDgBbEAtyMZ03hy15aPPSq3
OkWljIcRWycYKxzDdWiwookFcpQK0Jvg+kzZZOLoNLkGWYoFQXe3g9a7sOLh9AGY
`protect END_PROTECTED
