`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0JWofT0jpHY5f4B4xuAcrGtFgFaRmamdcGt299MCIEgdPud9mGismLTzwNIbTjsm
4Y7UqU+l0UM2Oa3sRd1E1wWmZubT7CFDRSI0VXzE4eJGjsW6ucd4PAenFzR2uIuD
23ktDxqmCS5xflMgw2mtZat7T3dsJOHiiOGP+AUNH3ajWfEThCA3S5lB3TReyaQm
eOcg4mzwSQgNBPFNVR7mU3i4MO2nzxLjuV7578LSAMKYGm3zV5ouEi+Mvq+leA/J
WSNU9lVR4CTcgH1G2rLWtNGxsOdMcUO22h0g1/fBgdo42Pvf3A1G7mdfm6cCEhl6
dI3kDOHUHThFiH+Ijd7R85c+6B28/TAj4DEskc4xLNRe9WknTRQnuJTOF2qmg0X+
gmzV4M/a0+lPg8AqcAB26MAwjC4TnLaWGG3FhDW/SLrtgcnUlTUFHot1xZQXcF0z
8S9DQDo0zERwiutkKmsGXpzMfgPkodfXWT1TQ6ceP7O6MvWtRYjdGy/Ryc2gcIOL
6ldFdbwIc7s7wAeXHObP5YfBUuJ72TKN4p3S66eYixk6R3ENsx857u3gvl9nxsWg
EyTH1HuiQ2uUg4JiPqyggqxlJmLqbOveKUIUeh7zBqhP7aTU5GlirDxSKdPa1b90
DmA8jcXh2PCNsfjEr7VFu9rZDroMVKYWlMhx4KM6C0bj/nurEJOtSIUSCYUnRCj3
+BZ9azmFB01oaLQYYDon27qzYirCn5GOij4aCF7M+2o=
`protect END_PROTECTED
