`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yc7uLpANz8fsUhQB5bdooALCj8TmycG8nPPV84+MTNRNrueHYRIfNIPO/FaaDXdg
jMQZ99bCjrNV6oR6Y1z0AbPIlw7Vs4MQLSZXUI7o87okB0OiDxX7Ytx3eeJtA39s
1LrWBrS2gsExxQQi3sygNoxdbftPpDTIp7j9yMVVCcvFEfMEeF9vXqKPkbeWeK6r
CVc9jb+q/uzqnWlZaM7oqWhIAlj45OkwtAJRIT9j0BtRsL8E1cgOtyGEvw1K1CT4
kbbduVmgNUPrHTylzq9jzLD0kXiyR/8m7QZR9d+VauZJxbhhRkJhVjeZ3jHlx0Vd
zQs1n/vef9mxUE/rLsxfvSUCDzGWPHQFJgwr//x8vaCRYdzKwHesyOpbuBnjxOEP
ngBINjlYZiHhSJSwkX2xoMtMq9MQ8PqfkkKMgIr/NfE96hkp8Pp+wvTnMGYwgA5B
pvnYU1vSp2SqrvfufRc0PL65bd+sh87L2M+y12+mAKi53GPb0+cyvwYn6yM719cu
2snMzNAmq/ZpFGJQrD/jtMhkvVKIjbCTpJ3WUt5jKnRNo4wFkXSGURqJbP+578tp
SMirUv6y3sCyOOVl+vi86CEfux94tVXGEdSJSGJMn6SkkcSREvnWSTF5cnNGDkkP
VNOXmYxVwoqhpaKujB6TN+z2o0wEHoYt+SeN/5/mETp5ysCBlKr/yTgFJDmyF767
Cmui1q1ZXDTzE0XzvvaMGjBTf/wXUoxD9Z0sakR8tdxo3KPKEa/ZNATwSQdRMKh6
CtcoKpTItwPiDjrrgX2sdcg+MK6VFBiR71NKGJCpeQzvc0eg2RaoE4T8bhfQZJ3y
Ul4H4gDNx6QCdpIX06kBi1zn5TwNxJCVF9Sow/+3Kw0IevAzlrfIiPUs2M5UmOb5
9LDfkJYpTqa3nG7Ah2cePGFH0lrsLyvaLbtqGuQgJYCqq/60RBlV957mUkB+26ks
TVcSGOwTSmoZcIVRm0ei4IRVFHs1uEP8YiCcueZ0KsliXgOX17j0uo8pcQTqAkhU
473ogven/bF6b5yOzpICbFHGF9k9duHQvBjBAQb0P+g96/CMaaUGHJg0e63KrvD4
5KwJV2OTNTGQ4bsi6iXlUxRyITC0r+6g2ZCPsWLyOeCEpGtgGIOeiK+85FuRiToV
KSa1/hnZyc3RB+lLFWTpbTHszwmuld/GIM44jjbMKc77Zn/itKa0NVykxFXaZLb2
8MpftIoPZRUEIISosRR+nfDsmTdCks26XyXRSSKYzmP/PbIYJcUwcCbORTKjT/Iz
NRMdFF8WpdY1aMjxUjqCtlHZ2Ku3anq9N2jSr0X9JRFSuJ6oupn75gX2omTiDAsk
c3Kec4rDXJ9SwePdiNdTzXq6mmDO7PaWUUFmt+/c8Tk=
`protect END_PROTECTED
