`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5tv0LeP+Kd/G92tScTGomq/K8y2O7DYr/FpvXm/RVXt/XN5gQCCW3cPdrJ3X5/8P
xpyttyLloMnogNqL0s+ZWvbDcm+tEy6+wChnWQMj0GQkZejGcqxup2IjBrGnLEpi
qmlq9vyMGfHJoZRBVd/2bdSas6rG/f2qrgvnGpLxCF5YywvUClVsYB+daoq4sA9V
cUTAgnkSeqg2yJgt+PxJPrdpPzxbDJJ1wZGg2LTnZvkbK8upFlRHbU/O+2mr3tjX
cITUtXglyeEU2VYO0zF7o7u0X3U2af0eNOsKAHp7HTAi+KqpyJQ0FZuDK4dWAbwF
2iMhEKTJiIJI267dBvSuWP65wxUWfwrtwlz2gWnLiO3LzKAJOhWi/pyounQ61Uka
Q+Es4r1W1ml47C+Lqa/PxEaapBzob7ZKeFP8tat8TBpfKEM8sxK18nKe++kdQz6l
LkUQL+7BNAsDwh2bCnDJZdBbHxZqmKlbGbYpclJ7NSSdwkrw6wx+D/Id9cDkM7pY
/ine8J1tt0aPq/wGs7L/7V8kmOfBGyIiZkCOoH/pCDtrMZ+n0tIQDF6IMUZ89lKU
jiUyIUYsQ4qfEnOVn9Bt2Q5wf+f3mrCOBdEMA4vMxllcFSf8QOEGQ7aCTxz37hpa
FyGA/9X+CQMr/Bw1U8Y2bIj2EdwTOfjABptDzOVgmW7xXH66P0jxViiovsBLAF5D
40miQQQm8A04l2GtvVn1AR1XMwxBWRCWlhbFss8ANeRgYk+mldKahwJf5CSrgVYt
VtoyivB1G0/PsvobInXEdIp0GCQIckla3pcfBnd95kxPXJHQMvnVAlJ/cvsGYFre
KLtfOnH8a18t7CFZ1HQYHXMbcsr9CEWBad4fGf6NtAU2gsRHt4QlFMUx+lmj83I3
USPVdV2onlAFnhyLZSDsMPhBis23g9LDeJmHaMxGNS4pkA5A2LuH6J4xspxL3X08
QgzKW31iJfCnktr83hHQAPnyzwLsOTZBXIXngD/hwkRYaxVCah6zAGUov5RnlOfy
9PZnhPePo5s1rf99e/EVUVDlrqdCXi6brSfv1OtsHzDPtZpCZuqnwbsRXbMdMauL
lNZTHWin61f1EHGkpAy21njSnpuZp0XLyX3mPYRomGrKwjLbYwhNQllOru3uv3b/
rweR2uVPZB3bNcQacogfez3xRuxJvMneRWluQc+BNKbAFffL5J71vKZz8MpJeY2/
n6JipWrVbkQC4h27sZLOChsRT6Ts7VBUzztbD2iW70miHBf0G0EXK4IwRvA1SZPt
i2y3d1pT7gTaMELliNRW2ZjdvNJkDBroLiJhP2UuRmoyaojTapnGpkyG+nTeHIIm
74c7I6SvFpHIBIh9hNcFFezSGg5yRmKSu0/NTd6YqwbipVrzTJPmECY1gwkCVRnw
FPRBkGxpyH1Dqo6oHiywGjlTm9rEC9X9cItRrsYFcmFPJF7ms9rR0FlqNTwZ4f2B
fx+qGaz6oNcmb0odRbKkJcUx+3GkcppYqFyUJwR8+YcmNwEU18hVKFyy8QUtVcU/
2WenwK0ov2JWvjU/2h7By6F5bHJdAK0sRyPfMpQWWO9NMF42I5WIXTeZKZd5xTV6
5dFtC5LDiEja9l8dzFTWdvrfoXIrxXPwfsiVyyD9TNw/SY0VLLsZCLGdwcUdi2OD
+snmGZzcvrZZWkVzpvhCDNnJ6OLKyLAL3txze+gx5Bfyca3aV6YgUfNVKieE9mNN
SG8BXNulVQgnM4DjcE7ioRHgaFCjPTNNaR18DTHM6Fgb3BuHVocWD6IvF50dA6Iy
lpHiFjgtkzymMvvBNsiA9Jy/l9EMrfpYo4WV6gkKiyfIiPR3u8lBHmVV5AY2GiJd
coT8sBs3eHs0TYzGoStawysvjOcXW6rMz3jfMEiNd2D13byCHQQbDBkadC7QzyVe
APXwddKn8Kw/3PlGpCVFSoChAebS5zslX7fveHRM0pJGHidIvS3gMp+cQry/4+Cv
bdznt5SbCg/o9Sxtbb01s05MF8Svv0ioXSRjeSj7JKDqfahnuyjpZ6fleBtWtXHY
0cBEbZihozrUONP5wIo+Pqw57wVhZ6Xpd+nW+l3Cso1vVZQp1mQ91Hhfb1ZFv6IO
i0Sl455i1wj13xLIQx7psS9z2zvDo20/mx8FzXPtQ6lljR7My2ZbbYqqrnTITbnR
mrlB6FuEuHJARYK4iQjHBqr4x0j8eucVJiYT1TT+hU6umbZqW58TrbVSjeZLF/vY
hdUPJOxgE5A+Rxm8v7BgOVITcgQoYhXjWOaeX9Pzr2rTRXnBp7WPG7EZ5T3Hbims
utFwvGN1UHlj4Bp1Nbyl9FqEB+PH+SPOZfanNeGPkLSqnSHFZl5LOVRyzcONOai7
24iKswGgZzsKRwBl1kK+yuJ0GaUr7FLMqr2J8J8iZFcs+R/lpftFtpCQhyrT42dQ
ZvYaAGmE7Fz9bru/srDOn23wxLm2nFdiAyAh4f7IgNjgWRM/aH5nRRoJknEKai0E
p/SUswJ9zfSYQe96AciGAtYU+oQS/pe/gaf/wMXKMSgIzxLPGupOVurAbMouW5Z6
Q5oD46cRdW75Wp+7pAsUHRWA3yIHTiajrkfzyInK1NfZ/Y6YipiC1Fs1GqiQET4R
ezQpBhgMzOo3LwvUyXA20pVOsxjEykRXvLjd7Bhf4cBhqWFQLsxrMmiV09dej0+A
8u0gI8n3SBhIEipWVjv6OiXUMNtcntV7HJdVpMvNzlCJo7zMR1eNloutcrk3N+Cw
yo6r35TcCtMrkMM2517M8O41di86E4KYYIaOf6kN0FTuMvUgso9Drl8J5dT6hjML
`protect END_PROTECTED
