`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CHgm0+K+aVrQb8nAy/RYWjzG5bJGEpM4+PVltTtBCS2qunWlrfZhC9AA8p15T0XY
bK5pM83zqfBHhNgvxm+/ns8oqh8L/fnB5Idg/MEIgix1Gkois0KGbb3+KCw4JG9t
LkS9pRiwIkuZ4Ibye8ebbeLX8Twu8l7lo4nH+BaSb/bV1V5z3C3NxTyQgwWallUn
vx9OgXVYsHwkhdZOLbeIKXF8wzZt2UekN7SGMFxZHq+hAYykivFAwm1XVxbZruOT
IBDO+Tj0vBnRYYN+w5x7xPih/i6uBX3Cmf8oLJKMnX1u1RS5YqMUZ2OENDpeM4n/
1BN0lyDFQar2m/yiMQ3950dE1/dsXRXu5s4oGYXRJjQkNbZLhn3jWyC111UZDqBD
gM6W3MoIZHGlDfmQAwVCaktCyXLdCVwlkIzE0o7rFosuvzTlNLKvWNdrVz0Fd4l2
xtnGHNnmZv0qdSgxvfO3odv6ync4ETGEPVU4D0+RWKDhGJnNUImdGNDjTHHbal7U
8zEmCj1AFLANP/HvCxda4uv0TOiBsz/cl+6R7kaXWDgaYAVdB0Bpqk9YMGKbqIaA
6PNl83ehvKr2ut6dZI6pBMO9zGXVtGzCRKhP9nLhh5nfRMM4HZyPL3lZWnglWAS1
nk+kTiocvyPq7UPqqlpngusgDmkkENeAuHETQA81GCmEh04SYOVm2v6L0OVQoQ+8
qr82LXaBhtHaIs62TgucLShA7tE5l8ZEfCs6DVeATwbhgxMivi9+2aUK3Fidc6uN
JeYLvYg+lHLSUBbF/vXt3iKLPtoPWiSU4Usm055q02DzYojNhI4fUIDt88Uo4QBh
WzlIJC3la2S96P0nAQ3/zavF9S1P4Q3wVwyfwazVn9/n0U5aRQkqgN9rc01t1njG
imFknA56s0lWfJ3NQoweuRiS29W/t1xbPix19Rerj1/wksuhdjdQTfsIEUCQ191u
yNHeXF0cqVTGeVxCgFMTe1O7miJveUGtCAfouHxcg1yTorCOAYVZd0lw2Zx+jWQF
7GQfCd6XtzZf85TlnYa8zTq4W4AKWRzYxpB+CvHfO8AvMCy4eUFuo/yZS/ibZ8lm
Toh2niSXiZPBaRU+Y5snX4M3iioGNJNSCzIzKrvMNq9ykGBDR5ZUtd7dr0b5vKps
4lj7pDBjEA5St+s157W5PAnQe/ITfNBL65peKEBUruWfucxTVG87xpnoCcpLgMVz
GY8Ml4n5rQ0loto71JSszYOcSz5jOelO6Y/TaRncTZic+ogIVAzcqZhvobIyJV/u
le5f/j1TZb8JUc4FYHdFC0Zdaz6aY4tIIcSjGER91aEmG0+MKC3mai0LBFQVNhrR
l5a/4+J/9aobaQGOdmB5zdi8wNcIKZsXmZxC2XUWWXcJSmt4DGF7sA7RQg+DQPOy
TCCBht4CXiY2vIX64f02Um/xBKolrT5XKk6ch6f4x3xNNWV9Pq5I58PcMaZRh+Ut
Ywh2Bhtc2HZZZezAv6oOZWBelVihoU8MGOMbQ1I1fJ9sITRVPriPzzsfWmr3XfCi
SgfN+N30AE1pyTyP+dF9LT9pvWMGqaz3k1XlxRfxMCcmpdrude7VIUDzeWmkR2yS
O9IGPhXoh9siEqVjjjjT/c5/rOFsVLT4rbmPAUaTA3t8gqOBK7mUR2AgmCOZBJwy
CHtmwxm8xkoH7kWfe2YNICBxpLP2XQokQlKe9Xl6dmnq48jtWEqYOiMMMnZ58kmX
owPqL4uG8CFQugx/YKkRICj4/o3a2IqF27d8jMLe1TGZBd8UgK3IcleCy3MOj8UX
a0m9Xfezm2Yh9+qdnZxkzSeeu8VixoxWYpOuKgMTjLTWyaDlxJFYoDSXo2YsqRnl
DHlU2z4vfSSVZYyvr9R6P4xT1rCTabU5lC4LmptvZ3ij19BnaHmjtZuzW3BdkIxD
f+CpbQ37gwtzdJnSWCnYZyYjZ3WblP7+7a8ZOCP0eHvN3ovgqG+LmwkvRgrx6KGa
LzvhI34frCXLjQk5IpIs+v47ndEX6WPAIDrdT3z2OmzzyUqRT7k+SyZ83eyY+WMa
UKZKKGJJowlbVnkODIBtk3q22vN6koqycMErQi7E4VKfujwEAZ8aIenXvc7m65hR
2Wf+FyPSL52Rjoi1k/hhUpeHPxEzraDHF773tGJEmhZY2DkpCSw3F2Yq6t3rEZC3
xwLN1+wg66ZLZb1lfWt2HOAU+/a885tP7pQj4NL40f8hR8PNstZGz3ANoXUIRkHX
R42j5fMucblSHbs+Uird5PlQZIcWdjrOinHck2nUt+4EJVeXpmA7j06X5RUtcfBw
s3mdeg0ihEEQKPHvkqzOgCeJ5bTtsNhx3RR0zIh0LGr2Ixfg0yborszLtzGW0bwl
0JIB228Xp6fy7ws0SwDB4YHmthPsQyS50gk1FQVDkXslZW1NZCJ1dQWhIVsBTCae
ojl+e3c3nfN8xuD9CYrXSGwR30i6gQC/iUwag7gKwQYQ7lBDSSuPwwPywXQCzYfh
jxqhUSgZI17P/r8oWu4K1BBY3Zg+Y+lC0eXk9y/VkC16n/i0bkbbPcpiFWGl7uWd
Oiivan1FwUJWI3WW7poHrjAnscjE2/Zo36IuUwn6cwdizwtQ05zD9rbZ9Ox9F/CC
OKqFsYTh66CdlCueWD9cz2rJMtr4jvqdIsPVROMeMkGO+9ILXQSEi8LKZL+cJXrs
PoOiu+yeQUKk692EmTTGwZ7jiySAWqHM8C5feAlg1QO4BvEt3e29AJox5Oq3syk4
OzFVcJEFC45rT1PYYa3MgIGGcER4dBpuf9Q7z1tlrUG9+jX0LGxL0ilC8XgWVKa+
HqAlxLFjN6f9AKESlQd0N6y1Zbf3LaPw5DgpL2/7/3/ajZq/T4QrRJv+WBNLKfr3
HLnxo70avUAOYYA0FdaDYqlOVYcxeHM+q4EInpX5kC9iT59CBI7NjeTP2fYoX+g/
7YIIZG9bboCzX4KAt2bA8XSpotEcz9RqpSE2lbKNYVgO/r6exh63IjPb7ucjMHKL
jfpBSMvEjv+1uTWuNTKgjMwx4yhULs/+yvRKVr4wItQxpdvGesnfo1jWofOVn6ob
0x4VsgVpiTrsicT0R0adyI5v2SyGBlhdF+8lVqsQr7fS/VNrRtGLu8haNu2QZs9G
rLsp5omnqx/6HpjghkFTxMYCOrgZXMJ5LgYwJTfJsx3Eom+T5+ImKIfKOOvn30uB
0p5Jz0c6M4KsnYSh9fWerFbtB7jE689OrUy2BTXM/2VFKDzOvp4GD9P3gdmEAOgK
ycQm9lHefgdECJfZy0+l1aVEwgWm27yzcxPIiP7hvY4dXcmV6m2Eqf8EC6YyBy3T
3mN5wLD1hn+2A/X3lsTemXbfpEDCDmcqFsiLMs1e3V67nRjgxn3hVsjnIdhfEHtS
ZACOQ17hN8XT40qaaTnVK6xI1Hr827vYSn/EqpBhBN/LsLiXE3KMCoHPBfG9DtB1
kqVTDJ2yRCuT2nO73CmOgT0qqS8Zomu5oQuUceBtKmoLrbbzz12y60vndoudn+pu
GkLkOSDWMMvUh2zgyHTh0XY4Jwfx6EifEokreup6OrEbqxri8GUrzcStOCWWYADx
CyJ2o8Q/VphmdVll5huaxbKtMrHSl0qSImv9OEUUAmkmPK41HYXUqUixn62Nx86W
YoqcXqAFOi+NLgik3T3aX7/gs+pb5jp1oSXZqavMmbcvive7LdQ/apDRbi76FPnr
Zj/h+Aj9l53AMZcy+8E9NS3MhyArO7jRkmQJkwTHiLbiiv7Nh03P/ZVMB0kbA+37
chiW4uNWI9Scf+KpZQRknM2MSoVVtR1aAKEX/8rAjAb7XZlbFhZbjN1kT780luJB
D10dlqJ6XvZ/bp9SGDHoNB9iLN4Z7BKVBfVbRDFGuyrKbiF/kxtpqbhMw5ChbD5X
x/6Q+0mJyUjT1VlTq6UoxU5SVLLfL6BOw1hy/pIenCjJuqsHKaxs9oT13uOey7q5
cIP/QRpxaSxCu0Lg79sydryF3rbNFSW/7slZ6V9rJPZQo4jTBPVXXOw3AjyEHAVd
7WjXT8yC5OuDxADVxI9k+B9EBeMmw7xEXrn/S6JShPzEGYZAeICL6eKDk51nF7R+
1x1emXMjNCHZtdy9fe8z7hmNkLrhoQQ2LW9x+pf+rvUdRPjDkGjaTiwfEc9EnfRk
gdRMIjfmq73JbZT23ffUVt7D5brBEF4gSsacJag3CHp4OTsuge7hCkotSAu1a4x7
ijPHqLYaM6Ae8ZZHRFKZ0ka8N86a9YUciwoYgBbXsbyXjkvAvq192tnkpCynJ7MT
WCefOD9J5Dpu/0XH2oLolKCY7zoXFeUVFIa28g/+nXXQMIXZTsASBAibQ8gKjuRj
Ot4JMWF8qb/gG3iqW+rHmQWe0pA8BF4x+Jqq9mp3GYTXkYSZExfcAZeXa7kglQsA
bhlos9LULoGv5wvNiNDTcADNd0/F5vWL/g29F9x7CZEgsnKcpWIkdlrlHubNu+Qf
c43ntNXP/cXHROfRu+g/h1xQyAoen3nOYew9NoyII2XVUHmA6jdMzXoQa83pJYnV
NJm8h6zyy6AXrOoX7wPPJ16lNu2Szl/F6paVZ8RR7Iam4++Fh2w2jd2EuHjPqndR
KJ021FFLb8CyYEo/p5PhzltwPuYC7dlF0uqZqcgFBegEIBCeJQuZggIAUKc5eM3C
S0l3Z3a0dYEyCU6Oa1XQ5A==
`protect END_PROTECTED
