`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2XyVO7EJJWKQ7YPfwC4Q4L4+3ydG0uOo4MP9wOtRtRYIKMOTePLrrVXwFppizC/P
ui5oRvXGkjs9/EY6qvr42EkgLjA9Tszm+WEVb6eeB2iLOpDFLMPoQTa1b6pki8Cd
lxtZoOmNINQyGjomik9zEb5bIsq2parwlt6O9dbyc/bWh+d282YihVg+1Qd/n1LR
N2nnW9ICiznLyBdV/U9myLGz0SSpGPoLVoBTqNsLfR4s+orY5QH0qDidWGu+cbhw
WNmpXV8O563vyks9UkLwngMMwMmRCINJHuZnCGcBKJzzI8V8IIgPiGOzNhQKTIbg
mYr5UxQ+moLiuyLtknbuXRz63bdTYaXsQMOCakduI3pKd/NizvnpH8Mxd7HBGvQO
+VM+vtyw0MRY4jwXzW/xtNfojogschSvxf8eg6FC+Zopk51Hs3yRBzDj4lxMgtJ1
YOfwJyXATbg6yyIqlFC54izacNJhXCK1kI2SFfjgqxQKQ1xtIRF+5erg8e6VDEVx
m3L4aFlPkl+XMXE/wJYuB31z2V0DjjGdxEWs87OUpT56gsjS/fCn/DVP7DzDSD9X
Xn640iRwE0LH6BjsxkL09ENBCJRDNBhO4tZkdM/TeD64dWMIJ9pV5hhhPDFaVSyU
oOxY7HzAWZ//w4tXOWILr5MFW6DO2OFMozxGyjvHlUwZOr/yqK0OwTZNTRYQfYx+
Lew8XoIyU/+9+xhIC2WGWVsc3HoJWTelrONWI75zk0R/+FH8PTt4QW+ubHS+/FGa
wBKX9AjpoExrzBWwYPgkNQGiRjYqaRavVcN3U59MMb2KZemcgLnehkmSQDlKnf/s
vTOnPflLjt7ovA7LaOO7hg==
`protect END_PROTECTED
