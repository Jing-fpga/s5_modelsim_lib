`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SHada/k+d025Uz9Y5TesDxFgCxtHfhDQiwFMAIPfn1i/A896lfFlHgIe1ct8k0aM
qBPMBXN/x+DM65b+r313fdO6LnVspPO4kK2GPADrKNvU3myzcX7FLfgl02XAnWfy
vMLkIKHsu2rbKS5fN6MyyOYMA0xxfPI7tebwCmuiO8QsgSpnQQiDAH1n4ckASqZF
9o0aYZZb7gauS1lz/AxOUQjDEjlvgKfmpYuwRW49UrjxyCr+KJQjuiTFKL6HGCZf
jmJWTxla3KihaVYsjSs09nI4LaczPM+GC+8kwdYEf9PbcePfFanpLov/b46op17w
cCllZowiXbPcJp5XQGvP72AjVpEhbJPFt2L2405R/7nvh5/zaBqQ7mF0vGMPFcBo
hoMmHZJPEcDc+MuhfLnTaPEHh5OdYP97cTigRBD0GDAlVXrtokPKChxwU5Hks7yU
Un/Ci2435MN5pJOfRb0MAfEblO/xxPM6ERQstbFZ7vsxg2Sg6cqgEtzpMHizJ/sW
8ZLoMaEoqlUtir3VOKiAoH7Wxr5++bFLbmyuHl8cWfhfobqW2vwqyGXq0qis9Vc0
VBExy9OE37wVVDm03VE2YVFbPSMxgzH/7kXlwwHkJ1aT5m6hcGxj8Vkte5XkJKD1
AvH2AhQZ/RQXKHMyKomJF5OXXIwqLaPqPDcJrhosReQuvBlH/aSzISJpB3GFhvSR
Ki8h4vXUqoHoCUCfcSxcwssAaPohF7iQHQc8auWN8gTsGiyNRXOOlnlbVYFZOaYh
6GmuN6bZkoBF0NbGw8uCYAjXSZv/TV4Cn/8HzACC7Xs70mCeulrwzMKc3m07Wbk6
dX8Z4d1uQCPpH8/7TWFFCZdOFnoAm+uV61pfGNCyt+wyVS8J3WpMMK9GczSuEaW1
rREmfLK5o4IKpy2YMuJi9FTjVCwlfgS7fVYkrlErjn63O+DrkqlXBY/bDNKAWmrv
m3mpzPsh03dyNWTLoQwYsgiNX7gLaW1eKmz6xz4FHTLJC0snaTMHH7bRUQEacMjD
uSAxCD2EzEsOKZf8BPnQTpTBP+dny7C7lNXd6xc2MF1KfBz+61WSMDY1cjleWt/L
dK1qVksSfoKY1ih+ABY9lsS32dmbff39cSM8oBSbRLKP3E5q+12X5kXgoxlOyg4A
yMbDd1qZdeefwJu+UDExfmdXXrpmKsWMKO7W+UJ9cey9XMo1HU1/4Cahg7zmd+ZH
5oY8TlL6vzMQE/6bL8iyqMI5tBSUTCu7nY3QJ5AWFjE2Ox1Dh6yzpBjPOqNJOfO+
vzCo/U43xRea0iVnjGc6L89u0Le8vWu5d1ffHS098Dn/Veo8q0oOu0XTo00D2Ot7
TFkqUfI1IRQ2nrBMlCxMjwxc3YQ2PH915wIDGHTV7gEmaQHWlBLnv4zFsvT6S5GO
eF/rhbRrXBi/RXQBJoOkLVx8GMnbYfKt3y0Qt1y9VWQcXFLZxLxS8H5xy7Kj1cXq
QPeauSITCWq/BZ85X+cu00XJxXlVQnlnPBVGVzwwq8s=
`protect END_PROTECTED
