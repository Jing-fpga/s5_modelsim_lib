`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ReX67+x6i3SQdSBTmhc2657hgE+UapaIlmZrYrzcWOwekeeH2XXcovdhQziv9ErK
IEY6923FyZNPIURGnXASxB6eqmJ6scRj7BqDei3y6h/vNuoii3mbZJGwdqAH2m8z
CGWASqG3U8BRvPiLAniq2Lg81wTwwjqxRyfT3Ja+8Xfl3/yNmYSozkQdiQB3PS5e
zsU3BhNrspw3ZiKDrXXmioFyR8WPphAy6TK4fUfVw7yq9xWZ5Rz3LZROUONbmTrR
lSDEn+t6iOYrjICV8WoYXfCVcjuNLg6wL1GkzLhRyz5L9QfZXqxLp/bh5yXS3A4n
PkYK2cYydtC+kU3FqYfBA2Ot06Fdct5FaC4E6M2+Fagl5SrM0wk4/ofBqzW85CjP
pdEMnLvNqdLatN9winsXQtnBWD5fbWErfPAdpdpEWJV+dfs6QA3aa04S9tRFXWZM
ckF9vhAnK4GCObpot+fUO+L/WyNSz2VyAyq++SIWQqZeElPjCFwKZy3p4hd/8Upd
0y6N//sPH4PVyHFYDKGSvooa2AfwN09BVyOZCJ8uWx8=
`protect END_PROTECTED
