`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BgI3ljvX5+ZmOijoLpJ8lbhaaC8bV+kFou00Tr21/Ltj/9LsBzCuXO2o2RXpyxXm
hFMeByhldeEX2+R5yH4pi47et+0HbMbmLSS3evL3fTFeluDZ7MzboN4u6Jo9HeA6
/9LVKtMVGcOsd1pR9JqGcBgrlX0AqqrGMbRVkL+PgR+ejT7CT1dTTGWmc0679gf/
7UvSsqikUmhRcG9hQ74YQMt1rTHp9I7rP8kEWkEg2XvVpGTZ4KPnGY5LZJlhhDgI
IHeFXc5zpiz3vDy+q6MnO0zA3scDyD5K34ksUHGJ7cYiGUYf7qp9Op/lBrrRgGl4
m0HBbITqu02OuXxR0Gi2l7zrhodH5P6LsYokUQDHvIqkvB68TCm7/0+Br/pK0NLH
iRKbdfqbKih3LdITu/IdLzvm7/NXCtfn0SsuWy0afyHQ8nWy3pkMHx4+GcioGV1a
yhQEm7RD7kLFmShRO6JxfdiaUAHnyOUureZBXrElVS+RZc8mOHtgX0+vkrYC6a5a
59HrYOBPUjcOxccaVUHGyLp0jmt4UrZqRmiIR2OZxB7FNG/Gy3Q491UVhPFeVJw7
+Q+W5bd7pAU3AFYV0OZlwpd5mC0v4IwKes7774JbTJYDL/sxpnlWRWMZOsrI7uYr
VSmO5IlocX/WVzYK3NcbgUWMGLzG3cJPj9+AN5/0daUiUPNTockJ7e7JGUZUNfc+
y4ljxeR8S5fTEPPy7t5272MoHrkvL1TpqiUfYBfyfHt7dlb99isGVOqUEyqMWiD2
xfjhvqUzBHdAdpsl++ZQ4IyzRplMtZNqwTsIqV+5uZnMau8mToiW1w+pEgb+xOwH
q3wMF77P5nK8xHK0na/NWOG0coNK1zL4TY+QSGuTyiQ=
`protect END_PROTECTED
