`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ygk/zl+qSTxs5j0qR+3ZEYeLDqSNBFrgtGqVvuFv2B+GnA4n1gdms7tgNHJ19Jbi
lrjH8jsUsRfrc6NZj2I73n12KSHaD1VcuautqXYsLXgYn5mpeJDz77OkhiceGkRE
zphk0KIoOxRayAaOtYwXoyvrq9Go55O+WMq3EXp0adrHYpJdYJNegraoGWqU0SJQ
T+vHNYDsP50wfHNM64L2frc6BPH9h2HyplVrGwtSCrxdYvKFxl4aQSq3iepIXj83
5m2ovCDJdXCRCLrtYAGaF5zkMzFoVcGAIA6MzJ5kGAiE37x1Yu5m0XfQobJ4u83T
+LiZKteNY4Z38/yc8n3eIcpXg+jF9+W3n+B5O0VPeIjqUPXSSOpeVqT6KAQMyHty
cYcUBgslxM8cr5BKiNrfKWr4hu2qfEOnImorAvpt8qN4vIy5U6UC6K9o4XZkVOVQ
Evh+TrL7+S9eYzKF0Xk5gN9daTboOCYrnYZ+FNwzOVeuODzF0OYf+7Bgfdz/OCF0
Ms3qvdSxG5bH08FNvtUda7r//3kZppk3O+5IiB+nYLdRprZmnFT54ZfybkRcsGiP
xtNU3bDLBLvXGNAp2peZ1vEKdNsxRL7k8ukXQ7NPKUZsBi2fFfOhWMPTaO8C6dv4
JM2etyg94iweeiNSXXT6+0nQsbOpioDFtnzERdC/FZl5vU4oMqXT/FA0qW+na2t1
RVLCE582h8fSEz6m501YULupPXnpTKaKFPTsy2qzpKTBiu/xXh+KfdJdVSovXyTO
4SnAizv9awjZclY/vKGUoz1QPTTDZi//CheaOCIPx0Ub9NawB1EDGckffRVYsr+m
bB2uhmfzhcr735VK9gLsnP/gRNPS9iLuZyTgM0o6d3EanujOc8ASYCi2cIqmBssw
eFyteyFmMXHQoQQ8E7rBjG6/vYkKgzLBwVeH+d1SX/ffdEYy0Ra6b7iNrjlsJXlK
acP5yD55U0PDLzdGy+8AlsBz6IvscrIN8+W3V8wTN+KrbclaLMkTpbQh8Z/XJxXj
nsE/8SJGX5Njr9AzNHdLj4XFeEu8lU3eIG4k98JCnA/JKqX4jaqUrnciOzaivm9m
FualbBef9uto5FB/P4t2ZS0QKi5p2zc63gw0Nj5cvBgGxzeY8CmgP9JGqblz74CU
MR+MtJHjy3bPEuleR0aXmCaiGEArTdsiMIH7mWjZ2CXHb/fcBta8036QZkuHXCOH
QY1eUxH3p5PSYJoLm6ZEDjUfou4MdFWqQN91gY+t+c/ABWkYof59xDT+rE4Xw31A
ZY97Ru+4b112yfBiQ6LG/4iFoy0xEmp+8cmbgAG48GIxa4mmqH8vhqIv2HV8Jzgg
SEyF0nf9HA7R3Mdp5dkpDsxQY0rKgjLAmowYFIaNavlUySbdhFLgsT3cuc3U9VU6
lEtcHzGMXOBuo8EWueequS6KzjhCioVpxPquQzbl07NMcqbyVBKJtr4sZJEWXy2C
tzrS6x+XasvMqqY6vlVHxQwglHUgZzNX68byf9GKNfpzlVhl+8WHvoWe4k0anM0+
p60kEWFJ4PsbAS3Z+Rf7f9tAGf7hNNWrJI+VsD4v6CDYPCF5jf3TyDTa0nl5zX2O
chFIda303doRSC/3mgRvqi+/zyuHn1/TBxeOGxs5zDr5pC5+lnEYBQY0MVN5au4T
h0LW8Mqs5z76WEshs9BAVhIhCoz+HdbFrERDo2Gu3P2GJJGXCWt3KDMxe5fq5Kt8
OWkz4/S5X/liAHDQWCEVb18nQc/dftIoThjiy57qJ52lMVlRl3zkHu2lG1ApJJgt
XAfd/DrZ55qMOXIhLHXA7lL++5w4ATWF3892Z3ztBL5hG+1aFSF+hUv1MgnCPeOh
1hy4CI4wgP0YUMgnynMim0pmU6DH7ADbFHVPQGMpfE+Duc4FovAwfGWgDcPd38we
U/WaKSll2KOpIoUoIbfsYTzJamDBD/gU6zIDEYu7LOyuo9u8SxQI46oADkuUWb6H
yBWlC4v34zfgt5JKr7B+3gCaFhn0fgPe8JA5Dpf3fIiyv7qr62csy4E73fYzA5w0
CAh38ERrTMoBH5qvnO98B79i/k/1DGXQgb7riR+aDL90v5kpXXG0KZMfFbz+RON1
IklHmGZpiGtiNRSSnnoCwmj/x27e0IkwQ7H7mIaYfrTeDSIH91FZ06k4aoymSPvb
CGOgmML9CIkx8aoS11MBJRZ0U6rCYxXl4SsoD9hwZfdfodXWE6JcXA8VrUFKhFkp
Qy2Wbc6S/t+z3615F7Ctl5P01YD975shqrG/0aQPub3bchINLKmdmKOhh9gwViYm
ik+vTXo6XwTVHCFV2Z5CI+zG8iF80bOpRIT6rwlx4peltZT3SkrlWA5CXlLbO83K
A4tjh9QHGd8/wQumfXZfD4q0KzSYBdVXfnaE9/4ux8wSr5HfEUe+B0Q/n8bMpco8
jtA9RIJ44GRs0rI7eg3xP0WTxM9jM4U9tqtkT9YqOVp55BgrvzHeS2HNNvN4aXbF
rKXqJBdjAK6InV/1LNz9XCgwJm3qlZVFK6jVjrOgjnC147onyGGh46dSfCfE/9J+
Imaqc12sl7/nf4o6Yg/pfJ6qogHAm1lDHtJ1hTAC28Zaayfey7pKi2duWyBvmDO6
76i6hXPoS4oQ12sLgd8TACKmaAZkJGEo8yHeUniSU8dhXDbJu2Jgf1hk5rbaq0iU
yHdYVI/tlK/3WJCAh7XPsNp3PV6XeWpXK3jN1xE8jiZcQrqj8eCfPb03nFfkh85J
wlZ1REdz8v8s7rIFVS6VMRv9ZEzYs9jcbirkbgkW16hbcK8ejN8nHS9bcAqLChUN
0FLJjp++ZM5+hOMr4VfTQEKiWrnvTgVgdDX1+BXByM5BuYjL3q439XUeLYu3dI8h
elqghID8vXe5CZHN/OaGlEByGhITV2bX/j5loOZTCL7s7qLjvwZiUPLCmqb8/SXP
XzuUf+IbvAQrDqFoRBPoSsoG3M3DBQVZ5wvzK/ClCMKU5fIMeBZ/ZTms1L7pUv9N
DiPkXM2mTtjnbWmRtpJszm/R/m64ZtKb7+u6JiS/oCIr3kxwpysf6tf/Q4hK2VFd
pQfT1nNL5rOt0FUL8Awhqjw8pbmysCm5/nRLpMQJq6hIddCc/mPCBHoAGF3dweR4
nH0Yfz/WMpKxiIux9xpWwjBu+BLjLBIE0aGXPdpBY5u93ITIi0vrL4kFXTn8ph3Y
VGOHBj/Et0n9GF/PndCYUw/6DJXdbu772VKkGCTRCEE7AixqUT/145sdSw/5Ef7S
f0tXF/Uz5/TzjxACLjsE7Cu9E/qKH+AbQoJgQOtxbEVc5idmgPXQRhUOSYMN3dgt
GAeufxbGQqctrdvJtF9pbsMHN45sPchpRRsU/eih4lKuXNHEoxdWDQIeWNSVS55b
PQGKtkpxaejGB6gto7rm8qKZfrdBLduqBVFDxXFecgKkCsHdKeZmXJJZGN/1Ii+R
joN4H0slHiEWNhhtDz1dBW4DPlDKZ/DqY9GJEO/7YWLW0XUmNFShoycwT67Fg8aS
9PshdrHZ2+qCv1pblZRXDW8HvR0HnlT2OMSTAlnFda1Lb0+1Flyjk7JVfT54P9kD
MGd3ZJkRTd+n5tCC6SlV8Xe37gsiP1M3E6pbVAZ3ZEhKq084lhbBP0HgNvXu7FqK
CbpURjoWweEiQoWjdqLrxmB7XPw5HOunqfk1NAVVWfCbmCu8WPIdl2sqVCY+xnSI
P5a8/wRr/JLUM71bASkbRJGlY4J0PkbxcIeQ+fvV4CnbOFiXlH2KlqjYzMfutmBE
GTN7e+076eK82NetZpM7AiQirfvlldvSoFIRxHo9qkn3+7Ej8ULUVypij5szBYPX
5zreztkOww8pdEMjnli0zvpG/kbEYyK5s4/CgeUrQ114vBHEE2EEJBIzYsaGdRGQ
TzswZjFT/D3zYAAKrhSWdgOuqq/5cQqlGyBgQDowSxE28z6Fn41V1o0zO+dcNFbB
6AFby8Hjeox76QUJSoDzvnDjj0LvMTRGNrhPVRqJ9/95PFky4K52KfxvfD0oS9JZ
GK3/jfJkgw/pXbHmH4fS2dSdUlNcDWHmq3mNQsN6m1uhMc6U16wpIpYGFhSsXB6g
jeAUYVUakiDXzJQ3O99MGXY8v2ODQm5g+RgzwZ6UW9RsAKCzSiQnhXz6BBq9GumP
5A/+ndOsz2+0ubnzj0wQvGQOJXUPfs9MfFXt5fgEnvpIQK8O5o5G6MsrRGztE5H8
eMcmdQ8Rj4YUROsAOWNTpDWQ6NoFduTIPeN2ZnfFjxQvzhgc93aZF1OMD+VXVDkD
nwTOAtKIkYy5PIjHQAAmSAc9xEcrQCWKHm/VKPn2/Uj8EaWCQWebXcqSL/0QlHgW
aqjI+stGLZTs/TTRGcc6oDIQaucddcUqOcitfCJJ6AE5Yi060OY7mud0YEQt09Wx
0zNQStKR0XjX9VS1HrCa3S+KxamlRnbrKrDntaG11wJjC9twYy9F7ANdkIV7sKfa
`protect END_PROTECTED
