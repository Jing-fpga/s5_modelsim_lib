`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XUkwPRFQbJy0fDUk2ZYTGV6pxYb6lfqdvsAUOpCfgbIsu3kjh2t+9BIJMO4DC65J
2O9eTLcEI+Lg0X3ryslnBZqtV8dCc9tF2789JCAPH/BwV/tAHcr4D9o+K/EXfqnW
1jaAAKev/fOHv5xIa/JPh/PHkfrScyd+FzYmogR+/dJMB09iBrlgsDK170FuyDO9
YPH705lUubJJ/mqEns69R5BV62efERav9aBAc5n90UniNtDmYlEA7aPf/nJK/D/n
WJvA+J1DK/u+FC8a6+1c3ia6BJcdlNZcj8rJg3WDhexNPWsxh+8WcK6gwOT/WOLe
aEV2D8s7X4tDk/ehm4iwZ7QaHIzigBFb80hkj4+wD/E=
`protect END_PROTECTED
