`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YDFnH4V27rf5v14AxQU71/GcqLSrfvisSTtfcDjZ1p0iBAn50LBUlxRI2/SmTUiu
Gg1A/YAbLb2UG2KCYxKhXxgFwcgrvRrrw1KtjQ22h+0TKH7tcue/JXFojh1uIBFy
BDYZofYZI5B1O64l7xgJmIGMwQPEwgsOIQw9m78KYaYMSqOz0DkvLPp53J/t6vlW
ODGqIShUCM5Dir8y3Qo0N4PYo1zo9a2/BHvsY0NODoql2aVmQE/AgZMfgXfdlyrU
MqmiSceQtwCDP3cXP3hI3Wvv7wv7vNABc1IOkAE8Ejb21T42nQ3NH7m+ReJheHcF
4F2hkd+RfpOs6Mk0hYztkxjGeMtgWpjy0MD7XTFYkjjeH1eM1mHgqPG5XNxP4t2+
sftS2Qyvl5bKPC3BM+pZZlVvo/etORPuZ04cWbJWrLeRaV/cJf2G/oBqVOOYGnCC
SQF7JHE6p4bZBHWKPN1FcUpkfQCsrvrPU7oJhmEh5LdlA1Bd1CpmvTd7X7A6WJdG
+L4ZSmyTL9ztu1mYuXZLBJD85zCDqBV67WbQbXI/3CBD1Evbcm8WO/jfoZFHKAuw
Ubb+1qd7uJB61IzCA2w40MBfVXg1XmkVvd+PeJWbuT8mJifQIDgRLhCIf/zQVRk2
usliZCZxeVMhpRAwTwNa4Wmnv0O/0JS3GrcxkaiFNTGM5n5GyDQkNoQ1rDQPkigF
X4AMipyT4S20Ei/ADNeXJPsWzz2W46Ad5V1/kWIOJvZOzbcMKDwz3u5w+bc7Bv4n
Gyn97t6HUOPTKtmprpgy619anAZLZlNREF8sg05XKWW1AhnlTsxfKkd+ntegFYhF
QCxRyImvxN21aluyvQfdkv5/NDjnb5c3m5HNkp8LTlgJVuAZQKrhi9OvaeU79/R/
N/tDIXUCe6azEikVQTiBAwOTJ9tY/Julj5X8uNVH5qx53/pBfcqm877KxwKWzhXd
JEcMq7S2zrz8NGkele1+AKOuIIdAWQGUGg8Zzl2eC9dSmKVVVksJHZKhBAsZakDt
KokTvmE8Vvq2Em4rQ1eEuWEbYMj1FGSIPl3AQtUR8wI3nsPUa8ioq2viYaZaDoa2
TFjxc9AAl+vMnix/H16R9pSar9Zhd4Y2PMxM7QJgD1H1jASR1I97Zako3RlUJRuU
WeKSISawO24CUPE6yIq7i3YC2rAUotbZo9cB1T5o/SFeVPDDPMQrbhDzLAFYMSFu
KG8hLI70BPnP8tNBDnoeg2beYiKmFnvbcc9XqPEfJipY3DSbBZGRsffxIGrcikOw
DdRu1JxmZc0fpXG5v344BlM0wrif9yu3uxPWLsd1sX0KBc0ByiGfd4AvsN/JxLiA
Vp+e+F8TUv6TelbMcV29c/q8rxLDxNxZd+jVxeniO1UjWzrW5wGR3yeO7McIGRsK
v/EJdmvguWPUqfjlyaN6KCb370LV2VTqgbvT7rXY8BujBL3ixruZtwNTf5ozXZfs
/9DDp/nnQQ1U5800uuZ5dIMYS3ZjvpoNXsAbFAYig8XF/zE7in0kJ4eI11hco4F5
kj64HVZ6Uzzxg3KjwgKTcwCIU8+75Hy9gNlWXONuNIih+HykqU63+OnjH6DhKr7M
YN2CTiS3kc1otF9FFJkp/NY6789OdUYHdZi4Yc2eZFkh+fSGLgdarX4RRRQWF5BZ
HP1SsrIdr809XIVHPBTeVwgAtoJSA9ZKGq3hX9aD9lQhD14FHmNHeScLF7YkANqU
9rFj79B4r25rGi0A7NS+vJE1raGeqHbhluPJjR32DhNKc4Z0vbUwDgPJ6u+e1iRW
ZOz9sMwlYkZ7jQV57ZrsHDBAAomqq2scL57QLFVRTsGFO2ms5lheas/bkcDPwiQr
AseAzSa7NiPA2bupNZsrmzUI7NSa6jYDKco6E2Gx40HIJ7vP/roOEi3EGHvGyFqJ
hOAtWpoaVL1qbTGjkUzKJ+xAISDz1MpHN+DcrUwxQ+cm76tQFTF277+bsJIQBiTF
OwcjX2SS1vsNvYmhSzzyTDxK5WQXL/AIHWKVxsl+6sytdsVBWRBgZbqp9xdrtMF/
QHUjRA5lX/uHDAQGv5Z9JgVcKE1CHfEcb0HKncZD7AJARr4ugZkqWFeXFt6ZuAO0
zFRcwDpMoQtjQd9bzTnx22l6+WpMK8KM/CnInklR5dLG663Xpub/Tx2YyPxbVFN2
8LPBtZGQEGjrhspeVhqzV4CGeW2oJpksXBZWbFVvU2m3iyYswQFky64ACIXljvfZ
4Vws/xl+pVIYFfA8e4+gU8OVVfRFxLahH9PP9S+HVt0QD1+0lKy7fVcJjX7EgPsH
dl7MMJJZ3QEMUknawtCz5WP0IgFpr2dnTTODqeFnchk03fCOvxfo0XHZnTkKMyfX
4k+U6InQ7OEIfaMP06pHBn/kCxkg2/1BfpY1rVSkVYNZHstHAEN9Y7SHC84RuryM
HeKthq+hZPRZP35TZniKp5S3zTreKkVRByTAcWwoH8saVB2uyli3dnQLefZAUI4/
PHZrsVHhJ2Rmx1UO81oq0DCCBaDPIj4c5+Nf3A86LoOeDcyby92UGdez/+Cs9TWz
qxbXjh8QQeF4Wo+TOlpZ4p4gYU9rnnnARROKb0VPQyv3H21CXDQ7jxBUwc2Qzv7y
BF1WvA2qYGiUAzWGJ8oohptMBsxucUMJDPrYLYTnBxd7R+FhknrD+TKhf3jGlrq4
Pk8mouPNBIdQSNXtkFkky6yaJnG0Fm6s1MtMToccOGTXHr0TtzRwJynHylml6nw/
bJ0srN8AAFhhgU0od860yhIOuZn0kBBKzekX5o/2RQ/NUzFqarr99AdP5TE6EBJ+
1CmORv/bh7p0XKgjqplGjbFZHyoV/cGPzxNLaIrCj8JoWOimY0PdbuyFRZYq+BcJ
sJlEGD0wvDW+eSjhMmRba5hqzWQenvwxCkEfziLzoOIJ7T5A5u7hXACq7wJzHOsj
Vs1T9fSE/0XocO0Y+Xn8QNqVcEZiYVFvRbov3ZvywINAk2PVPn5pFnELOMI5VdX3
7eoV+HKEhkaKoU+hdJXSorWlfnhwZhKkQKctLcodsu8LGzYDeskqB/qj3wkIxBWC
HnEOpFY7XyJ+zggT4bM1b4VIQVnIB648rEh7qtpSPJR7lgDrJb2EUiWNZQqshxde
bO+64F0IMVtJdwQU2llhi8juG+I/I81lTlnWGtsmfWorJ7BH1P2/mAHogfAIaMHb
cuEnXfZQCLOymWMjGIPSXeeXyxLNw5uSM8i9eHpaOsZSoVNhRR4XRPV0EmDXFazp
KhBo2Hj86Jq+6zDQGRSbcSoLhRLCwNVyOGBG7jDg+vbQxP3gZ75ZwiCBp0UGqF4g
z8+fiQa7YPIVUTDD2azyUm0B0+/SsnlEWtWxfCBz091TQaMPRJwwirMgu5HuAZZM
JEc6QYCc222qkBR0QpfszoXrRZS4ebnJbFukZce0ijlJzm+DVEK7c1DkPrApQ0+a
IcksptT6acpKFcE+6lmDrJQ1hWQsvt9EqRJklDswcBpMbKesnV7uDNymLtEuQAAL
mOsBIbd+gbHrD29UQaDD8KuQIM1UwIOp0MOLaaksDPiOWeWF9AELY4kB2xm6+Whm
XGP1N+5vgUvKc77TNbcoHtXDMvAr5cFNi0zU4Tv7myXQlubosvIMQcwuM5xIHXqe
yRVG3BQ1dAwhANn40eo0S0PZ9bPQEXkn8qnsETVXXnrMfMw1r46NBt1ImHMYFW3/
+Md4IlVjcO5rh58fmPAp2ikXmLP3a/8jKd+6ZHbT5xuC+EoWSxUoqzSrihBH75TQ
949jHhFLF6vKnto9XsgtFbtxAmKbDRQnpO1KV+Wb5qjx67RnbmgziFJPTsZ0ywX0
g6mrBBrHBOsuOFrEFHA/c3wt8qglar4S1MUIKXN0Db7GeeSkY0UBaAkFCI7W53vW
NfHQDaalIrE9/oGQ51j1poqCg/lpl3bL2bN471yPvoQxoMuOrK4tTTNbbSL9713k
rZxENJ2Zs5msHzZWqwtIjlQ0F+cddkdGrHgZnWm4AdrPxV/e8zh26PX7He6tPgHg
Cwlv1nykyjIaCqOhOCb3rbyPnkvJe8fMY6S5onMxRJoMzMNPig7PsY7Q7NBaBQZC
WpZSn/JZQBeh2md9yoUCS+wAsKVt8aSRSydovT+c5tAkYsAYp/X/aZmbZnFfdRXA
gwlgkF4n1NFoCEsJKAyO52EMm0VWuMkXPSvT1t6YRbbolV1yHizRkGIJwC9uJDC6
4DP1f+rxC1w7xjA+DXFmBL/2xT15Hhflap1TBvBxdwoiJBIVACa0Lv/mT9uSa0Vs
vExvL20glG7+bKqdz06hoqAb+AzKOaSCumAx8uwcEYQCFuVVBtuWE4I5ghQtEl4y
PZE6nib08dY6w6lsXz8o6twZVhXIstjczFwKQIb4+4+MwvvrT34TagO8t0gOVMW9
txh0x2WvYFUXi56yVMPhivg0GRlc5ZKdvW6i+9oheNR1M3H44APZjUZfv8807vI1
QP/+EC25rg8BzP6F+2ZFvPzpto9zwz3dll38ScJ/wTgfHbN1daRPgjieT5x5AoD+
lTtmcS/woJqwc9tMAXltGnPSTGdUWpHP9V61JZG/H/6ue2FLmcszo/TidGR1yanL
gf1gisIU565+xtZA00GyTliZrmXwj5zeLfX3iAN0TWNEj7GiQzWOrvqvIAY5BHLu
`protect END_PROTECTED
