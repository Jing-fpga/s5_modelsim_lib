`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XJx+KznVxkeoDbCF5VavZf1Y3p88JsyZz5OqCrstMgxdZu3JmDUU57uFMka3caD+
/7cMdLqoDcJH3fkHmqRKRfcQf3ksU6LKoZ8hf9gL6YK37T8TeSSu5Rvp+uDVBADk
MvDbHAWOPSJZmwYWQ1L26GUf1StV38zX7Y78gNfApZ9nDOeOzG8c/mVn5wLtS2EH
5Q9yFDuhAla3icDTAXuYGsi2lTMX8QL8LcKegfGaRfKniNMNyjojJjxcJTv3O1IY
TdQWNA8ewL16JcFOCKEvoF/rxzpa0knAKGkr6yet2Sah/xwMHsoJldG6TVBIG3T5
xwP+CboEeWtgH22c2XyEkLGY7EdfUFR6qWotuh1LctyWd6T9n1eMA/ZREJPQ7NES
L/xodFHdINtSDI2Gif53AAIaq9i0QvWkasaoVygw+uCM2QqtYVXKEkQQv/EMX+wy
rBoMFQNX+llGKXshe9pRnCLicjmR6yLeXpv/f/qNGR2SQt6yqzzkJrIJVkeiInK3
ppgINpdegNMywTmYQY8KCeXeCCSZ2vEg8Na8dzn+CDpuqRLeanKHUI/sT5FOafD6
FCnlJ3FsTvUIM216ZFsRCW3nqjhchTfmV7bKHr+YiZJRAPQ/htbgsbeCImXy/WF0
EuHFqafYgoLpxp57x2T6fPegOl36VQE7cP4y6mFuN0E=
`protect END_PROTECTED
