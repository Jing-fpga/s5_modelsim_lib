`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CBqXEXDIigQ48tPdfCpGelDQVvo2N01j6WW6MM4ip33h5QViLg/YuOrbrrBT9PrO
QG2ijeJ09flAY8LMAccf5rvS/X/KgdXvy74aStfUuqIbF8GoV8tJr4AvpklIzmLJ
xop63pT+SU9B6wyM0F3h6SkKwkAE56NMBEG9rxrqAlHaYE79TolF9dxImqmbPikK
SNKLExFRQi37iSIKopBATxErtiBs2XAxR6aNn0Fme9JFfmzBLCKzLhT39/urEayQ
Ow+aNGKny0a2HitOBISQlbUc5/r430XWUERBfNp42FpXZ0IgpdXzl6dxWVnwm8GC
uI8cE8Twybknl8eMFYM3F0cOp/k992M+44XeIKVXYkh0DGormOq/CegSaNx3SpqO
sd/auNN/gtTKOLQZO369j8ZO+bY15qY2TZWyDhMu6WS/o20ccbf8wFIhG7FVqRCZ
orcxwQORBpMsNvagQF2yaWTsSY4qEh6VpntCGC7JUpG5vFKY4NXWD+6iojJbFjli
MaYdlvSoQKl8CkZH8ahHQ1E2sn/4wUb5C8a3pV9KRa2Aus5xAHjSOrkwpwzMwEmK
pOBKPhhDlAQUN5RRc2G43GRuD/Y/CmolHU1UaKtx6CfY6XyxJEjoDTjcDz6wAxUQ
dA1WeV8V1JZDHcSlJC1t1BcnuYX57L9ff/QWgOLVwuORUu+2YWd/93l2oRGRzb3O
jFtvQBXmu0e/JtRhWD6IPp3X8WCda8iUo7ls5zJOrdT3DBRGUISw4/hQ8rBXXDCo
88MZwAcdk2oRigFl4zfH/0U4/L27slxlmOlkZRDplkX0Y7FExzVWA0gw3bhQ0ZlO
x3LrX2uC6Uxyr7vPM7qz9C02zEUQWhk+Vd2n/XDJW8gVPmyJ3xIkZBYq91ge4P//
4UgvFOSFXcxPkRjCr3l0+DAmSYy3ck5J0dIXm5DaCTW205974FZ2hg0Zv195U9rU
wJer4C01zxYWOEBE9ZapUJwPXFApe8Cs/Vh7k6IQ0j4oHEnAnBVj1+H20JUn5Zko
Pm2ogOMVmnGq/aPYu3np7R/WlpOM6NbGwAl1ib6Hs4T1n/O12uIwV8khmhGTxSSm
5H6OA6H8O6plVQT0L+hKMZmjTC7XFVz9rjt+ukJYiwTtSuIQG+elrL8X3phb1sfu
5xeuu/u00ncbd3rRHeCugg6z0pj38EjOa2JwRcxLdoMnSQj/DhqBQGsAp1X2QRJB
gme0bO+QZ+14jlhsyxo0FHyJRumEhIaLpGB2RvGwxm03cqLjonL7bj+PkeDruwFd
5JECzlEBwzeX/6nPG38xFL+T7dAc3FHk5thBBxlkZv038C567Bo9c407AGPZMLk8
5uvrzjK5C5IZ7HacwyP+JRkljGmO29ivR0NbAMPTZGVi5lDvQ2EI0Py0/RqMouEz
fPKZu6/9q031ZrxFIGlulJOoLeNF6cGjDfKMxAjqxwyOFtYXFaHzVkiVnESMpcrB
pyGfiMwNXcB87Dmmlv/3nZHdc2zjwD04kXAa9hRN/D4DvDjxCZ09ioTCXqgspRZc
/8tu+Z7/GXwJHlZXckOvPPa++D+G8E9pLdVb0w74sBR58hwxKKlUPEfuuH2BaN6+
sBv7GhlkT7dZjL0VFE4flCD6ktpaY2Fdu4dU+4nUbnk1UVnaE32VBgbB3nMpY7q9
q9AOsaTOULijbDvzX+rfcnu/peBgtUm8ZLGPQJ/AlddlpYmZn3QnWEJuXxBOoLds
2HZlAHzs6zXJeU5HwjzQo9bK743hI8uWlW+nn5gy0cPgqs4WJEKOWjxdOr5aPSIz
e+TtRSx7eJ1OiigoqauAtQf+b7TwXeKRdlmz88P7FMGkrbMQF8bnQ9nl8yM9bPMG
`protect END_PROTECTED
