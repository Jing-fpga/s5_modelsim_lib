`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tA9VsdSey+yE4Qb3dJglvyfuYHMzIMD7JENVRRPuUO9eMtVDeUAgF0b6x+3Uq3CJ
NtU08+fInbnrreoqPIC88KJRsa0BZQM1tDuQ/OWW5zuc6q0uJ3fZGmAF3X5Ht+19
fxSHFIgQCsbp/BvtVg8YEIeX6T8BVE9RkukjaHVvQAHEfywj3tBpRmdLwk4sHU2T
CTt7x9I4Xn/mI4PmgO7qLHY+mIJOCiR2gTuAQ/fPayqxx4OdlwACU4mV+yvWO+8p
P2hcD17AWnEhu/P1rbooKvIHZ2Fs58kYxOLsoLWCRh7BE0ncY47tPYnPhhHj5jV8
queL/rSojQyFCyY+tYS1ggmnafVdvOW3BMMMHBvShHB/mpo4BpVn6k1xHLsV/XSw
UNxSpfy8JSkA6Fi2hYmV4VDjxz1njrLxT+JAxf/JNc3cXwIqJep8NH7g4qEoOXuA
O/UyUNx54Jc/BEQMmKvxml+U7mCZ4beGsxyW7xrr2Abcr1We5KY3+Js+4EZA5wCN
ZifAqRBDyVOU1K08dz48DInuVBnAiedJ4WY1/Ul2AoICuOYV9RiIzjmKbg7VsecR
xJCPsuzZkollvLA/KRMXr7zJvqSbkmSA/bSGQj4dY8Ivb8kZ0SYIUu6ZECyfPUXg
VNGb08hiZVB1ebaMdKW47fgfa65BgAoV8fMqDj4ZMwkAcWPWNyscgcTGgt2WAIPw
`protect END_PROTECTED
