`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JuIBkbgvjwcYbOrgKoINIHalIOFZstd7glDUVEO9u3g5es9Taq75NHEdNoNiPXgw
PhvkNQgXRl/Gl3oa/jpYSG5n5TkoRFvb9XPhngwUJxsQY9mkVX8JiDZw2+pgSPqR
qMLrH7DOIy1DJpO/jtG6FsfefL9ZkfkPpJmo3urVMywTb52bjRXGOGdkLOXQ06Lq
jd9CW7Z1XSP8t5u68cDkiQijrCkN9SaeS+GS+wdZ8U4q7p0n49/qhu9DuuDtMK5b
vTiUVTmW8oFpX4B2le8nA+FCCoL988jkfxUyFM+fKz1vm8t6eLM07Xi4HjMojj9c
8Gfew3071wqmv0i1j+LPPdQL9aRKWiaj0OUatyfS/kWMPUgPKabj94wHAbgGc/er
DCX5M0jgbLU3LbWGA3PDNctlNBtkNR1RePEo7Z9S6dAol49gfv4dma5WwI1kb3Nw
K+D1VS2I7HauoJPZnZ5grHH7UkhNr/0xHDrZDodnzv+ds+dcxF+1eHXxvDeNKgz9
GN2i9MYzEbS08FOiJaTPSgzg6kbsNBwbqhUu6RuZUv77jb3rQTVMyr/t3YeztMjl
Gl1A08+WvTKwvr9sA367ZQTVO1bw10KtYswXzyEnau6TfjSo/EFz9odUMVIYXCSO
UpVaEij2q8MMY3H5Wlc/B2C4aUA8/raVLSP9sinT//OgbQTyusx+vNAMYXtMM6Rc
jg8dWqubuEyxwaEoB2U8XrK4GDpBZsPCDMxkdTlxxyOr9Mi1kykobwAhGnZQ+x5U
wifjY8Uw7HMHDvJzvBbZxGi7cDcnMJa58g54/tLHBWn3JDyb7Pg3ZX4y9cY+B1/6
LR0k27rUNJN1ib/ur/XZrqwYG0PHf+jT1+I48SM5cWQcBwQmcGKxzOvzUqK4MRr1
bnXwSNWa/GA9ISRkox+ckk+1Ed4Nf6vcOKzNm+U4ZwfT2D3kfoV1HtaVM6eKV0K0
y3W1laTyGpcODOhcwltVwuunr7j7MJ9IFV1EYtZsgSkJklKE8OgJ7iRRZYKu/ysT
pASXHUc6rGjwjQ7Ajzv6KhS/9VE6CFSM8XUW9/eWSy8sJcn+fPhdwU3GViikbSMH
3DBwhq26b5hEfzI0VCjzSugGn9IGHzefho56yDFYXFySUlR7DLFhw1IssC/Gqr9I
4mqNvCufKuow0CtKxJlhNx4hqLwKZPLjnSW2yMMTBP9asVR17QtCEf05Z4IjvS8v
wtOkEZqm0x/l2KmIQmwJ8fpUguG+GdCCpfs1YnxS9KfmQ6F4XhON65J2/VwuCgdg
xEgkzbb/grjEg68SBbwZLHYVRArWrIN+MpM3BNnjb02vaS01rc4TpxFGgc1bvYtH
hD7sn9+jf3LRzu89OSAN4z4HPSXyFpcoLZSw90hDBCfEulUpQRkOYC/TPmRIrYX4
9i0hFOKWj5iejOx6++ziNSo/d5uDsASVUpIUFJ5t+pPPvFIh4sztZ9nflEYsKM/7
m+Gw4pOiy62XgNnjXfd6dTb+AE1wZ0fAhbjulZXxOavRKcY0aIw/SIySaxOYJTKy
ctUQa3BHj4TJNHmvHP+ZY5Hjoh8Pz9K5IxFB1f6cZY+QP4mK/6AAgtsrDIBIAMSu
Fs5dUn/1vltW3Tcb6OM9kdBu0PFC5h+Wez28E8XFtJTo/jMar0bCw7O/qzBcouq4
BC0lPBaSiqEu+/6ylvb1hB5kI2P2ex2SvvAmQVTtFgq5n8Bm65A5VleusEBErKhm
oDv7V5JTwgAY3Zvp1SyvWsaTR0ZuWfXc8OvEY/7sK/z3GJqVicX5G0HsgDo6r+/T
3g3adrz/1OfKhCwgMYXAcUAgoiDhMqvCeRRy1xMiMEQFKuswKXOuAqC4ZQGYBqvi
kLJOaWHgK847YEOjvOVMKcvQVfxycD1Mzgwy+dhMBa/Ha/p4/Ib3R68T4L2c5p0y
i9NYOndkfdK9LtotZ0rCzvtak1W1+O0pDmEoUesL07MJCIyEHrpI0YnT/XbvQdKF
g6jMluBTZFvFT+nV3fjTZdJ3qR9Cvj/kA+D/Yegdo5HgodlTbf6MkbW0MoS3lKCQ
7WgfBjVxV7mGBI9Kqhf3eDsdGdMVoWNUIixx/BURTXMpUUikVzPPnyKtE36d/oxF
+iaJg0BRJFGErpDv7fLm86hDjfplcljhiqDMYd/LqoJMY2ER5ENzE1ALLoz0UU27
dsozff/F82os1Hor2wODzXYFqisrUxLApXNGzuFZwgY0O6frdfZKaFWDJI4P45mD
zK8pr0tMDjShvRxErXIrBaTFwdIorPHs9bSGwkSBi2ZY+A2TCASbyYZzRqv5KWJf
RTZFenyDMVXeb9sjYnkRdEyaMKH/Ne27YusSieFmSYIm/riXSZKD0Nn3rljo3mzU
7WZYlfYHCyrvjlDCE9rKszmpjaNQ2qbp3lzdzNZV1l1sFMwY6uGzucBhdos9zwCj
FvFHd4rmceBJxjPObKRCGkkwKImZDPOJ03xyGENym9E82gumSX+Qr1QCdcEmyuyW
t5ZBqoICNI/HO/JIUKO2Q2cT5O+PzZtNK6ucMNA2qkIQ+dyIrvy5Uo8OhaGrRcqp
rv5+S0tD+vQXylge0ut3Mx9q/V1QDHuZM2m0h7+b6EE1Ul23xQeD28WNysxJGxhv
reem8fqap/MSS9w9LH+nqmiNpJjohL06pdW8v2G17tts6LdOdxRLB9B9MBIHleVp
DXPExVlQXZf0lLM2EWjx1r5U30Y7WLjJIufSdG63CkFpnWar38yd56X/dc1ctvRa
xgWG8eTmyTM8YuqySXAv+2jLKDXaGbdRByWUSG/NLMGd8LNJO/2nyBTNdlO722tJ
Wseb0GPLCC2lXpsHgsM7t8bhdKsKa+WBtoxTU+IB0CJf5jZgH2rY3oNEEmExjSf2
uvGob4LxWfLi9KThnu1LPElU2U2EUuLh5Z+sJqmFHEJCbRhKhHej0NzDL2G1keTU
auNtsn/+oBqMmgudGy/XPd9+Kda617NvuMxMovGWSQYeglJP0qYkgUiL/Y86d8gC
wj90oJO8ZkwPQFY7gpeRheAJ73hmmQERtX2bAl1nNqHy+6zl0rbyiOwBYz3qr9WO
VZquPW2tLeI7xPMW8F9xESsQ7aKinT8dxa8jLacprz/oYpd7qIUM/nMvM8nkpHgT
MNBnzc3LSj8IUG5urqhSdGzsvJlM7h30vVDPyMIolkE9v8+jmmAHE5+X9ig3IoUB
6esmFqqyjr/LBbdjIn1kz1np7gq2xxkPiNqLtM0wd6C7Er1N8Lzy4d7zpISqNZaA
T9l/ko8XAuiOUrrOVW3Iljwn/2+dyG/kjPQGt4Q3vuq3d9ORjwInGQTAdVDfv4Tq
JmphF7El3ED1j2HQV5Z4o9Xi6zXaeFt4vTh2giSVhCXGGKGi2HELaO5RpV0hkMmU
zBYC2qOaS2ndIpGWSQRKwFzaeKt0i9r5Sq6HCtxO0JPK3cqWpU4V6Fc9905Q+Ct1
hf5INZJ9yA7yqxBjNw19gwrFkTcrn/p2OzR3T+Y65418wCJwPXgXFpM5rnoUrxf/
P6YLCcxhU6rsJgolUG6hXNaM0nl6OPGnQV5/6skM7KiUNRcsazEgIdHQtUn4wjHc
TX+StjkSpFnmyrZLcPdsWhNTLguFml7yiaR0VXCphaKHfQt6G/DTODKWnOFz9mKV
mvO03ZhxdmN8XctcM8nAHOqDoaQblrR7Uu4s9ZmEE4WakRH91wOs8Tu2Zi05o6LN
MWKICusd4OP5DDIKi5F3Th5RUhkX766U0w/MupPvkVYzV3qiSx594wMhUdb3Wx3k
L+hDw0X35EOp71SI9nEf6LnEzHZhgJ0GePZ25RQrJKVRad1bczvRpdHu0dyNKD0D
FSm/BDmm1qkWg4ghMdw6O6RFsAphEzvcoPJLbTN2SP2fuoqNaWDQczRSjPFzVUJY
zVq4q+O7i7OuXby0bCKJxqLZiVCDZxzmp6qkoRJogkj3k6U4KYEq67EZVMt0T1B9
NU76iDcXTANKJ4goJVdBknjozUpbnzP9nNw0ra+BS/7Es06EuldTKbAT5WvjbaZe
MQoA/IvXyea1XBWucRDtc3PUgq1n0ZhZq3r8CovJqj8CdGZmleKeDCOTEuJJzwKJ
FOZ7q40XVEzVft2ze5xHYvDa/heE1CY/rvqhoEgvU03RHjIsa6aEkXhqc2Tcfj9v
yayr27FY66KYZofA6e/TZpmudeXEO797ww7R2aqfmDrzPggGo74AGJ8q+Xlcz5Um
VlcUC3/bZxpD8yyB9TpokqeGotasQ0Zh09sXpleTBTbtFTwzhy3ls96633GwHLkx
uT4T4cMsqDexY16dmbAVurZYT9R4O8nahgdGnuY01zDwWX9OQaakm52IWPjoef0F
tizV8FBZgK0HO+GBkx5ydUZHbrkiY+AD1GfIbRvJYs4a3ZaAF5ROAuZsjfc5i4pk
H0kgomdnHaNi26ipMLrUOjLYqlUxoVLMfKCG0gOXgaa/m31VHiJaa9QZ84Aeym91
cEdKfTgsKsdcOfpNRWfQHWeY/P3EIGzwHmBBnLjqbw/1IV56WDyDPrK5h9OOH31/
bLXju6eYPNwW2dkRqYZElSHlhhUxIySH8ocgODUuVi5ysdlgmTcmRdpMeqQBy3fv
EMyWjcgEuS85mYnASuCS37NiiT0ql5OXNxrIB/nT8qeaaylbAxGdgrvF5CBs+lRO
uXgil5hCzNCQhdlbscHNJhvNIuIevj5PgYmVg6Q30iCO0hnk8UI4bwTsoIvF1jhP
8/oMlM1Bsw/wLcN5Wg0cD9dQMRWRqOZZw+TpgCc8oHAgyIR2oOO9A27kc9IIqe6m
cRSrfTKJf2UXQ4IMBanM754CjuONd4GM8VBGHMQK2/OHNNK0UwElCLnwjIYPOmO4
MbaF3EXSvvsalGc4InvbyL08okIZT4yovKkoQQp+/N51ZgI1ioKS/lzDQRB1ZFly
zFYtdKvdOPS0xPZhXdMHsTeKTBqfIkoBv/CGiLzoqAyTbDNxDUB/K7yELahZn1bP
Ewv2rXf4NSazj+k4lO1CUL6KolQXy3ty5vF1rt0LbPfpZOVp9RMo6m2eDXRueZdw
43nO6za79hKH+EIfGKGSVCprP4nRCrn6sAajiALHxGK2RhQwLQHtN4ZjBbL5rofj
MqXa9S26V7OZHWfEmH3V8di7GTKLt1q41jg9623XWzxhn66ogiUs/FoinSGi+lGR
sPpyA7rXWE91aDbJbku6WUcR76+VjRbjJgRdnZ7LkiDNJ6YTaFP0l+TsqN8tbzN1
qDv8IvZSePY86GwHmP/bWWCJ52YQhNjtzVd19RhINGVbMcs+sNteTKxrVTvXOjlj
gFIOsf9bH2QK5I1tUt8yiRMLyiYYMsHYOztqaQrdqSd+w9Djr8n2fwAPG3dhfyo5
k+cQMLWDy4JqYwyGFpB/h+DYbEBqV2SLbekI5autDW5zspsZsZTWIzhoDTj2x7VN
K7P5ODwitSJIGFmygjVMbaq40+bT42NPbovcClMWxX0m2nvyAa1zI2jvO6NPtwM0
xTku2LCf9zawQzuWJeO8uPvDROVXJ91NA883IqBxEmCfJ/QpRzHEg5BmuRQ/5wL4
wCfNEQIagZo02Jjvg70eaO0VRPQkK1cmB/bqOdGi82PvjKjjfWtwA9KlWP+Cj7Wn
Uin4IHFvGSEese6w/bhCCYgYnLHTm3sk9fzuZRf6o1D1hMXvOUhFljY63NVTleSG
cC+3lXFMIhEVOCponvLDZB07xrMgOCS1Q4FBmAUtY9SDP15Wk/O2En1Vv9CxS3gd
BIZAXRP6Ir3df5NMPwL7jXmL+zx0D3OjuIp7Lab9c44lEqwF008rxQzVCY8hRKAB
NHkm6Rme1zGHZSMumiieeAFPeaGTmYqU8MgwHdKunS4xJvTyV/o4P6UtqFTliy9z
iRKPT7NtitBf4n86WItCBDM8tbOAFzOEKgSsFIrFzlSndQonhG1ewJ5Ztw/btTL8
NUOZ5n1F+Xf4LBAvWG3d75zipa7AGJVzV2MPSKlX6lBO/dO1l7YfnWGLfgJDXmVJ
lRgTRfbFHoLX9evwUPNUxzD06qdCPQZWHcK4gq2WNLVBkUpr8cbUfwBvIP7xbm6E
Fu2kzfnMt7RLVfJwBlut3LRCOFGcRXehlZknQyF2xh00+7ejozxWAsggY3LV6wBw
s2ybPBy1mzwwV/g1cWke7q8xMNqyFcEmCNJCzaLGPCL8mHK8KVMsEFabaU/0bUgC
v99kdKcrF0qid9wA8e6wun95iRKJejlDvTxNW06hHI+K9xx59++ytIOoGlGMJlb1
e9yBaNPUsZomGKZ8OsoOGvFnsJShTBbkmf2yxNPRmaYvSH1AyOOGPQGpO4/K/2Fc
dIM9FZD2m+R26pkKf0Fw6ef4yiWsC8vb229oT7fMZsKGlbjfx7k3u1/HlQ1bPcOE
zWWo+XD+11Ts5sRjr81F7l5PA/M6ozin/YTNb+gjeWdRgl2MqtAWnB+VbS6x40K9
zcixvAdkuzERfB7YnSQy5B/g/AtAn/Brgg/eLz9DcmwW71XskgEuA/iKZ7aFzwCW
bZMtcp65fz+ssfMd2A0WI6ClgYvmBDMZ8stOVh5yFWMgSC6pF3Nmp8Usm49V6j7t
n7xEG90Ig9jHgM5ooNcdiuBkuRxoDNBy/puGe0+t4c6BzLK5J+LZ5d1sYIzaJpAt
1ahQIdA4iOLhXTWhaIv5DQXSBIzV5/IoZ0haYRNucde3gIeQWmXM84ARa+g3dZmz
FxJPE2WR/UEUZPWC2rdSaf0ktoM3UM8sIPM0K1XEtdsX3I5BRvBMsOLfwv92hLlM
HCUntTC5q6VwJmilTHyuXDduxAiEgUDRgPSpN5dNfx+m72GYwjQypRl6875eWVCC
r7/A7Z+N2KhqmBfk7uZFrdz8HJnz4FuwP059NupN+ZmxtUDa43KgrP7MEfDfyJyM
OERGw2rhzjhIV24dCSpkwu+ENtchfcpOuxlw9eemnadH3fSj8I/93dWZ/vAsCN0e
wLx1DIiLn5z1WZzrWgwNzdbu77bqvPvgNE8qFO7lUfqAWk126paCx50RR6nee5AQ
MwycKtcGcFZ3L5gDwusePLjeZMbs6MRixFmahGRFQ3KSErlB8yPlgU/BfDMZFVE2
v0+zWLCsdcJhXT4KlND6zsBXHzLQwVpscncgJl+U6dNaNodNojPe3s5PCD5LxS68
vHK99xEvrAXG7dQWvmxX1shvytZkXzMoyfhh5jEW/Cw+dD0lcr5s26Mv2ilAQ2cz
gDlNtBvzHiiGXRUlHBy4/uY1/8VWFdJfGBY7YH1kOpJ8GKSZ0Mgt4mjmlWGnRKCg
+/8i37Jrw2s4tenU4UqIMbJbzZvaaZvs/8nJEGcFzI0b+HmLkK+FSjaYO1LfU3CD
wSbPIE2zbxUKhMUBLkbcMUETN1j/AP2zZrWyTqUJKtDb5+5NVamZ46RpK6CEKz7l
aIcxpHyxeCBaiUkVvMhDyv+mT3c9KCbw/lEc2bCRZqCVAW7GKiJaWwsWCXKVgWZu
JQvIkFBgMw/4fHq67Gv8HNlBwR+0WXD53idLff6ZW2lSaVxxzK9CkRJeFco2igmt
253pxCaPNPrTfwi0zLnatzOyUAhSLO8y0iJih+QIYyk0Nyy7zBAzdn+MHKOEBTkj
jF/ZfTXv9tiNusYoRpui9E5MWbnQpXB4PEpr6Ki1ZWtMeHLiCr/+xF37oSA0oQDF
x0B4KCz8SrahhCf3vJ2Qi9Iprpmwv4F/o+34dFeerS0uYLw5AJABt/pMSxkEdQgo
oLFYL3/5dLmoeGBj8XIeMIA0FUvkqANg3iW53IUoKRb0xfSGnl6CBc1QtbRbGn9U
kk9oeYGqrpa9hT4p99Mf0s16LugZlqMT2dKkupmreWQxsAJk5Bcjp/wKbu4UEl6r
zeKfYPXmzeyNP4EsvBt/uJZO2IAt6poLt5gptFrVR2Kp4Te6wXaHAL9tWPXGDKAX
oBvq1JBTCaTu4A+Y6jO8H5Zifu/tAMtip6GaeCOmnyTvxtSAYvwbry0QiPE1sw4s
/YG/LqNSMW2fC25+R9lSjJ/8q0OO25kpzt1G/nZvcKkNjlBCDmk09J+87IZz9NFl
cLktPq6Egn2rMx6cbCyrURiTtIqyWw/1psYn0bJ4fgWi1VcxqfhHnrb1Og6aCHzC
dDNL9cdrXomn8H+XZkJwJfW32XxSyUS/Wx7xNdTwX05+NKJNN727G911ASSNy1uS
l+IL/JsexSGAwzmGeU8cUKh7/Xu4+5bYHZMW6xi43N496E8BVQHlYMfHHyf15lB+
ilHcqRbp4kRR4B0/fBu07nnnVYlNIqixhV9BtS55AF7RyHutO/5PqArU0MsaTQre
ALYJLwNuu2OQL5g+aM05eYEaSsYTpqUKg1NLQUlctBjFgCMkkAk7z84rGwsYc6dD
+y2jRX+c4wq2aqWvtafFElmfF0pI4zkDm1v6sRRYnhIv/GT8vIKHXUzE3NEwpc1k
BnjZRsHn+sYwh6yjnEgqE6lC9xMCgWvfUA/uKmK3MJfVJWJQzTvFgU99cOOa9J5b
8GQQF2Z1auCl+UrCwsspshLmZGs4f5o8g0zi7YEn9UKIS2ou124vXrtVysFB7Tb7
OFzYHWYOkRnddIC9p76Ok9tNQPVjQAms551N6Hr9IjYUGmXHFgIX1dCROV+tntaK
Mal18PAavzZYCC1H+0yVJy9Mb5//u3vAxOiS/E3seFbgPPBoLVC3JJNGxTrYKb5+
nCFiaCCHh3aE9sG/zsAjFAzEpV0PoK8lnEeQt3MFDb7cBhXvUnWeZEpR2wKey8vq
cdDYHL1m2EtZLJxT2X0sbwIPxmL6QTLCAj3f+bgS7EEs2096ZJQy8H4lp/t6XmJg
0kY3D43Ht1Tw64YVZbS5Kbj3bWrhiI+MYDmoLqXFIMLDBquQe4y6rlxkGWqlFApb
luKX6CvYKDeNjdEVwVXXWsRlqp0AkLMlGnlPpxM2al6KnEeGiCVevgiynNoOMz89
GIGgjC1pw+HkDKyF+Lze27i5REf5v4AAMGnBaRBEwYFEOBabnumHYLaM/c2P39JG
DDYidn6MEckCuMx3rbdylaGmflmag9TnbxMqWzCLq64ajyrO6jN/5CJjAYA2uL3W
VKXK90aWCN23KABpaVdCFXcal58scL5eZrixGeypxU/vYj8VE1WJURN4faLqdROh
mJctdNNsw48q12SZaDTMT3vAYLeJv0dOLpefyqzNC6ADUI14XMDj7qNEfpwUUrBv
dMfLp96Gk8fjouaoZNmTr+q1GYav9UY1YlTzU2eFNZ38ioyfuDRVZ/yrFp5C33aW
NecSeSiVdGd0+6Eg6vnqcD6pFxk5gv/6wEFxWuQi/OmJrtzPglbEXgRfAcjOPoIn
HHfdx5TdIxEtodQFLc2ZdPqdCFlf1clyAlUTE0PL0IxjUCqhaZMuZyqELyWkpsR4
pPrP7K51p6Tcjh8OQa7KVOgx2MObUv2wim68QbMcBNSWWaHovns3kwaD5OE+Yb34
Fgz4rfBUXI2WdOZpLHo9oVprokFEiaSNDxQRaFAAwLzoKTYpLh1UReAZtAXIucSV
7khetIiO1ZLvtAtJF6WLVhPr6EgBOuM95drCWxdn2KXkYK0TatycBnLUc1dGbTL0
8GBzXxvBsjE4YPcki3w4X4Or3mFTOaZNx0KH5CjjPXFJdVuopsRmENn2oM55o/bF
fJjekG3sxCwFzdzeBemaRmdLYvoqa40PxZAt5I+GsY2m8GecDaFPrJ4d6C4PMOho
7DvKT73shdUCfXyreffKIEYk+BhOyMi1ru6R+3y2RpK2FT99vYqO9xC6W85aCtC+
Vw/6I64dDZ0kMzLYuxlZHA6IW7TEsbzjsHgc62pwsC7dExOOsKuIZs25KmbSAXm0
npcCGO45354FkE42sf6mDcLTZBWmBvAbqPuBpYqF4wFu4sALawPFAQEv9hwZ53Uj
3xaBBxjQHnYgI3SSQcFakg9Uj4igunf8zd7F9kjp7wwv4g4Ge3buXU5oqJJS4Dfc
lvz7IQb+K8Mb0Mgl5jl3KmFAK5oVPGsG6vpX5Adn5G/TVvOUvYYsZtq6Bisekub/
0/ASI0NYEv0s3P/Inal7aVTtOb0Klk90Aw9B8rLTDkndVbY3GRXsdYb9+QUwV4fU
cuM8QeLm6mVu+U9+op9Z65NMoxFqDNxS8xeO5ghAwUk0v1gmJMfudm4NuBgZAOOO
GhxROs7m1+KHeXyvZ8RWOSFlakdT+7LaGnh+XUa3bHFjQ7Y0K1+MjZRTcIx5q6Lp
zoS8C2LEnBButlfxRDRvWoo19qooeuYP5AKaG0aNnLP2KBgVOFFq7i5C50VaspMn
PlXi3pHBJTKHgXfZKO16438cZenO9GBsom5UfOcadruk3aLbz+95YtbyYhrnwxsw
mgQ8eR8hTysFvF9FCXf9F3q7CLoDQI2wTh65GwoggVoHYS+vaAXZZxXYyr0OrzBA
wACpiG2tz66u5ypaSYGmMrCH4PS7f1KmiwcSg+CF4Hiu34iZHN6buN2IMcNYZsLF
PdTxPBDWJAnKbu75o/7DkHoY6OzIDg3Z8SDYbHxGdUmDa4r2TONC+GF0d0OaF893
GV6ZA/vbXi11TK3DEXYViNwOcTtSu+fhwQURu+03QEp5BY/lsK28BxV5Mcp3pqxh
okACXePRnYov/sCVeKtv73q95pXZ11ldeYZOAoJQ0GzPGq/iH5CnaAFNA158VdQi
F/NJH+X808oOB7a8V/AystVDESHvR8v0n9/iTYBHsEA=
`protect END_PROTECTED
