`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CePVeCvsUj/3d3w5okzlZslARotHyiZCIL2pvanA+LYv4IxZGO8W3ozIKA+W3XPS
FJUw/V2ZGkqFElwXWJob5T8XAz4KMauhFeI43/BT1WJk42jy2lIM4SCmaMew2ufT
EpMIYT2lBY8naBBriNuFB/ykHlFdVuhZryS97JQGHaR1FDHWvBxJVpS3xr8aN5AE
XelidicHpqtNpcnDT96Jf29WF1aKZlUWA0ZNVQLIRkpnz8jY6h4AC7qsqsbHZhSG
I1bXmnsgtzOPUF42Cl/NwEtY80QDWKaoP59kgorlplTrwMndiMYcwkzqvvU34vJE
ZrTKaJT2jS5LGDgwT6iE90kViVnLmGJZ2Ye6eOtRNsCKFjrASOMq7280MEMXvwrT
z94vN8H6MbdLBzmKMVecKmdF9VdtF8WN68my8g21CXqI59Hb4mYLppHebkn0t8ST
5vRfKbxjMbV+Rfn1ydIxYRb9yeA1fHhpSSXMKI9WRudPjU7shHqEYlXsLGPk8zhz
TlA3rRKK8Due8sxvc/XXIHg7sV+zVNUynCETFMqv6VCnocBrWiCDL2wLyWxZn2Xk
XKvMHGGQgjJmKo//4u0SqbxaX544b63C9hpY2I+SrhbQ0DWMoFajEpZKGvvfC9qN
l2GFwVZsvYR0t2HauWiF8gHt4x3Mh8lX2C6qwD05OhFgrXTJhXEDQdT4y5nGY4xa
Y91FkQJZkH/dSD8xA2UdzOXpqJkUiJBw/O/QGGQ98xTRWoxO30CuvHEiSoUNmgBg
k0eeJPDVlENtjJyQmnCrYbxi3d7ebiLhS6s0P64H3+yO9/W9S8Wj9Ja44hMHvDD6
HHPAYAR88z9F5CtNl5JCz0MnNj5wgxjK2Y2oWB1WAxfnoWgG0+RC6jKnDsstF1Kk
Typ8y7JFm3d4F1YP2yaO0ngtxVD/oa89VXs0N0Ujk5VbJ5oe073XPuGF0HkAOubM
twgCaEECNhmQE9qIV+3ICHFhpjA+xegYsb0Ec5d5NNkBvmLdYq7pn517Gd/4P34p
OS5o2sK/ULpJ3QOU4ESiNZqRs3asCI86ARrlLh0BE1VVWmk62xHJJNqS3DRsNPH+
LTrQhnezRukYTit3JSDdjxgLvbejk3Jc3JkgfhdBGh45e2SD5sfy8Urup4I2+PWi
MvZK5HJCVkOIB/p3j3qYTVdYxwhyYWnAfrZrDkDqu1+vXDpuNM+YxkXaFbd3RoLy
r4tEqZBoz7H9vqKUZdElNoa++LPcpBkOFwTduwGGU/QM393xb7eNbuDxZ50KFyaT
urJK+0ajeIG8JDip4vs/MEEV0kar52tN64FheJwrpChWZIGWPNr4nYJmTJXaCfDc
pi+PomZJcifZDHV6xKMg/XeQf2kiD5iA84NR+Tr+n2YaXWoJdRKA7KkND1Ro56Sc
yzVfyPMjZPnsQWAny9MYYoZfcX6mq0lDsj+lBsShJie+/G3NmUafoeHkp0AqaIll
iqMlNgNwOU1ugrWcaIa/sXuEqyNJWUoKlms8pX29p/2iPrCxstTDPezA6Cj52YLq
J6pM9G5tvv2F/CDZTz+TSkPOS1072xArnKpHFup1lfuYhsxru6f9iHPbxybT95bx
ZRNDwCvshM8yr/8X5rpeoMrEwlbNj03pKJdtJt0IKrYe81KvT2C6VZuLyAkaM5BK
RFW6e44C7Db6Lx20hENlRMp8igE3rnybhTFJR7QBKcl5MysyeZ6XaXGr92ylfDpU
DrbZK2AWI+D3D8EH7ax8PUcDqV6dBYiiGNqdhEWdALyvy6nGUb1beH93srlSBH5c
m9ube/1Rbthg1DtDrL8xNzZOoCMlSR+xz6i+eG3HfrKwHeEcyCfiRGGDHfTBtjYa
rbMwpu6VsELIfjKJFEGCNK/+OUXzlLj7pquR320qLplT+tPNJmgoqdsKLoA47jHb
++0Yi0Ra0Egrmcv60wMkUb09420+OxdJMgN2nAD/EVlS4QKG4lqRdCeVoWNgCEaZ
XJBkyjm5oeqv0FEmjt02fmBnzjh4VkAS712EGMvP0JsttNv+uqE/9hHXXRAUl4FR
t63FwMeMTYlK4GYKqV/nLF0splUnvRiN9i6zx2pzonRF8Ae5V7KhqDHUKRsmQPUN
bnsE+XSYmxVDdryYKGvg1BEWdVTFYJg2zAOhYRbKjz2TQTF+ACg+q1JgJQty+h01
wUEOxnuYl0Yw6QoZMw2WBvaJXHpk/3htkCbaOcSC6YvcRDBSfzMlanCHUDfCx91I
2D4YMa+vFN662skXIzvPmGBEZDmzWVDM3flmz18C5swjO+7GulfhncP38nRcVB6G
0wkDaQE2kfJLajCZSald1ALn5ZKSLNEJ9C4KOZD4yjNaXeih/QSyv7Ep8d9Psy4p
UHhM2srbQmFzowKEY9NJ3UqG7CBTtEF5t45/m+yW+oWPNooSwSiyn4MoJiVPQ94d
no7BjQgcWFPGQv7gRB52LJpRX+XpcCvCv1w86VB5vKN+LQ22kNjHWDDE/rkoqEDl
Ni2TJFHyzbVuUJaX+Ntyi8ZQ4w0vGoG/PllgGwWsy9j39jPwYjIPoBt1XCiu74xF
XzVly3iIbC+19wE+8ZVcO6wZ4YvGNUiS0XbEj1E3yBKK5Jn0wWQ7D7cqy3FholJ6
Rbw+SzvqDdXtkw6Sog9ILUaIFTKPb8DqRWzO/3aFy1Vz78JeAuJwjHxBvRXs+iy1
zQiVS5dbmAozbASjGXtB/b9NPHG1g+B8g+EIIQpBTNTl0u1QrV+66chXRrXan3Mi
HK/OKlYzz6wpH69rWX/kDpi46qEB9aD5bRRHLTj1CemejAuQntaLfbhT6tn96WfH
17VY/b2c53eg9tSTGM4IMM5nxIqyhBfRNKat54691eneVKhBWaGPY/GpJebFE2tR
9DYWAuS3DBVn9DnWYBgORJ/snI0Ok2MIjpP3FaiuesYwy8QKojnSK8k0xYTvYrP2
OfkFCv4wOCTcdQx8f697GFzsi9fcubPuA/jhBlbKmW35Et3n9kG/DlCadIfN2LdX
elHncW4brRRrc25Tt92D+B7wMhbvNoXtOP4S5FWhMqtylgRZM0FO4Y2UPEIfxKMs
LttxfSgTBRSZ496nM8Q/N8iUKvg/M6R2dUJcQTdUx8gefdBakVzq0s+r91/p+b/c
29wSDpeRKrb5/oTrp7yow7NskHde9iNvjC3cGz5z9m8Ux9hTZas0X2du9vSo4x2U
R9E5CGC3jkr4svn+R+MRYSIhdZqFsBU8byQd049xwVzgZAnOTxPe8ayCNGtVJHBL
0a0IRLLoPvNZLUeFN2PaH5P3ZAf76EnaNls7S2KEgDMfLI2+mUa0Q9+asCXfycnO
2fEoqJkMwv02tOV6sfxHBaQ3HyrWaKRBGZIDx5oIRdMneEu5WDj2BbUKPThUVAP4
q19BDYIV7g/LfhkZe6JrJLKMB6Zbz1++rnHhCmjnKTOio3nkqpk053DmsjOIfnIZ
PksX1lTF5z93OyHKxLWcFquWo6P0HjbG/5zg+LZHevR5mTmBERTSuPqzwAt4zk4E
oHa2c2H3RqmG4EY7dr8AsdnTWM1RAVWUxZdVNReRIAilpgLEbXdhaAMloH0LdKBj
dRnJrJYuOLFcyM7qMrPv1Q9NqC7vdXvP/ej7a8F48zd/++KW3Ca12Jb4pXvj1qtA
6IS/kElzt5vBoqJtYUeZRL3TDIXVTitW8i9nd+vB9pWfdRkWqN5D23hf98BsZifJ
Ja+i+e4i5w+Xag/+pshbEnUl5oTWld5I7rXBKx368lkqaI1DS2JOEsM8EyoXIdp+
cSXKmU1tBOuEzsu9Kv0RwHlTDlZl2w845wXKlqk7BKjSTVpGz6Thob5He8eAB35s
eCWimwgY0ij70qDlQk1rku9Z+LyLV+ZDSEa/9a3gu658uKJkFeX6XcECUXi2+3+D
DGcTm2vP645mZueCtO2cberfXprSOGkj8kXCXVVxgAdZt9kxuCsAvwmi0mpxaYXx
kuIm4sBTAMKQ59A6sYRXkrrWqTDFQzv8Ib99C1q5a9ynikSlWpZK7njpP4ckoMRi
d3CXyMH7ei7YxXJfaRKjAImpqRCONJahpcK4UT17zmakt3xZv2eUqSDwKLfWmWPy
xSnrHp16npkqpWUpYfFVsB0vFxvMbO9vLv8TcEHrPsQIijgtgfm/FJddLWr7dwhp
CgyzLYhjfd1QL1mhWzqrEXtjBZQqv50cD02sgIcrqJOaFDAJYnKs+DoUAFXU6+yz
nxAH6lwWNm3iaYsyPO6YQBDgsA3IeHHnkW5PlvSxDioMNfQUKYNUJerNgYbHiEAD
YgMF0x22EkyxdksXhz8npXSh5CPErrGfGSeTkOanRyoMs23/Z5UvbU5q9pCYlgFr
wyXnBdZsulWoAwaIn2IjDyTo+6aD3KOSS5eYdOOqma7qY4a5FGrfGlKJjZhmbtAl
P+mf4T4vvZ2qJO79hgtAo/b4Z+SyyKIIOa6XJUsLUdFjlvAjrE5xFffM2VpwlWAl
XEWEtDtTdc+aM4Z7ftniVEwLNxQecE+TxzMTeCCNPfxSLj5CvICY2MQcm6wYR8jC
dePVNoZUrD1PDxQPDyoAqasFrnUcJNiVFUYKQH3D+Pg068MDLS8xpzpMXVPeDjeG
PNhrc+FCd02OJ0lu1bEK/sEIsv4FRgqPotvxzs/dhezxqBzMpkoOewvASNOnlc8Z
N+RSJtqNJeUM6ZH6QmBnhGA62b7OPGQg8gO86jhF6PGaGuTiGOf22B8AmvkSnGuO
E92cyPmtxZ4uhgD7rFzQyDBDyifbSBypL/S60eTMmr3nPEGhexmfIU7yY5FXAhhU
HkQvyAT7hxjYG4wI5W5mhw==
`protect END_PROTECTED
