`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rYZuR5pmfA1TdUHFqa8A383TByN8o+8cjdVCTKP5bVB5Mb0mI/Ofzh/tAj8JSWdJ
7bPd5J1YLEu0WWVxj0ChCh1dDEl7MiehKLpGky2QSZvbUp8JjNA+k0po2xZvqhsq
KY86KXiA8PNBTDLGO+QYtF+UHDKXIHGdYzZ6g4/+sOAmH/q9/Tn1y3PKpNM9356a
GvbG9uhudTiYJ2wSpifUWJitAqMXtPlw3bS071MRo2NrIfsdqH+Up2LkNo3slzM+
Dp7PiYuvJxUIV0S3zLbmJ82yg1130qjnmgAIoh++Tvd+tYSFgOUawA5wcGbAZfPy
0b6554MUHEm3/dGWPoZV6Uc7IFhkaeQKnBgzHM3IBhTPdEYaVzcPjxwR1fcL7Uem
9mjq93S5zP8HdfOqxEKHxyaBmPtjOy9Q70krgGD/qqXdTt/xuj0Y5/RWjQtbBezA
8oRca+CKxZme4EMrK113f3vhbS/FKQzc4KX7ImKtNzkEcXHUtLdSUHM3tMPfXLsi
suWwHFfYD0BBuYI9KQRmxAaTEqGTSqHCwHGT6nvohzTAaQ9imzObmS3sDnVfx4Lp
EBYeuh0/Ltcydkmelh3KQMYtwyPmgsPvgdtqpgv2qoqJqX6YBq94Ha8ttORsyKTB
XY1ZqZaD25igsHWdh8gglu6Si+XqVx5LAIA4J37zPPsyckgxbvySvpGPZkiM68bl
3UL5k/sgzkIQirzo2xnNNIfeP2chPwg9PxhRnu18faHCuh+SPjIOwxNzw5O/d7fe
JRhfEq0tW94TdNUvxTGcz3SRmXuU2Ybgk5LoNtWGeHoM8kwd2g0JPkMynBGPLpeX
bRJCIGsuWCMprZfrxnvL6LY7FRn/y3tsB39B8Qkv+LSiVrRZ/G4Ut+RnKpXUJrxo
NoRGHiHENjJH/2+9ZVdBWyVgl/yfc8PziHDSnqOcIaPMrayOnQ80eUsZ+iUaVjTD
/DNysdVu/kM6zCx/d5xVrCQtTfr8rZVZzRLr9ZF6RDYqDHzMLOA6Mfei82OlBkRj
zmKFZH+TwDsA0883EjMcWaddhOrnnN7zq9XkdL/6CGOBs6L3vH7j4mWtghFoco85
mWwWN6lLsYCX8BHD0yv9voh7KIu7VSo2O+dM8nil0ygrGfsDeFDT9nxARpyYKGdN
nxTk5MJtl9QDkER3XRKKzpNlwlMCRWepElF6gMmBOzmV5sQkYZqi+NaDGBhqSvMf
DPZbfVVdrjuWt3iNrq+KI3qeeraqooy3YG42jJucZcAcOg81j3pJiC/slzzgYl+v
ZU9/VS4iCTRyqMR59TDeyoIdEVEFs+j64+DtqZ75NJ1DVaSTD9B1oz3XVzIJiZXp
rzUkiDLDs3L3SPQIjdxanc7BV9kkve4pKpBsv1vQWp98REk2guG5JMYGoaGbesqP
YEVdDkEqXw2DBt+vnAvoSnkZux8uzNa5pP9z+VR4gMSTi1QCJ5AzJkThWUzXVr9s
I+3SZoWIG3yFsNH+hQchBpvPJz/QxVzWSeBeJa6FUJK/Vxt6UUNwV7iByu5vnlAC
do9op7BlUQpDZ2hxpPtVaN27T9S1+0O05e5IOfXwQ48+PF/2v0Aki7AeWbAsnSW+
bLeLB7Ta6H5pVPnjPWwVIRYjrbdYt4ART1Ou0LxkVGlzAZHR6oftoDh9+iA6V0mO
aBHhFeqmYOf4zc8NnHOGi2zHpKgPgRBBuLHZj0d4IGznOowUyp8gaF4cBZeveKir
HSpnL9FpqjrUWY2iO5TP3fnevxLvID3CLZ4+VSt21V3egPKNdjbREenfsrUFrH+Z
OS/rSdtvDd5pCKdDu86IdQ/UpTIeUonsk4na8/RYO6KHYVpMyzKKYkx3IiQHQGGG
ukoks6TX8iYc13JAZB+mk05rF7BDuFqrDSkykvaJ7IbrZm2fijcn5TKnplD6ZUmM
ujEMP+bGt3GEUgVMUM55OZQ2lCr7+jsd+awTKmcd7uYiEruHyzSRtaVXVYPfayUi
ZgAT9FCRvLtmEKx3zBCt9WewFnVWRPL+SmKTEMFOxTeikFcVJeiiMgyBgX76Vz2k
k/kb/DK/85NBmiGS7meyIIYtjr+tZ7fqtYlddUYOvHMeEq3/vXRg8TsXkTF6GTxl
/bhpbTxf0K7dZo0wQYfo2PUt64Ssrsd80hIShjCIKVyNHUbJ7383MLgRGOwV+vcR
CxPMrEocCw+wBMqQ4rVd78Y2B7PVU0vOEaMmg2vfHsbI220LQXEkhiY6Rfo2cBdT
TSeMvJLL3aDL/yy6xNCu1T1uusvrI3PPkuCR+Je4toilkAukBjWqeNwUPopeeqQT
UM8DisE9tdeL28z6t7rFG+84I6LOtzvM1yg5IuuhpcoIfr6M8xChe1jJCxLNdQ6g
A5KoAseTf8SpCxiXpEZQxxB7kuEaHzUvggteX4ZyMzaR699zbhGM9brDa7VVtUvM
7RH91vD7SYmSrtN4pyMxrG8NaY9Lf+BBKShCjkJK0n5Fopgn10VR9IrkRQU1qqWj
XFsXQ+H9cfCCuLJs0gA+9QM9Q8CmK5RvsWD0lEy2PpTlo3AlHw1Yw1M+aWuqbtyM
8xINv865olkGUIqJCfoyN1OiCaB9IPe5QG5PmU6IvOl78ULgWwr+IUxBGpRf1il8
HFgOV2yOSB8p2hSrT8FBIzNwRpgtKGR+O2+jNYzmDzd7RRA9TJkg0X8mG4ZdhHSP
KzCxI361rFZ8g7wTMXdlZ9vHaidWdUiTEBvqLMu5RpgrskGmXnuwooUCG3ZVhhu7
JJTxNi2x5OmTSZy3eDXra3e4/xmvF2We03Esg9oDeNYtaTeMQRt4GqBN4Jf6Ocno
qXjllXIy7bVaDwlTi6DXFN62zkkccGKOqzTnE7O2GaA+LguFwZMLEsrzI6u7951u
5rM6iyva0LHWQsGWxxWNnBbvTdnYoSTE+1SlDK40XQvVo/WEJWMRENFvTysmXGSr
+O5kFAqhUumjTdpH/hi23RoP+UeqflD75dxOJitc6D7vLgvX/qD3GlmTw2Wm1D3i
6jYcNqK+E4PZYUDUY3+Jrl1jxLzshq1U+qRpwMA3qZr2GXV4pCBXb/Mqjo/ddD37
ihp31xvhqFYZFSlPa9fxznILVj7j4pVpzLtQRvJeGzACxNkq0gYLP4DyxUF3HGSn
6Y1J7xzeA4TVJLd+aPh2hXTVAYBdFfpg4zQgqcp9HswSm90nQl900+UVyhOnbCjA
yph2pEZrwiJygPgx6Myz9bWjKDreU2Q4j5/p0sDp4d+tQR5TleWKnoRlRqYQeXrX
RXi1q2fxbe4Kxhl9alYksA3CgMatlAGWBWEKqiPmr5DOmdbg2i6z78EEhZa7CWI1
fyTQ2LMWTC6BErbIfpvbYYBq2aqH/nCroCFhjc2q7WMmyTGJ52Me2y+U/dyy47hT
D6hTHvSOiRYc089dindb/rCzLziLX9NKiLS04HlYqvjuaB+i9PsDtQy/i2CEObOo
rSloh5jjsjTmO1Cw2paEhOvOwE6gFi9jhWxOZx3qFCzd3d66jqZ+3fJILTKpfVN0
JyAQYDc/co5k6lwiKPIqkgjj7g1Vc+964z2SDKvmlJJvPK8BFbtIlysBebTh9VL+
g4GJuY1vBaia/cSq1pQirHHxVx99eTbq2nw6C1LpgXu06XO0IcR/rQY+Sq6Lm+nw
hMr7cwJZfMrJk8UQqpqiUpMpMzv20wtchzlr52GueW9w3ufabb8INt9bs4OAIeOG
2PQ54nhuLRF2WbVAX9NbpWSvHeNgEvQY0w+eQmV0Yud/a+JxMu0ApTaB8l7ENNfv
rdHnfcwsv50KiLSDtmOD7rAlg+8YuCTIxzxRHti8xZB7Qm4wT8kUheODpDLi/gl+
w4+Fi9/w5jYmNMov+iwMVekXCh2IaQS2LeX2U7694Z75L6Pu1CbLAslfxUNXjIqw
xTKcktBMWyBzIWoOgZnXrOFd8VHP2OdQ97Cx0hDj5x3sRDN96nOnMOngDxOdfAqt
JP8hBitCc+UzaShW5tYSmU0ybeI1b4NwyKhVb6nvIXTwELnpMIJfnFUdJNyQ89F8
PcrVxMAo+Rdn2FlFXAUr7ttOruLM3+ZILCbn8yb4hwcrvnd8VtEY6RgW0QvqEYYO
5qFFq3kD4srPTDRVZ9prJELRZmnnQpMykp9DQYIJtxRs05EdP9RLq0RCUMvyNOL5
NPZtN6lNNoKtRHe3cEXJZvUbNn3Sr8ethFeAfJcMrYpp+KAwDVhiua2eftpfTtOb
ECqEXG9jQ+IoQdHzKhB4FNBCU2o84DJItrfajVa/ObOHYLk/ZzcUwVXgePwDGZxH
5+Wx8LwitjoUjSbNoqKCB07mJa/mG+yimtF3lBa/HPcDNq94//UuKMCTIfNBCiXH
YafXhYf65H93OijqEMe8tbj8Se/aiX0d0a3GjCxgS/v7KY9RF6Qea0x4ljvN7HCg
ds7QqeroQw64ia9gPIqhzbVO0d3OwnulGsThzOs0KnE1BUh+O1SGURzn31mIfgSJ
FCNYdutz/5hi1UnXLfN+yYefLDR5tiLX0FI3fbzsMjWeo/FZ87rlSCL+yypDxB4D
FbELBrBQd++DbOZPzp+eo0dCYHKhgDYB2s1nPlkABt4kVIPNqgznlmod0eJJxyp5
xbimz0ZYvl9ZWpCqBvQki2wV2e7asa29HhKm7qSx4VdX2HIAABMRjbbSiDwF1SSE
rWL3Ey3osCeQkUBo4XKOdUDwkQaCD7OAxNgQ17ob1nZq+I87kDywvbSl561UCkLK
iKc2MTRXeJnhnmNt9pd+BtyxuwxHYsXX2ziGdnjUrlIJU+2/65WfnGgMUfRyIwcv
++ZhvDfWzL9eMdbKH+GyAspc5NQOjVgjaYjNrDoZujNZ3AiRVkqVEihLdX4qWAo7
wB8P06uXfffBETq0+lFxPfTX82gZKbmflk2gPvb+/GawgfSUWxVGzQcdbscApyh0
L5RuxdwLfqaiTSDjlAYtbN63ms3YT4H1cD82xZJkkJBdZIjZzCPkVH7fowEpXIGf
lptMrURFVNPogJkDPaMPN7pxUnK3ZKMYjx92/i+MbrSEy8n8e8RjjP3l0oHHF6X7
EADViI2ro0Iih3xbrdDQpXC8+G2nEUNd20e+bPWTBV0Hjx9dNLo/KzwuQVfiUcND
QZpfuf/eTsGonyCeuCIrtaoL7rtEbGe4aAY7/UNq89MjFvBZROcoRahn0ubTsHgh
l79JR6cfHMKX1S0Z7k27kR/2YFlG5apRjbFyHFQUqyl5Gwqur/0nchDl+7Fn8jdK
BiL3MB3Qao9YwZ4g45FI4VJiRUHfdNvHKSC3JmLU0dkDIK6zWcWIsZlTSnbeIKn2
EF6SGy0BAg0u7de7XlNgFA/7JeQ7tqtKAPDKgDsoVQCPUQZnIST8X6qPtXNdVDdj
VkvMCNXwC9LMdGQ/2Bttg3nIFQfl9YpnKY2Vl6MbOssYF1B1dzz5emAscyjCmHgA
WlDCLM0er9ehkzgTKUQlUqWAldnMHtnzAAHIpcoKKwucDB/cq9cKtKGjwdGPdtMQ
hP1KCGMGqOOmK1Rjn0wzerCGbAhksLwUneVMKRsRCf1qOqgnAzx5IvYBxC0OTCuL
uJygsV4DjHFywR693qZM2sncGYpYYPuYODHD3YF5nQ6Vzw5tpnJPYG7FCMev3Nxu
Mw+ldqXhFR8HJFIAGmKKDvXQ5TPLvnMjMmiCLYE5c5wT9dFXpPkZuAww6dNULdnK
7/k7WmrW/Z0E+hWEt8Swzij/j3C02N87IQLWoroJMRUAQykarNWXzxAHtchllhMQ
TEhxOWfuZ9VywQ6LOW7rpkbe9PM/CLbVYMCaDO8rQpB2ZXu/byfU8F5Of2xIF96q
L8AAUT4iklNCXTg11Eslp3k80Uttl4cKmII0zhOmaRYnVFJV3h3r0ItlKYGVraaM
DtRJDVBEV7xb3+bf8MwRs9vQaKg0fwdeNHzHl2ScAnS6MCc2XGR7shuymXTc8lCf
FKXW4DvildtKSIYOAWuVThK5ux4qQDKo5PBLLUoKf3KqlkQf2OJwjzWNW0yy6x2+
I4ZwIshxSUTol79lD72gVWvY6AH8TncS4lf+9KxaTtpfhc1MDzVq9XXNONmGfwV1
88ZivqJaastLEYz0Zpy6uTsgRApWjjegQvHMyiUBlflZdYS9senKyR4tLnVGrpIS
/3jUeC1OSun8ZYfIP2DzZNxnlbe2U6SjA9iiyVdiKcCjgRex9+UEtkP7E2V/q6EO
BclBu5DLIzp0of9NWrpHbw8xWsbZg6Z0B70zZCOsbm8yQj2rKCW2oct+dnOM6Q2F
SBo3aEbkfYC/2p5+gM/zSK0n11WULeIUnaOpV6bZZqahlzLBEJJP3K+WM/SpWF5Z
R6wo1hWgUTpbPSShy4VpNepV6BmEIr9wzQoR/KF/HvCREjC6ZnfydE9rm2HkTU2i
RLJk8GQkimhwuSrLC5NgL0zuoJ4keVIz4v3cErT/YkXblZUojIFK8hGoV6lrRS2c
f99pV4xRRBr8egJFEtxi/7s3uS9FfQwsB3sSDaYv+DxSPe6FQK3ov1k14H2gUaEL
FHDp1+QLW2zTsRZ3j7JHYApOsnPnv4HqiXtWnjTc6Au/Cc0/5l+FvaHOqax1FTZ9
aCtH9l5Jvfx4jNa3QqVVnLvxkxm35SaSxkjf9cOW+WlTyOXIgjOmw/MLfJw28Oow
AK7BSDbBKGLnXGL8TczngMtPQ0JKCOx+muxi/j/42YsR5ullADnWbKX49ocwt0PW
JyXBqTWTQYVV05bZGNR9aRBYkaOW4kuBSJ7pe57rZslaGh1UAFwLRIN0iEvJA2QU
FGMXgElun+JyUCzMrM2svNhhBypj/Sxl9MCf95sj/6uoWwdslpQ/v+c5xOtnAlys
vZ83qF3nJGIhFWi8weTTHvMA0ue3egi224UuQkSY/URvC4SaixQBfPXYr8SMAFfp
ldkR34bNefX012Rky6K+DPi5UTDjzo/GtFosWIfKvAlgU+DzQf2BVqVK4vt9K/OS
v0JZynEoz6nMPkgywdjvT/HDaWOH0SsY8fJLwEf/Lgi2E1Ls0Ld+HIxMy/OVsi1r
+HN8zYYl3GwKSSZ3KxmELoX1of92/uv2QavjUmVX/584LkOG+R73mSx1ngY5/cbN
SXGf/V5U4Tvdx+ztvbjigCPYNWeuNqOpVG8FIv2ZXXJeDsPmdQpHvVMTBl3EQJXD
koV+aPjF1U+raHWao/cgtEtDN4lANpzpQjtQEtPcP1+OXjN5/F7yBeap5Xx7A8+W
hggfwrGLklMO/CZZpe3s4lLurM0VJ7VHooKXluvs9JUKCnPBur2ZlkjtCd21yBL2
p+VEGBclrewVtiOkdT1F56Iqk97e+vrXIkpfuP7+j4InjwRvtaACSFW3Gcz+jcYk
UZediwnljCT7PkU+g5zcCsQaY5h1d9YN3/K9kuv5aFn+yaHjj5xHW7J/HXP3GSzB
v+Ot9wJ8SWf4h9J+JYyIDH4htBgBlNeXhU/apauFJaqpD5F6KCe5tbuRCxFitrXo
A2ybs01+FJeIqcWvU4cATEluNh7ATX3tft3PrXcaJkh2CAs9nRPXCHmOdn9tB7kJ
rhf8CFOa7wKEVLSsZswb8T5GNFVQb7ZeSbGwR4BLGdWYvWcYXiHU6dXbwj/S+21b
mIZ9c3RSGPubrInvnoLgO5k5gNoCegQ6QRWYKR7XG9xgTFc7jY1Fdo1knzhEn+/r
veMnD115asElcj2LETnc6Hahpgv/820WaIrn1vDxT2zHn8ci9Ja1q2sby95hqYPr
vxI321esMQwMhRi60k7VTkx+K5Z9vLSpKDhPmO9+YsWXlJvIVfLhRRUHeUmXADG+
+kS6Jzum4QELqbs9guuITVoTiFNKVXcz+cHYbt/N+BopnEgy6EzPfc1mRR5q7Euz
XMqm5zll466L91A/mxUUAzUK84WEJN1MCAeXadHcCCb5QHoXnLZCqVBejoxtaph3
CmcJuz5KlvaB5HRlByIzL+mTdAYBNvfpbKyjGy+kniWFjTD14CoCmBdXAC7q3DhR
YRTh5e6YXC5JqIcfO56MWW+kHLjgAMHiiX2/Vf0lOkL3Pbt7U4+gtlle3BDYkG5N
4JHO2lok9dEJd6W9Jh5BAPPPEbIgxNg2LqpDHzcIvVPKgZqrBzn2VreE0s4Ceuyv
Z92dWo9zkLfPZDedcI4wt1fTh0makCHsn1ZqZ77rYA4w9rt56X+5Ei9ZV8GEX39R
3M6vf1A4IfesyrxxGecYtcBRRudZ66WN/WT3tQBtgh1h1rxx5GnqtvKua9p527Yi
nMRUNrZEFMF4ss3tyo98JX1S8JKNwf+u1YBo7QoY/B6lIiNyjKRKH3Z+aIZoF5x3
fcZM/olKBQEquZD8S5vWhRWLUjnU+D31JG28B6IaKurutU21jKdf5ENes203vhmc
dkVEpFHK5dPBtCIVwQy2jnYM+wuc3P3pLTIdUTnt5n6I277TyZnGUlWA8NQp65lK
J8/ajigN8s46KzxPfiCVwb3YUj/kJswaGZ8n+H+pUmKuD8DFe4AYcoHBFh+Pzrwn
y/qfcEffmO/tTlVmgfbnUJ/GOyaHGQYhyiiLZQVEwhd/0qp7EoNtKlOFNduOK5FR
LzsetzbujnTg+wFPnEQY+oNowNv71wLwMxenSLDS6MXeDchST9tmOwrcNlAD+g01
UKmXJTnvWP6U+1IcVs2Pw+2ZMjtS8YLidx1l9jr6i0RnRGqUq90qZxvYy4zPGEMY
QK9hE7kCv9Emm7nL4d+OzIr7bAxHOy2dOYN3E3LlmU1Oz2mqj7SEZYci1LEdjQNS
7gjbud4gEkqM2qu5rHS1UQMvk46/FRWE7d07xk4io4OjVT1QFwMhCUp/is35WAnl
16PFqN4nHuTH2NlvngSyieghYXiXBu9SGZXswzVCOIcMuK9TvFnr4TsNsrHk6cDZ
uSJlv86SdS/4HwZs8m1lT2BmBaybRbl0sS4aegtY6b86NWFxMUkmB6+es4UsbEHQ
uC2yT2ID+X0GkgaGeV1D6MwYcq9DmxH3zHW0gftXc0+5FE/nIPD4sTCLhpu1pDbB
SC7jNq0NDmb0SNbv+q1KGbQJywkFwutzpjfsmmZNveyDP17wat8UdaPPcXNvlZFY
Ws+yD5ENak0ozTqQetIkiJvSQxKTG37mGG0LAVjI1E+A9p6Tyjz8R/w3oI0D64v9
Iny9//qdpiLmrOzS4Acvh8lDusHYr0FknbGGoXNSrHjqnb+R0IMLdBDv8Rwif/9E
2jU5ffuDt8Iw5h1TK/908ZfG4zSv+ar3P1LwXUykMUpCgJ+lcPkK75ruU3A+XZIF
biH7+a6OHlrqdD0bfZnjMdWLE8+Tb74l5ZxSxtQGHAArfD7VfnB8wmfmnU8m3e8F
2GINwtWYmSUJCTbt6l0DyjRozWVUJ1BzePjeHQ04EZplIiG9etHACbAVYUMuw3fp
UiABIkPHq+dv8BagnVie1dDo9b85iswGML02PzEdZX+3jQxQEayUEWwDwixX4ouA
Ym9qfHnUSPt23y50YCmVkwqe/pAcyXDoL+aEFZY5L+GeGUBWpjDReAjr/j0SEYVC
nm7K0r0+759fpjFsaLQ1cm1b0+xp00/Am8mrC/ziSFl9IhTN9FkBqtxfvqJ/SZA3
o5Mg3TeMmDbbML0P19hVT+jBaYmDY1k9Uo1GLjBC4IQtHXNwm0gcEr51EQKwHYRy
JOQm34HGPX6V/gAiRmiXhkTUrgvteJawLfCMtETOFWKTC3+CkBjie1OeYAZBj4iy
yEUfvjYnyaX+yUtc6N3l/plWkwvNlTU+p3XPuSLmcXZ9anAv0VTIdbID3V7VFS6H
/UR5uNhz21HegKVK2SmP886QPhdGAnL4YEcKHhUT/kVlGGUhWJlyVuFecDuxqsYU
esUSX5qW6q6qgmFnZDLisBV4+KzP+eqWpAzANfupdqqSeYSY9kocGa5khznQN42U
h2yCwmq5yETE0it97dOM3aVZb031tf4+1AyvHU5QfEXNWmD8+fE6shI6mALYcX/P
g/i8MmZZ6yKwjS9yg7wtvBUICj5jb8hX/EpNvgXR3vmG2sYDGvddd9/4Nozyb5ZL
iVyxADcWpGU7zHPDJzQ6J9kOu8kU/GOh1IzoHsgbegVdgjQ1nvRYsuJ7r63WbbpV
Id5FhqXxwyjJ4mB5JOLRu/wrUDFtiLwaaEe55QFWQr1pbcF6oRiPvlxdkQd9FV6n
JWLWtEvZx484nyi1ROd+qef1S7+G7sEplMvmAZxrrqyX8eD6n0VMtilafCgGmwpm
c5cZPbPsHxUKZTb74qIy5Z27K+Cx6u44xkBilt1C5T+ZwLOvF6H4J8f9NNkf7lPt
+1lWt1YiQgG+xFBre8EF6pzrCT3vhFD1237/t6zbbmzz0Zj9+QVYbkQxknZvW+ZW
7SUdB7jU8irJmjrEKYVb/wLjsDWga733rMXosFAEgIrZHKyWeLz1W/vdAGOzbLHn
zzCfWfm7t/+HZpYnnRXNeh7J36DzuDGUsPcaZ3yg2Y4Pf5/GkKD7bcHAgCVeI+9W
yJyCvzBPoew6mKG0Ib4nP3N66miYxjJd3c9YgI3Md3TmaQoZrWUVJdHx64UT5zag
rm6Tk6z93nj0ueHpcp8xND/VKSj7RqyaDl/oFdtavmZB1FwMJnF6dGlVmBQpFP5G
L8fsgRdrAmDMJ949uZPvar5Km+I0avXZmRwhGDzcVChmxs3H3+MAvQpScT1j1YAE
F63Jt8IbYuO3wUgB78HjKJLxe6bdAKVWiTJqJWAKeOV2EHGcYYFdAktfyXi2K8BZ
1uvoXhynH/fndTNx8pqwZEUZEJuzyLU7SHaz78OmnxHoKq7iKhBvYyL8LxtocMIt
+SMLlUq378RpdmYIuO4yKNJJWDmWjr9BbsUSw3O1WCc7UL6h0uB3p4uCMAu+ZSY4
IaRztSOJwBkqTW0aqg2w/x1VdYnAhxE1HxL45xwh9cuVyKJl8KzskqjlsFl4HnOw
FREDUEogL3jwaa1K5XzuzvBbDCdvfv/CCTDbEllyCPsHy5/ih5vOZ2dCMAOUJawj
PhbwX0XfPH3Jt1mIpoel6IQ1Swp5WLdlOMT9Zc9qobUhLuxNsfhKtWzUy3lWCEbn
LKweWWfptxMHBBpbm5g2//XBkqA8YcpujtyzU9lJ8EQRxkw7W0SGRSVgKCs1OTK7
jbvU8LmX45nqPP6ZWIi1IIwmhrdYoCC7FC9zYfC2PoDXVH2f1AXGiqD9S/+CsQfP
7MEZ6qTmQPDwQs+JlYmCu8ZClkCEOsqu9bi4voR6Djp9bvGx0wJDYn7a/mrluzrF
toq5/tw6VYQ7cEuN+kroE5PduF1mZJZ+T5uzs/oR5xhOZQDurX/8yd6XZuVdM648
mpFnRlc5FX7//ste3fiz8MsFo6juDe3WVeD1tbp2GAv1yr63l+UHcReY4iEFWmf4
eaRYioDL/KsSDnFHCeYcSMMZjBh3NgWscatnOflhgtSYnqzQL11JKlaVUsPmUdJo
sx74cpmxojFZBWqU+0gZfUx9k8j+VCLdmP5rM0j0/x45TSXEKmCWBrnR8MYYrclY
C6iC6wvR2t3gt9w+Jq+TjN/n5J28WOAMNleJLhgIFCwaJigvsv18KDxfha3yMjy3
3vLn6nqr4nbWDcTdJ5zZbV7OY2qIb+tFzWgdL4XWp1x6o37adU1Uv1nT6FCGvW+Z
Vtk/EsVlZHNWny3eMb2gGn47d2ta3XrKy3YB7ssr25QPCIfEQX2o5zyGn9rqLcAV
1ZIV56omuIQ8Reai5AjTUC7Nqw2Ahc67atmvp61esi9D41F6C+Q8MVnjarpN/zqO
Po75sINPt1ZUZnxaMsirESws86rf0GUuljTVZe5fqsc+bgG3Hj3HDYR5bn8iXSdA
eURDviXn/anoMO8er1gTHBAgdMXfigcPrHj6wyj4ffi6IhX00/y8601BD/eu0XVC
DQGWGtqzxIpOZSQrLxRJZajV4As6Zqm3wuR0+07d23NQ51gHPqpOeDvn4bLXIFBT
Ud/zoGCMZdf6g1C+9oXXset45MFprDDgo7PwbuZ6EULmaJBctuU0cN+EjNAk4I1X
C+9+sDpBbqUazvrhsSXhpA1xrE1A0xoZPw0BrnnE4F+UKYVZOsq4jDGgz2Iyy7yj
jCcRNeecdNdT0o1z02Ftqi2XCksktQd2a+LpywN4VNrZzf/3nZYhKX4ocxdnm1hm
MmeD/HlVlH+GE3z08vDzpwHXGuPn0rULU5eHcaWc0+MPM0zvmDnBfNDUrFaNY0B2
xg/PAKU6zyzkawyunSsiOWOgzD98RIc1H2NncR06finqnXW0MbKfx5LhCAOC4vpk
D+9m/qfmcKUeU+BDeMMFqvTjwlZGAVMyGrmcCaS8nJex199YfdxsaHmKio14Yk16
y9eDQeDw9k1eJx0EWar2kiqKuv64B5NChfiOJfTfoHtq7Va+LUeutIlskaqm2iJq
GD5xFPf7wK08w1WY2ekiM4VISfCYzFDbG6ZePzZJUyzP8TYi82n4abuZbiTDcCv4
4atHK2wcLbp9ucCENU51vDbwGBS3g/A9bTLrPh0Vf7WRFAVF9KoElIRoZDlJyhzc
aN96Ry1Uk2Jnzxga+Sdq7j2b6yGeDuTEWP544iRzeNV3r2h1YJ9h07Norny1wJGc
DhXu/qyxddedW2eKTGjDt5WrkDK1SmFAcWjqEie9jc2SWK6rrinWz0ioaBzv/fdM
Ie66pUS/FxWVarXeYDNDmu1vp1hGqT6chYNjiIm8SblPg5xLPeT3asu3AU/wII6c
PsKzd36FeHmb0Tde3U57PKqBWaGVs6P1mi6o8BY731Lzk7NIH11WgtG5e1jLkJSN
g8BCQUENXiwu5dciLcQpfvr7Cm759NoYp32QO1uQJ1V6zBy0cTEHu9Z5J8QcOOuc
/+1BS06LZHqgj+wCiuUisjaa78WYLgqWl1pDVFbuGaDEk/G4AvhUigwnHJL3T5V9
2dLJ7yzqmOJhHymINTkCVPh/m0Pd+As+NXmH7SuwrL93QVCURD2FIbCVuC5htaP2
/QMiY5VQKKImLrn9kUHItrkBLDQsBYfbjBUZNtOMk2O93oMWQKiYnBPkv8rslMN2
Vv+ST1Pe4LFiT3bJSrfFS6JOX9sEaJnZu5udk06skLKAZEBlBDI2ZwX4e/19bjVY
N1B8nbJZD5Dwrr91Vk201F2OV8Iw7iU7AbEEpqYXtqnuVj7vUkqpwiZulnYA+ZUc
a9zHnoL1qtxwBrbi1cQdxZTuPhCka8X1WE2SIaI5EUs=
`protect END_PROTECTED
