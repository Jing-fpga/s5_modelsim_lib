`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
04G28qn/iZlKb0SQynHRJzmJVEktV8LZexs1L7MpcM7yaDTaahhzzu2B4a+/7K2s
i5qE3oJAqF3plVGNOgycnrnjg6cfUEkCC9CZnoG3iT+JFrv4+xHBay1Q7uJuffVa
K/6/FKGaUY2ZT8/Oe3RTANq5hCqu9q9HIyguRDKZZF9c/U3yEf7HnYSlGETNl+PC
fCkctADmu8rTudZXk1sZTMnXBfdvycVRqkmm2QrWzoNxZZor5GEZTbwl07Gl04q1
9RNPoCWTLW2V+e59ABL7jmRA4uxqyH5ilwx6aO105FnFlOn6Uwy2NfsjZtNjx6HI
Pxo2RsoFYXz5+4+e+nyPvCw1LSCaEl/iJoF0lIsek4w1UK62GnPKXWpVdVdng27E
9Dhn5omkFuK3Teunr6Dihy7yL93hpnyn/M8I7i2QqemXEQ7XLl12Yq8DpPgahZ2i
5ZwjRLQ8t3MPpAE35sEZkwoShMf40FcRR5TZiJNW6/lcz4/s4SKY3qNn26ak1iqj
xFltD1abLcRkOGv6yFdJHWh+Dzrp/U3BB5HDwhSL7KaomJJPa7i3o2uEziBHbSKI
7uansoR2KdLXSz3oZCAJYpaFbt1Gd65dmsUw8QkjDjwRL9S01ADXE3aaR8XXBEuG
ugjL3TMgdPlQ6sQZtkFpiL7n4/4YspH46DDsQ8bVn2zsbYmGOtZqYZxoF8og7o2e
Om09LfWUCjSVO+los2R/uw2EkjDj+gzYYderI32uL35t5mWVcH5hTUaj7gfpL42V
3z5gsns/Bp41RH6vLJXP/wY83o0cdcf9lkE2fXIFR23lY39bzpU8bY+0A1Lv+4Wu
n2RV7F0QhDUjmvoX+Qrsok6KP7iSm5sWiYS2V4oAGytUtBjcrJH6kmyv4eJGlq/N
/R26RNwSkFHjOSLn5w6HUTLBhPCZ+lm0EGXQ6tENOkBidNCRy8eK2Yr6pS+5fkaB
Cu89u+SsLqinkMrbI9Iox8GGOoe39ECNhcOV5DYssXjOcp9pfunvjdcO7mLxtOj1
EI4zTQBc4XcB8h+hEE94HB6VQFNjtskgPvHZ7dVZs9rK16X3AA5qbCIAUCkR0bpU
zlgsXPZx3GQDPtBZW0tTiZAXbKCtOuy2rMXbwepeM9xTYev9qXmjMMsA8X3kj5Ja
YT0xr0T0vIJ1TiJmqpACuP1zQSnc2Pr8HsHB/NKVt4u4x4ovs2sO9vwfw3FHI+02
Cd2AKHCESChmMCTGnE+fAYqDRK9nokoX5kP/YrpRzGk=
`protect END_PROTECTED
