`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pYDP9VcwugbCcVTHfIyns+6y/l22KO33PMFc87XuPWAUCIhcAWdYfg189nuj1d33
eDVlXq0/psel8/95T6ji0+iozmV8vVT9xTK1x2wetRLr2E+Pvf60Skl3hkKYB/mH
VnYra/MZm6w+vnJrCNNKCnZk4Fsp6WZ4GgGfUP2LuDXLAEnyzOqKnW47+GQQOy21
AoSEZywQ9aANZS0fYtmzWYbMQNw7aTKrMqjooa3o41ObThDXymXLli1RaL1mEGdT
fPqpGCpZDP+Pvwk8l4zB8WIilVCZopSZY3BWExmQ/ZMWvIU48YYz0RiuXX0aVKie
qnbHivD2V3QcHQ/lVtFhdi3RTICuGRxBQBnosCiP/zVmlyZASI8XsU6ByAyKlzg+
TY/p1AXYZ4bL4SKOmHLpdPw1gQoQFqGqQEQ/eEEd83s4roDXpII7nJZTFdCe3E8U
jzwMyd532Rq1Yy0SmUb1vbPSjQ0yJayboPVEXAtvmT3uFW0kFqEl/WvyjtIOm346
0AxNhEDCxI1ns3FY/9dVAh7kxKkiHjRqBVQ82zCZ1H9c+gTo47NTxk0xP5KVPLcY
8LWAc+9QwnXrLy93/e19dABb1/tl47WTevbukcQbwxOWz3axEJ38jk8RbppyXy1O
5gUOY997nGBoSLze6GOAh2wGq5kusuP9GXTY8gVnZXeNtmhK7Z0LxrY+BJKYWYBZ
SDGA1HTY+dFROEKguArohfoHRpdpM2397i87D+nL09fgVZ8eN7SNXmo2lKFi7fly
wNb48SMWsG/HRBa1NHfdIofzjxVUq1egatWkYWzh5A/W2eJyvubQkEIVLg29NBtC
J146KohZY3LwUbFJPI1p5kreSQtZy/L4CJJT7QX0Z/MKQ6RyUcnfHRAHWhuqUnNt
VLsmCY80ibzuW+qDrAaQhmmEMp5Mw1byJEXpCa7yovsrAQ7Vm/X5NL/NLJMckPUw
wPdjQvTrORSwpQ/5MeGOxvDVs88qNciNdNBbkepacC5bWHMKWgPZexnQePCzONyO
kkGYtjSQPr+cbMxTuQoAEGGW1YhYSGyP8+XvKYQyet1Mnug/Aq3yWh1FgmHr/V+E
OpUbX7ejHyeC7Gf/oVS6//Yg0r/ytzdDUC8+T6Ys7q+7NsuC0FwB3eCumbBQEioI
spU46d7Uxj+CwmiMKEsJjQFMXA+o82h0M/T/dHoRyJ31MERudR2mRlVkxyrMNCsP
wOcZzA94GKO86ws1J6ekIuoVuquovJAdapcKSplpfEDnV3rFeGONJfB4IyNp9kNh
HCciSpRoZEFBXXZx2CzZuUP0Dt7sfPLG4HyPt6PW1aYdcfuMkcE9oGh1WuYJIx0w
RIkUw1I9W0BuctlRy7Evt0iThXP2PksySdiBRNy5gWaKttpDbrqxPlRFKJNNX0SU
IgjGthhgXmZD9FZFqvFcBHWEuix6mn6PLO9G00IJtJXjaI0ELZn4zWuj1WbrDvM+
QTw6dtYxXX/NGTbWisbPzYLVZ0gagbQOFDs2nHfQLK1dLjxeqiwlpnSvtnWngmZH
U6rn5FX3oqwBVBJmGd+sPmlSNloa9SGbXrdFkTQVCXNNu3LztDd8uDqYWjTDp9aP
irkapLXZ2jkhncXVFZ95B4OBxuubhc7oiGnNiIQ7N+Bd+S/27y65XmOcuVwePwD+
/AsGhjbtx8cstp/NMAFmwzMfjYfNgFzirwQUeSfr2iByd9Urhx7s3BdWIFId4m9w
mIpk3cTBkdJDzDtjw7A2dA7YFtd5M68RLAdzwDwsoFKtc8ejTmvk8vXsYA7k1yVu
jHyvhF+WK+YvUktWmU7Ham53k1WYTbMdmfO/K3nx2sdMhnTohcp0K0aVT7aI6pL7
jRkSqYclmsrRD8wYpo5yfeAy37/EjzB1hS7wAGKuO63MZDyDlpLGMpbHYhdxDxCT
ZdzCzxNC/8bNZqJ6riBNzIV5rRi76b/wtADD2VX+bxzLBomydskLNLOEgD49KI4K
mRku0D+ocLuJTqQvQYYezXhtKR/d+7LrfYEmbwfCkCJwAvXwO/hXzY5BLSE4E94K
uNxFdAi3DxmGuunMJwVUD/zE5tWq9FrYochmYRteuLMBou4ma2/cU/eVa5i6kDNi
uELzDNKsg5JXjsqi9SlWFHWW3kIJmtlBE5cls6UpLY/jCwaStGDY5JKnwK7q/Kvm
vYc1UJVXT9TJnowUUQtQYi86xgY/YIaiiYxIx1y0Myso8eLQV2oCs4iAbZyVW7Qm
Bn3fq5y/CFQkj2mvsje84iKii+iKReqcyn5CaIl2ATRMpVuGF/ivv9d3RCP13of2
SUK7+o2TaiknZwp1R0zgd3MD7cEvwPMHZLuCcRd3XbXJueKUqyGk+LEIbNDNOaLl
LAgkdiIbxlw8xgmFNUadv7tyJCB1KLshT2K6lv1GYowrkJLAY+N11impk/Xi6HNO
qbVLSmoSStpc0a8LkYWyVqtjiPHbOznA8mVqRBoEPakuj+LJDq5KH3Ou4APNbABr
5/JkihYLv5H2aw3XE0IWr9VWVueUg6UOxT3BZm+92yJI/DZfuXd2nUR1X9LUbDzG
sFpL48veojEsTC0gDsGNuH7k/YJJL/otu3DaUpkbZR0IDEzBLDZzj4X/MuftDRsi
+t9bHToZRPlSHZ7WyQrp/KOTuTqxefRF1pkUotpcGYB5Xwl5z70Hw2BJH7mbfrS1
adwXbqURv+I2EMvOMJAh+OBFxZQcm2Ffv5auLTR4pbo2L1q4R6knxBpGpFQyfkYa
Y+x89a7ZgXbwdwPlrI73QIZSXD4dDDYzdyBp+TPfdj+7gBVBeVoGGE7NHYtO62rJ
wf6l1i5jJM3DxUKQ1oIeyrEEO8Xdy3uBsHF7XqqxO8+UTeq0IGgR47VqX1Yjy1I3
TgjusbQ2ThIRCiC/jBxtkDqHVfpaFCIg4/viwstxHtedwlraLhdIpQSO68cCPgc2
L4ji8Q87dvQHRKVhNvKDIRRc5hqC0Fn/UbhyB7O8PzBIhLudUUk1O48eAB2OgjuQ
VXztuk+GtJTsegf/zDnEwGjRF3kDtjvaS0T2Lj4QWldqdpTTmMqeP3nVczXJh96P
iMs1wg4CWUIHOROmfYetPqJ6cjwVPkVAZZe5ybCsi2RVLsS7Vevlz1hlU4mpEUg4
T+m4kmD9RVRHbYcIPaDf1eYZndBjo1PoLMX30VAUBAZoEQTXMTyz2MT9gyCiQF4u
wVtXtHIpbuUGBPjXgCv4X96J3TFQz90LWJDy7oYAlX/9P7VgRNwd1rrp7P4fRuBN
iwl34wFhWIPEGPy4KTk8lTf58zBK8ENTK/Nl5oJaBiwstvAg/pdK+3vAfMjzET+X
Ea6z2KoV8PDiCj1sG1o8VnVAaEJ3bbpQPVC7+E2UCiQ=
`protect END_PROTECTED
