`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LFtFNkH28lTxEFribyjzl5Wt0Wkb+ppjfUdelrmSOqua0cjableOkiaVjXnCtqWF
WvMp0U9RJ0TxzMA7nHBZIrg+mLIkL6LkTIanOMqTxGH3tHsTzaMVyY7McT0LsHst
ucAZEbo91LDVgZFOjJuqzahO2/Ku2Ri2uRFcQtELS1VFDy7CTPpeZ3StBOJsGsax
qQvx/aNEV7jpyK59lgspVSLr8d1RHvNh5gtzBMXwb3o9DOycP6Y37ZYqjKU+rv+H
9SKPc2rlI17M3sYi2mF98+Ky1fcfuVlNI1myvhrsdzBGnbz44i3X2b7ruiM7d8n3
yocDMlY8YPvmKfecL4u487o6X3HY2mUK7BMzfiO/HhjQfPcTe+kng5iWba1jF9Lp
9OCn1opw1DDTOpj8u0hSV+Z1qGcqJ6VNKlaMbbSTPOVo//OvkyUGigaDu/X65WeI
bAggq65rCBfNVR0Gcitx0xddzz2OrpYGMTfi9txT0raBFr6AykZjxsV2sY60NPe4
5RvbQ2sgLrEDDR2oI+2VAJvFazQEw9+Q6zrJFPpo+yZkiQDGsOoL1QLhuTUtECTu
Z0d10ItU7TDCjebCn3LMyAo3zjXwjiSahrFuzEwII80obK15CpvbaA3nefFyTQWD
VF+EIzq+NVCtDYbcIhvNjGJCtaEJGKNtXWHD8faooqOqaIueAYbFc35Ozp18D1g7
jiO9cPaKonQQBFVzQsPErvA3qURmrXj4XVOyeFy/16MA8ZUYxAk30bUE1U8AhMMH
bgdW9DSyYtvsJqMuBKalxFQlRd8QL31fHjlzoyOqJC340zBksQlFZX8CcOrp2A4N
vHjJHdUmvOqgn5v257PwADB1aqz1ialYHcSv+sqThq+VNTgf+pQSIdhTqcOehE0w
nQhObCQ+0Vuh0xZscW8EIxAsTGeul9xlZaUvJCMPIIypDWSJGf8Fkukq48rRf7fh
lde/yA780kptPSF/+d3ZmiuXcZTyB0KS16iJG8YNvZbZsUapfhl1EO4MINPc1cRw
mSc4llFZBIeL8+z0OpGp6M1vd5zrzfTxBeBonZ7/bmMF9Pe4z6adg9w087XKR4EJ
yK4WViOXHlzhXMVgK3mybkk+yQJZqnXoc3/qUmhOVsc2mHRdYZ+9sQ6kRLR5M8jt
9K4gz5sS+IuacYfuyExoBkE1Dcslb8kCEcsBNHkRkAN+ULUFN20aSc3SWR6C94/H
mbu4IzcsyltshuNmVorvWcoeQOI/1BKPWPslDcDU/Y2deJsJBJ8oy/ZUmToWGyaF
lvSvqWjVydfZI2U+Dt+vfZTaj7uIZpFwD2SRKifSU3VGddopyBkDa32b+fspC1qc
WgFqg42V3ftmgM09BO3s+fHG8qzn/tresSzrJPSscuFIMa8r3SuKN0/O8Do1t8fd
O60spG4XoQBSSNMMWnt3ZK3kp2tXifeBS+3riv2SH5/B45i6jCS5aqLlvgtDzKZI
BuUCNkbglnrMhuXfsirSZRAyfzoWqU9nSytBCMu60vxEuxSZFllH5UkpJ59dVEQg
OEysnejqw2rztzs7O2MZHA==
`protect END_PROTECTED
