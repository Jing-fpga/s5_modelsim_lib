`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cvz693TxmNCYCc9GsrottP4V7SKymjK65gFUqubVe8Rg69eGfy7ZlSJYwxKYc90c
aRpEnOXT3bIaIwB+P4nWcYFVeYy4lkD6BYf1r39pnDoA60lXBo69lJKokvbsQWf/
No7IzYeqiGk0lksD16436chH8Sorknsytpa4lQmfrPwAwwAAxdlQHxe2CtKg4WAR
7ZueUx0yILrWuueUlH4wo1rN61SAbE9U+haUG50fYm6iHLVKvW9Sh21Lyj+o3yFT
//XciUM9C/Z00OGlvuklPJNVAu0CEcVtn+Id/TuyQ6lMG0qvC1wS7HS4/FPxzf/z
HdLnpQr4RNac0EuyrnzpmcGsuwuGDGsv98t/AdZSGa/JHyQZNwNGGsV6GAtiLThE
qi8AvJowCdbbaD8RmQxrNNZ1Nvmy5jwgUdIzjuroIhbZJ/xN4G0ESQaF8c8kVA2g
5l6pUxxLKN2D4BcNtm4W4ZQ3bluoDz9tB7jCM8nAxPKeghQP0yjvlh4/5HcD/5pM
98Vbo6hJgrzWPnKhwT3jl8g5JdCNxNPGHUkmW5qvJ1nvixU+/OOVpYyWgHLnaWSq
Jxo36WlRAV2FeTWB4qi43EezrhVzp/Ej4BR+5PJ7o1CSC2TudBvlvnV4FLA6LQPW
8cRmN5T4IcFARJk/a6b21enHzXNzz+QIWTuJQMNQCLkAr+tM4baOBhamtZmGt6fq
qlqYlBhGPeKohAxlaAiTvY1cpdlA+JucOS2hzJ0ejHY/0lyukhGHQGL5zHZXOukj
zlg8k9hhoQfyEwaHGtzpfZunfZTb1HQFE65JcrW/Mmo=
`protect END_PROTECTED
