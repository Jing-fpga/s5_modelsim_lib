`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F995vDOCvmBFL5TRNykFQoyAgNH/RBuqNlvxnXJ1grYJLajqjDD3atea1ugEsNYs
mTGyhr6eydeH6h4wvD1ULsoFqE77zFLxXeLdRrhNqe3qB+2kOdqRF0k77baXTInk
ByJBhCewiBvezIU8dqcuWQWq7eFwqGbSmJRcHcFXRnvzlRy+rpnvE6w9zOOibJv0
4rf+g9RcAr6Oyj3Or2FZogbDzwaTaiczUG8AkVRGwaKiDgWS1NcMR3dlLAOrYIT7
stRiV0Sj/BVcIi4R86BQj5chgTvVqL8BS1Oxa62KlNOxYtbH4Oi9P41XvruGl/Go
YtEJ2bG8Kc6I7/aVJAv7UR4c+NMHmMCujlDuRCXqK0s+thOf2OfWyjkfMXQNWNBG
74FDPAu+5pNnkytl8hC/F+7wMwzODZpPcLNddnX6Rkcrkk5FGItFILAIGfqoFwjx
2M7PNy8YG9TCLP7ht1DpprTlI9ax5HGpk6hubklibJWfFII5qcshRJVNXi1uDPLB
saj2JNWRAxVr9y0C2Z4+pZ9c8LoTsZVHwOya94B1OiM/fQqgvTj/mZoBL6lASmqa
T0/NvxdG3CHnQULctRgpGAv5TboqJoqvNQwSZoMNozRRbtKfpD+e0AyveO4CQETt
4iJfeQOriG4cxi1DTOmSNf2k1IycklNYuMWT+cNrTnrb6bA1BjSL5wj3FhxjwDB1
11N4H40r002ZuwrCnz98AD/+Kkaz/3YNp5dkzAv7tAbBD//9YwYFDsS34tJpz7QT
zu0y/g3H/5p4SPt/Vuxw1ikf5pHPcIUktIOmdIq4KQu6oaJSgOcFBKkytoKBGdTr
gGHzDJE9whxUHjy538FDnxAvEqsfiq2dGJZk/Uu7Du6bnLuggFdWoehtBLu8T2AQ
tuON/onabwiYb6Ndm7UShQ2ZqwDwRhcoXgNVLHjMjEUJT63eg6YXzMNBYkthWmFd
tfKb8Ep17TbAPUFd8SQ4bRkBC0MJQbW38sgjPgHbeoQgdrSag2xIAAxqSMdJ0nce
553/JGOyfqH/pK6kYF8HmGvoTYtvo3VNk7WbxNeRNVj7ILfKPyk0yYp4OQc81SAu
9cdvwDtEz4SAt1qYoadlHgp7tPL2l66Iqw6CthLlN9r5Y59cdCWRggw/6trqpXr7
yNe3WhRchS1G2MYNLDfo/WU8UsLzhmKXNrLWUEzECEJMIrBi340C2H3pjN4RjbD/
7PRy88qKWNxLuU2DhvXuzk4VyUWGn4gio1ijgd1xA0ZfdEdxKxVhf4xOJe3rL/C7
poUbYgVTgHv+Mj2TdiLdIjmVExjMfzcz9HetpBhDlBU2ysEEkblEESsZ3gcAefRR
uzQQFczlOcMxRophJjCW5lUq8F+0L//AFIouzyaEyWv7l4/6Z4pq2he9MS4MO+yu
DL3q94AIX4UHQqSvlj6onLH0HD1jeIZZMSwvz62mQLRiDawqIHg/MJayIPdwwsOM
2kYpl0y4jK87a7O7ZNBJWQ8TtEb6ZQOEZGoAjmJzf6fqXrUuoAWaBInSHACvZFVg
B32HezbTKYbzFbOA0WWyYQfmIolnJb3vcX1jEHa4/d/CcX1dhsmkImrbOLq3vxVZ
IobDvZO/0QFoO2O55EZiZAlLsPks2naCDp+KJBlHexvQMniLXOpxjubWK7F5Rpni
s79NgpCucOM9nzXlgt0fiVxYi2IaSFtxyhcSH/rQQOUWHCwLrUOIOIDne6hRzg/H
Hj4uF2QX5FeUPmo2N7zUt6bSHqtrAfgYAQD4ezSLk/e7mFA1pqpKzmLwbTBQgnXR
3QvWlDPSzBIP3mTXkT7RNxSHKhC9MxwVftZJ0KIFWAkXoNRkmb2kBKt8sxmX5krf
NzYSHiunTA5IeahvRGnjd8wkBSZvc/6+7+y2fTPmxG3lWISzoSzbger3U9wkhD+y
CKB564FGeDWukazi4fvckaji7iMtQHXtU/gnmsC22104SW5D11882+EshvHC6B+o
v+a+g9N0MtGU7Jx1tBy7ssEN2sZka28sVhSG5Cb5ZeRf3qd/cgzCZ6F9qcjfodE5
Gcd/g/mtsAOAUWVAWucdOjCmaSTZCbPEnzNsnzbnlTG26FE2KGt2szUdNXdJCwVp
vj37HzGWSdezMUmiSbfMHRYK/1K7wgEgyLmL5v9qUXRmj7AKlZyreIuNbtPFc8XS
5dnV/eU9z4wCyKhR26cxFFEBCUD4HBhpWVHsZ4XeIR1BoJ+asFoJITW/rdWZu/8Q
fTnn4ZwE+gIbK1AO/8+MZ9PCWBekptFAXRo3Tcr521C4ukTJCP7Tl7GyXVZeZ822
vILxM/LBgME/T8pzE+UW1WPqTKpUoXgDwo1tl1aFIiMEEJewgTWSO63suFQaEFY5
osYDuIalaSKsDQO/0/ktc8Avj9CHUq8zMph4x4bkZsX3VEP7i6cUwl7EzeSDLQH1
CCU2lj0bj4RsSd4L0lcb/lJ0oVLCyspoJ8iWUuj1cN5l18CBKyBzOhR/ojc+upiC
0tacX6lrZzH1qymdKES71UBzISVfNLs3KIbu55LJd8kEXDGKa2lsIGLeT554GIW7
B8zxSqyCfZUTY2bJaACmkyIG6moOhzjfZhWrqStEMqipppa7hfE8P7tpkTtEsw4Q
BALKqrVBilm3zSqlCy0zNBOi8xImpMmniHGcD8Iazz2aWSyHjKhHpWI816zF/5QA
nSoEzOJhtitkH0IMyrh6L8IarK3KcEwEkzF5KgwmDIX8yXWG+Dm3ceL1lInkcU0N
U0HHxBzDPERIpnPZ7Fo5d9x8z1iQqnWBSRY/rnsN3nPkY+XRiAyaLtdlXMJtZX3Y
nGtUGzwexdg5a0Y4El7qcIAFHFnVPAHW2gRFdcolESw0jNYMjS6aeHYt6nHYLZpi
CQtYQXAj9yoZwCjqGSQxV6V19femJKWHEerXKneN/AzkLXT8W6fMjHvvc0+cTzzr
ZvLQJ1+XDbhPV2g+EasdQ0shBTik7uSeyMYv0j80gABC86ycvIhsEb/zTCdZUmnW
LkFzrQj4tTnbfpMDM4fgWyzFLDIqME5oKiRTHhAdoHyjkbxwbcWh/Z4BWmS2sl37
FGAaceCB0FXWXTSXXL5Ao1cUMGDKPSjN6uaINFxeSQZeHSBj5nOxJ/eeJESEyKQC
bN8cz8QIrRz0pBQIHo9b+px38k6YVu/+c+lHsw3/RV064cdg6+Gj4cjfVeJvi7B9
+xJM3w07gMD2AkzAcNdbYsSfxURiinCllmvCkdfv2hc+JhS8hc76XuRfyehJgSRl
NaPRf1QNjdWP1K26yPvqgqCr1sOTGKL+ac6noJBrGlrzSRGO1ha9oxGGYC/3u0lC
MPIdake8p87i9cHHic1m96PaNkUX/01TJWBKnDdvm12ZkUVTJnK+YHR7E6Ou6nx/
zSNRFoFM7/QMQTXiiKiBG0ZLEHMbSaiVXpxN9pfSYjxAUW3/aknxjXK22AFX+GA2
GK2JQonhY1H80n6KzLTNXtH6+o2H/cFB5XytNzxGRGXY0UDcgvMdFFj1cqOQR5Mr
N0FmgngLM50CCbc1U4zT8uEZAmKY1mF+lNbey39KD/FhwGVZQ/JRBbpWZZQWB/3H
WpVRbAwZ3E4foWvXHgkDmFxZVQrqHR8Oi41LmQ1zSDSLNcZkU3WLRUu2TalxCkYq
SJisWS9CWhg8v/PCP/fP9Fqs0vYdUXV3kkiIfS1slVNNB/S7gnm6yENOpc82qokP
OXg3HvrCHMU70e9SRkKqed8AnynWme8EDMRIozUq36bRh3jq+kixi6l23n1B114J
mhBJvtQW8YnguJ4dEDtmP2Nt41NVLLKxI1SVm80EoGJiM6GqAqAUTsidaqYdDZh5
INFgHBFVnk+hthXpFP1F+nON+2WhM2lzVCH6lMfotkj8zCgE1p6b6HEPlm7esq3N
j9XxgFD467BnrEx3PX+8kQdm+4T8290NPyzQ/KEGGGmTfjIKnly0ztABxMriCO/a
cAAMPtyufZ9ejad2KKKN6X0GES/M3qfN8oUXQS1LLsUkk0bLU8lg92AesSU3VNK/
DWJm6ktmrGyRTNB5k/gxRBCbHBRacsg1nyh3wChH98D8HNtWNE2siGU6KNyZVIIS
655p2PzDrsVqtjsZEbi1dEdsGJMrXcKxGTKu6LLsipKbDHJbHswZWz/im2HPkvEL
tRB+dWdQBUt/uXRpJUqRr/c0EqWITLUeYQDgPszJTjxrOrsksszxnd/ccjF/7r23
5Ngs1iAHV4aRaUGSnKuX4EFWXrmo8+n9iyhDhLdQxxFqbfQ9Tys/Nfe4Y5N1VukN
`protect END_PROTECTED
