`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qkAXD5FY7Lw62/FYwcDqw36bTCY8KyDhIi87IcPw670uaS+B9Pco06FG4lnkt48X
PJ+h1AAvvyyd/mk6UwI6xsXQQj6g1liCTiDRHCtXlenjKp1O/AXFCYE7u8i9IjNA
R921adJxZCts4zQnJF6iIWV74fdqy4abwg/Em8ktIo8wy/vY7pMdHqOBIUz0ck5K
N0VzQWJS5fONu03xJQuDkfBOEMHjA+NWKcVStOr6E7vE9/7P6ZU/2kCOLTQQeIGw
BH5s0ISFD5Z2TyHr/VGidXTwRI/jX6iokOapIvZWctzp4LalltVpDVSb7jXwsI5o
Zz+fRALkuqgyk3/V0d3y5fTbVB736xfDjPz9YdqM2E23KsOpGPvxhSXpPQD7kvxB
VarG/I3X1yIZOZVfd7JxksCseAnsSMZnmEklahn3iw6yie4KyiyP+DxCjcnH4x9D
v9w7TQZ9URrrkYC0ufLMCmj0LAuZXwMyfibH9BaH7qy7feUn0Gba2H4WkoW30mK3
MNqF9nQsGUC6SwQPRvFV9uYWn/setZJOIoNfgI44/RqPoDFpRkAZkGF9j4qt1TDd
0d0OWXLL9IyTwzOUQHczP45+msSrZ93/bE1RRfkpIf8U/+4qrNY60pqZOQBFjHH6
a/TBVLjrcvkI06i034JgLh4XdJpndR9vNHPCm+G5SEk//btwJWGV/OJ6RtfGwKho
pqdrlAdxGjcq1kqgJcb0R85g1D+37kEaqQSBylqTrLla0ly0tQEnpSmnfiGFkZmR
wPQwyEr5NV3JyEsvyF7CA8PVZ984nuESrT0YT/PkUiz9FfxIitNzCj+ASD8Uq66Q
bO4jxWFHv+vaE2I+2NnF0kshNCQPHAAgqR/zOCTHO8SxuzEhwEeZgCupXjmuzvXm
LAAP+9QUkXe2VZJRHHJu9tRHcL32V3iwhbHIGOn+6o8d2oicUcbrRjqkzZ31kiTa
3zyWBqFFwVyNzJfeZgRHXaSjeo6z153pfx+30PQVuPcpoDnJITYVlX7wALH9nQs5
7isrLUnFY7oWrXW6RdRUp7Lh8ULsXXdUsC9BpexQ4dQxo6paNGpvuMy4Vr1E8asg
ElVsY2ZnIVMhr00ZcjEprodG20CNbi5Z1fK5pg5yZxBTO9u4EMqJQHdYNfBSvXaT
mtrP7JmzPV48LGRFrCRcEaBXNXD01DtfaKXjB5O3jaIwUV+Q762/JwyeYeyn8NLr
QBda1x7W5J/qmaOhmepd9Ceu7VcokXcBNzH9uCrt83EpOmdXH+SZufMuirpM57ue
pM31+lBtteh43nYfvBswPQ==
`protect END_PROTECTED
