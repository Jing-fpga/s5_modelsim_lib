`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZrYWlPmaWSlGmxs++y1NUa8kBD8EpgxtqkL4Wmd1c3YB8cfIDD6/PpF45VP3Qle0
AR8/wT2jYFx36YoFgWcQ0xFTdatCo3CL7D7ZPRZC4yNsc7JpuCwtoQstuTvOPTCy
CZdsyKlhF/hpIWyz4VZ6ixM9x0ItIFwvYs4D4p8ynOGppzpJ026DiARh7cD4T/Ia
JpcNsxBRd3+f7zrrcrtg+Z48ZpG2wEmlfhh511vazzthhDmNVm2sR97dMUcSiRCu
Gvu6ZoBEalW0EAtT72Yqn3Vbxjjs42oLqsZYRFurD3fAc1DlOq4SwIP+Xdo4Le1B
9PhP4OAZcGOqo0I3+Nhqf4Re0j3nAdxikl5r5PycxUm65KQ50W4sukMRSlHbEH56
Z/1UDah4Yduw4mBHRvtHoG9O+63YNvrbryXcnpaycu6PuGKlb6ob8zCKv3x7c4QJ
TWrmvG6k6W8h9gLbWRW9RlVzs+2ejRiBujFlndgjHfuzK3aAmtS8ar3NvsJZbq0V
X9I0vIBoFIohOdIdnAJMAnqNxqM9NdE25sKGCuWC8mVQQ5qze9PN1Q74//bu8iLk
lNRI1fXldJI8rd2yI9l3esXV3LSipXGBpw8nflh35vFc4zMcIiUkEawttZECdisK
W8vziwA2ApFyS3llC3OswF1c8HlkCRa+0xXToyMYJPukbw8CuD2nphvMNw3nVD62
Xniu+weaUfosQ/VZQ4qerAuq9xR4t8z2bncFo3pp6T3Kws67IiERz+BDNAoxNmlK
5Hf/vrUNZPQEwCVaYrzH9lLAGF7I9/vR0uIMJtX6n2yrzb8+SQ3xFezMtvYbgC1X
dv+5PLhK+TaWZCez2xPgWB9AbgxR2dzg8dRn+7cXl0ob1GWOKztrTh5wv7MZg4ij
sFEaFmGy8eGipjVXvJLuFTJrZ/9XBvSboQKwRQRDKgm1+Awervs/2uer3y8oEkgl
zqnyc74kYmsFsKIWoycRlcgGsAwbDsyu00VGvgzgbJZa6sZMgB3ISJCg8P+4MiN4
mb7Mk0AZE4ym+mcEl7bZNfrGW57ZbMwa2s4I1mPduXfvyRjPjQTvEyOvLdBWXKrd
rcim4Ayc6/LDrB0jAX7g8kdxsbnWVBUqURA+gFaAsx0ENEBdLKUgAimWatVczOhM
b8mHgShptU1eOkPT5oOxdcltDeL95jzTP2TwCKV3+oqwxU+Fvj2qXNW9VqRdBUPY
/3C5tbEY8pHOdonNTyao0vOvMouJK77w9c3FxtUTFin9rd+zcXRLbnujMpu56IpP
`protect END_PROTECTED
