`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mPan/Rmbh8M6G1NP/JVwLwL42pN5vNeq82QO25v0OXJHGG8sDr4BgbqreihVEfYV
HKgZdZ6TrEJzf5rbS/AJCpKPVCOG5GyOkQCQPHkJDPcqrYWaosvx/FCD2ZLAxLLW
CzNkYnlFdBXJsr7e6CWfvuu5Xw4Xbiq6WhaOJsYtPTIPshL53633PhNPsVip4KG7
l18jl8nyj1kaO6+fEGsXA+U/rz25sGuuvuaVUoqxNWOGJ0mhZ1x6mGhjDHpkRolg
eC0utbKVXb+d/t3/J481SE+okhLdO6SzYyMTctBUCeNZapQfZMD34vcFegi1ONnH
UIwGJGCLwQ528REDEsGN2SywhFlLY6qdmeokkOItyOQKHK+qX5VCBWIXwyLU3Pgp
okmPnYdfEk+dS3PzflzVg69vlgplhaGUbCpdOpv8YwBqmFZHPEkkzwlif7wpu3a+
dOoWU7zEI88hRI8fSU1NbAVxXkPNVvWLMM6ZK02z8rOj0RuS6ZWXNDSYpJZsWWsx
olCU4qWl+2z2ssmxVK2hyRAjDAJJvzJcXRWLVy7lm15pj/6yZbZUYe2mtKP4GlB4
sCZPhbMzxOmg6eHXhSzMPYKbgMint4tYH4PVEAL/uJicmugdFp5wdEUByNhrRxR5
ajBRKuv8I5BXY4ndBX9d0l5uaPPBF1m3ilpnWA6SnNbsi3AjcluTWPK6eC7l8Qsd
`protect END_PROTECTED
