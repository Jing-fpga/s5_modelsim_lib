`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QOdgCWDtDMaCqA3qOACCq73uiFGg6yufVq8+IOSPKOVZVgCHvUnM+xGapeRnONm/
Cpj4iWFiliIIduaEMKRwB4dflyUk6BzvTTYffCoy/sRzOML/QsjDeL0GSbXcqTP5
nJU7KkYaAOK0hpCAi5jgsOmaQ/A/svSwHgReISXuf6Xwi7mBkA8FOShsGVdp6K+G
LuEG8FnDXnXYFBS6U3eszprTbfRLfZ/euwm8S0KHPVtQ78Kky5pjs1HDlByNiIgK
Z+9eYJbQlzsGEolAvPzlMh0jIQ+X7RvRV5VPeQE0an0+MgAKZOAw8duILwDkatpY
nplZ1aR4qfHjR6gFAE0ZHG9/r+YmsDeX3ZuQSxZXh9F0Og+4kG1qXhY+iB1vt3jE
FLr0FgSHiSdvrH7Lm+Ib5jNsGw8Q06Xw8Q8zqJ93Ecr1rMcwdFxLk285W6GDEdh4
LqOoxssbdQFxfIAQLTeuKbE69kfA4ELI2TBEPzAuGItbo7RrqvcGRGuUhBw4X7Vv
Y5H0BaI7dSRDYDHZdMg9grmDPGg8jFRLHr3azMf7OJ4=
`protect END_PROTECTED
