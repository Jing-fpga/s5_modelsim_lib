`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JeRw32/oS8ihbIJMH4ygaZei4r7OcJogY0HzJsEsQJmpw7oUw5ukOfdbLWq9MjOV
anz6joKa2hffYtqOaSMvf5v2QcHe5cjt9sTiLrrpS593czqa2hsWL5Eb/z/woBcy
rP/adAv6LJ65pX4NRHsdHoz6lHwoFOL9vLgQA7yo7UHz1Up88cDsouOz3Ia9udnU
jJw7G3NDYDm1KieF2mlcYjxFe2q89IbI+BaDV4RX3scvecvYTu7N7A09uur6svKw
7fP5U3RJ5RtdUtaflOR1BcL3hxMs4yjtyZ+RhuzuLLO7Oemh34BqWwqqPc0Nr9hp
pPKmtbWsNcEcZ1KcJxtKaIJDUdJuLNAbasrcqcsYAYIfROcmdVfSRhn7Ce9TG1HS
z5osM2SXYC/eZb7HMTdVBfGPkhNSh8HsaiS+r7P42mCt6i+wbYObIwv951AZsmGB
dvVT0vfVfMuy0OznrCuoMFhQFHcZQI6SExrx31b3w0mAUV2QOzhMR+5ZnPMHpSr5
fRRv/sWXDbjaO2IBDWd9XGpMeUSRuyVndAQ3a3OksToZg383yFudvqREaThOk5hx
pYT0sSQ21Ac3tRNKY8nnlgfD6vgHcrZ8aZYAwtwWS19pu21W7930F7APD5O1aZBN
ZGQ+GDMSqFiCav/5fX7TXcYKlIcBH3UKAdXehtsv6Spg5VPU9R/J3y9XkldPxiSV
95vgnna4n2nAnAz2U6NdsQ7L5fz7v8MXR3rbO+zJQZVgchVviPZo0baC4Tx7nrzb
TuHwm0TPUM5fTyg9tKTw4tGLeVtskx6+f0RTbZp6uArbwnLY8hxNs0nBTtwXQHzZ
wtqkp5E3a/NwoGGqXy9RUG798H4d1i1q6cEum2gle03YZcl4PoJ+dLQleeLYJqg8
UUMDnAVE3Xq1s6HljB12QD+megl1/Sef0km+Zx8IHKR2/MTCmMlGCjjhw4Q3/8Fb
w/tu8bNu8FY3h6xDEEm0Mxawb0oOxPXTrvY2sOGYbM9cV+0mh84nL9b/DiqmaBA2
+e2gu32Vq3ZBMexXenm+Gcyz8veoN5eti14zucgK92nX507wLA3w8XaGQcKA2Tre
WVov8bwDHAqptBdPnUXckJ+XQfxbHM1y4C8vu1ja2Lgg/ho6hiSLCxwi7uAq3/XQ
LkCQ3Tn3Tdj9UIlB7W8bVQVfc7UaAmo9HoUP9MxGSj8cHttWrHKiQvyoBXjwGihM
sLO34d1Hw8cmnPU4cWhJrZxeXgFklA+9zCM2WmtV2IwLkmE4sXE6Hqlh2qDpNVQ0
X8yssFMRYtUEI0lhubbyQTjDBFgXb/UdQFzghPvH8hRWe3HxL8lQN8+Airbu3/ap
Q9+JvGNw/v3FjBiSkUQsTkPiVQBBsoYEjG7ovII659ygHh3an4/HOGPxPdecLIpR
Am6K959jCig7yOyq6JhTOQ==
`protect END_PROTECTED
