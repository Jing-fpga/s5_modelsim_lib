`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f1rK4M6ZbSWIQ7YMbmvY7UhwsHCMM+MQKOZ7Rh0zgdo1GVYrPd4p4McJxcnRf+kp
a6oIN1VHsJsuuC3XSo5P/2rMbzAkx1dGo7NGNi8O5uVz01n2rfQoFndZwvPgzLYb
rF7DBTk1dfFbxFfyXyS02vJMOYMerjwCC0f13XucnYXrm9yFTsvB1YBFasQOZfNa
LogiyVCSHiKkx7OvZ5ln5Ci8J4THDjyq1TsdA2bP+MFTNJO2lja5y4o5vaSWs1AY
QfX+urQ1L8gpGPlPtkpLcaA71zS1umq0pA/GumwRy+8drEmXeTEmVzLN0Hd7asoi
YmYV/zoyf4Ap6lOscIGodNRarInCEKNVAP/JL6/Oi5YQ01XegGpN9wB2a3VryMjJ
GEoXDzTY1FZPxWc1NixqcxITROrOwm2tD3ar141y6Ph+axfkEzn0cI2YMsw1DUbL
Pf7uiJdTrN7lrmiJuYm28mg8Kvmd1xeJ/nJ5Tw8RU8C0FhOOrSE+9UxizaWvpmje
LYlXmdfYyp0ROfqri+l9ASztuK0AH5BDFTJRlOXoNxCaMdAfnYLtw7d5luwyqdnw
gl5t3gswxBFoq+LdepjY0Zv37XbGDlz4YXD9WCAWD4qFoIdrTc23fwjW08wbQdlB
GnNw+zeHbfqejLTemWA/TtGcm8/iWnnMmyQvZIzCEUpSN/1EGj1l1vCgJcyxU8I5
f8uAEcpqv4HDlkT9CA5EmvOHj2oUbNeD083w/WcQm5BUce4MRlpcuDi39CqKxop9
VWrQWDsvDAsYPpQmXa+R6Ik4lKBACqXJqfTV8p7sc6mRmxSwScisUVVXs3jn9EZt
Ys9AhgbfxqP4IgDuM5nIoeDNXbP6Qw4uCkLW+FzZPZhiWMAZlmYjVNf2TCA+Pyt4
vbOkBVFmLtoXP+eiJGrNiF9gh5Z3BHN73diBrJpStsFaCHNwzswM7Z61F/60qit8
qVTInpXBwFfrO9jKZFV3/wgF766Shd261Ce/K6sqKep2KtsXY0wp4WsqsNuACze2
Cx8mhoCf/w9AhRLbfKkPfFlVC5JO/L+Nxmps2DVRJHCKlc0WqiVcPc4QXli+eORk
zQ/wwD8jLFP7n0vqFlRENWvBzRBdqT6DtaQpEkaN50jB9QZJO9U0QQAdJPTCO1kw
u36VDJfbM6LUyA5eplxH1i4XBPMW62m4jBzd0YaqYNVpx+pdGoXlFuZkDWe1GX/d
rUYtpj2wTGHBIkLWUgPjJI2Fp5i/kXarexrzFOuNbKAwYQ0EOCVzYiYrNLz/CgN0
Mzj9jg9Wz8uK41sr/7v7HnFMWJE+eApGncuZK0SK5WkW9VbBN140VcwmTZJlwONH
T7p+SI2zb0ZZAuL00QCNiGE4P0u/LwrqVAdd0TuBVI/o6VcoK9PLEGQsRXZOdeZ7
EBWxOkhOI0H3BmJSkJ/HHZcSr3mMG90wN64JES6HgmboRtpKS8X+IwFuAArR+FXs
Pr2kVNOFL4yxMf7nesn+/pya24tiwB6CZu+bjT2nl2IKKSS82HEMbOsV0Yqmtj+y
CDKc0CEstttF7WsLkRZMTRk/LJMngLTXxEIQMRlsWEq+Nufywq6s4+VLFr8G++pl
fINEU+guooMF5nIlJpAZLND3T6SW6plNBY5DauNcSWoXQzr9qBiRx9XPVyo1cwlr
hpFLEUbPjbcDFvo+iRyQ0GvizZZvr63KM8mJfFNaezxa+ArR57rz1Zh+GuKN2kZM
RklK4HiOLqf6y43S6/vo04UPU0efZ3uhrlmeLFgq8I1TZQG5Gw4gwwV7e3oZb+Xw
wCEJPhUkaOApBN28QMQFfRROQpcOoNlHYpdJ4NbAdmGvRbPTxtp8RTRtDyg0Y+NE
7re0TeqNConbhjmm0OsKMfTdQrE2YF5hZn8AXPSR7vUX0ZIktMw6Xb1BXkrt9efi
PqMj8CW0rC8AluTWwikz+IFJqfG8DDUVfIBAbltAxdb7xcEFsHWZuNH/RlMvqTqW
45HPRXgg2ZsWVVt7VYZP/zQC2F0vpTKysCG9UdMk6VkdlGo+yY84CDfVUT50g8nO
9qZYSNwGQzwhcUXwk/8+hhIZ338YtDH9Vw1ifXyOrqivCm0qVmhd3OumKzN7u5z6
v6JwPoQJ+eV7S8LRe2i/dt2gp3dvaOLnEsZaYiiBnck0+HPH1ZNNnVLFTkR+JFpx
ogvE6Cq8y2cebk0yrHsi5UIh1yuapOUu89YWbXyi7NevHnMD+lyFB3SLwwjDcI5a
uL3KQ+J/0L4phppNDdOCuYnaoNV95ovOPScipCjQujeluUYNWbGpR4wae156WNTy
cLkLYfD5oEcGl4FYq31+z5NulnX9aEqNTwz/IO07nt87aEEpHvuUP9ndl9MNQ8jE
T6gcptkZoblbX8NaW+MhsmiHevAw6XMOhJ4kGzj2gTNF6DEkHmtF+GFMhlLMBtbb
NpVMKsNBHULU4zgv3RLKWgd0yfJm9M5I9xYKl2AZ2ctssRx0pV3NQ6qJ/G6kyXgX
cr7ANf3IHkUHJcYK/QwiLeIz8uA4r4357E15+7kEOwFd88PRjGHTZsQ6Pz/8xFDF
n7bHmn5SCzTaMOrYJxCXrTPaTpe/Qt5zVVF9E3shyhlDNiE6isDCkAexRlR+fDV8
NK+sYVUNe3eDBd9a3aesKDQEh7UwPTWEDdzztfajPYSUVeP8iA+7QkyMdbPSWqgn
SRFeWtgrlpd8Xs2KjD/ICFhLd1h3kgzcxeC2vSjjPa1QfvAtrIW6dOnwxFfyPXuS
N8Clu8Hc81PAtgzVeEjxeiZVJ2MH18r53R4YeWD6qhKctmsPjJ9Yjo8WyiIY06/1
GIn23uDSeJ/ByO/3jlVHCNQGQC/5o9IpnM0pq0+2LXgMZ5IYp+l+1MNrNZpjspcu
yGZorqAkrCev/L5WnujRt08YFMGgCjkP72RwtzpgTgnHNkLinp9yWAX1EvEeVU/0
IdBGkewG4+rN3usJXsherxLD9Wc1y0Yjkfq8bRXINH5y7xfi4eJVHvhoVrN+0abL
3ADnvm431chxBfIakRyql37leWOhXMqorYItg9PblHG5P8ibXhlG9tsrfLegickj
M+wLXgn0nUyKjfdFMz75E5eoT3eTXFPf2QSP+wdbtPUy/juyjEqEmlzBAOZvvEBz
pK7Ocixg1sJFnOHI3Gz4XLDovb+Coc2R97NgfwIkBIkeibooLSToDIwDagpHuIhj
dlSh3PG4v4i8naaqhgpO+IuEUzxsd8vto8DSL3jEwBwpR7Y9En1YtK16kRgxa89s
+j9Cc4l9il5tufaHOHw47ihFviFajh+OkgjJr9S3y/vHGBkQ1ZMtQvO61yjhXFKA
7HLrZWm9+KRqzEQ9M7nSu92HhPBSbGB41XkvprbpVq40Su6CW9VH1vnrhhph/kPH
/o0LkBPi1WnExJJxKLIgK2KK0UCtzxjsiWe+UVOWnqR4DJSv2r4KTmIoRY+e1fZo
0UkI9KpvB8KosLm9iDBz1Z7UyCW4dGiuw4EdscStSH/D/fNLhgACaHQsHoybmwVW
5KOXUDBK0pUzTVh0LhQtpRS2uvyTrDkCuEztQrnEsRLvE519FhgvuSwtrKTyZd0v
ue4bK6dNw4KZwHjGB0XIPbLg675rLjHzptBkKbQTOt+ES7DwEPqrptI3mFPXk/EZ
EoIFp/BiTgh3GghCYvMmVLdP6Y8cZ1Sf+DEEwwH+ql476XKg2WEnjajxLWn8jYU5
qbYhKthPdbOr1tZS5Y8z+dGOS7aXbwyJWNy2VHLAGlD7TlcXq30zY14hI1WHpwPS
rr4EaLHtjJIVWPd7lOWVGhszAJvGXyZjp4DxUfqJp/q8nyASgFnvU1iwQiP1k1JX
KPUtdNc+E97JFqhGBolrppu0MjD7V9tm9a5tJR5cajXiVkYQHbcg/zVJCbveqlXl
AsEB9/Rp6gZuKYGWXD7z+8KDplYKWRW3ee8Eap8htH8TRQnmPaHjtGsXzf/pN/kI
7d77NWs5BpR9ypFczbDCWwpibxYi0M09egVOR3r0vZ0T5pIqNfHYtJnAjbrgr+Lw
gOP879jHo3uMMPm+1BJNJPT4mMznr9uhuBGv+mudJRxZx2g2JByZTukGKj5pDQE9
hqEFdqfzn+4JvplMeSFN0c2j9DzTKBhJMdW9VtUAW0yaouE68CnlsQOwELqVW/gJ
AggW2fssHNjiyIVXVgHR3b/9sUqHKBFpZyHmh0aq1JVhS68+fw1ej4xw3BIxZPBe
Q4VMeHs2WLN9r8bQSo2566Z51DYNbN0lBogQOGPmvAMDygvsB1OprI4RX55vDaXI
5HDnLC8CjxJ/XORs5O0SKuPSC3qj1xW8lRQx4/xoGk2JUEVUujsjprl+Feeb02Qm
hVfpzatSVqgW1/TeupHAghTqpFFub+l2h07pGkaFRa1B3Um0n5ieGGugaWC+LF1l
ypdtKcZowVedDfapq5PTTSZy6uZeHyDRDPvGWuUj6sQGTj/fEaO1g/sNen4suE/Q
9tjDGe6FQlAqJmkiEFgjwaGgjy0xfnXLvU1QCK4WDTKjtBQVzi2Jgz8gJbRv6PbX
q8QmNEQfYJ2WQsuK2ns7KL1FWd2DdZeyENu4/tJs5ziZyH9ss+nxDvi3IPe5PkyV
/VqII90ersfP6QDL1UiQPoUSOsyYwFyhptq1+eU38eIg9qC3VwrZJiuhLQxvYB9i
UqmHrj5s1V9qFuhbThvxQTblj995SzICHkFosswpvhfdy95xlKV8KPrO6JB7peoQ
ESy1DuUs73djoDXHrdBiL/wn0RQHL9XTYKU1HkgZNkn1bBQM9GmfFWKQwJwE9mwf
WTTt/Xi6Je4aYvrdPQIQqMmMO1xnnfzqPbaz91ojaktPuSzzknlpFLHJGLYMXUn9
lkoF0mhMc885XCg7Kv5iIMBWOi6mb/0HZ3KC/utg/A00zqWmlicsxoa9wIUEGObG
uhcYqFUTV9fV/wlAZ/HpCmg+w7EBlGCgyKvycZawtGARuQmF/kN3YJIx5PqRMN7c
kZkvqnzKs9KRpl4uLd+yEc9k0pGuOcoobPe40zp4tTVEB9BSo+Ws+bE67zfUp2n3
lOF2JMmmgRcJlK8Ae78VDy0Ud939/soC2DWO+WUDilOYpt4QTviTvXKShbjVECk4
vgJTSqNv/Pc+6hkKdOcWKXP3khospwMEqqsR3S6FFAtO4USas4xl2pXB+buwVdBU
ew4lEq7ggbkTuQERLhVEM1AH8kl2R2plIVNUIyUYJxzmCcDRAhe7pLT+Mz2uMTvb
tX/Wc35JqYeXRR9n85XpEuFSaCi0kz9cuJpm5XUlfyCD+peHme4rqfrSbmXVh+xb
yOAdpCug+T7fcgieb1EH/AlPzeYZ7B0DnI6DYWtvdaO7mOXM0MObYnFFij7wdmMK
BbduKxzrNlKeWrJLcSBEVBBVMQe1N0jbh43K8IyZOD/uRD3o2wqizp90Uwei2alF
iTZbhXLRQ2auvxve3inQbdJDPvnsYh/TlJnD8e9Ma0FtKkyMNvO/k3OLrUcbjxWt
MWXD4jxCXMSbS0Q6QH57ZgGpUQEr+YXw93NE4oUrJWngXHBfuKMVg66bi6XN5Sik
osACavqHzf5uKd2B9kzS7DXqqNBO4vS+8T4KmJTA5K+YpBDIx2BfWmQ1rgoC3d6M
h1KOPSfwlenVRVmdqoHnQ82VzgBCdeTf3YTKLS2PnS3T/F55KM8YIuK2sFB/A4tj
ZpmoKk9nAcCBD2nrqDcvvHWsI6ZQxl6BWcTqrqBkE46KyjqOJDN9O72t34ZR9vMm
yPuBi6eJvB8Ipd5QjQdk54pm1Ivgw4zZjLJqBBFJgVrV6SG4nES90309iQDHZoB7
TSO0Y9ObTAK/Df5u0mC6VRBGcaRBZDFfY701e6aOIf97Kbs4WuZk65hOA9UaEF6t
TAzVedJaqJcTxochWs2KcHX6XRT22dd3ViYxupR+pXGtQRdKgkXqq65qjhhUrVby
2pRG/EFJeEQyiAYMvSVS4/As/AyyIyKJ+JjN1iRrCDwwGqWWcPFaH9ydKT7MUIki
uAh4vMuEryrPSjM74uDUs9rB0ly2qTLtkaJw9/xI1cCZ8/+y6ifgDFgf0Eah2qzQ
mTZGTNUBZGddLtXwqTHyJtWSHf9lItq1BDwyiJNWLDbRs077RSkLTzDkq6rQuBdx
5XS3vjdaQyiEWPkuRrJdvs165jPNOoEIY+Aq2GdIi5uXrz+FahwQ1Q2gvI+7tycn
Mta0LUmvF9JdRnurRGVF59X9CVNAcgwtZvykKecrUdVvdU+82wrOhbq+yJ1qzwk8
8azsFNzXfEmJ7iuWrb77kCDqdtNfMg+cyRyeIsgDh3pQ23VOdoUUZ3oBWjC/+ll7
f17MlejIo5+7cN0LBdkKKiBdMYcDFRoqv93sh7CrtrEmFlxCqkIs8HjLA+dZnRsc
A7fLP0YAvBn3UFyOfgf2NC9Aw4sJ7zNPueGeT80X/C5b98QctCevg3BcPyh0SlEn
siRx5U/mID94M9oxyokqjFmArHcO2n5g4QxJtxYJTN+2RhbCCvtRN8DR5KPPDXs5
+MmANWOTTx6IQ15uszi4tp7/iVU/HxWj7ZkJHzbTrI1rqKoTBQwbt8JGJFl+g18m
SpBOrkEoC+6ovmEQ1HnUufZm4GWyAW1VgZDquju1A/fDa6CfSJRLlMLJxJnz73Lu
W6IajKrWTiF7yQN8uRzJcmx7JDX3ydKaF0KqMYDkCE3xLNHC9uYNycUI8SM/U6xm
zGqc2QjfOEs+nya6jRJtnIaE55tsFt0PD/L0whx6xk0G3ZNORx6j3cTFyfAZsmVx
DsHRd0lFDvY2nBOctY//+GnuxKi3NQ/2Od0BQDE4H7lWyIn7MZ6qP5zFlEH+fkgF
bLqNAm99cif54j7KERtXMC3+LCthPCN58JXIpd/r069BQBtemRhAm5HXpldYKcfh
FtfZjB7CHB8Ow0MADPG4IH7pzQjCLC6NfhoBzeNtBvW+jp7d/auZ0X7ZvM2OH7lr
sq333oKfEGQUoQpFOjHsccocc1pqEX7rgkCpZJrogpW5m9gTh+HpQCCpIjulhlZy
THPkCXqNIscFU67PdaPjFpYN02L26wh4cYVOd98Hg7ZBye8jeOP3c8b/PpuklhpD
1W84taB5+S4XbdmziF8fVJWkoB/iWMq72X9K2YBcwHLsV4K0YTNtqCJWsK0t9LOg
V7eNpSXONQ+BLksymYiGtmJUTbf1lSPI3KzznxkShswNBX/qyG2IQq5TruP3lAL7
0wR0xp2RdXuiDEUsRKu33VifUpmSXMzVanzIbDd2IixJR7eyfJJL3KrTq+RRS3b0
Kho7IqG8VeYs10fqTFhJlJ7C4e5aQ3VnSDvxv0i+lx+opnxOHcUfy/uMDWbYKChe
9PKc9VSaA58dZUpuZRqfCUpp9nsh/AsbiKl8houbGwu0ZNbYUMq5AQ4yHUMqTRNl
LHN8VkjJh/vqcnYeWN8Z5wM0MCJ6h50qMpJTuBp2Fw1vGwm7jjFtFgUfYtRPyOZo
30XgiDUUxpmCqvYfTwv4ouaWL9sBUtlIZZ3g8DRaJoxep7E28A3FNAS/MSQ5n7u+
PIOSoDLBOS+lwQtCAOBXqsKiRxraKSk+gFPF9BVuNmb54ahEPgpn09jv9hIGD+JT
snnWnenrQNSzNr9xk/wYrFq4PuUUx6ms0qYmfMVbFxKd3yq+geHyP7tR9ZjfGr92
xL29viWzeGSv2gzx6a0C061VV4tqLjvUOMvI55HFEcxcI6KNKslYq8Sd2QRJugfz
SkQxZfaTirFkIXDcDzpU8FnUl/XNuJR5wVR9vObR/avrU8pFqlYjgLcmtlyhddwK
w8QGAHfoVuRtYXzXsckTGLhjYjwBni8wX/8E1JQsikRdyui90H0kqTRdXiAmKOGk
BN7WsBgu4xw/bhUw/SDZptrwUUJSsTGWXH9mLPV4chR3meC26zeZTWiLI534Wg9C
ck7xPLQiCntftfKhIbjNWBLV0Yl3qt0zQTi9zGeLS9/OmP23v2b6xaSqWbhZWoRi
SoWbmFl2yQLrgX/Oy0Zqpn4wphhfuhQhx6Oa83Unr1MkA+IOj8+n70OblhfJfO4u
weUmSxDJJNSnRxom0B60GtpEW4QsozVLXF/W7twcP83Jmco7sNuwGFnV/uqPKwzS
rVp5gNdBC82YPGj8aW3zEercNaRbV8i3IhaIcwkkJ2JLaXduZC8rzoj9cHy3fWmB
eMLkC6ci+KoIoZMTZCNKdAZ1/DCvMV3ixUJ6H9bhgDIBE38k2AygV3rvaQ9f1TBB
P6RhA3oL+g1V658tW6bgTrobIbNTkucttwWjhFpRcXMDk5u0V5EcbX0OOS8PWRj3
ARBKftlz4LzhnGFmCgxxoYtmpDLplCxkVLvOv4n0xnNqPLH6Qk4ofuPqWGxdHy+B
P3IokTWeUWtgCTx6jZfA0pPhoG27UcS/wABsmMAtf5euKDmePVUgSvSJh0sNHxyj
Lb4WWyHtTq9coSXfaIeLClIJl/2nqKVfbsGZlBl1tJJoJsw9dSSodj8gTOi/JsEm
L0ku3/H4ErPH2dAJAsPYqMRpPFtrdFSrnGuX6mEJdCX1vTa7gxupvTdSNW43XXbH
hjUI0nx6n30K7xmqjMCkdqaR/YNVgepyoZLVao0prD845UAgDH4eeu8OVIv/Z6OG
enTVMqQChteBsEjDIkm1wUSC7QrHidel65jTQDg5Ap7T4WtvAfYj9WlurANlDLHi
4J+GQRhhhzAMcYOcYTPaNKuN/0vz6ZZolekL4Y1ByPwcpQV0dp0sNNato++GxTBi
rJlKmPLCV91yA5KkqkgxB6RdFB0Bv1SBSuVSKfKav7yK85L4KSgXwumeNam1OaCh
d4ZPqSqBpe/utNm7oG3IJSVxJhTSqnUcIFHPG5IEZ5nWrUoCPym/tb7Q4Cl5UqFx
LTj0IZ324StVjLzZNUHOtvPvWy7CbSFZ95d4aN+nibOPIatDeK6pKj8yVUdIWPLE
OxUyLevxz2zNz3/vgYsF/DGyllF7pMyAWmNaf1WUTnVoTLYPrHdE2DeuApQDSage
iN9lGkRG8AMIq1CamAYQ0bTIpJUutuMqTNandRSgprRn5AREaFOcCqzA2dUN8rex
ZvTYVqW1gM5z1TSu9hytkAPbcMLz3eSDtrq3w0RdhohH3eMqe80XlQSYz32Hm0Yp
t1Vk6vPYa1tjtb9MT5DCPIQEi7OxG+WvaB3s7ipiItDgo/eE8Vrs/3DP23LBvx4E
JqTLdPu8NI7YCwHKp4AAkZFZ1XadlywFAovvFPylNWqARa5vY+cJzel+a4m3uyBJ
R9Eu8tYXyZCs4q+W5m63ci6vmnIgV0ciPFM+dQrFcWZ0Yl0NX9wN424aWS7/0IvO
snV+XCypGOC9BVCAg1FtNk26DVMG2cUdZ4CRsoPZ0KuwRfb1HEBH0q7QSY1XraqC
Kcolozk9Zcjqv7mKXjbupb6D8Kv8bEOSUvVDUrjQUl56i2GDoBnNkqsk3jbWcNtm
Zzci8J/qW+S0HbFcyzZMN0rpPWXREcbxxaP+ek3WBKCUpIrJ/Ho+vb4xQ6c/BNGA
8ci7YYKIJ+tKZ7I22bDi9OAQjOW7AbiEEvvvRY8nBb2lJXhFFatcCiXXeitPLRtH
MzITD0rxEpuMqQXE/wXa+UAwz6OnvFLxYdSq28Sc2M1j8OsF1ZLJUcB2fyo19tBF
l353i0ZEHUX0bHClEveM3/avN28ukW673hc3DBZ0BpeY5PHWW/WurSyE3JPYvziC
8504rgB3kLu3aidiZ41pZq6mTh04Rccs9O1lvnGgLcix0WrtzxLU1/Mahi6tr1cI
GWHO0pKt/wLfXjknwhEgS3+Drq3jHaLyF0VqXl7tf4p1dlUx/XZu7nQqaDlZ7NCq
N0XyHN0gWgH5tJH68duf2tQ1M2g1pq0C4xhU94wZ2MmNjLxO7wjyIL9QA0d3+2bm
0qO5gXgqziRKi+/S4Vm9NkYQEDupiM9lv3xiwWXS6gvPAVWQ2B5/bnohuA2Bt8jy
CVXJcCDZwa1ieeSRXGkYxZE07XDLMIw4yHO/14WL4Qy+P5ocb4vgf5Ejx0fxDHZm
D+6L7LakBA/4vF+3ewFSjBk0tz6W3+npZ9N5Z9pWvItk9StZuSjlSMAo0eKjgLzS
jf0W7o0HlNr+oUOYrLz9NZs0ud9odrt6yOaLZVJlgRRLKUSyFMH3qiPmwi3wyNGE
/gPuXh+HPKrLmXGGaPltXf2eDlkogBWWm/NoUkrXyYX0wVq+8wmRPKKA9rweT8oi
yyYSeQsbYo0P95J8l/bIeZ5HRvyJ1v7//nn61flmZUZ/3BglnSYoJxYRAD1XnYt6
KxIb+Uw/aIludDXFi0kNPs0uPNIRiGm7seIRjtB23Jj/z9xYH5A8mVBAA+Q3S1Dj
CgmxpQY4uQ/Yzo5QoeCrTQNpAPJks6Imf7qZWstV/CwAcaBxoNiplusZzihfpfLa
KkI8fwYmiZtVOPpRjqldDPxxEvjWtJBQGi4n2JjTqIIJzv+EgVz4rbHnA9qe9EW2
0pJQgE/sLwasF7DXgLshpCKH6x1uRdBbXlUjqp8TeZ/dW7w+FZVNxpKwzpuahXR2
k7Et2L1pfPJSJE9tivaMMARXGSI9Tjj3k8DrrejJYLGSYlYuG4Vx+zjkucdPPK5/
e4kqNcQq6BQbySJNDtzAg5mZT61xmyc2zsXPn/ArpxbStF8gbGQGZt6QWQqhDZgi
aPV7I6/JtSMovnAch4UAdH7Lr+zSu62XEZfSTlE5Y/bjZjjn7FwnZxDNwJ6AL75m
jfQ6VZ2X70r5cF3rVXxXkqcGin/rEaK6ci3kL+yTf9A408wy2u4zZn9MM6cP9bAG
X77BuJbY0bPBJbr8ZFQyxFXdf6rf8XtKR2xA8G0TohFxM0aUxhRcmmxXI8VUhLPJ
1tCtn7BOYFI0RVX+jdRZd429BPlWNemsT4Wc45lKzdvYC7C/lJOm9ezcRR0IGaNB
08PHc5dIVWN5Yb/gthYqhxl0EZ4Xcj8QNKlzUKdDguFChmrbiUV6HldN5t/sLX/9
5mwV/QJLHRqgTHw8mb7gpppRnkLrgw5yj8DCeyvgSIuLWfG2hd5JZJrBmrYETc73
ci4ZRpiNAmNunlY/kPzXa/a8c1HVVY6xDFazZMD/uKwA44wyue8icDPvsJqixTcc
Z15YxGgyfkxS6FblLb+oef1idJJJqpkIp1OkvZ+FU4hROB2UXjqgCyr/ymzD/xmL
dYd3NSwk0eOw6MUxw+1zlBpkYoaqQaMPxfekhWFxHq0ktdjtXO1+Ps/iARCnkSGr
22RoVHihy0htAgeA2+aO396QAFZdZ6d5Zs46RYG7PCpFQnTzid5fOg0DYLG8HGKJ
hky7ivF+vv8pYLBc3ATRyljx7+a6H0WHcCKt2Iqt0ac=
`protect END_PROTECTED
