`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1/apAur4Y1kM4vv5IjHfAV9N3PSvjbefQxJX3PsS6a30Gym4MQwpIM6/yruAdHcw
3TSObAmwFPH0GEg6/XWiINZCZh1ETuV7/ZpNAMuJohyMM8lAXCXmOQN74cZZ4dk/
GOBAcT+OnOdYbqS9eguP4ntZwml/prEdCfH1zao1AI3Oi6GcMipSXKJYdzhnVKOK
/P0DFKNShvFPlKOlIZryjb47WJprn4POBdtRx4yiVcXECJelTIpkY3wXeHXEsTx7
SmXbcNZlrWMey/xvgzswSKo69nMxzPFdnOPFqZMha+zPs6wHOhjIhK3ezepksFmD
t+OaBIdarPs25dRoLDmSacYQO2Lvujw0icN5naB/mSRQdHBd3e0T8SIFI7Yx6+hm
ayE8Fje+65JLTunQtXxJ8LKz9jhB3iI8rrODjobSs3teADlIBJ/TMSjNJLdMtxkz
FH2cOi+3gmfEoqhOHWz2mYEJOjw75i2PzdbxrKO4qWyMwT5emqjOPoc9MpV4tERP
s1eU+agBgY2pNWCCfMQewea1kOQmIayUWMePb9ah5hoOQXQBp4tb0BQVgG+8hYqO
phIk/F8P3+IZX1jVBCfZyogSbqY5xEv3tDN3BWbiMo4g+PsUCT0OCjRMNsExaKSv
I8PzPGlTTFoc/RZGxpMYR9xhQpeKXrEXmNpp/mwWM7d8C6YtonjgMIaL9CPuQnRg
0aEpzaCHiOmrGf7QcP7qSac6FGmPBpVyYNwf1/GSZOIfylFW86crhaXpeE88Jb5d
VhrcRingLUuTnH0+BY7QSgz5If5j9mLl5rYf9cW98RuelgsyxdWALoYR3N6HE6Ms
cw/H+eElunM2+8PrgBJ5nGS+FS3KNL23ex8wgptvLgTFSmfSv8rYp0X9N2QbIhUn
IB1CpfhItxlaNyU5MIz1H5KDsMZa6eA1IFi/s6liTyZSl3r5lgw9M37DUTioc7wT
iMwCbj2u9mtS+mRL6WI7UZ7PdHcWdKFzbGX1AmKNpth+NBrhvm3zFmBOcPrmqQ+S
XdD3isEhUb9gjiAesizQTHiBqQe+QWjetrxu6f8/DymFXFh6qXEBaB6FO0Zm4RO3
PqGO8UgwWT1yIT06xyqCXDE2VwVghr0uVX1/F8TEnEAggW5oAKXcZ9VwBxk7U6KZ
kMGyLfwa0Xv0VmdwIhhtLrOEl+Q0cpAj04V96T4N5pbfDwgd3Vl6t8yF14+CC51a
JxFH+H8Lh5CcsLaaYap2CYRmqPEIbS+TwbX2jv58t8SfTxiRNXeeXuIhxqVcZMTY
`protect END_PROTECTED
