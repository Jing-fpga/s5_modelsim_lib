`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ESqhq1a9oLRReBh3XmLemS37zwloE0Nihl3CMQU29RX2B+F/Hh2X722DdGmZorln
BC/RKZeENjtLSyCNQDgdQK8ILa+qjo+laDY3dSSW9rSyEQ5R7dmJiWkMZUGi7l+Z
ZkXMvePqOLR6WwPsGlz4+PisvnNEodoUjX+L1B316dH9++Bd0eTF7pfFKPO4Oxy5
WtOP1VtA0kuE/TJI7RVvcrdwJv4FzutHtTUaqeGQwhqNQazVRWYLBB0t6mePjn/2
0KrF9IQVFPG5NlMWfk17/NR8cNtNKbpSRRoKdilcNTv9oQkq/Vfo1tA2xPLa9Fmk
svhkPgrwS+d7da3e9M93P8y8efql3qmLRy3oMmmdwkIN3Cx/DNuQzkRa0c4iSXls
ItUKW3thqfkz6QTcpvTNNLsbiMO+748XyiqZ6wxDH7IKZkvCsC+CqzI89M/DY0jb
95Q560dxiRqGgJwokiv7JRvX2NA4//QaW6icJM8c1v0f+FWeYxEPMhaF2HdNEOCK
nXz5F8aQ488A1ixKeg+dN6bT0skyrnmxyllWTQrWW0/DnXgcoccWE6iQaCYR0Wid
m5anmNxRfyfWX6hHKFA5KK+ECNgnSpSvO2XEZyYQTSDp6ZZpRxzYzUsFRNlXDJPo
66du+3PX6/+TgliXeq1gmXKDMZhKLzo42bfKwdPBpGm2tnlRguwxDN5f8j7MwAQr
mjNRcplPOG7Z4G/INbDy8X7EMbdtu7qRS/b4bQ+W9rSeq76+DFWgeUYiqUnJTqyy
MiiI4siKjqvBUjSfleo1fMkEN13WdJV8+SidVKCUWfAMiMPVytOtnUPh04N1jQ4f
MpXTuKlL/AE6TqDlCWqbEvKvMvj//kswLD7dV2SuBLceObJ37fKcjCbNy6EykKGE
URojeunel4j9Q1rCOGLv/KrcTZW7duDvhmyX/77Xl7kjOevXT9KElT6v84d04G2Y
HszECL5VxSLy860sSPuyxXXuFb0Mtc/ZvBRp7XQtItSFnOX8SuOWEvQd24WI8bh9
`protect END_PROTECTED
