`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
20PuZrfEVF98ke7loIQRfSH/3UmInD9iwiByTa0V7LV1fkKHp+Qd21Q4MmtTKvPR
EqHX8SiI8dWsXpQVaRHRijvEHe+CLjqF1rSoRg5274TS8v9vacPKh8775400zO2j
H4JvEUk/PCHVQgpvFjuA6hxb+aI3VUMHxh6DVY5c0bgb6CGb754kk2tUPtoTgub5
OTEiz1Pxm7sb86Crc6FBM73gbLH0C+bziwyO/d78stm3YkLtDROzNAhuEuhM+1bU
32Q7OfFQ2OWmeANfoyj+1y8+2XWfcexb+BSXoicY1tVwoKXZhnchAfXATYmdZjq5
hu172bH7yW+mHnFm5ej5SRAyA9tUz5AxNBCFnrPk14lgdzgxnESGmAIv2PWveZQw
tKnEXccERm03THXNw7n6qPl6UxzGGjBheW4t39O6eeW0L66Qby4e0XLePeAF9NLq
mcWX7UJs2p0KAxa5IngWz/5u0mYJTfjyVBKb+KSsQIqyarGft1ABXtP2/MOLqvZR
qUwzgp+hJCYVPzbaDPP51+4WH7w4Vkg6nuq3beEy44F0OQxzJFLvcdVCI7ZuipHh
ptu8kGaKMQ7lS4+WiJvJpNnGFb235oEJSM+n30iQ4idYDsLlUC0IAE/l7fhVh9/Z
T/zKD30jlHOcNbt6uGER8ValkLTbZfepGR0a+hJqCGEee0JUOGbSAMsKrfcSaD+Q
jgkgY02sJVIf2ZSW/uQEsW9zE0iKiLb0fWsY0huouf5udiJiIE+rPuXZ86CczBmw
+i3me5KEiW2HA0ao7FUVASAIG9iHL+y6Sbmjj+Y9SoarCFprx1CHky/tTT9246ho
5BZbZV5yVJqoZppc/3CiJp1Ymc7/uTswzIywoSpDvMBQHbdQxyibQIhLPmNBs6Ua
ds3AALDi5jRmn3mWGx2rh4Rrq97g9+8wY2VUyKzVqo6bBeYJE6qDAE2uNdcZdoe0
3BHU0jYI+rpTbC+si9U2FkA5sOJO+HShulYJLQ6arsl6IImnv57tMasfXHfWe3Yi
hZTFZtVxvyVppdbYvPyZeoHccWtWEwfOw1g4sa5J//DFsiqaWRRCLTBAE5PMK41e
0YKKLQKEXS/KFh+Is5zlvZiTDa94FhCBEwgwtGJEqiN2mLeFp4zq+x3AaFIN9ryN
Rw0bb5HGtNdTRP5DONgv4Qx2j+wlEhoeshjxGI2Zp1nfBLPzTMuDp/5dIQ53xTz9
vwE5U90HuxAwG4vYrX8EzO8m7HGtbUG30oje6ckDuyVwiJO7wegMiFNGWNyl7Ma7
71jEAPdDCeAJvM/Hh3HoNgOkgeBizoS1yQ6Nql44XAQbgELQsOmwvYnAu7fdzVW2
BhG0nr3ZJQOWnqkB5aBMjTkFJ9NtgGZyBFJ6FHMkry4=
`protect END_PROTECTED
