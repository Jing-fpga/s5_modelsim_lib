`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y4Mzj5xns2GgorL7qVjyNYxqgeZwz+OrPsdwsbU0oizLxWXcXshAMaxu9sUAF9r3
adZRe77khqt155xfu5Cs2NZ1OzeRDlcP5dhfJZmrCIN/bcDxszjN8v+z3Iwomn9h
hPsUar4NCSa7BPATnCE+Ort4AJQIypsofTC3ZAq/nyWF/RwC/P29tlCHR0kh12ag
SB3KPAKo58njItJQgyhJul7GQHLhu7klwEhPzWghW5QaTZdjByUdDdTTW0GCnA7n
XS5/ZXzzFKuqZ0ILnLTog02xW1gc0pRF7IFTn18ylifNXVlBfrZGsZ7AQLN3AQYz
l+7eGNFl2D2es2H1mTJu8PHMwAqcUjXcpWIp5uy0Ls0HwhqPWviCSf+LTqSGMeIv
9Ia+Yy2Q4May4UC1sybD7tGL69hZAD9e3jBhpwuOIAh58LeOdvFENvH0cvWzfutD
jhpaJXOOZwOpK8UnrVFB3lzKrwwoIPvXdDRibXCNONdIi0XGuf61Wzyip6XvcgvI
QAyKxD9ZGp+G3icW+U5V9dJuxImCrYDoaA1mg7wOYClmNJwFYNMizLyY1tcSQTZs
4vrsAas1XS5155t/qkq5EJtnQ0svh44lvVeRu2nVz259A5IIyrJehwjhYKBPiIWc
Ptg8X3bPXCaBX4ca3qs/6D18//p6SfDQF4tQCaWnenV3viNO0moBlJ8MFjClZPte
G1fZ4UIEnewp/AUZvYziil9mxgadYTuaWnKCFWdZLR2K5PsTK5EcnpX61IYI0yWV
rhepea+cB01r4dQdYS/X24o7fo1s4wUl6mCtg6dVQK86z2crYNhDWnchhj4w3t1H
2Nfr60n6UlXPrvBjBcpDBDr2A3SMD41dGTDN+RYQCLuHOQseh9RjGOq7+C+mDzlP
f+jZ4LTaqvlWhd4WJi12K/vEXicLuPFx8NT2mcumAsTBg9Tw7gyHU3dwvAADVyza
mJS5uJvQZNczlJahOpRpk9LUb2OTsS1qFguxFerud70LxyFpEwV10wHnAa+PMyKv
sw8J8neGAbH3PAtQfFqgUuy1fFmbNGj37mRWBDzvRMO5jcW+7wjXaWh3mEpApwTc
OE7ULjN3IvfaxLf4H2Lmfkqj1Xh3eQ6lwJ1YTaNL8cG7LP14UN5FdpgAYNnppi73
0EX33BAkkgSsc/AZn1cW6qStffhcCaOokUpg6emfbYU73A3TUhALVRbbBdpiXsRl
+e59fL3oznisgzsm86kHkuqx3A4+easCDqu3hUAVpLRsYmxy5y8TWLpRaqXtn9rm
CNBFqkuMY3pZY7fJS7m3knt6egnXqpHOhrofEm3UABwt6NoZ/0l/ZGrx5r0SYIu8
PHcLUwknPVOMmcMIMp1bRq4nwKYDRO1gvtnlptd7sf2AfBiqa98Smz8YiUI45B4H
QgtVMVXb3MR/RCbweGP7BLjEiaunrv8DmGPcczKPsHkNmLzSYRWAk2jqXPVH2fw4
9t4k7kcuA0XJ69xgIIeaHmTqKPTAtYG+nN1klBpMMRyQFjB9HQJ90QMOzgQtuUjL
5Lo3SO/buqWSavPdoJ5ln8oEnS1TUlL8JncejabqXGhEPcoLnpHgDlvHdA3zXYPw
M9dCBE7aK/Nf/pFR+2PDD6zUkGeurNyexNQGcplo+ZVyrHaIwu3yG0/lH16W0NvL
YxfUMotQdWL5RAwhggG9K64ROgfRouwtB8x8sWC7ZYTPA4BkpyjWj1VWVBcYxOV3
SO8OGJnMpQalc1u0trfQ6cTYNQUFD6+ho/HA7vT2tNuh/2JBj1A/GzmP8Yy28R8H
jJ3ATU2XJDYFD+GBvLOXsLHngtRWliBoRpMOKiXcwUqxptr5uOGkNFVH9Km3YEbe
rFNrPjm3vZ65MZUsD82YSWMYI3Tu5kGPBYvg/WDfRQExEansY+i/jDV/Uehcf+fj
00FAmOBvptbST9YPzV5CIj4yINoCoCWHfeDEvgjXDQTCSs83qex7W0H9YIP/oXxx
dDyhOQEzpo6v46it25ox8w==
`protect END_PROTECTED
