`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Xr8SSoOTWpVvu7gS3paAmUdZylgtXCejPbmww7KTDHUEvnFVR0s7fJ55qbuD1Kc
btgBvOCTl6QNjJu6nIok8vWmOxHWPIDAbekKxjxRl/HJ93y5kRyve3Xnk8xjTFiA
HJAAi3dkgTy0qnJWStzcaB+UkA+EJBa7OegD5mb3eG5oDS3BwVTq+riem1Z/UIKo
YjND/Hn6O7tU08rowBcvE/uhZ9t6rn2WsuVw4UsUKiXuYWA4DV0HrB93ETKAPD6V
uIA0zDw2baPUEa2Y98mAHirTA3MfdCtxrPNRTgUZpDOb46XPr4urpc8Q9ITAoAvM
5a0sW1eCoYt+rAWHt4pdoDhSmaUD+GcTzPgOF07uJEZZJXXO8AVU9oLATiXKyzjk
ncrYixIycUzOfR8gGi8f/0TSenlbgwpnGavLSneiYvXbCX5EiSoYN4qlxjOllFZx
XOtp7tN1x7wQZjLfn96CzUe39+p3Ub+YEH6LyoDObuQuUP83w0EfyHh4A1gYKBWJ
FR9I1o1oS9vatmfEtZNXaFnosA8sO5Mfc217M0fNP2t+tk9nSysgl2eTt782T9oj
rWHICbnPritDjRFYdksG153dkH2QGy7/t6DwHbAjS132rOSrynjPWtwNJ8fa+cU9
hf/G0x+DwRGVRubQyVQbjG5f5kRL8MiLCRi1BsIlIey0q7oPA1avU48HUDDdW2s6
p33EbXzI64mb0Xg3n2oZPfHBc4z/7X6W8XUFgWuOmiWI2nQ/a+gASrGdMDbTM9RN
DwnVQLYKipNt9n3YdAII+isNqxROGY6E+XQEB09VUSAM/CDFhUE5gx/rBv6HcUVF
7fFNU6ie2WFi4yBwVrUxamu/VB9Ufh1wbx1N3eQaASibeO6JLa/OkkoHQiKlGptQ
qhei9j6h10gc1vV09hscv2pTpdSsepy9AhYNMqu2gnVDnFN6SfHhn9HLswBt9gXX
VvbGZD/yT58YBkSJYUySl/uVxheg4VfBKzGgZjxVZAK/q+5/LoHmvP3Sp/2wU08G
tWE57QeG+rbSh4t7RkGgt2rgXUuf6VqPHBPzxWxitgJuZXmswlEFqQOhvnJI2mdj
7AGEYokpgehbIYakybU+A3vV2o77IutpGmRfcfYCYySD0Y7PlNhGt9WvG5F6PK6M
wUXlTnkWKcENB+14JDYgD0ch80BCxRO1UNsSrITZcyA+uFaF3RSyQMhA7jzfOtRY
zm8hGB479JF1aErphSKumHI+iRNPYVThprzpc0MwDCQ9Cqpq0TfSsA6zHPhPak8H
iSxpwdqF+c2QpktXGMTpXGOyemmwyrbw1fgjyMG3VaqdgbRJA9dBw52VDMFaw63N
+io+g/TbOSyUOMTt7QwpvzCgfeHsDrlWBnDeYoCzxhKPKMLmQAwkRr+1qVmtC8Cm
2BebQqlAUjjZmsAkvd3x4RpfmeKBjauAodkjkdq77fC3m+/rdkRpVxAViwGZqfBv
GYydxmSGuISQByLH4BXELbeQDqiAcElobJhxosMukjMhwRbqoTVuBqRlQP3+oVTT
cAT+eVdh+iAPN056xEKdugT9iqapSvtbpizzMmF6lJ+cKGY1A2HxxNVcbwIvxwf4
kEN4diK2qkzGtIeyduZHtgPhO2TNcjzVrE0Cq1NHp8b76PxxBpdsel1h7Y+bAoOZ
9Mm39xVjxM511/hJuI1tp5QF6oFYu3HXlwAyUuJ1dfjWOgJC0LA+tuBgLh/wux0T
AHZWWZcIHqjTqTjgXxGHY1CYbCIJloivhUtknBRMem2kvYHFzstAjVoOfefVjtK9
krNAJSHpRszRsnhWK5AE07FNCK3OKIXDep6Z0XtvesXneCtebeKc/mx/JfpbZ3x2
DvndTB9t10NhQCnxSc5RlMOE1LDm1BCGBoxvDDR6qhkkktBS874hvo+GUPQw1DUD
b8c86sBm+sIgE7JKWlATQfOgEnANDxXO4Ig7QNTg1FpPeMye4QbDyuNJ3Jx24YZg
xS8A1QQ0Ad0YtA3RjGeLyQ3V74gSqfONnrr+jX0/P2eqLSMb4ZFyl6ANbYGWMHIJ
Hm52X66XDB0iOcEaagpZqJgWt5Ke82KLKRYORl3MqqpHV99BYzJ9ck6QoebMHEIp
kG+uDe16tDgbJlQZQMnYbOhbLptKsxXXeWzeOgbNEhsnFSkC5Df1NY+p42CezLvO
69UqR205dFqzRzUcEjheLH8Ym+2m7RFaDYBKZjZCc69RXXUbk55Sbgl/9cg82jcB
n6zReb6oxOB8AQPtKW0X0mkrmsbJy1u12C8Z3PSsukPlmQhCOVrlI/dFg8HAUzXQ
hiVTkbCw4+L4hx4Y6Fsst++KzVW1P/wX4PSlGegXqeuzaQ/Mtm6JVbYIGcbtTKlz
mpsb855ozokYmof1qZBDERAiq8PmWglgUBeYm3oIun1yDTKcKtN+k9sk3ZFRGYu1
vFIvpMuoBddC9PUJ1+A8lrYOttP/fyh+SsklwE9yjhrBoH4f9Fhzr8NkvbP2R2LJ
vEJsr4wYAkDHmmlDd4uhMyz3UroWgBeWDFx5sOg0KNzDLakUdjS5ZLx478oqOmil
c2aDoH0BQ4jI7fVbgrAXEzqm257alwHJQy0Sl4xS+pZw+D41e/hAXOyHEjuOthLl
PX/cVg2ebIayBJl9ysHvfcIrLOLoeI55yExUQegS3rhHKtiXld1daaDAXurZwn99
uCq+/l51l5+4WbSlstMyUf5wahrC9uqaLcO7MfnHn1yT9Bu+ZT3CQmQEFTO7EUKS
Pb0Pdv0o8aXp+iYK3vVOpT/Ur2sZJ3zTZAKsAS4yJPnltsTaW6Ve0ILaeYLZ86IS
qxoy3+M6J9J4aY9vHFAm7tjSEAiREZO+n6U9k9Gv3EFkWLE76RaM17T5mUGFa6pQ
YPONvKTlldl6lNLjmSt1nrCuVjfiiCnztGNcjAyUwrQ7b8TMm5q0m34CZqPrqm6Y
nNVQNopwZGPBhNzgE2NSz/iX/rkWrijExKZTCyDBgR0g9BAGjvMOGCkaHpMtbpho
Avwgp4FjZporraC3MHFf2gvBTJz5Yz7VoH5HlJdfoAU8r3XnEb76MQIp4hJsi5/Q
5FbTpau4BfnTKsSMCTdYIBUKpEJr9A/t5/aKKp4HOT5LnjXAvYSfUUeKB+CD0mp7
lD5vGy93qGGe4uKwX5BSjRbgTQhIYijewvC+cazZULqWTM2XuW1DEDgPytLcR2XB
ymbhC+tB7BUKQSQCBEMj4mco4K0b93KSvE6zpCeYH7ZEPq22BaAZm5MpuZGDIKGr
tXHFF+qtnapaYitJii76KBlfqveQGDUBMahbAQmRwa5txMVM9fz6MnwOq7sPujN8
/aHUAlvfP4CdhsJ0QCtBy9c8XTvoe2Hv6HoGw0Wx9tCOrBghuMgSQTR1kecGksno
rFOvVCrba7b2CDVWbviQZTWCT+w0ZuMhPBEvyRZYy8IfrIsk7zOq9kUBgT0vavJ2
LKCI/lEbrWIfz33kLkh243iMYZZBDH4eRX2IlFujh0LMm4JjgR87KGLDIiI5hVii
Za0AvXWx4DRCcv3uY0huu+alxA2wTs2RpMLyx5MswWcAOKAORPohtAvajPemkUjg
exQ7c4NwQ0xoYEuB+yiLLBMB9Wh1S83kn4bj7kWVi1cp7ThGqJqSHeDM8FUKlIPM
nAfAPAgVQ745UieCVgweP9OGL9Jmal/BrepcQVFo0fZs9DiyV6JXpZILtnYefxrN
JP4RwfIOUEsPQRsYuHXWbxuhXKwhJNMM8FPxnRoIjZjjpJbXmuVDBilNHERSpJs8
jBAZcHIsi4eVZvG/8Qg2Krpjns2bg6EsmBR4zR8AXxHB7Z2V4lVg7cnaWNbtJ9Ht
DeOH0ITx+1O6yG/+JNae/meeB2g8rZGWyaZYO7UnUs8hw6cGKavXaTBQpuas3XZ2
gZsNqTvSsbyQu2JKg9UMTEXyZ6CP70Ob6Mic4NTUk/MsJhkXm7eEpJTqm5XaAFy6
AAghAW0JB+0PrqXdMb9+ft3XQMlo8tw9MkSFnN9iquxoegWL45o3w5GwI+auc2A+
4rJ/1sG6S5OF1przaE2AokNeSFbB5PdjPnPmrazLg7pfxkNFtoiTNS7L/q1QYZbE
kEY/SRY0WyDk6Cr3ENAm7pMfMNQV7NKfPasVo85ONjI+vsvRE0nheMvlq3wS6Wui
tkDOPIOk/MatDPf1D/5KufamC7dXv0U1EOISYQ5WhsYs6Kmi5/ygQ4Sjp2dFUd4/
qsR034KKZL2tSDYYCfRv7MlTn2HwZZiHDYx/msIRyt5ToHx/wovolmKffY36EqfP
MnFJ0FHgSK+anBDq/N6qu/XA1HWhocI6UjFy1dfRsDt7HzAvaucgFHB1SDkuL36v
j79c6tFUaDa97/axlv9+DEIckBALYijlIi90pOBbIF8jFnZ9WTD2uEROfh/ZoevY
jtPTqFN2903VS9zGk4tnhrRzmqOA43bRkZxly2G9RkGbVB7bze0JeU0JT9LPHdu2
k0WOYhl/eQPJa7x7WKdQq8YhkN1fR4KneznKItXQPulLu750/P4W9JnwOyzEpdBy
3eAIjxXgfCITcF2O+/cDuWYcHba65FcaROGggImTYWEDW42WW2vIl0ZFph+PExP+
1kCCK6yNirCpMP0bE2AQk1NwBUXTeSR4vvRW/yDvtfZPV2Jg/+EFbsa/5PUA0xTC
oBNpNdkJ4vr2dwx2bmRmbztKg3ZVsCANqSkLitHVPWy/U5phkHqu7cluSPOLvj8W
ZhOIhDVQenWjjro6JAcGZziBIUNnk23YG4ZIC+BmyzSytt43DUJgZk3/54EhXld0
u1H6Np/RNsTlRisXW8UFKDxocIPK3IO/Hs2Tq6ALu6hLt3Gh61PkdjiiHLY5jklv
thJ/WAtSeLEnLxPCubUEAjQEnBh25Nigljml8bYNJ8nPyv8PI54ZMjbHi2UyPMP5
w5iH0BBlCm1e9cXSfKGtbo2ytsoOUq25btWAgtIbBMeQqHT+SFYpYqZ0mQ3irJbB
w2fpwCPmNs8+ahNyq6Cmrd402/90HqxeLMD5KkH3uc8xaWfjkkWMi4XG1cuDLHm7
q9N17Lodymw3ogU33IgluxFA79NR/PrGD1nkSM0TQ1MvPniqf9wrnY/KTlYhkr2u
JlZgKgc4glNHxE37bnnJmLldObBEUmIQbLxYH31WcM4m03ByrpSN7R/q4xpma0/Q
2W0ta6fFSUlDLc/fmMFytfr4JjqmUrNryfdAcq0LL0VTa96crLRRYlMyjVvDp65T
xoYhJWIv+SUI5/NlypET0Q7M/uU32ojGIRpTp8FMwOxsPUVrIPZ7xwZMAEw/7FVs
PoZVLOAtD5CfMfNlg6M+MrezatqvUyozKQiXpbtis0xTDnwAGEsiuPExYfRg27n9
3xugcm/G0lQ08Sm5/GDU8wLyH3KVN05/+wZ3hO7npn8kSpzUhB6hLgtHpSIqOcDZ
+7EBNprR/EWb3lKaQAZIkpcH6mLXZUGjDhxWtR4Av34XMmlE0AfExwsL0TarOxTM
NUUqmyfF7O47vWIg9Vj/IGMrBeD57KxiO84lXEKsqi3uGVCPQZ5q43+e9LWDIqfh
Xc9JQNyKGLepZ4qDXKatLKJQGNvrRHKDXAhP1AiwTao/Eva2J7AZxlj2D0E0n7c+
SinzOWV4JZPtw0hLijwVVJCVC7EInqhvj/3rKC/arX3yckNvb/uJY8k3JYGFgMqp
4so47ar2mEG/IiK/p+yvzPCnu7zkChlFvj+RJqKRIGReU5Y8NZrFStFafQqmgJ28
HRwfaXoH/n5+l3Gf/SBX9kAt4gVVuNHuCmBbq/vysED1zeCMXNjqpEpdb436aQqZ
6suOtYQHHBDSAGDg1QXq8hz6lpguBnVL+bNwSIm7VrFUqEGfnY0vFli8L9XfqU3L
Ysjj/BKGweaPgg+g+fxomNfqwabNNpVtbGZOOgwY+rQlhfkaSZwbwVUAyiBxWvwx
MJObqI4UGEVOzDStBOWccd3O/5zguAU9+0CIi7OoG02VimKztCOIrKS9Kn1swTy4
uNbVV6mPXnv1M4fN+fUsz3eR0HClZXCHOmPq7EEGMFddb9OdcI0yfKJPCZPl588K
JyCVhmtzKsFMeDt7+5HnT/wKzH5SpfdSrPL3n+YGlhPizjOdOt1WpR94EoeVYwrW
6EbcCLWUsFptGUU0Ka3HxW+TGBSTe7D+iR8seovV6PhEgwlxbRJczBADZMTTwgay
mn194pQYs8Dbb80pJGI0UVCnx8zZI8ELKES9n9bMAUwNTWIsrLno7qGcUkUD2Bk8
Peufhiq3CnCTUhHWvVfW+neVmfUDMBREQNBv7v7saMqYQmuGrLKMp9PMWTlUi6Cu
4gCeRIxIvCNYZ+2qz2224ZOlg9ZnjoOrsbdT3eQefW3H9si7r0Y5qZWiwHNt+v/E
V3VeV6UiNq8LlvHJJfcKi0J5bF5NKcc0ZY5b1V/e5BU1pDuIIabOxhAm/rdMzOhk
nB3jTbfxC78cOLdOoXobvG4STiW0XX+jyutOIjXiyFWcSvDpgsQ/JINf3SIi3b6X
BmsdJqjGNSJVT4nxWb0Dfl9zNUOOq1eglzf/mkxMMs2YuRadjQe/DMpwiF2Br5L1
OumnlMY0PFaBUkuODgn/wyIb7Oxlckl5x54ADNHQrGmnseqxpOIBMYwOe9RoXpgC
VQo/0mgNxBC+fkZpAUmwgYp2qohFzdoT64B5WhC61LYEpGQvNOd58OjFX0bKR9/l
4oFwbKZvK6geD7jtsdsK6AyIpg/asO4T8Y56Sxj/1gc2t9ahXIxX1y4TDSfBdbUy
wj2cVxiZkVJizSBYRaVJccJ9nGmiYCCnF2NSW4LlrsFB0NTSAH58DN6IdcCDu571
Eja6a3YQioad6M41zOOewYI4T7aBFjWbK2SRR3Qbnxioi4YhMDNg4DNFIHbN1PUR
PQX8TtAzxM8J5Wox3h1S3sAXXqCvA3ab6mWvkzYM8u3ZDLaFBBh+0PLs6CW4P8sV
MyKw5oLRYJzlqcJzpBHLcxbcrurf+cgIwCbTawhAfw45grjKNPNYKq1Ao7KR9URD
pB1XDVvAAcfq7DWoiueSb4WlLWA+2IHotjRNfMrYsrn6WK+ZzeQyt4MQnGz0lwNF
XR7lU0VTXWrdSnEJu8M+3GMrhwKa85CIKUoKye/Tn6ILaM1vbhglx8bRg2CkDL7t
/noUHGjQIgl1WuXCtVcEfODQMtZUalSWULiID/szFsocNHeLpVwke4nkiD9Bg9uD
CalAyxwRo952X7HXQFeCf4YPUBGtSBNM5dG8RqAQENbIj2dq69K+JvqfSvQMRhct
ccjQ90ctExstLHGiwfj+w0K/Fbgz5ezYbntB7fT1uezazxcFVipkWIDCNkD6eFfv
E1v5HeDjHx4aPEaCF9XUqeQEBbhzHk8S2qv3vYPI9gTveYBTsNdox6zgYFpni6/f
QeJdKH8sr4LyubqaDLQzgiX8tF/MQf4bun1xmdZdTPo66wTxju1y6EUiluNGMD46
ix7avZifah2/qQsamXVMMfZqpUheKcUwNTBxZnilwXLhMGILpLV/pPVafdtvlgUD
JndjdRUI+O2F8dtvQmMmSTyXFuWHMZU41lDNSBXpwDRz+ZqTW+w0lYmBd7uw3JZf
Q/kyh7JfevCYUdMjgkNoSdeYvih/jnvLqNN6ZL8eNH/Sx6XZ2T9Vzz4RYzozymZZ
mkCXd/lVKZiEE6A6k4GTAk7XhuMZgatLaOJxGiwl7XG49Q1mBqnsrK2VVqnoHBr/
CnBrm80z2FRwSI+6V9Mmihc8K8IKPl7kNubQgfvtfU2A3TV2jr8b871W5u0U0em+
2b0anICOlUMf9Y4GR0H7vcSshGdABN4H9CKe1Qphceg+G3Q8nDGGgFS1OcA9/bhR
2lauKJLiMV20vyjeX1dfCIpFFWlEfxA8UUSsbSwXwVhQ2wCQAa1xPlinDl0LzUAp
xYQgLIRqqUOjLLT5OfkkK4z2wsV1b3QR/Ni+NjkMbHsLMGUKbRhfy9SA9EB8DsD9
hZDqeAc6yBxsPI+geUWVuCH9t8PKkZMoS26QuRxBmj6nS+ECnYJ+vGNK1XCWZDQ0
uBLEkhzYdyrZ576MJ7NsUEn3QXb3AdvPZ7uHkGQIyBbEorsoFPjJoNirqGB7lvXp
BqopjoWvLIY+jTh/Ttoad+HjTsH44nhkK6dI8OvrT2BxHYitNd2+WvCp+h8sIxs/
EQFxPWj4ocajUiPVDXLLnD1zfHx+tfN/0kCMl4uccAOVb0mbWRjG0fnIfn/ClbJh
LwepexHThuGBVb1ptK0k/kDS9ir+ICtO10FTP2lUe7YCwIu28xgemXe3pdM/Yi5i
/yhs4gIZU9vO7Ju6CV36a5vcmSBpFsFt5j3PVmuzi21+0ikaUTr1Q/QBkQAY8/Y9
TwN15NGtEl3YA7WFD9hVxnxN8jSEqRGVmhbvmaxFTyHjLUTVlW4OGYa/j795xS+R
HM+ODRUku3XB10X2SsArQd4a6PYjC/0wXWqZlm1fVJ/Sv5j5eUdBUkLFMj/4yQ5b
cIpIgy9ejVcqv+qGU24nbHympJlTg04Ldpp/X+sVNndvo+zkdvpPXDMOQHQw14KF
mDtmRNttQxf66tUYTxsj5wITQVpr4v8i/y35DEAEU6Tj5O8dhc0hJ+rh33k78NkB
79oJT+qPt5/vQqK6qxolrC+skqxgeSNsDrd7u7Il2HLbE3lOJAJe1eQFPWAOo1oP
RVCm1HhTFEYRygJ4XYrFPBL6cfMJSu3eDu9g9iAtJe8MICfBVDMt/SdBvDy3DhXK
XIZssHRCPqyyWk5k77LXeV4yEEfBWQUt3Q07dOkCgXE1heFIfI2fCjW0AftaCnKZ
kHQvr5midhbXLL+z+RbK2oIvQECc+NPo0hTlWihyhpNAFLHyODyyXvVM5RenQtVd
3TiScBHUIntp9okqFeL+JGDaUKZJztpKSA5DlLcJiP9x3zrdk6HUR7z2OvqQq5bo
v5AYHQs9vSWyrF2O+rmdwHaRNaNdgTTIBtCh4gAXAJ/N1k/QdhEy53u0kS4iJwxd
cKiKnPtWvfwWxk1bftC94z+Sto9a5mTZrBdbl8AE8arUJiP3DAgshAVweYTvCGvI
5jpbjUsJBIXuqqD+ywuJzo7uSCHD/GDR5VhyOS5/DB+6L7LObbAS46v3+sqy0O27
CfVLTbGGGjGInCPIHP51K1HFxiuUjHqdr0RLYR3ipEEKaCH3BCYOqTeWyQUtOWIz
vlRFNUx3eqa0GCajUk87M81pTSzWB/aZ/2WiztuoDdPmX+1fowC6X+y4RbCbbHht
gDV7Y9u6vJCcwkZP0i3k+SUrArFyjgcPMcY9hxrayeVBqX4bDQx4qKMoe7dwGOs1
OS9MuT0OCRaKKZoXxZQhqKHHrk/MCOw8xz/BiWuh2+jPQm9tu6y9JqsxzBh/D0Br
c4KU2NMoxyr6QMasN02dd+JBrrRXCCdNZkNRF/sg3K0Ki9FAqfFABIPaeiXJPBsq
3eaZRk5JA3IzQClZijh1aGl/159+PvfwiSlMT31yvJknfNk3MUjyZemDbKmI0AjG
NgvNzqVQ490BqrTVNf62rxhkjTKb8iQnHPUlWLmw09WxOhN8kYonCsQhNArHxCv/
ANNyMipjDjinvQ6+WB3xkoF9TWUr3TpRp+7wBWXrlKntGQII7u7BdLSaWRHWqDiJ
eU0y6GqE5GxCQXQ8V6vEfCSBSDaxRQAzRTLhIn8LsRP2cKWIyQ4y3bD53TXBmSaA
2HCP7qJ+/YzfJWBa/YhouYOGGr74/43aiJvvDjlCNdcfA/Nc0tlY5UYZK1BiD03n
lGCc5kwDLNJ2yVC+J7aGSZCLcNiqlawtTjXHl1jXI6LUFF8gyzlYh7ieAEzjMBpE
8Z+Ag/yBc/so2bdQrE3CsQV6zsBmZFIsBwN4wfDI3X2rnMzJPASsGzEM92XJFrjs
VsIy1uKzza3GKa7btr/sgAVU2070KMW89Y1kRSplvIuf9pmUcxdz5lIJY/z2yeHJ
GvsGVJu+YCqevmu1lSvg3Q7v7GG8V/3n0yZPCVXSq/DQaot7PSSnPt9hoJV9Kahz
taUU1lrEdhgCZUMML+z/mDD4Yhu6MBGeHxC92qnsGK8ZNmlPR93ueCQuyPwldMm8
my8KQ5KFZ8F3tpxCfxN2yOgzM6+IqUDeJi4dd1pOlZ+jJIxV+wDhgR7TS6DWrwyG
hYBTUFgcipJvBsuu7WIJYScDIBQMtPF6/Nl96k8nVi/DTHCXcCgFvZLnYhmSY1Em
O1i88VIksehav4w4UNkKtT/zmGw2baln2VD1JowqaA8QHunfeXDYqKBkXJzas2Zf
gEhj3i5dV3zjoCzqKuvGrqdzrj/0guDwIrJu9XhmuHvaagOF1t+vUDihpxIv7zL0
7YXziSb0DwuXnYZdmdFHmcKF2BkA8V1U1vlWRxL7X4uDVGft87Mc4aBAMMJhk0IQ
yCzHOkcc3fL0fNm91sbNreSMVJ4SCUd8SkaW17uzfmG9M3R2yPkkVpLji6u0Qp1z
sJtHNnPaY598o7dVLLWOeeTi7NMIoHrP+s6/OX/Z1ViaQf6anNXT37a8Cdf6vG+M
9K6/KX4JRQODYIcpREV3wSvcW8R5+BrhgsH1zDiooBIeCizQuJuuNF6dDVt1VA7E
ascHduCIHML6fqCqyXTqcbawN0+DN1ACSdkstenvLBGT4+ixJymM+gnOlHve2owN
vBxgU6YTO3HUzVvX0DY+e6AkvqASj8VU61casZ9K9D7X2B0VSJYbf9K1lT2Mpr8k
xU6o24RNz1bzxcAfuAe1KeiwnjuCp5z3UVmymlvlLC6RsN8pNMMcFN/Js03hjV4T
5Bqvy7B+OVG5XNkTCokYVXRsfguo5FBmg2AST5InNM/UCmGB5gIgBMegYDeZfNKO
4EtIZrrrVA2hL91iQGSHON6JUtRutwwtfqBBLVPwnkhCN65z5Uxdl7y3VVPOxG9l
XrhBOFS3LlhTJa0GP5DpCiturnGir92Z+fBFtWuWdv70NSbyieiMIQCjvBWYyc5k
RN1ps4PWoCQENP6PsOXRb+mmQAwdojMyFhW60n0YQBtnFqQM0AZVD1AUmrSkeLVg
RRVbXSnqv3Ul3KhtfFptJDid/Svn4qf9BQg/YqV/t9Zw0YzcEdBcIWyGMvBl1qBE
2L2A1C3coUqWgEh33e2dXWhBBP7icog3NI6M9iKlNOSkbSQcrPFkRM5xWUqHih1+
yx86DinaLgU+rk8/DlFQiQ/EJXbfkQB3mK5bmPeFmfAeVfA+FZMRD/3BOytxSbk/
i91P3lqazjynDx3Hqyv3uiwC8rYSmM7csnIZOYYZQ+oKHl/R6kC2w6fQtAQL9/Op
mE8+VFVBw459pYexhjst0oLC4E+ZJvX73IVrqeuaa4kwc5V28HdxYBvpKWN0+fvI
rrDeQQyn2bc83uOIL5aOMnoZKkHNRDDdZAD8DkWdhcU/O/h9AwXRdIJsO8So4upz
cyGdgohiGiD3N0sGkp0QCUwP756tPi+RdcuNAXFIc5Jx7bOo8ox4tULpEvuf+AZ/
oVe5B9hPd9uNeLnQDctn+s+17+0vqSXfly98elmF9DPR9LchNUzuESxj2OX6rJj3
Du8GtySTuC1+kruU5Y6RC9aVoLfPgo0Y/X94WIyxyQArb1ctrjdeHlt8kcht8SvX
D48RarleKgPAGJMq8I8irnX0+OMA7PLpdfQKjIDT1YB21//6LFeRbTocEe1yGPde
qj/UA90mQUcjzPfS/gHLsQfSNNgGP2Xv1uWVqrnpFJ5YKTVNU1AM7MhmYi+VpYEn
wwjSFAPne+5bcIz1iJWi8Hu1tSraJq6Uc0UHhc8vTCxvr8+Y/H1Vw2thhNvnpsOc
h++XgYnP/ei4Yp8vKaEIKh3NYbQF3VlUo0W9Kukv16uMKzu0NVXFhoi5p/IGOSFf
iZ+8kv8UsB+Kefw3FtkNRcHzZSMMRMSy8CKfYP+kePbame5U55mJdwZJBL7yEiSp
RIpq6t/+OOZHUVTcLRxaT7I5h5mELIr/WzfxB/DYYwYhIEwrbspwf19ARErjI1x3
pxM0wEU8OY4kpDvlVrCbeJhDOZrRLgmb3ULfgFaI0wBoSJqPA7cZFvsm5gUCBaBy
vKsMkq3ym1r9zfNza6WJGtFu0UJxTZxeA5ifMP7AmfVHkag3qMDM+qxEbzMev+ZI
EcuionmTavTTlgAI9dW666qEPD3SfZuyMOjFnnxqiVYUSz7213OVgZiRzdil/Oxo
E3OoR1kVAnUSZDU2UmKQ7mi49DJTmLvPSj2yJ36OIrIQv9qku5UmC1iPr/5fZQUy
qEcZmnmtE0AATRVATJh3iiZMJrxbC57im/d+X+SGfHp77kG4MXAJdk4W9AZQX57A
dkGvW9+W0/FhrjHth9vvcWJynG/tGTIULzwmxeFdRFwbrOxV31i34zAHcvCdlrFR
Y0Ebqvjp2MB/Ks+bzEq4+PqjdjxuKwOwNlk0N0dei7/Ao2hejBVnHLU0vPGH73OU
tnIFwF5i80dey9jNPz7P4eyKYBQI5g1Gon5MDneLzrSGcW9gvOxKofvrPNiUo+H3
EUi/ORf+5anR6flwWg7BQtf05COyHmI1rHgO/djqjpOJaYUvZN2D9gYcRzghCyOx
/kn7vfrrOhFUk/3WNbMdpTPHlp/aOIdBT5kQ9fLiYBpjehqHlTXtofEL+fgsUWmV
12B77fdJ9cyX/KGh4idVVC/Y17AJAOKmBccqHOJHicAO9MrElyVBI9gAvGekgDam
dg62xCZydAVfwFmJ+chaP5lml4VNvtjScNyV1gs2+w9NFK/xdEhiJBfvsMCfolam
YLMbCLL9GQB5HmRdF3PgdW0hqHszcish/oh5bqncchAUZAxRaXFlpaSFu5MRE7wB
nMl43hYt9F53HoVZtjvJil2/Y+r3PJXSyaqhmkGxniLwJFRtx8I3GzvPEl9kLGX8
CXq92LWrfuW1vpgzopRXqNi2Ps74hquyzAoEew+MwR7ekMWoypVVPkbAk+8l0WfA
LWi2Kbos9HiWU1qR+AzarczqfiWfqtBC7fY2QmmkBsyFujuYyzuyQVBKaWhG6hek
Z2nFfRbOA/IqU21d0dzEHLCp1+oCt54PZOAobRSJbmAppN/n1pogTfM0ZErj7YTI
OvZWSzShumbD5alXm1qDTNJKgki+UYbYVxq0Owunnpe86KduQxNsgK7D2XigytXe
gueRXZkmTopjswbGdniHCV+ShajkqA/GP/dij0LQmRv/Iwzw6v3wy5mJOeYNFov8
5TXKztzMf8oo6mwmN+men8OKuVQIWS7CG+5UeNVLLP9+cFhLaESA2hhG5lc8ehfq
/KYegCRA2kRXOAzr6TqB69I3wTMORorbd2EDRCsJPwiw63zDmRspkuvNWKgsAY5p
0qpss8qyGi3uPkagCrH4ncQVyaUiq9HuZmVzNYjg1MuOyt+UlENwHQc/cXAjfHUq
+9JFAWRG2KEGVh4LMnFUzHrBEXAF3aGXfSwsscWmnV85xrOv6yFvrFrXNLNG4UvV
HQ+TX6w1ZlryDgbl0KApMdi+dfa2bbnQ7GSPea1g3VwTKMMq6+tBSsRxQhQ5l4V5
Xxo0RrkoT2Ypui8qhVVi2kwnTGRAqX04n2agG9i7xntDpnEpuSnBwrkonmnhA0n3
mvjL8+IIfi1CTWWR6W73Hvqj/KCHr252qN9HrLku4h984y95H8L6hfCgqZ7RhMPA
RXxIejckSJZPGSg520zEW5ZOv2BLKm4+xQ1nVgyQ4qfojI9qRuRKFiULvuU7CIGI
q1DFfzRAilWJ52zu7MscgYEbJiLhgTfElAxtr9PluuMuBGLDFiGCmOgXii/aMfaS
oYu3F8KkKYsVBdyLKM2NVjEn5g+g1qBodD+NLLqqo24sBVMeFWu3l5mXbRA5602Z
RBU5sUlD2zE8MS8TqNR9bkgqpTJcgVZh4V3F4oK/eGiN5Or2+qP9fCdGS6E3/+3/
1mEOWQSHtR8GEHevLU955JfDkpFn9mhrbuGHqLPAZCFsfB6VZzjy+MOUrxy8lkYI
70H+RYnYr5iIlhtWwlNbb/kHAmAsVaT9r92bDrZbPRymIxEbdAOku3ipVdR+L5ol
6TZ7Jm70wIikG8hIOpaMywgcKzuaifEqN4OU3NcDVnhf3kbyMi90RjRmdh4cY63u
pxB2r6+vsNjguzubw9SvqMyQB3eiyCcRFzPmwkbijbfKUxQHpSdefbLF/JQTIHRc
OsLGO+9CZEkUw85r3XIS7FyPqm3Cx4BozjEdIm3pAGHRWFqMQVxMmr+H9GErhKYS
+VVw7MlcFebw7FivUBrFfPNBBLbTLPvAPuu7BCk+pSo1LiPdV78BpHoavEvhlCtR
S2M8ErzTmivMjD9A47OzvUIWCPKQ+5Ny3cLbzop5yVAfDytsAmEjAsDGNwU1q77g
cqD2Z4gQbktfJPIdDzG9O2uBcQkOLHtsZZrm5bg968BBdTg17yUjAG5Xt1x7mTiz
EZE2A3TvNdNE1MOj6iaxHUUhAczTBh9lIfuPW3s22kSgC3+NP1LFiNGqRyupKyqU
SbDbNrRt4atPgjayZdSOIlFPrnIUNqDDmxqlSM6n1ErEDhBMn+ez31JYese37Src
9Eammujl5Cg85+RLp7Bnl3v2pYKkrSKGQaXa3cHeJ/qBQn5il7/YP9qRusp8gceY
3sfi3ih46sSpYOnz8qbesqpYIkrv9RVXIlqJNBbSZuxWVtwnjRGvMBXMoNHheU0b
kV5Jr9+n/1cwPPIbe2EEQo4kMaioRpEeWzAncMorc1xIoKzEMALcHTq4k8726kt2
nIn6BfJiSfSLo1o+mMq2ZH/HsNPj0sI49NzDQljtvipHa9M+8YiO8HQkGpB+FksI
ZCbs4MQu7+YukWwudaIPuDnAL6UDbicZ1FhjSPBrXOK8EOWW+ArI8HV9R8r0MXc/
c9iPFxQQ+dIjgvGtTvN1ZtBKjqwBtbzooe9GVolOsqk7TpGWQQa1TN4gX4GfJjeB
ZeIkp8cXb5zNjsfOQvJ54JEoD9rTu6zEcVPTXLsvh3CHtAlJZLn47Y1W1SWmeBZG
Bsjwguw5zGK9PBLTh1raZy3KeVP1LwoGGsXEd1rkYIoFnzQg2dGzPCe0qqApmhza
0K6Yc/QMSwWDfZTi+B3Jo+i+PIQAPsHImMK+lWesfyDaNcYVq12ZJ023WrIyrj4r
WBgWck7+qZX8uIzAi05lSTjf3dZJIL+dfhynelgO44RNGCwFJvysAH+/FaI5ziIW
cbCg/Sqdg+VJdEsfUnwiX1dgEzClV75fbOmPsC3vOxpK67J1jMSIS3bCl7jj5Ic/
NHKw2+Y4vzKilVZnrmSoDMJD/AVCmxh3kKbaTvc382TnAOGLr+TqWLqaD9E4dm3a
HfGe1pVYwv2DgJlkuNii6bw6GW9F9/MbHGFAzvqtU1vTPVgixYCN5wv8hygfmMh/
3cSx/mTeEKqnYf2Pawu3Bm6Q7L0cLcICg9hoswRmoUjj6Jd2ehc/pKVO0U8oZWN7
QDmJ3vBwpVpoEEyAgdgC3QCcyK7FH0IdeDM3EdDqoiBkmj7uCkAQE63ozro+uS8c
gPSYetiC3Ga5uevDnHgNMa1yWTyEvqcescl986B2222jQWQG3hIS2yNmEzbpBWsO
aen0qjrt8ocSegnQeNJxQrr9L9YEFFe8fdth1GWIse3biFAbUu9DKDZYM44gGdCh
2HRjoevpRHQ6ssE/PvQK9o5hhPTl0dNot9Uc/EPyhy2dUjF2qi4ALpfwEQ+9Bt/0
CgW+w/kUuws+xrr9+igfaa0TlSSCxsWiL3HOdTq9YpxySmbL748Jp3K+9qFBumOb
2eoC0pImtt9crbPH5g4FWHS2jugexjkuu2qzU1aT2IWMFN99gaUclzSKPHWISG91
zsj55O7ubn4Y4mxwD7VnAzfLQnEiPimhWVraKrovqPFuGTcxn0WFUlWG46OaZIga
JjYQomXbQZigiR18vyqfytOjOLQtGsuvDgjIkOeRupNM9VmuKIf5M494sca/n7mq
XpOWcIxUKB3ZcEfevwOZTG90Cg7UIPXAyPBYoxdg1DiPW5E/Auyp78CsiV1PSBBr
Rig6Cz/9/tMsjBx4P19pgonTMYsmFVdQs5rH6RnIZr6nUnL31J11tew2DFXJBuMv
GcHlWBVe2OzL87f9Fj6eH2VGIpiwblhoaEPURCT0DhQLIU+d8NZerOAPN6SfVI8J
/z6K6PXxfj3EyTrC1+OyoBK8wKuUtibctfKEj2ssPSe4P9yOdyNAoTxEfoJ8BzTS
c4CVywLLJpUkDxwP6onpsNvve/FPU7zf5em6ycTKn+f/rEnewL+CP3m4CgicnySR
tCKlv4pjV3ECZbuWRNXTjxBO4aVbJPXCKtwmeY0wB7geKXbP4yMeFoexx7FMfXAu
H5C6Synx/CQdRCOQM5SqAN6gde1ON/c9p5LURpE6MmXku+8v5dyxRJjebG1WyDZM
CUdSlvwDafTH46Ho672NXl+10nar28XwQfg/EJDLQCXUhyff6Z81F46aw9oRamDE
Mf8qJyLMdxPhegNN9Ykq2VxemufRJLEjYjuW8oBgVkJidFUNao5v981oeNT3CQ8p
Hm/qa+0cAdbKfsSfxNGAKCKeYBqqO07sgZxVd2fXicjQcW4/Mbl4f/bYW0SME7qu
Nsx595W6zK4yjlO7kvAK7L5uDVH8ZpLcPO1VsYi1R6VPMbb2rsEUOeKayPiWsO3n
7gVWuOjjtR76kCEvynTeUV7+IG4FtlT49uOBsbSx9L37a4V4MvJ0mFQhd558Pqxr
hymAkuDicuiGPCe0GILRosgtTcL5/GyNu/U3R8c4SQc8G4KasUoH865RGKXtjewl
Ves+ELibYLeXFfHN7Op7kYrqwFuRo6MumsUoC/gwp90Jj2+x27hxSvQIcAZYwWZ/
u3BBVe3mrbk5Mo/NkOQ8FrlApXUL5vjbQ8PGx+42FSSVZRxqxANQjGzWLdP5RYgR
PSoWl6HIz2dcjbUUwX+jbl6KKipqnLQ+jBC7/EEWfDoZKtHQ5f/FBQZZRLa5Bggu
MMhGQ3QkdFd3lS8JUQnaqh4pm1bskWBCv5Q9aZjp57GyPl3hZCd1LUV79k4GcpJ+
k8x2ZS5qQPwd/2hBKlMo6P6RU2KtpTtYKAhrwJYvqaIna+NNd3ygEnJ1VROHjGin
1zTQeREdBMQv7q83mWZv7uDzFQ9Klwk8K9vK+GH9vUxbYA0imJd2jZbXZPxASdfv
i5bc5RnnAwhLH1f0R7FTazTpGVezgT/hig5zoxAJxHTn7regieZY/BMkEGezTXuR
3wWIHV+ik4rgPkFcdMQB8JbXtCkEJMAKJBwChtkk3BlH6LqsyTlY4JUNTR+PSDqW
EeBAt0E2yoJaq2TGeKnnAw7bvL1DZEbRDFgZ30K3lSMNIy5OBvghMZ98dTZDsScN
2zMXN+u4KmNyBFmrqTGsMUufu6XuiqLeoREUBBlvZrdnGf+5z2LqNPQiiu7CsOUQ
hUPfUsgnllCalchKK7ubCnUKcdwLTWIUzWaZvWhhrhvevOVQs4vxk+asDn6vablU
aIljH8ebsNf9vtgrjGfF0gbz6oAH+DHuZk1R50dlQQXIflqzPY7/dDYlFrimM3Of
V3TxYTIY8zstGCN0JEfaysAdQtxbDhEaXOxh//G3cvqOL+aMwJkoXJo4cXvYfhCY
hR7MyqR6n33OLmwstuB5SJMhm7gWrPVQjRoen0xNhXPLHn2A0KkEt6CRfFJAdU6E
91TR0+nBhE4M3+i2adJlrzUp11qeNBZxRLvjoMe4oT1jPoGaegI2uJ9vvtdWGwak
Ec8p6tWdjkPH+iy35N5fBGWA4sL1mANKaUJ9IHWyxZXKHdRiKfd+uKLl6+rmk8Kt
N3hxxdAiQG7S63DUqOfiXBT+Vu4k/lZQKt8vvPuVx6xst4nYPiCISbTgA2J5zKHT
g2El3PJE3XExhz66TDVohotfjXNJfIbUfmcHU7QWkv41hu5TkQUMYZaRWxE9Cv2K
+NjU2agvi55YYfnfeAl/Rgl4NC7iTjzbs3iiwUuXF/yfrffTJb9uk6R90K2MPCfI
2U+YyZ31iNURF2unNlwZai/y3fz01tMyQSrFAUHO5T3d2aG+Qr2WsMJeM0cheFkp
2D6XVPurOPvi+QwlvD7Jgu1panNNjugG2b1ORsdEqiyRcsp5C9VE3ZPKDkLwvJJ4
+21/wK+1P3+bxpFBeYXug9xAu9iDoykSd1c7T+fHhyNBLrCJXfiVbZFOoqfIv0q8
fSgJ3w2MKz4DRgPkmLsm1VUAu5eh9HRR4S9r8tfGbwTpmCQXFIQsszuVKK3DswzA
WcBWLxjwBqIkuo8d+/jr3AvtcBZJk4JHuKkhrI3qEp8GoyRlr+cDDS9BtuWuXMbp
cagchPlLc4P4MidHZ4R4uBfscSRZAa3Hm799QSg4A0m04cp+6qrlzMuugQyXcR8o
ddYrVW70XemTiN8K9AZx9hdnqeW3sVZykJaRCUB4V3VLHzh9hBH8qGP2w7c2LTZg
0NPVsWEm0c8nh8stpG/6oeQffkwIk4+mE3xFYv8UGn1hgjiV81goBFM+fImAR+QU
8UGLuUpTheMRpODRZS3Ms0/GG4ArdP3LJxM2qBE0Ok2+hqe7NSaJbYHVw3Oq2Nxz
Nkc7/fFHySBOk+aI9x/U3HePRwl2XucMF+rewkEsNDwm9lvhLypw9QJzMg0NRXEv
Ewgb1PIsy1WeMPfQUlxDrSWG0EpB3H5v/bXiKHjuYAzhZvulAltKD0U4ea9HGOdv
kIOjw/+rzerD6sW+iNqiRDmszw6l1tMVTVlpQFjIQqtBMZRfr1qHrBIYB4LDA0U8
4IsVCfZ7huyMwZoHUqjOat6+VJW74oYIv2FuvYfuGn31nbfB47kDqCXlL65GMs/t
4BOEbipjXqDM1b2zHeSsYbqPrJwf2firSvgkJwJoOFNQDsMqUOSHHB880tJlTajf
EuzCQs7N3ltxZTqCnuxqk0xu87sK7LHY+ABE+EFPs05dWDncZU6jr6m9oR8JriL5
svGUsHhyS7rdFQgbI/YPZkSQBkETIfT4ANXpojbPhwpdiCrLqq+cUp8qJJHNsV4/
98CEOQaK/jE6C0qiR7ul8C3DOJgoSlQLWeN0svB2b8BasU2x48NV/Sk6VTnTBJy9
R/NBZZiPfcZZPWfLLN/J7Y0PeZbZpFAhW5H+41KYqPfaTvw/yicIcZ14kuQihwqN
v/+A3yhN0S1m6xj4DMUMLAAXA3Jo9oLaGQXIIj2L0k9j72NBmj7H0EclLA5Gkk7k
GUMpfMvoB/DHmoBHI4D2dBW/JwUHMW92fOWsIunuHQqQxIoVmKIGrzTNfcK7Xntc
SvoKCjLiqcff4aBWVCvml4ZGRwUIdevxwwgKyzGVLbxIhJ7FXq9m7/Ym88NsjdR5
dLijYMuN89Gwu3Gt7lLnDqgUMmbpAEf6bX0mvHdh3FIZ36tmeTTb4urNs9wmt95h
n47+/CPEbJEcT37HOLb3Och+yiTUkanKLmIGGD2O8JNmx2Pj3Z1n+kqlfYOyyczc
JP1HJLsB4w8/d+tcwijsNJCXxaj5v2J5XJxCQ8/XakxBMpdGzj2gT7lfLU9PkbIc
bNiyLvB58w26eE7fQgSewel9/JVTG+tT1Yy7AHr0ycPie+nhCRo5WS7jjInUBrkW
4EMBEh79pJGzSMNeKKGiZ9m848Vr8DFWuCYtW7Wolh4DHgTCTrVmTxXiKnRl5Bv/
0q+fLcMdosLYDEuJh+XguO85l0fFjTdV0psR+zQlMIjzfsw1rVN6pWVNXzlrxis8
hXcEMjjTtM5p2CjPWFCHt5HN2zwFvuZnTUhoSMLOqeFbGlX7x5dh9dqG7nY+fmXc
AlWoqBXXK1bxAf1syv7DiBAhvqC4MWCdq48vxKCqDe3XOOjuUNGZKA8ozn9l/oDN
cCEmIOUwB1xU3E3W+IzU15meNpAqdNtzqD8u70KATyhQrZDxUYoYHMKlMw1bs4tc
OcChtGNsIaZZ+DkPjKlfzcYB+puYj+AV5vpP/e/inRwxffQM3tgF7s6dgmGDnRvH
InVnm5TYW4X7drtvTA9w4z3qKBOg4CqML0aTNpFDzVOqs+5joQU75GXTC1EEfI6e
+vj6x1wjGgbNMHh1rg6FnUsvaoB7X4j8TiNvTydD6R2FZjbJ6WTxwq7GJjmdguJA
QCpuqhng0E9MDBjZ1eblHMinYAeb6XSRPM39K0K/b22XEakqOZ/VpAQk0NXj6gBC
b22EmnIOVSNzi0WegGnvtxJMxYJr2MAULlAQlz1WDJciMV2aifR5Whhiwm6NISYq
1+4X2boAYIqme1dtdmwJovUG4JLGuh4e/56xtOFBB4F7A/njbiWoAYT3Y+S1BZt7
KPJKC9EBzt7XITatybL94r9i+bEp+bdKgqPp1JBgCaPWv1Dgauj52n7VutfzVeeR
RTuiCz3kDOsCNw/UGHdWDPJji9KQdiEVEL+jWu3qU/HHM3W49X0dlBZMyRo9L2V2
3EGs7HeZSwGVhSVDSj2fvZkVWfIGIH8+x0FRIMpKXP8htZvNkJIfaE9Ciis6FVfD
drRn53x8l48MirQ4IxzybcwQ6BPAr/VF26hTXKxaO36i93s4H5pa2kx5b5K8h5W6
lJ7+JOGh2tKvIUP+3kumoif4t7RyqBv8YeDAyIG9f8YY9rwb/5E/4UpKVeq+MeCG
3QHmpTtkpYkegEon2pyzj4Gtd3Z/pv/sdr6fFd0hMsVnreEWGusDF/nKH1A2h2on
CzqUUX70vwiLkfzVAO663Q7xQvlWgztvhV1OFEMuUy7E/GFQqr22vOLsULc3mlO8
iqwc8CeJkdA6L5BKmUet6oYUL4OAF5ND/WEgCjm7RiOLSYtEKV2OGG84c/MBXkKA
7VXXtfhM+AAHYtwbLQnWle4cwCWnEMNpJiu7xt5yuGU5tlvEdGxMiwiOHjTDl0K2
c08SSIHpSXc7C5Y43ANVj+U6QFvqy946M6drgozphHh95pwifrzIMUw9BYcUTp5f
bvn18q+YYRi+ze0ZHzsOgHWKJI9d4E0KsjOG+/we9/5KrbZKlu80k+twuX5rZTDT
7Zz717hDmdx39uUOhc94pcQD84ctFRztg4cIsudlSFf6Es3r+sMye3zByfSkJWrt
pW4hJvu7ul6SC05L5spMsDpXLopi+TjNZd58fh90GTc9Qo6EYlw0/dcL0etANfJK
gdxSSP1dISI/D5qMY2X2IkXpgWfOV1YjWhWMLf97dLvKMmgKtlJ8PCeeVW14iYyZ
3FdIfL/PpMFDcaKevQ0g6ak6KOB4UubD9qu2G6gV3bnuZWGyiY3VLRdvXirvpkne
kdB0BNZrSL6E0+Q/nSLtRbS7QPE1WRKabNPadLsH57cUGZrTjbk/IuPujyU/RqnI
WKBMWb3T6VPGbJ61Wuor0q4IlYtvboLU7uteg0wgS7v4MWbazSDEffkEkQwbq/xz
8cRH4ff58l4aJS7DfztFgUbAtbFIcmwMH03rvRNeQ3sI12G0oIsGliLXsOMq9mww
H4OrcS44zkAPO1h8Ua7bLbV3RpE3Eg8YP+UfIbOvojyLaUaQH3Q2ZlYLikUgOgCg
cDPonZbkhy745TFnv8wc8ZCkqbBWZ1lN4ZuFpCIjvei7+RNSQjp9T/fh91ojLPq/
`protect END_PROTECTED
