`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PTskvC5v+WAv5ILtM52j6KlAFPZokjuFBKWqiwig4Dz5Gz/zTJgPlkcJWDTZmti4
JmlZMCnLJaYXkuc6yp6aVZL9h+VtcR0Rzj3iFodS9zFGapDnOQH87Lrj9Eub01B9
FaFu69a5PIAZQPy1mKQ6HOEDhGFxskV4gtiH3hD8Nq5aXqSK1zmzS8YB91Z8K19A
zVxNCYW6aT2XgKw93SNTKJB47Uax4BLVgJErMAxc3Z0M9ER+0WTcIswtkTQdYrXZ
B1eBVnfKGg3fHXeeM82MHglNJRjiQ2I8wPTf7NbLbyPoQ9O+hthusfmJ4QwhAd9w
urPmhZdOKUzuLi719tw2mFbAH6A+vqHoCfvDZn4hAZuGYeyei0tIE6+cnAHyytbA
6VPvzIo3f42vneFLVQBUdxIH1wZmjOzTjmxZ5B/vDXIuj7HQjbFG9W8noZLVjFXZ
0ItjLjf55UCcOYQaAVWd/gqCV6WFMIA4NV9dlctwODUhCTXxWbRtnY86XdpcQCIG
aiGQp8y3HfkRhi9EfAJO93coOeGfrN56ztjLZwyvLprkhHRiUtz38nrtze7IIf4v
6WuxhUE6+bO4wsFmYf6jcphhzNpw7TR65Xn5X6PkixOU6OtjD0t/1trQMeFUYB0w
65AblUnUZJ5r5qCIgIZBfV7fC3pfk6yi6fuY99M9i9dYdWTCxPfcPaEKaHu96bY8
sheLuVoP/dZsQWWAuCCTacbwcyYZViXwB8/lg8iUhdKz2r8ynrSsmk5xNOprBXTx
kt7IFrMjIkLVHXjJJsulz3YVw3C7GljCw2Cil2hzOENaMfvG94Q1j1QZFxvEj4g4
2apHzvLz4ZDZcn9nU8XbE6xaNWl4NIj09y4YXL87oSUL6GGpXEqbBBww0PAwzohm
iLf7KgCHC3J2lTeIUsPfz4kUFeCufi3ZkYafu7VKOpg0pot+QxfOaDtXzCHyk13E
OJI0LgkgRbxclz2RcEMdTJ9HEvmORwC0uVhaTCNuJZ9ZSJwcOpLB7PvaQcOeQk4d
`protect END_PROTECTED
