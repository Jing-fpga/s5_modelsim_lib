`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K//0R71M6DL8JKVgYsK7qlrRtfJPy0nBpObOWM3sSCeDSVCTODU8FF5FFD9+YqLy
J2d8gOBuTg4l/f/g3CJgu7gneK6OkTMUOmMATrb2CUh5zgDWEuCC+G68YA//KbjD
/v1PgXcluqYoKg3Cb7EAT+xGx1eZAs12OVpiCyoWAfEm63Wcj6Val4sfYqyyXgeC
`protect END_PROTECTED
