`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3e6OkuiMgFjiCP1v7bHNoYzRQdyNenaT32sABzYN1fx5ZbT6gSjc9l31/i1oo7eh
2Ez8F5D+cYO6rJdVhH1u/2/f27zICRBwMDN2lezejjouD7jueuTo1hADBB6p9/D2
vq0lrknzvIugvphfu6rNe79KS+qjwb11u8C0sYeW+A38bK+SVGe5iAtpK1TzAe9e
MW8y13fSrL2NkzFRBU5rcZBAsuyKSh1byezbAEkcIwlehINsnTGoAL+vUWW+sW/Q
2k070rOjMlpIQin1bdwV6HANcSJlQs9Iu2jTHQIybM8TgEhFBl3+brMMfsCpKzk0
Y1xlhBUEYsnovZW4bUTsV1rFQHPPAIpuqh97gs0wXdIQxB+zMLusGUR/QQ4zAGrm
s9+fRqzC17Aa9U9kN7pp5nG4UnsL1xQDOu7IlEEaUEHuKafHfDIckNWJZjjjPNpj
Yoqgw5Jay82OFhbp9x9H0Y3OkIqJstZw2zzkmkJ+awrZ7ThRlEHUUM9d8v+cPGAM
dP4O3n94UqAa22AmgDWgrqh1+PIYLNoQ0mdO8SVbr+/SqiK+dJBxIb31RiQVuhTZ
IPGUCdR7K4qOcDdmuERGiYlwCGmyEVmToioDPeaKPwN20sJXf2+IXwqBjw26DGoo
e4iXXDTK/TElHWdMIjI9NK7Lsi/xYBKkXzCp5tViXB7Sav9eKQxMCPVazZzIn17D
kpkQofdQEqUnxul+sYImFi1Xw4MNwldNhr5EciUsPEASdV6QhtlERpRXvrraQtqP
UIdc8T1xpwrORTB5w47YesGQGF2MbPph9B7DH7HNreTteSMpG9V0uu+Tq8zjl1Jo
dPe7oUdxQyLH7+Eesfiy5Ft+xkX9Efoc9zcvr6D/iZXYFeMZv/NgnAyhIcLz7LH4
ZptSOFitheqZgfMhFEHnVaaXTQ44Yo1jEuRaUpMxvR3asomiuNAPHYKn5O246VGj
8dJLU5qiqKhu1jdiPe9Jzl6eorQenbeJGa+P18sffrIuwHoF8zM62a7+oQjBe5xH
nuKCbDsErwfDCWm0u8mlBOBJF/VHfJ+QvFJeNHeqWsXg2is47UqusEwq+0hA1FJI
1La1TTVAfWozWVyTLxdFHzunS6UFpo6LVLd00Bc//vg=
`protect END_PROTECTED
