`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yjU9QbbIRhXaPiZTnA2xUA+mVn2+3bU4eYnahzh6skU4/0IuXN7Qmzsl5+HIXrmX
2bVZgiSQPT60UjIfhzSkh8MAvQdlItDCWQ/oQOq8UEpQS39glHL/BnWkU+SGzh3g
wM9YG5EoDATYxAnhYvmilFKMYXXbiRLwD7cMG79eJs3o8cGRSYCB4h2Awjz8RpZu
5WRcF0CQL42KxpymE9yLm7uA6aGFTx8wuccZWIQ3Z8I4xVpSrq6XehIkyA5Tf6sV
q0qNL3HLF2asQ+FDoRc3tXz4tTM34+AhXYO5NGF6GYvMCZ4XmDpS5YRzuQj3CD1J
EkmCiLOyKeyaXN8VXRZSt8OE8UcNJHYvMZgpuPrRMoaqWByo6mnhgH9NKJFqAYpR
8O8CGHDTg1z/6HVyoPaevpdfL/kTKc3Aemd7glmqxIVZbJybW9Y4Ma6t9wM4tqVK
e6bKJRE4I8yFHJm4VAmRdFXNLmbVtDoC3quIZflS0xoXM+i4VI67DV+eudP1JIgy
Y8HIYZHqlkuVyTw78nk+2EJ3zzMnTr5IcMv6HBn/Bdd8Jo3TXksfaS3HIPYXxkXL
4MMUpdTrwMopNI56dLlNQ19DOqQDDzaT3ftRlh87XS6iNUsjxItfOKAfvB+xh5c6
V/9IVkYcu8xJUZ8mMwoO8lfLo0kmoi7QxMKXabnCGBrckPMqPs6eFGQM0fy5xEfL
8eNPgT+1Z/xq1ylBLZ3U8CM5Lz6NvYlYAned7wer1SDMUN4fn21yzXYMooHiV8Da
d2CCIwKRddyte/siZUqm2H8BldcZadq4TUfuwHlZ/kSrbDjZl2nvqbaWDwRgseTw
k8HkRb7RJR8ufJWvN8rqsncxJUabXdwd1yj+dkjJzLPYzpsfL2qKG/TpX81002GI
MClJNTfyMmPKkBUOcMPvFCFujz4NIVzfl1lV1P+08ZNfAzkBITKll8jsJLKCbULU
lS7vIkpPA3Qb/Yvyx2r1g5FiuzxHze+me9aalKwJ0+3pDWpZCtuKqYUkYFCVcTtv
8fLFciGQ/CDJaCNza1d55gIYJ5CUonYOIIUzDa9JqrgKI1lRYJ+wP8ttXLBmJhwz
nCz/voZa8GiCa+dUAOtwEGwbQZbCdyS4tho12nosJdgYNKC5sMY+/G3xtmmtI9rO
ZIpJEcd34o5mbFwfUqnGPLMd78DCOD4NSQCApFh0mVsxNIF7jNPzcVGkAdP6Zpr2
7o/HV4ty2ARtKGxEaYVd2tMaKQsI+NzWc6IyjzP8gwECM9qpfr0ptGnsWgrI/7wa
TqR4i2uP3PqvF4uLE7O6L4d14waLHXns9Yco2SroVyylUTFH9nkNUyJ6jTr9LJRE
JcB2CLBkpRH2xaOJYj26M2V7zhl3KdSy2aNoKOT2osxRj/tCjecyxCz7iYRjuALe
`protect END_PROTECTED
