library verilog;
use verilog.vl_types.all;
entity shmkt_tb_sv_unit is
end shmkt_tb_sv_unit;
