`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Xc2JCJm8g6g0N0cT9pNNX2ZgxW4MxdUDar4cdk5c/sS3uMyIpJ9af8SUz1hIXJf
qdjN/8c50AMGUd4dJk6iXonmTsn4kXSFQugdq08a5YZAJstWC5YwbZxaS7LRnY6z
3iHQwABfqOeQEeUeVeP314iSmdWpT95Sztruy7I8Y5vnpEiYCNVouqhFcKoalswf
zodvlatFZcc+bgNkcJJI9jqLghXUW6tVMzFWkTZVHcKnDvihGJBoa+vPvY1s6dhv
Fux66udyVURPMWiwKKLSpIqZkk0EkHpNSDAoGnNJ3WA+RMO0xNiIN8OejKewf9KU
5yHuAuYJ2BwfdEDdT5QQtiE9NkiX49BMn6ACl1kypErKGh+O04iyWEo+AITY0oyY
9289TtdtraxBmzfXjgkhBuueZFNLKHJydtOFelPtdzuPX8dRfSjUv8xG7isgFTPG
Z2UsPz6acqMUcassSLsP7N56oMP+UaWI0xFN+XFNn0XkWon+kgve6+c0S34Im37S
ZY6v/9gFUyF9zz14lN3lFhT6wkKg+SYBooCQBvtOj6eYJJ4LQ4d9DuPRsL2VwHo0
k6h/ZnwQiR7KVHjzvNGIN5gzGFPLbjKs+PdG30re6ZE=
`protect END_PROTECTED
