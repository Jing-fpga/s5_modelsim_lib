`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D5HpE46DbxZG/Cghx9iUULFeIVn8whA1UIVUfUlIemTNRvnFvROJThyqss12HVMT
IxrFd+E+ZzpK5KkPJyCZqiyZS3snSfysYAJAiL3Sv/i1quLmaIUU996ngSdPjZpE
1f7rTe7rzhbT4Vxh2qa+lv33XC9sAD0/oyqHUl45LbjKrQn8a8Bu5e43cAQcGsmU
Jyw5EEog65Rj4RRmWxkCzbUNTr980i/1FnGU3Wew5huMTHN85iCNJkEM88ippGeb
zZY9upQg7B8PJMMMxJ7kIR8A2VisHPilqyO2a1ju1kDPOxmf0m7xhEU5eQ0U7HkM
V1VanTXUS7hdaXRyjxgIlnAbzhHQKlxEEyMiGfOCdd3xql3fYWOslSbfKuVZ9jaq
Kv595pwAkgoCjNb3mkWJuo0z2VuP5HDFwXZTj8Th8I9/gvzzRoC9hm+IWcwW6MzT
fm6hif5CQZjiFoPm7mN9DmPbRYfNIAGX5HPbFdmZ7yiFIyMWLTRqYjuBWYtEmKcF
dYaCPWlsPc40viNqujr+ky3s8OovxSBoNs/aD0wDjNE1mCZo6OP7HlsmD9t0FbNG
joQoLe1NC08Ffp3DTyPRZfG02qetpNdvjBgREYd4s5ts8wHpfwatAthIFSVsvXlv
nyBteUo2CZA7Sk+M3+N936/y/uKWhf2UhlX7fSVoyFOM6pAmBhup8veVXVGgY4Xp
Ym/pDgi6ysE5XMd8csXXoJkB6DHtnt9Y44pcnsoU7yt/3Kqi0quT6AzUbqqAEmzJ
AjbtbOawaqhPoEZqbigR2rMIrHMf8a9lkyuEqu3d7YQkpHmO9jFFVKc3nTwEdns5
c/rtMnvAjvb/VJ+0LYrrWJYBEsPXR7GVc3IRExV8Z/iaygnELj5YJHPxy4bQ9wvo
kD9oJhY2wa+FNs2CQ8yJbfDQkhf6goHe9fy74tyopUhqRxZhnMVbV6+NAbxeyixT
Br4hsfMnpi4GnK8p4VoOIuTyPWXF8bQ4vpI+PkXvn3OWKo806JATnWTj0awQT9Zr
pCs8prpM9pyScykHbcXPNVPKuWt3rxaW43QhVJquvOD5TBix/4JhwGQr8kpAptY/
nw73U4EX+xbCe8qWCyOQ1uNAZfmy8rjMIlLJT1Vl1Xh+NvNNAF0NggMCIxwycqmp
RitGLP3Ah4epTY1ZhzZmsQOyCnUua0oZg6qPtpOMDbQf5JG4FDmKhbkg+/QJpMuL
Qh58+V4s4w6tTItLK4DrKwz4WY9FmV6L5hxKQVHG07FdKjB+RkPcuZPTXXWRrDOa
UlBQH2OpICPXLjJfqZ6EQjrqHEkIRzU/MSm81sRZVIS5GXZkcZQLqnxpcchoZjv1
QFGCURk9JJtr9Ad6aMUggiesCBkeuxwaNl2pAB3WmWaIesIeosbK0/YSjPva33IN
4g83HtMLeUgozXyDTyZ4aGB6fb6GtENXCyR82BW51eUaBOeH4kqZ9q1Nl46okjdq
4OKsMGIsQ2RI3e6S1q69bqAI37pyfl9k7DwmPVOipMMWUCh8bb7CG+bcrdu/1L8E
pRUzzICuLZt5869H7nJ5mYzBGuhOhCR5ckNwaYpnrswuiFkHrwdyYwOaLhZJL9y+
zXkzDz/Y7wz0WI9mJf7VLfWsx6ELnEN0qm1ei6gwILtwBxITWmD8mIkgyNFIvZ5C
PKRmyfdPO4wgxzMzQaRc5UNNG+z7OMToyVjOs//DkzJv+1f69RKAPRHu+tObsHLH
TD3mf9aguiQuCIacoPjJ8a2Tw77oR7DMUt1RR2yx1RovXtX+1PSvI9J7soAo/C56
a07nXd2En7nOkI5TbVfvUwZapBuEQMVllYeATi6yyb/UkFClyZbR5ZMmlhZS0krU
DefENOBy1GroxTvWs/U4O6Ub5I4eRbCYAy9BAcjbAuoiZktNcssVrMhCe/2Sd+3V
WROT95DBkpbFFErETr3Mq447mSPB56mLXqdxXeg9z1qONhwe9QNV49S5duU4ikpF
bMHpdXK/z64mvehpGESIDTVwqSFaibgI9E1Ls3wcFjqxrQoAe1dLV1ciUznAo+d/
6x5GvMt8n+K1G+0VaHHgQ4vJEML1ApqDMvUqnrQA3HM5CxEgZJuBGylz2aL5L4m8
AdPdYQnwDPYBJB3SNkyHElUJJrYz8PkySh1HS1eYLtaUj4wooXA7cc0AeqcCTcJi
H0xb2cmz80agvTvFxxd4zJQJ432TbN0TXbV4qcivB6s7zUgj96DzdKYtOUuSJjdy
MjR1sWnnMPrFNVpqz24s4eQnL4zUEBaBRcxYsYa9oEGf1R2ImE8b7eEvXRZ3d6+2
T86qIeQGkcMptXWXjRvEdXL9Ogs7bUAD1K770hHsAGbDeNuy1kfAEUDCJ5tmdE9K
95bL2C7Bs2rkDMlt9A/6wp3xqvhWBWQJAzO5tQd7eUGYm/ksya8cngrTb1r/69/V
TvLdr0ZXel6WDAwNwXpSSK16WY6rIBryLi+s5NtmDQ3mZgdRFHysuG0F6l/0KoOu
fqfSwKp8WvmRJ7ZfhxcqkNWbC0GRujCNnyNaK+0wGjs=
`protect END_PROTECTED
