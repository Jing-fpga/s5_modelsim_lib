`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pdJ7LO27C4Oq+diK7hGU4wmm6SWGrSIiJoctQH4R9bK0y8BndlR1FZPIhz4YEZeH
RrXQU2V4UaKWw1uEmP7Wk2WYAwvURsOGtM2WslSEtyNOBttZvZEz9Zv+GM6Zai00
iJO8rMSn2pdhbS44crjgtOchfny3Y240R/+jkZmVOvn+/CKameVqXuxPib3t/iJP
N68tizrFJJEZ5xE2tqoRjghGsulqTpoa/buBUa7X7KOM0xfYGf4+jsxfAcYyFycg
lptHkGsGU/stj54X6SvCzHjg8mV052AoP6dTronAbzbVaePBUBdNUoK9Kh7onuRw
b9DeWaI9iPRKrdoU12TaqJ1Ku+ev1UI1FzjwqFACIbmKQpq7e0qeqYJyf2CQ5Tg5
/Nh8XWQLWZpWtxAvO9KZeGPowD3PP9U5wqhQdWmJ+qmETk8F6yHZYKsu1kwFtcUo
k3yfpySm20W+wFnz5IC7+2pSwX6nYpuptNOD7ywg+8qFezTNsYb0505oeStcaPW+
Hb69xjzlDt4fAEfVKvq406EUEqdhXVr/Bu8q/q6bnW7A4/fbTeH8x7ZASHWzW8fj
9JZ5DkMnpell/2XEvmAl9ZeawfJXsZ9oAxt2XWwH9cX2LkpQj1t1orWmpjN3rGGd
emQtdfPZffVwejB3MX6iGe84hH1YzFQ6Hrs96DF7eyOYTpLBr1X225FEx3CRE5vD
4tUZ1PAoPMg08AhfMZPRB21p62BUVH8+wYogVoLz6fm6xTl8V5yzAo/tG7Uxa2R8
Uq/5J95iNdLVfn8fx+wLIi1zgSw0kEchn0UnLTMORhqGf5Y+d0pTz0NRUwP3zoU2
sj3sYWyDFmhXRtj+SDYF9IiXHx3qGJkskgX0k0vab1waGG7yQ42mnsckSR3WOCi2
I4g+6SsXm9Yzm5UGnloeKUk0A+RqUCi2RjtHflH+KFuHSInG8GVSvb/ZHEy6ZsuO
hkjiKTqiHwjuvCTibLEfUCl04tpXERjbIC58L0SolPXCJvqXjdrhvI/tQFSq0L56
PImbm4Ig5mRb5pDmYN1Vxfbo8rx781TuDPyEdIyKlyMPRMZYs+ODrmpS2JHWCT+8
PScnJy4jsMfWC+5h8lrAiRbsqe6GfiMUCdU5VOCl5oIFJRxdDgkRy6sdlmhG5LIJ
AlqF5NusxwgOoROaeMktH6Vf61ohSsni5+FVfIcMQz32b9KuybVgiEL0Hfb2EA9G
gAeYCq9MzKQMPICWSrOSgv12AwZWZ80UUjoejU8H4XBIAuqd7KCiL0EXJmN8djPg
xLhPSFHf9e9HminsNd3pGRc2j3AlTJC0OeHEho+hB49yADRMUwIpWBKSLT8N5l4R
P049buWDBEE05zVzh6ZQcZcoj2wxKvLtoIZ9pgfULhGRKlPJmOv2SCthlXVbWazB
tA0tdmyicLMXsn1LfQ0P8TRRfOoeyRQpWqfoMHu+aKZdW3kw+93gYt115fSf+YU9
4Owf2nauyQoqFTnJHKxhKco8rm5b76JGojgU7vJtxyq/su5ba7KfF1aXGIqetOa5
CyTP6Mz40xY+JiVBL7L4uCeZK1lsxcP6xp9Js+GlR7IE8EEN5t2M6D5lZbUNcw3H
Wje+6xwM0jvxtS0noYBa1LtF4puLHGa8xWG9sCKF/R67fF8ct8pxgckK7XSGwUJQ
x5hOWT9p+Zrwcm2cbY9y3X2ia0XXbhq8WWmvwc+5+HachZkGr6Dj/utlWupYwXY+
518rNT31FKeUkjDYl4xohwx/fSaKSPPDoweIAWn6sKBSnkvSsIGaj+EQa80P41VH
tt932JX+W1W3l8Sh/bZMjPtA5izj9Fj3v79GR2SybE/DISdUSGdYYMy01XtKrhH2
kipcJiZjHKqEqRKNhTNYht+T7xRmfb8EZFusAzGLR7DyniOTrAoMBQzlx9ycw0xC
t8lUO3fp6dkxgJNg3VT+zSiDB7MaAj/oy/ILcg16vO1uN37N0emznArm0uCAP24g
gdCUQ0qidJ3oSAXdH31rdlgIBT1/B3bhCtSHfubfUWvOV8MjUvDFpLRqNsuZUIo3
bNhMsRv1UQM3PZvDXX/Px949t7uBU0CFAJKSfAcI/e3SR0PFrEpl04RABJk4Lw1B
0ndu8ug67k8Koxc7MPMazGpUpg48F69OkB6J7EG6evP4/XnohGlegwv9fAvKbl60
c06gWZLZF0VGqNp0ipnfXOmLbyGNzQgiS7Nt9hnJq2JMDNTr1lZh6ZCpvUtgNAdL
WOyRu6QxdTZciZ7kXw8Ha2yWbkTq2sH17fhrQZLqsNUtAlLOl53RSSw0Cdif+vt5
cKj1Ga186AUPlWWO2O9E32TUKrt71wHoHB5ZV7d7Bmv7slnaH3zvoC8m5UsuKLNW
ogwEfygT86iQmS61866vmq6V87dGtU8jUbJotiQEv18qA6N6PxrI/EktQrhrXFcV
CSSp69Wt8eEiTiKykLvztd0eb3SXcR+wAeg5nCmlm36FsfJy5hPYdZIsFeDTZdC8
MkOOixjjt5cPM8aO2LQi59QAlPIJEENGNW2G8G+zcRRQuKjhaEomT+8DgEflIk6d
tuyBO8E+P1fW1rWtIDsVW/WuB3542LNokZQXsTNQK+c3958+Nz0C9N8tg+tmawYg
0MCcIdN7xCSvhenXObqVz8ON9foZLX8aAB0d5GJZ5x8FurmqX9JpbElkkMmApgPN
75uUDFeGoldMic2o5Y3HvNTwBMzs7ZKBL3TNoBl6pT0Tu7glJQK5HLr6UrwkrGaN
XEhgoN5wV6n+mteBp1sRfwlRNBTbpG/ULvl2EWQR8EIthNyAkXyd5ejpE9BY0Dz4
FSX+OFzJ+KT2M6GnX1OnzL4K23H26YPyyt+O/X8gC6/ltY7cwfb5cYbxkQFy3vUk
L20UrNoVmU1ZSu84vWrWhMmQ8VSx0jlNL/pwvv9f2GkO22x3PRwEoBU9baJgJ4k/
6E2ypX8G7Eep1rHdwZ/YGjdSSndkWUeA8ykG9Q+Mxq2OWPXzVjDAX/Jq61SlK4U2
RA2rHB6GRVxNNSFuKpplwpMNN5ljkEFb1/oY8KmG0yn9b2OG18dnm74rKct7zFIj
as/NY+5LuOTOio7JAU7KRmkuspkjhoubDlVFSMrSd5O2jsT+ZBo5j5boqV3kfqGb
bJA1WB698Nw+1NGYgVyyuHTk0jsxndjbf/Gx3nFRfIvvvQZPNtxjoQmJKRfo3B/I
xIaT9vf2xSRav9ldFOB3UoYttBWMT1Wy3ZICx8HLLlomkv3SDwTgjzkDPd2a+tPz
H+iul6Y9biN82K9gjb43mr1Rd2P9D2sHNOj56eAkNasi1+okeSi9O6HR2din5ky4
Vjv0CD6PjTlNl9RvVvPNDh3QY+xfMpHb02DCOT/kPZMg7oz/sfLik1c507nSZ7Yt
P7rib9vvr3bUwNPBNM5j7SQe9YsRzu1CBLWft2LsPL/bNb0A5zO+3hOReuBwB1SS
VDx4o8sNQs+y1riW9zXNt0Y+AimBz+XJ0B0ryDxRd3OhLwmX06j1J44NfaIpqcbE
nSxFRiGYUWY11jTUm5/I4F8EZiKuuIZ/JdBqQ1FpWdiQVo13GcQAAjjYZrbRLMCT
9ibs/5l/8zk9g3WsdlA0DidWZHyJyar/7LVK1GCT6r5DavCjuanNPCN9751hr4wG
86F9Zq/zbedCV+eOKZnty+X2EWvQPxJKFmC6HqcgGadqRn3cmzQcym6GFTKwuEDd
G+yPD5yv0WR6sfFIn5ti6/nfT3+ltH6PQxc/cDP/NUU+bsMAVIkD4puJkq+2RKGE
XcCO2JDBVc7EwkET6pXfVW4Cuk1lQL4vLyY9VbhZBDelOYmW5Wn+o51IrqUfob02
fcHL4IxX7fpPp+xb9kykE/0XOQ1GDiHr6NytmMYLuMeB+2v+LQMvqPtVlIHa3wzI
zlY+fUxmLt8Ngb83yUVithxNH/JpkC1ZqutAkqfPb4Q8l4TkFUjVOYWmZwU9JFEf
8YjW/cVE6228Ouyqc0aJeScZDnWq/i3WzWhUnquuWyzJC35El1hHI/MrH3pucOlh
2iYU3fqEzQW1rylDTiLa+JgZ8nTqP0RtpQlOlJDseu2OUo5mExj3UjIPDNynZP7m
MyJrKoGJCF9k5Vkvok2044IwYrxh5Y7NMSc0tIqnp1ji0fN/WflzmyAWNTpBROBR
H7nad5HGj4qjxHgUXWF+VbhdUIRLgjS9YVZ7l4aldnzXvo8BdI0rbJSRh2BlOyeF
jBe8dTrRFyE3A13Tasx61CZDSas1l2B8Mc6ujYbGElFFldiADYss6cluJ+MiMo80
QW82QIYUe/JeXVRBRkX2Nnb+DFAQSMrRNgAuJ7R5KQkiyNLIAwqY22JM+gey27Fi
/UwnVvYRMJ2Ry2I7YdtINIdDrnEXmx42mIo5Co5Bm+FRIHLYmkCbM/ZdyDrVquAO
LA/b+mhxFd3Dyux2EXGmvStzuIbpLzddEq9aR9pnQrSfc1KVoiIRRxRDrcV1BEg0
9Eiap6tq0NOwu7Jfd46aE3EnYS2kRqzgyCOLPPZh0d9Axhp2DYqDHUcytBF1bvXi
LBEhDITszNcH3UL5xLXDQgS6JdfJedImU2966+TLUbKiRfkeB0zMIIj/Eh92un6d
vJBpf3wnh3zX8NiMZ+VgCHsDytAtfJYNp8xpPCD3Q0V6WRWJgX5/C0RhJ18SUWjE
cOudmNgWsbXvTCueWiMNGY+u30rK6+Yi3rTxZ8AiBVZt9BFrOUV4vmkfX4rLxzyX
XKmcBiinESUeQnZZ8m7alZinQbD1cfUWLuBeOpmdjVoTDZNJN3QtGwNBvV+K0MCH
2Xq6ao2vcRKS4J9ydeWCJWsKYBX0Oka8KjBPtHlou5l4Onx4QWSN5cvnrU4C+5lg
aa9yKgp8Kbxsldmx7Rjx2wDz+apAI97gY1Yt8SSBD/caB3SrFVpkH/RFfLYDU7b1
wiobsrvDn3XMI6DfW9Df6S2wwG7XZErQdP/Ae0idOa5fhxb5glc3SDZvy8PGj1xw
bckciBCnppGOMXz726pURhSyyZiH1XNBi8woPLUMNfnIcqJBktSECgkL0qWHcXzD
Gop9PpSRjHeaEMxjCSE7jvXaUjSUcNm3US4O238l2m8tHcp9LNDacqSoMc2zqcSX
rcgGSCU4Ch0VeK3Xvm+052GwWGklkHqzb+LK3Bo6Iz1ENj/KBAR+ZC1CIiGpDin2
1N2vXzi3vig+y2wnBd32HQFthlMK7C0cfXVr1Uv98Z5JhcIz5Aw5a3qn1CVem+Pg
d0sTN+700mVxvru5B/WJEwzVJvBp5LQcgtS4z/EoExuhaVuwUf0qJPg9F+bCG+fZ
vyFk+ILALp0vMpvrURoEwwqXxIn/dZ0k1tNs0VXvpxafF+pVplf7/dbZ51Z1XXxu
HnXfXqohtZxkknx/ec8l6qCgrG/7WiFIr7nm5yHT95pr8kZGBKtbiXpBHCSLMS9T
p3UsqHnWD4sxY1V5qrt/pWNOnEYYIk7+V2j+Kdk3eMCfEZc9GvXcycI5oEXMRzhp
9rTnG8R2KckPeKxa2mCkCquzbAaqw1Z958mRhK0+32sVC7F5uoymcxhbG09z+g1L
MFCvu2VCT3Mn3/EgxraecpJUXZQApTx7c1x3UBLeiPZzb4ZfbOoLq2t5tMe4EWXE
AUFCsHQI2NSF7tVTVF9pYX8b1usqhJJ58sDYPF2IofnsTo8OgxEhKaMLJ3eqcfju
kRVS+FV3iJulqeX70Ge1tiCbfufyQ9N+GbUtVX8G9oZcymai+jwUor/sLfObhJ51
tUdBdiAYcfO1o3yM2toUI3xFle1JOyvArOkF704E8yXfAu9r8bnfxIi52f+pMDqA
Ntc/FKn8PLlPyhtq1HI6Qrk+RJXQDX1RkgcAcDmUwUE10ULO6JWCoF9kSkB6mnFx
UPUTUSnKxAtnzkpB/Uc1IVZMCjZgNGr7hp7eJ1Kui6GdDNHBLazX34vw0qs1iXhT
U+zDpJfxRs6kYyDOB5ALQvlinzaRbT00sX5YTLT+eZ2B0ZACgUom7yrksBN9jhU3
JQcTZVqXTyHuAIuMaIEuA69ns9UbxJL+D0fFhJ9J+n42Bz+MVmghM1YZB5gVIpcr
axHml8GGIgbyFcPUN78P1IbLqCMQ8lry1uWZMHtwUA8w498lxxegu8BbWQfzV3hL
TgffQLuq9JFlnJk8nQfjaDfKb9NSw5p5anpgqT/7Gm94jn2yiY8dGa4L0KeKkQ2V
I5XOMJqEDplBCMoqMWfEUGBKzYxnbnwHWewyC9aIAi2WLPFgejZa0/hSkTe4KwkH
z/TMv28UO0FLe7WoyCRygcmgx7da+a/U5fC9FZGBLo9of1JD+ifqasCDeoxkC8ve
AzLFLqne/CX8VHBrsK3ic2a0gt0s8gVuPGv0uzg6QvDPotkZ5l7li0iu8prgRfr2
3HYqaqQYGnWOLyrYsY2YXZduk0QwCQ+lw/lDJ5d0UB1xdQFCuUXOTqNvqyRmHae6
zzF+XI3he83YHk22VXdia/7fiFwA4Mo2EPipzmXcDouhEME5Pv/W++MvzP14gSAn
rXMeWR3CSTFnpeO1TnoSMb+EQkKe6/fwY5OH1I6FiLzWxAmomZM2thxi/umS/Stx
/+d/mU7YwA5L2wrEgyNv9j1iyL1TkkLRWhfNGsZhFBQR6obEc0CODb1H5xL5K2CP
6UQa8QO9mOJ8mX/22uDC24CcNlModBsxSZ2dttSQvbSuUVar4dQ8pBElsOmrMnFt
YoDb+WYdMdQl9zyD+heiKpEePeCxAB7lz6r/4Y6RvlmeZE1vtIM3MfzZhkOEN3oC
NPAeYgec7mw6qOZQ09yuq1Qh4rNcTdvKjL9wpEXyOgl6DO74OLPjyVXPP17uuFEn
QZB6syqeupI1q33D9zBYo0owJ0+aI+5F36+NGpbMCpMfSvy3s9vU4LnujzL+JTUv
x049xaOEEAZihp6Y7aLJLhALwRvwCvVnd3HGcUIDnEgJ0hdv+T1EG/nB9k0L5aQ2
G6RS2NufWOWs50iyr+webE4huEYZb6k7YgbbWd2zX2dk4R+SaCNMC8Dz1Bw8K8C4
NG4RftvaVor2SDPyl+P6Z3lXz2N2GHAECXffrptemVcsonRM99dyrXaO7Yumc1je
3Dj2jyxEhvjcE5VxMVWS7GSHuVlK2j4Xg8KXvSXdvmIhxuawjTX8f6h+DL3dL9ce
joHK76eLGxtaZgv1XO7iU1bKWCWhQ/hkRxmu8TKV+VacHIFOIVXAjnNH3eHSkcU3
r2psfKh0Zr7VEwDsea6GS/7ZoUmrv1puQ/X0nl3V1Vnny0plVxqv3vlz8gOpL4HM
UWYjYT22nFoeUwsh30xsF20p/l0sDV0yFPgUZTu3MS7RpRIpbeZ9o+F5YcVex4wC
rRTfEzSVEmlJyOWpRbvLsUjXSbhBl2mFZ4umF4Sl0as+E3dmSNHuy0GwRdhwlV1G
saSTY6OJPE8S4soc04SVAk6Zp3DrTN3LHn6QzQByV99FH89IaD1okkUoY+ikC4EG
EGVeckorgef/pu81d2IcUytsUy9MuQMbpEiNyKatlccYKQXz0jRQMvqrNbfS4nFc
PaKDzcvcAQH1wjvRjdOhAcCtZd7pvKodjWCpGvsWbh0xg9OV2l6+W2LXPxR+39PM
B02M9TG3m0DtQHfx8UJ3+UZU/FbmkZhU5E60wJyVcf0xwxw/3/LLkrg70yCx0ACP
ChtPlmDOZlMreoIVGQ8m+Rgmhu9wKw03Gv9bKCqTltoTP4AN85M1klzFhBehFhjZ
qIA5sxpTe9g1FSZyAIWGQEbWKf6rHffOe/W1h5hs0lekU+Kxn1/BsQ+oK90f2q3i
efb5z6xNb6/3L6lgtmqQyNlUzQ97bkHWX+6HgktbCMazDngGejYIveWOH36TamnD
pQ0QW0+TWNTaxcHlKA0UgGIeeC+GLe2M4J87Ri2GN+4fGESwxF+rYpFHPR3vHsJ2
tpcCVbbrO4ep+CptiJE7H0azZhN/Yuje9j+BuhH+1ZFgNXz1I2f4dxp1u0kv0XFN
bxypvii+VBQr1VETl5ZsoLoASdQdXSFHpc/Dvj4JB8pl0ZdFz1iV32C/hwTr43VK
erb11Wrm3+Xr1eEgmQupTgd7MnLRE5wQ/EPFF/j5eUZmrJna4tesneb9YPJmz6LP
UPn4yg+a/lRiPFzFwRDBBLFyIMtE8PRnRc1oco2mhy19L9sjCX++BxeeSL6cG1tH
MR8+CKEParTq96akMY/gCGvxbJhBhg90BcfEyIwMxRP/Dr8o7M/rCL8TfW9p/1U8
0Lf9BuzEv6H/NTc2VCU2NuoDPfUCOWmTYhMXCHCB6VglsGqfO2V/gtKggno8/mbm
J0JgN0Y91O9UvhnqlSAvsXtfhKCw02M6wX9so1Y3djHyDzdHM2bsgn7KgFFy6m0a
/8w3urbw/V2NXlsx5OCf/Wyrk0C3sCpvEyZZndJgrAp6LQv1fa1pLWiqdOJ9lm/k
VnLZ2M7Vp7hr1KNCewhgdKpTb12Pue9V1jeYyLY8NSLKy4VDkpjiKKkeh9/mmtQt
3gl6n8H9X3Y0Djn9Uv7KR57i938ZcixQlDBG8j6XI1CKPsUeTjbrW1ZhLuJwygFG
rnDzgc9IcsSHTD2FehDwezmBuTznVdj9Q2KLjPFI3zqXT56X9jjF0gY9QC3/gS9K
sgasO2C0oT1lu0WsBI4Lr2DUji+8Tatw4N5synJ7vOw2DnRMMmwwE0NbejX+qRVd
YB0toQ2wyIUgtlitx/nWpvWakYkuVNBMnkmqdtd3Vpfs0lLhlXJF96ZLhW7X+CO0
7TXiuPJ43xoIMlGEn3aWVg==
`protect END_PROTECTED
