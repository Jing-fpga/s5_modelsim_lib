`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rl17ldPgTENLhvWXlfgHzcui6K4cU66OvVxvnSHuhWs3Pd8zUDIxl3WXPP0WMNRw
6YhNrt8QLHdb9DUHptkEuN9Bp/ObRXqIIn+2U5pn4XQTV9qNHJrF28FxNmLl4O59
nxRQpb4RU/x/f4k+T7247SJ0U3maUmIofzGGgTBfXWvHEArtKWXjJ7PM3zGcxjHT
gsqcwI3MWb8BeVLrVdq0+W481mAgW2kNSqXEp+m5Vk06awtDddlRlNjPDJyMyZXQ
ZtXM94n0FHIHd36W0eprjj6aMZGS52TUAApmPA504IhLCfq0lvJHo0WeJBaO+JVE
6KlVh6EY+pTOXZdzK4dD8efMRwqg9B9vj6Rzkl8oYi8d+uTWiGzvKqgW/YId/whf
LURxexfeNze2uq69FWHwl3Y2KLr5xUd51tALLiAalBh/gzzGpD8cdh5sPyBfha4V
5t7qcjg0jNm3NnoCybj9RrsKJcyioefhf0DHy4xg5b869STfeNQftn6G9+RRWAW/
VtBPdpQc9HCAG2ngkoTz90kIcwceBxL+AVBesfk8a5bURScW52wGxE2nzVvkwIgf
Moxn82kuKBsYYun4NfPyk+O9PpVGhBzp3/mdl8rz9KeZkcvjn+YV5CyNV9tQYjXt
Zbp4flbU2p1ELsCTN8EUaHnWbyueV6HqdruwU5Q5OdZrbJGc9kO4K7SIdtTBIaVW
zK2EdDgg2rXrTFIbVriAxH3TDWgwsFV9+sJlMZ73eOU3yv9DiPQKCfzXuA2SOLwZ
D5kt6kLtxajjPCMWDLLjZpN94feWojA0TUL7qUIrmhrh1K2UdL2LeYwiS/2KSPk8
8JV2sM0oJ7zi79sz9t8ewx5DhPo/LFztAtlaY4SC8na6P6j0llEYHlO26VcOk90o
k+z3K5uTu8HbGK4Eb3b9bLix1ayaSBjLqB6dlY2ba5EVgDxyUaXYwq3G3pXeoLgk
T2utir7G65DBn/Md8BKAW2dCJGwCro6MQlULxT9G+62K2YUqfCMIzb01Gt03VeFz
e7PsesJsjpoJg8C7n3ZFD34Zm1m5AdX1cqsj36YfiGqvu73MQ1FlKxRuFyH0+DtS
PDq3b5zK0JWpvk7uzggVcHiaE7IXA7NASUC8JL7L6WWhiX2+4LITsVQNX139Z62G
MpE2gQQXp6EZtpCcUiLyz5dcoeMzNuA7Dw12rSOOWkotWFf/qrmqhWa8m16D49LG
40REzEilFmJ/ESoJJbG7iu2roeucKFGm1j4Fow37QdCksq3vZS1tf9qO8Bf3Lo5S
aoJhTlBD0xGKEsH9WkzCUQBcuC0pdtOr5als0Zs/5g94oscscGNY/+c+aCZq/tDH
oa5Sw3udtFDEuWTu/v4Y9qwb1oh3iN3rzJgZZ4xk65lkeVYfgR1Xc7GLRbve48OG
Fyw2H/MYlgXKdjApQZTvoS+0ve9QI6XHkVsBZmeIr+tiqdrQmDicTsPbTce5YJd2
K1TdkMAQP3UTL06p9GPsrjuu8+tH67/+PahBvn2AfaR7V2PlXkgw+nkYSmGYQRto
QuMSR/efIjYkchx8Y85pxkLVhyAXViCbbE09rDIPWJgM6ctmYHohBaz6v5Hh4Qga
ENpy/A2pRCKsMQ2N2Qmvmw==
`protect END_PROTECTED
