`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YokaReIWHxGXaxulKafy6aQCvyXRWZb0G0DgqO7QoQVWlHNQ4n+x9ucx+Puf7KqK
GPh7ZpPkzO5g6SIhPwGVxxrMufb6TN1n+Few75FXepMZ3U+bOhvNr+IxWGphDLJ4
rjXmgWLHALee+9icuI7xxYUQDtOlKzmXglEr98Af1aSaowd+7uFM/pKE5XhNRg0D
7dy+AZEm4Rjo42xU6xKImntW/KoGwdxYlBPcYFhpR33lHwQ/AAzyIWi4N1COhjmy
NEPvHDy+fd6H5VaysHI/BWHan05T2nUmYwjbku+vY3nBG+jNeZTHKzCAckk/Ard+
uKP4rs7CxwGnQaB428aGcmh4/3Lv6Q3ZV8Op097yJ6IO286Hbgoy677gJJzqzLPf
jexHDNtLPs7BoeKEkaRIln3ILGwLnXc8FEVxiMpo9SM7THEK3wPLfCgc5yxjYcEC
NQGEEccthmDHGnBK3roEUF+nMUL+Vme+Lxtkyddk74nIRQbPpqiRfI64w8b9F2i9
CBd21V7JKm1lcc4eNWfbdnOeunqvvJPkITH/FRkPMljBfTUEdKZf6pAToDaonLSR
RuV8LJ4n50c9colV2Kvu5uq6tm80WYC+fp3T8DcoUIn340W1HLubCJgHb0PCt9YS
6RhoBFdHOglmVc9rzxub+xbbBpqKljDQv4Xf7tLtyEYiTv2g+FfCa7XmCwck/pcP
0TzFztws6Hosb2xCtlx0pcuktG9Hg9pKc7SqPPlAzXLu4m+Pd5Lhk4W/JKvs+fR8
K8t7F5ooI30oRKECnAYwh6rzfvix0R7vXLAg8EG5KWSnN0pOuKSNEIB9qNvDezGq
0kmkcrXzqGjTrq6ySotXBWqhTYxAxUtTE6IcBfXTomwwUPUyrNzBcbhPiHdHtkmW
e9jnFoLs/aE29vdLHstXeuB8ulmEf98mqlw1XDlXpw/TnSR2iq5xIlfZXXMSKbro
9a6TPE7uDHNLDI3kOfNdJu1Z/Pde4UU4mERqxLC1tpuNCsz9okyU12qohYth8+M/
x0h+POWNmNwWysSrltYvWGXa8jUWcxu2x11lLrvUxSw7ZrAxH+5Iz1LsHd/8i2RO
LyQ/j3NK2VIHvvT92StYMl6D9+tMXmOAvC8CW3nRwRL+I0imw3tpmu3AFKxorGSh
8BBMlLoSK94LSX1lGX1/Mp1+kXFg/6lBjHtG0+AghYxuibpGtv/a1dIyEZUc21kd
MVOM4ld7sgSAA2Fpfj/vQs/3htwbM7xPygvrCZyB6tLBCaecHSM5GFi32urbInYO
E/LmnWmaQiaQO6rvgHXeiyVJZmnG4KqFYDf5VGlVZd1u0vPNxrikaj/TbnQeXsIx
5r/V9fszHjyxCxWFVzN2v/DxvjShYyf+5xlHrtEYfq31Ixks+k36iiC9fMcJz0q0
gPj8jIyK78+IFR7WYyZy9MTmdmsKnKwHqd2CiI4U4iWozMLONdyjV9tR9bLI43vZ
aBANs721ap9wECwMNERevpeeWYKVkyqXZdM9MiC2t7ylJTI9l0dKj0mMLUqCuAf0
vpH8Tx++rRvo/mFuBc9I4pGWTxPhs1l61pe9rtuTD9IVIf7p+CmveZUSeEKgRvKm
AJHNICVD1T3VeKrgsjri1Kwn4ZfWwvakciS/SNyF/zPiE7ApaQPUTcgwaQzBdIG3
uv42cnY4QwIHzh+PGQPZqJCZytrx1UzpOXGjlfK7i731Kw4+iErQf2Xr7uisxFUu
r7to4bD1T1juJRWz0oFaaAYhM4cfZTtVVZgfV4qDgysfT2ckz8NV3+hIOnBzz3f8
5PQY0R9Cv8UNWcoKRs6wInzmOl02nIvJk5gxV9b2qM0VqQBjoJGN4SEGLuWMdWF2
P1ufSeLRXMCQVATGWGqrf7XtSCb69DQ4QFIM1ZNIn6scGikoEJxkKiY4wq/kEE+B
VzGVaVlvVDnLNeDXdU4sieS0pV/2b9kSQGl3MOparBDJT6Ptwwy3FtuUVihAPcHo
5LpZzpay4fjo2ExubsbMuBaUDzeoQ4oTKvEg+vHGwRaUrCFFzC0VjruGmFT+h3D/
Sn5ELu0eaG0yuZmXwngekP4Joc2KaSjaVmSzMXaNKOlmuicNXSz2wsM3N24qbl0z
iQU9jPNrwpzaN9R7ZU6pKrPns3kXP7m3vSWFoHQYgqxh3a4iSQH2gmrU4YJgLXJY
rkbsPQEkdiJX+g2H0EULxSizyzWjiYCotGoOfonBM2+XxurepRtPQpsJqKbvFXdt
n5MouDkyIDR0pCH+WkwdapQs8iGFcygXyGdNCII2p4a3O+jP/Jw/5NOT4NbXejY+
34dewm2m5ghth1SJj3oHbZTzGcLApET8OICQmHMv3Cm9HFuTyCxA7bJwy7oovNl4
h8AStqZZ+P52ekoYpskkf2hvUST4DAW8VIbEh8ioJypsu9oxhWwiP0nXWHU3zZGK
O/V2krAzMNDIpYuIkszMCwSvjsbyt45PbRzpikLRHD06PahUVnombs4pRbaTEvNY
G8vQQsrvm8LbcgnQjdrjiHpFZntvu8twons14a4793pHUhFXHY1kdAAWWnNezMMW
1s7fbKnWQzXjQqiZKghZPOW24O/4sxaXogX+m6jbTocp9NObS79S7iT9oW/ZP01H
4v4Wb/NnNDkk/6TuNbDD11L9BSghF3wlCDiEA158gpTQG5taodrD8mInaPFc7dX6
vZdbX8V8HNck0Nxqh0dtyr1gxIG0rb4X7BzzsB79LQFrg+fSEstcNo7VqrvkgMmY
8kYEx0RAe7gjMlDXM+PrFTNFed9+oxQ5Zl7WYNzsRc6pM8KWTdlKyD7uqoWZmYIi
HXp4+lpWesippMymSj2oRe7M8XNZ6ANXTdi+JC/zO+uVI4A4GXzPIdf25uoC2+Fy
0voS+D4Y7UZNX4EQZPIyzAKfLQ68MKcDx4KpLqRbq5eG4B4YsrWH1Pf3GvwgskHC
7hXpTvjlttSdE3HEE85MawkLmVJf4FfYLCRUgZHIvoa2Rf3INmIZBZrzRITrNWxw
+471L6lzOer3jLQyhKZygnQk/SRhAzgatRTbgJoBh7vv3m8tD0XH2vyOBg6xF2Qd
HYtchuN0EoY/bEDBlDwOZ6GIyqDIF+11un1WD+mW9fvKMmyqpmQDkq3nxRpV/QTA
ZztQae9wAbiJHXg+HR8UixPvLvn3l7OcKW/YizfbGu3iPY5hNeU9dWZcES5jgKE7
HsVMV1B4QQgPfxyOTfMScpZhJhc724pZbHNFfelAaB7zJzh4WAvJPPaM9rEsARgA
cIdfns33zoZmLvF2TRoqOI9mKQvqrX/wfCcrEFgxvT1BVgRGF8PDh6r47b/3CFPK
iAwxuAbgq++538XhkNZJRYQxmrA4mpNAG+uiNVK0eVVJFLdGcHpJCZZ2DqWNAu0+
qjkXn/+w7Eb2EnPrYtezOBKUFJcHQz2CNtNnZlP2fQR5ogGGlpiy4LAhC1uuJUH+
4dW+Hlwry9yU/ZrGyola5qjLr/v5JiBCBdHNelM+p6fhrBvyrnqUdhMtVu0d7ZB7
Lf9Cp2hbVkPJDZ6lRZXDnnV5ZVOPuLH5l4nuYk2x0NkuvlTqHCT2j5umavDO0k+Y
CjCUeAIZ1mD5L5oqfQABbX7mpvOQ8sCB34cf9BzDhTRAYjF9p9HdsQzEjwjhKpN4
7Bg2FUQs2OSiMiB9K/CvUHBCaAySijzoGUyPferGgJIGG77l+sDM7CDA1EssxtB2
39s6WZGF1ozyCCvmf8V1oMhJEhLsoJPBGgc6wcctUv9YSL/CnekPf2FvTLUP/EtE
2mN1WVuB/C0mTdIB5JkbCeKRUSfEvxBo2kgAkn+k6xDW2B9FT8lxLZbvlEUI+LLJ
qNI6aP7uzFH4pPV6GyxhYRUMvnDhaGrhH8O6HToZ0XqXqP9iUGVwZnqPt3uT6nWM
4PevKlfAD3oIWb0doOr9+aehZM2eecxqwrw5HJrFMhaHELV+ShD+ove/+52rW+MV
3WQlWWhtV7nirKuGkESFpNql5E8PdM7g0jR3KeyFZqLo3W8L5UXRRH2fsJdybVPU
MiXtfN8X3w2deX9t6ch2ftnj2mM6rpTMAugvp/BqGVzz4wv4+xOaGPcrr1nJ+JVl
mOxmG3mA7qG20U7ilahRlWit7VNyB5ZlSN+UgevDKW9STJFHRVfmoQlO2BMsBW7a
dc3jxvawE29NFm8jF2VWAaD76pbgNXCvw8JOsjdO2Ldf1sfhwIOSVT+siaKug2ZC
Tx3qXCwzsFdaUO6QMJZX9mSeh0YGQbHdpxeqKk9PdMWH0k0LsorCkg37kJaEau4K
5Tj2eNU/ouTLgFjNSRZHm1mvFXvSYiCiLGs8SBjRm/zwl/sQdThQOUeAYKoRUz6x
nXR97qGNhRzQ+bVs/vE7kmytqy8XESprjEhDFgVYXUKX1lF6heJSmNZwnESQx7YB
k/oo+mGzauBx+3HKzXaYBcS+3q1VPe+FGflpDc5z1blemN6BC3SnIvWWzTvB7H8H
UOUpJ/z4EejZz8w67KfbhwYGcK98bexxyyqkZsOwoEQDd6nRcwBhRqNskN8lqwyy
LFzxqMnw0TjfflmlsqhpCiRFCeiGt68LNye4GIm3smmKQLpcRU0U2ZL0xHvTMUB/
aSjDVS9fUiRkUt5Zfvc4US+GpY4QUBLSg5nPhnzfj/n5klgbaOnEq4iAW5QeYwoP
9ndED3pYVHzyF3P2Lqx+VCCm+Txm6BguuBoEEhSoUaHAVDDeyog4KBUlonslK5kO
tFlQRw4AhihMZJECYDjtZOxDfFTcS0nyXc6ywcePgvSS+pwE0fILHHUrtySfdyYj
S8ZiiMwfxWvICiu9VqFkxu9NESQ81HBhR7LkWbl8NiFgp6wglGPS0osHbqwza4lH
vC2MIOx90/b7ODJDYJMqDpIEDE4Hn8uHWXKp71jeW+vEnWO6aMVxMm6D2s9WqNJJ
SDvrvvzOIRlwpULeJ/2L0bR3vTTNzSV+uXJ08vDlOzSs6BrtVMO3L2UNv9AbtmDT
gmhTbafs47AysF4mP/U5FgM4gUdota4QvW4ZIJiPU3aXrz9CSkcj+sJdCg5TjGwq
j8pROxu61c2Jv1smEcF4TGOyMA8xfcZFxJw06jb8uCTNCnsLz4pmFfVF9kJRW5QM
xJiaRK9i1yKHuIEp1/cBXB3yivHBJ7XyW/KYsCMIJ3IU61eIZUNBJ6vTy3m/Fu/S
rnMWKvxLZ+1xwANwjyjeoK0B7D5P4euEqr3skFF43Cc/C/eL7DQ+7umb12rYQbt2
OMW+1tH/I2ru0BEao9ak0kMFKsMDGi986/VBhm0D+5+lVRvfwpsPGmGzh3krPetx
nkpMtqQFtSo9FvmGQmSj1mMGMYgDFxTBhyxpIoKSqIZH0l9xiOjMqYlDWKDqbBKY
RiP5iYYzO+p8piDCZjyRDqVXPz6lO483NedNIB+3Dq4dtRPV3nKsBvC+l6kB0KhD
DbUPhT4YsOf3tFt2Ztz9CHelHU1sKrre9WZl5eOal4kqNEfEYrav/cKSO1xBYu2F
GgEDbz7BFpFnNs8wqiA3WpUC8mkIq03cnNhwDY1owopWh3cz/kyxvGGbbrNG/85E
m20xwWQxZGBEE7UlgMqun/QvgOXX8m57EyL1/cycsfC1v10Bg3AHSEAKIoz2IY9l
ejm216f2lLM02HnasTh/+vuWlHjeWJbQi3EaNiURPBawBA0WF9hdrLPQTmWB7sRl
etWsCeXPLkFHEsFw54d9+oJ2M0XrTbzKBOg/P1PeQTdDe+9aTVDGsa2WOUwt+IHI
eAOKDCFxZNjTr0PBgl8LvsPamdeX3srtERpu4v7yvNGHAwUJlwHQIPELzPIoq5WU
70kj164XBxjfFROpkbX2w2LRMr+Mcl/ibD4RTS9dDtUaqKOcvivgs+06L6yrXx8c
F27RSHqDUZyU5g15vc+kwnD8N/Iwv8SEZF6ugK9sOytlkqUPeAwe2e7HBOz5pYik
J9akpc0wmXURLBr1PlD6BSlQpD3iM4AUZl/r8JCIKiqDHLqjA1P8tEZRfCEIRqqJ
RwUDeMouyd2KgKMm1uEj7kbo2hrSKBAistsAJjvL7oqPdilHgKJri2ClHnQUqEkE
75SUIqZoBP88++ppq6mIAqHEYeRTh6xq3NfP1dTSpQsp7kd7ICLu6ziEwuMXgA2s
Yuz43E3dQc8th+FJGtvuMsQ7auIfj0aO51buSJVoo0xmwc0fRuTR9/gSoNPK72yq
DitrEtDk17WVMuPdIBPzM/yC4a+dYXwvFDaA9TDpua0CWGa2THbaALrhk2CSlyjm
UtGuxxhJLHEsKIxwa7P/fDzX9QLorB4CixwwpaMoAHSpZ8bu+ypKceY3yKsb52nR
L8xTqx4ZHyp2ZjBTgBo3uQ6ryP9ULdzj3jM0uthV8MhEP+5FUIdrDbx93xdmQmT2
F5bk3VTDl3WhlPSwUjf2OPoxpmHZv2IgH685+ffx8Q1vvkkJLh2J248F87pCcnNk
FjEJmaPLGVV/q7QrL6BFEyH7GxOGFpb5ozCG9mFNAgVgpACrrDJXMxLmuhRY9qoz
oVxxOEIiiMeayhCwiLcsQLUaWSerp5WNokBxMi1URgAiVhQTIuHqdwVQimeRKT63
aaDRqFIUG+IoDkHQjiN8LNuGKFh5BBDtmzi9FiX2MgXXtKkMDjCtSVkW7ltRxArn
GQtsyDvj9z5aYva99PCXTXacbUXHtNezGdgWgnP56iqiS/YSRZabkmZ4HHsQ5uws
sTJMEJ06zmQnkOw+zSPA+bT6x9D5Gd6q1UcB4eaDnaQXTOs1fg6190e+9OS6tZc4
NlyAVkZTrnm1zkk9WdswRPBFeTCFw/b9ai6BxW5/Yi+tJAG8sZtcKHi7Gca3ox09
NUus+2CFk7xzHbkx3aTr7T/EYVhstWiViLvszpPcaPEruenfgYdz7Fh7+I34emfK
7GtZnoZFAlYxctykn/XM4+zOQjZGooiH8zeOT5Tp7od8j5EMqKWJmTnJ7aahuQOw
2e14mDERMEGlCv1vHvJcsvR21lsgKN2LoadSwHNtJvv/4NMHAd7jwMBbCZMM+5rU
1BnH/NgK5rodLlPASWarD6G1IKENBLscRXYpfPhBMI83BUZTsBLQjbGEG94PE8BI
JFyRb10X1hbvbXN1PY/opKeBjc4VxKjQZ0QzXOA0rE+BmLWrREAK5TFE9sl7PFiR
vJX4SyMcSk878LugosNCZPEp4fCTdafnK/v388D9UD3+t49tIVDIeRELrUiGTZ/A
lznJKDtLmlvyUtEuFNjZzOK3o35wyuUCV8T/DB7Z8gMK/a08BR0AYb1Y4SMypyuk
+7SyaV4m2WQJumfsjjtrNleUXIEpmV9zPgNUzJ2+rcFM0KAoJ1oJrFBi1bU+dpHi
JOpaPyjEIcEC4ryvWrwpa310HHMqhB02cjLF+1sEdSX6oR6/ykyYfb8lvw1g0oq0
bMpE/urU6NurgzfplN4w8o9eJRYGKc4PJixUngYqYuHZC2GfkaqOa+rO5OoXhnWv
/8AoA/tBLMzNBd82Vlr8GvMeG3lCls+92n7jyVKaknhzDmFhg5NRl6l5FS66oGxq
CLoJXHZKM3euA1v4L20i1FVsVH69qmUsJtrZwe1ZMq3LNPi+7aRgXn4qDEMb28jV
jBopFY3efazmxwM4pmLlMwKCUz7i3P1uoKuDyoiQncRr6cnZbJ/TTT9pvQHujJmF
XvDlwxRBuQi7kx0lq2sEgBNwye6OJsSZGhFNA3Ozx2d4TPwcQOqFBGfS9EIbBL4n
uU2E5w6BzzA1eXSjZ53aQu4QN2IZs/LI75k1LLENcDcqr744JpCEv3RsveQ3q+ah
gpFjPEYKSIY4dRKyUMQ3raKSFbLsqFgpQc1Sm+Nw6ME36bI2ge496w5y3mqqad83
iwR9OSSnK6/9hPwCEdEmMSNylf5HpdinUu9GqD+rEmWfBXTsaD7Gu0SdiIRBw33Q
cCuoxLK2/82dvs+6f/8bmPYWuS43UUsewvzgphnpE48FbMhjmZu32XHKRtBFy0qQ
yzV30pXz0ujiLIVWyk2RkcKKWeTbrY0Iko8ZFq/+psiSsc0qnkAY53zVWfcEXMxx
rRuFEGfh4AeBuACiFx84kJ+QTGwp2g8fi2xHDAa8M5JegDxXJUzoGGrAgJL1ZNBk
ew9JGiDVWN03OuJflKICTST7hkCZUMiwjQjOJppUNXuCqM2lcpBokEZ3m+RwRX3E
qPjhtYJVh1ncVZYgw1VHjkPheAjBSg0MyPPGADUB5qce9vmMg2gVK+88d4eSk7CC
h9DXM884J+lGD8e9scygBxV2B95aJ/Zfl106izNCc4ZykH5HRP2w9kdgNNdLQgJX
jp3pUPLxycekX7lxDRR2CDEID6p9Yxld7M57ulhB5f99fUFo8FkSXS3/Qv67Eq2P
w5wX96u6obhMryVZN2Wm7JyFeVBfQ9tP50DcMetzSRunbR9oPT1tF5zgf5YETHke
nJmbhVCL+MmIoQCNNM/ZtDq3djVM6oq0tDv+TSKYTot4uAfkoUL/RmdDRMSdgtV8
pEVYCcOEcZfi1CQSv78dPKzE48w6wiXJGHva+Y+SiWCbCXqWozh+l3WOYrCuGhrw
XI6cWAlDO4AIXYtxZTbJ5KBpYVHTd+ptEoCTcZhCj0ONQbnQTtoqqPIic0Fqzydj
hNXs3tUsBtnAb3Tm6xBSAvx5VyCdYoP76k+KMV8rnCrXe96r4x13GLg6xuw2E1Ir
D5m2q0OwRgqOMHRrxnFGOm+JR8vaF8iYsxCimGtLXIHGQik2d7tPei0xXHGpDbBb
N4fNfcEwiPMUWOyRz7mY6oZhjFwdDAG+yeHM/AqpNGZDmhJg8tdOReh5w9d55suc
z/TM00kBi8mP89EwRmH61XxmOEIhLB1Tx+lXq4QSqyjJq91Id78qeYyfBORe8jzC
`protect END_PROTECTED
