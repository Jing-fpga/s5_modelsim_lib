`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8QL7s02QjuaEMIblh1EzCbuhhPJqB1Fgqkg5JKjG/xGMJEjHmfXhswJ7j+g1wkLS
mnaMWbCBODocZfU/dN+PKpQfS+/6sKLXk3yUhM4pG65MhnSW/S/7yE8QO63gZCUy
EGb+5AmSdjdqueZW800ux3cbuROGGfm1b+5G3QmSZlWODkT2GXnHdFAY8MouohUj
eGZQL1OqR3IHLkPSCgMQe9PBcIM9Ren8g5WDum+OdqmWrplhs8EC3yHdAOP5pyZM
Tj09z/YyIKsgEPi3U6S7KkzQ2yNi+QcDcqLWvVlQiZnrrzgTCv5TPeESvk9jML+J
RDIIg7kM7EewGtPsOLYhNlDGpoPwpaV1jdTLhSb6syIl4F03LqboEZ1qGQgk6oe1
lR3J6q5onhcuE57qbL4XFDdLxzLFioYTiNEOB5kB+npl4tWc5WtkO2sz123DmdIS
c1DjHqu4GiXkJtCGRQ1vO8nrkYvgB+N1YJ9oNs+oFMKGkz7OpwowXbR2Brv89jt3
OMlwgUhBow7IuakHzhwvBEFdaztTkWgttpWkYCtDgrpmUnbO8xtHaXR1qvxsKJ/m
1DklgCfiWHOm4qe1uesMljg7FLW3bUC6Z3/ysjajU36a0T8SsIl/NbfOUWMRWIs+
0fAiZoN5F7ah/rwwYp9khrjDVgytI53kH+O79MQwpcytG3gKBZcZDR/+dqi0lu8q
L/h/AZmhiEmO+M86TAvPUlj8A9wEiIC0c4DpIQ57gkDjNy25JiB4X1XTxZoLpOhb
scQE9dArOFq41jWGV3paidPFKoPVOHBQy0E3HcBme1oXHMvqGbRuI+QA5e+WZ3EM
1DNpZwP/PdNtZVjE9PTD8Wg70BoJjBWzPI6161t9YxpOQIHdu0+Rym+6LKkNZG2c
w79EBh2/kPxecylIqoNoU5O3gXIWgpHpS3d7yexgAxUFq3eJ6gIYRlgB5R0rLoRE
hWfkPCWr5BSB+aa/Eutk875jtEdWB4jQbYH1QOh7H1nF7NWS2OP7vE4AUd5i6sKd
UdBYo26SnSxXFPXiE7QH+PotwJKpJCvcLwWC03skYTlnN67zH9rxSQzA1XUxOhCS
mUXdfdtY3OtUTSGO6iiT/E9M+feII/XM/kiwssw4lKZxDE/LKTQr2ryNU4Lw/y5N
DY653uBykzHIobEzIJNwWgTha/9owAi0d01Hbdeoo0wLp6cBfTAQPl86Km4dzQyq
q8/FLcp+FR51VvPkh+Tf9HKuj/hcE4OwJPijlmOwYIcygpklGm3D0l45VjmWo7ks
VEOSB0NYvWyzk1rNdChzUeMuMACnOp86WJexRf05yVczw3VmP6G8CVGSPJL0i8+e
T+W60f9SdU7BuV8JDu5iZNT6nQSxNUulxGg1xt95+1QliTEHKvZsj24sR+PBY5Z4
T6UrVD/8qzRH+uYg3S9LLxDrHFcBt5zs+q0YQtfoPb/i4mqkdMam31mVh+KaNqlY
57SCnkQF0GmXECrZPh1PG4ViRXZsx6XVgSqQaJZXcQzpKea7GaFAQ8FsIAxxgjIa
MY9xjYqH1PqHMmW5W+Dn4OsYm1543LRTQTGrOdwY1vHEb3iGI+Q3KrfeZJIR5+9x
rIEGxGuFDbsgyi6+t0LoHfXvIVBccykicQxc4Y/3TWV0ikqFeejawhNZxsT3sADu
OACJWFEJ1opsUXIwiL8aht7uPYP8knpwOlT0OrN8O8asNbaTAT8W7L51rBzTVVaJ
QEOzo7kb0URhYodbsT/iCQ==
`protect END_PROTECTED
