`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
irbUNW/jFte0mSVmBDMwp7JYtWyIasu7Ci3kWvJrtVDU8g47We8TyFs4X140218T
j9Fo+zWYQLEOwJjgd8fOpPQbp7x6DLUfLV31hkgzcqlHpnehsBxy2PGtpyLc5iYL
lnxaoDTBXcXsEkpY93HQsu4A4w3JB98S4X49VPAGQ18x091g2Wq21QmdzgyfviFk
pxE90j/PaeYSdfLqr8G2h+1vJMte1F5v2KBxR3FiHMPwXEhemlVZgD7GjMTwT1h4
1I1EMiv6CMhgPMuAtlCKKZXB77iP9WVxCd5RIleTE9KVueH4KSr7NSGUGV176onS
TzpXK57vnfTiXvr3hO8tRD18fQHQ+MqfC60MxXhZexo=
`protect END_PROTECTED
