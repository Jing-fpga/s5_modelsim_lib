`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
spqyzhsdE85n4p9Zr4AaVkCMkW/hSPUDfyAP/qFs+hggsle8ztaR4MXyJGHyrkNm
RkC42Qqhvqldl5aMTIT+PvIJCF6WPycuTs5urbwLxspaH373AGCDJvcvTKP2muTB
GYhrjPtwerkopHwDQOFQQ/jTI4c8cLnMwSa6lzTrK0lNEZhFeuClBrdCdSIWCo3j
4KM3lY7Ft2evx/bhgXjbYhLOIiVaRJwgCi63rh++shRs+HKmD5qqz/diMZYnvlH6
tOr4bcM4DtO70oSCTFvuATRtGwmxpKO5M7g+VJVeeuRiALH/c1buuc3UhqWl70RD
xpN2Qx3QqAOYZFkybhcyjGbr8uCtuo4gkFnksUGtycnvvYEEwvJMYcG5yxGnFo3+
99Y2HBaA+HD/N3S8fmBHLPKDJBt8iuEi7PP/aS6orRFj2ESn/Ab0+CA4RsCOoWPA
PGQEaSwM2CRleSjXCPI5zd6IbkZdInxe6623U9nnRsV1iEPrA3jOgLaPbgAoUsEF
sxOU3RyfhS8EgzmKFQ95r2QeraS+dmhnpWZdfsmfPcVdlMEIY96ou/EfAMFHtpXY
+JDaNXXk9XlTvp0sArrk1kr/0lUadBLTMqCslKRsT6E5waHtE4DWoVqgU0ViIPwq
2uZ3iAqi+bnnHzdK9MMDR+DEcDohB9XSDwbmsAB3P4lVR2PqThA1av/ABgzrAic4
7TkDbKbhmi3d1aVsTffIvn2vMqDNLMPdEf0h3PHWsba7Q2tjEo8wjias9JoftKmG
LEenk4jGbNBLiEY6cgLWUNRqnYMfn8RLlt1YEfxwwQJQkTiJFkfYR5/SaLcLJFWC
WJJd6lF1eeJCsCj3trxopIgXg1V0zECC01VzBHxGW5akhzYWJhBCBaoygSQlnMRW
dT4Afk3vJfqoJHAohQxwlHV2l7nWozvUlD2SDGijib+Gy8PnWKdlP220H4mQwQOK
CE/UMyzvKHZOYBQCKFoMIr4ESnPpS8MiF/usnsl8aVxK3IDm3Z5I2NBS/OF95T91
7vA5v+eDS0SsPyqvKsLjHRgog1k3z31udzqAs/FEqWPaGtPEQhGhKr4BAyf7aw8d
Ith0IxfSmMtGZPs4qgy8v7h9+ixja9wbePln+y1VuN9N+I1oIY/6PtcbssMKHqSv
FYkGDLzMJ/X+nOUIQDuGEtHhL8isaBPMUo/SMsG1bLNXf3PsjGX0s8dSMfoGVRcf
xIbQi7asDQYIFfbKxXnajyrMZhBj5KmIcZ8NCAuaEHqSOaNUZwdKL+A7VzP8de19
+IXNHgjYHs1lZLo/1v4dCJlL9H5/ALpLkiUWUZh7EIahvJpe9RYNHyhxQl7sKg/y
NA2Pu1FXFXLbN7PaX0py0DK9rtREoPsLpJ9hKZ07X3ksV8wTxHMK7AYXlerlQs06
8LoGKKk+Y+nuozrXkc7GtaDEk5opUhBYh2qM1Fcjd1VIgVLSHOLDXy/gTuatLIrP
GzDn8L9mtmyWQeYQvtlswCTsJsun2skQt7utjPgzS5R2yR0ydaM7wYO8GEocV+Bc
g8PVDEIblCy4F/guuiupnlo04sxfg4nx/dFrEV0RZ9f1BhQJCAc9z/ditM8A9zNr
8WYagZU/aGTmrOb/pynYStgMSMXXUmfgZHJOXTUEGEJOlTVZ2prsgwFJhKmuichJ
OIeTsI/JfKhNJYsndYT3vqkesGREiGqEo2rCvR/alHtSIDg8dtW2djy7MHCFRHIT
yBeJ/nDJH6gWuGdT7I2q/0a+2OEICnVsJCHpdeSHA3s=
`protect END_PROTECTED
