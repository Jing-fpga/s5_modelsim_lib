`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zKDT4fD0PYFKsdlDXH2F8kWIoUGYpmTiaUpKKsXv09lQkLHgV07gt681cSj52e9N
fOFm/KnE7gb4E9X+OF2EXYzUBtfKoQTPZzstgBRIIOT15Z1c1ryDc4ZX4DkZfCOw
aW21p8QKr+YjWQcT+oRmjj9Dkp8nFRIPHq+wjnHUIpe33MbYiHAgYiIL6kbAmMeE
uP8uTW3Cgb+xGDWTogEkaJdsD7Zb/AqSyL8oU4EHexF/uKzI2TtP1MuXCIUyT1v1
0DVKJVU5I8UJMaSLswvxuPRMvUjA4C6lxBTJOQTyR1eNpTpc+gKgPDdFrdiRFWnr
8AlLjwSYEIYQTAUdhwz/KAgY4WbmpM37/zk8bmcCi+rRqTizM8yhAT1sr/bIO3Vh
n871w4c05C6UDejQaY8MgAgU7x4tekOYCbuUKTdWWmoG5n4EBl1sopddRsC2d5is
i9+3gfSvTMHjMws5ACvg+RIaEdVUJExqA1rpmtzv6eNX42DE5wi1lYk3tbgpkLZM
RO6mUxS8lolDTZZ4iV4+zXeqowlIw96Dyoe96pyUqgzQ5ZddJmm91568+wu9PG8m
Q7R6ZZOuGSjByV6QegbNnEteHPm7IGLScnKjkZNTwwyI1SUERNNsIUy/s+gbFJzX
Co+uW6wbv53cFq+rHf46OKck5M5lbqm+5XGNnaFn5GNmPqTF9jgLL4ZPH8P9hN5l
Sf7lbfWRs6nSWxppaUD6iWmS3c3XE6yLrb3eToyXNRw3C6kQ1ep6zx48UW4aTYBE
Q+uyD52R0Mg0j/xE8qkfdo2D8is3U9vsQbRVVaFTNtFxguIFiaPhcOxoyllsqD75
pnTYqYg0mKbRnZ6ZPz05sR4fsondeGurqTzFn+jubljwZRtTBi+uBr2ggG4GsI7C
aygGjAtLhpjg/EojlJJ+FBXQ9NmGKL2YfkxMyeH0fMOfzbBwYQP1tIUr+rc3lKXB
iFbGctD2ruEROtorU1oaW3b6xCLg37+M9sJ76qsAwpAHtvy53wnMUomKNIBI4IML
1yKy0DlcAhcnMYNzWSf3gyufsY7s0qt1BlOR9UZHSgxhFKMpOuuLQcgdJEd0CeB8
KM3QdZSjIefnZgHHdjhz+SUtTZ7ZLQwS8clB0E56ewVfRm9iDgAwOA2LVY8niC8E
4zwZqHVS6a2pSQcEtPf8yDqIWuph7HKYVZ69qqcEAw/E4GEexrEog6mgJyOq6MMM
wOBHEFhTF85FL38m0g3ZwybsZT+5FoGNcE1+JTQRWfhFQKme/rLc+2Jj2XsXQPv5
TrwSX1pFwV4RxmoGMaiEQrcOqzkbwILcbvAcC9wlquDYI+lH3aWnIdDuzBNBnflf
FJJNYmsKAyc2XmYkeDE8cQ==
`protect END_PROTECTED
