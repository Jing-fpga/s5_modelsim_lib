`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Whbj8zlcjiu+qARbgpii1KIRrFMyYVMv79i4/AwZR/tztCk/TA95cZWRlWgOCTX9
p3+4LhOBrQCBxVn+GKzEpFyFrbkdW/lImY7T0ePwRCuT4wcSByQx3VQkle2oNaLx
EMxtgHMPf4EzqinEh8P9ox7VHSl+Ik/i6RY6e2QQK0Evxxrz0gvfEayZxBW9Qlbp
wqOv4JlGwITRK+Vk1sZeSikAV8AcRAuTBK8nBlZHxWicy+jjLuHrUJSbfdkvOlZd
Bmwp2kD7dnw+qaT3pKQh9O/b9WD63bKix+F+UUDqHvaOJ6j4u+oZu4C5ycwPxyMP
68gCkp9AfuINjU3poGmxl4MN3XtWHgKHUf2kAX7vGbwrGUc/Uv3tdYlbcvPBgumt
+6EY/R3y9RTX3u842mSv3Ov4XTAkLWangMWaHO+tGD+nGYgHoYcgaB7wPISo4L7I
lk9A8JYoPEVcxd+N+SDnqjdABSaDDY+PVqkheCLCO8ahAthNoHrDZZ7aE8u2Jk3w
ixAe5Rw6m7smAX91cupBkzB0F3pkSF97jb4nwpjmzrsjfOlGdXzetelQaVYpGM0g
tR27CPdxoOwYZVSih/QgKFopDUPV8hMkmFtmckSbmuQEEo9JFNm6B2OXf44vBD6o
vXcB6QhwMoI0CWk5jXIVJ+w4ryVShoxwM6imv/8S7h+s6TIIflECPzy0Tc6DI/xh
gf3e9iJlW0BAKIqC8U6FTymgdj9+rg6mQLh2MVN7p9UK6GKuyo+tXZQeH7W+Fklp
40hg9ewKdbkhWrTmSc9WeYVOwZMz16ssgBCjf+VsEkn47CEkViIdlj/z7o+F30Rt
Q43JFfhnNQYiw4ZrG5fOww8u93qSk1RxVMflB6UIqdpsrczejdxtTy9lrEuVvyFP
`protect END_PROTECTED
