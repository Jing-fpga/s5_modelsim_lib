`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sdW5ipRx7yglugu6w+Pm5ceqGo+lmtuRqJH4CJRFbTjTHCsIU+PFNwKqMdPykZ5+
5Nhzt5LWPICPxOEaWF+9e1BUtzHTR2pCKentvI4jGGY8//qFqbbA8vi54FYbpEny
WiHUxTl8OvbUuc+V+KDXsGVF4g17P+YJKIveWR3idq8X2MRCCundsXZlOpAG9MLK
XkDnlkW/ib2AfMQ2o4KVQ+hw9jHb82s1mxFQpAaxvJRA8MRXWQAQEE/kC8WGUxCH
/mEQRvxAuqmyL3NaEkb0GqDDINcWszl2oG8mhGtLH63Uy5X5H5Z5MDUhl4YobLSp
agPZpBIxQ++Een0ihAq2O8vn1HrBSlepqw34Af1kF0F5oAjdtEjDcMyP1Mi6oUR2
OQzwmQV9MCBxO766V9IX4VIlDJcl1m32UJI0IlT8yxxZwI5bF9lRMgRGQLtUmtCk
ZPUvrbjnJQSa0IRk0Crov/pyGWx23LZyMWYOKUYl81tj0GiToTJaQpsZ0oK4DRmY
lrOPJPA4sNe8003k/Nyn7nUvJWqErfCL/MFX8nXLTg5tHGlM6lTgYmPTMuawhRa+
CVDjLELIiT4wuaQ7nmQVdGqUbp1YlCWZ1uCEyMjO0xwZN6jdwYpFxlD+bOV8Hv07
YwZ6hTHDDCKyDYwQrdJceHdXfG92xwzR0F35glTwA8Li/wy3zcyAMkUuWPugq5f1
Wqxz8RFut41nglLqcleT39L+QcUHxAunBRe1XCzJMtOJQSUnkKR7AxuXzXFZvVRg
Jcip4b7FSVOEAE2JsHJCCo4k7zkggNR7jImvLSx4lT3WLwqpLwkZ6MJx7jHUVxjM
tqfudfCSMCuM3G2N6bU+i9HdlgYdjpHPQZ9D30fpw+ti6SlxaotEf/UBVMMjMkPq
kG/GLqpYfAr4tX8DLUQKK1BA28XOY/wVpi0IfdlcwysNjyttWcPepOCQBKnTzsPN
hfa39eu+KDLubpGaeCO+dKIHj+WY/SH8EmMZFROpf7s79QYQSPL471zD4roS6oZo
EKSql7rCh90Fkc66R0DAA8baMZBJdjxJhSnNsX1uebBU0QqgJm3DIp9c166p0gWD
JASqoC+2ZTNwjq/E/eZn3HD6q8T5oz/XTObU+OICJz8Q7KZYCurw7C53sfnVfZ8v
+5uFY1rik1C4PhxVbGw/QpWzBUGN+1h3NY/NRhy0tMGCev2+76Ve7ErVPkTNbyst
mKrkItIHVViua7flYcqZxH34HsbcmDCWceIVV2XLohqRBnQ6yGKndY4w3VTTbm2N
7iIpOWXTmoBzMMU2g0WThpfi2n5N9A751ogDYSz/fQuozIASdvNB1G8oBkf5zGdl
wU+QhtKjt7SwzvwfYWhXNjjbPqckoU9LG7lIMidvrqlTQ3eFGSpY5bCf7bZb+Hnr
cLbGv6IahU0nzYPNO9R7xhN0TMqVhZSWxDc+gc/rop0eW1JebfXWs75Hejr4LQRx
L0+Pw3pKyWe2a+BkylOU2Q3e9HJcP+QQjNZ+bjgViWSYjX+Ps9g5+qTfp/Z3zf6f
699osudOpP9UHoAbpaRMV4oYBIhHdekGX626FbXDBIzXTg2mV2X+o8DV8KqcLpYI
7Tor6CMAj0vb8SrWq6sEpcol+QOFpfxRuDnVK7qfcX6c2nx3dZMM4mDM8Q3Eey73
Yf/rNNDYKk3KefHnfeMq3CoV40b3L1UOBg8A5Ws9Az0rzyCX5+IuaZ13DAD18Vnm
7rzlmy8nVTDPsj3NnhZE+gJ3LQhlOcFMLFjsfAs/8CcwIFdBxCIC2MPoIzFbdUum
WMVyWpLbMSwldQTnJC/5VNOnT1HB/zAQaFXiuxN9ujnPVEkj3z1EqnAPIhsXl2zK
FPK5ugl14nq/kQS7YBXpHHaavcQygTT87ihOinO0YfdMTQECj8A0cwbnmJk1ViK0
zMTRhbZ29RS8pzhk9Jtdxrh0aRgOye7tQej9M+vw7r9fCplCcGXuBqxKkxey2Ehd
ZGaDc/7harTEzZZ/Gu++KKx4R72prApL+f+cunG2ngfyWuG0kvLwW5VX5FCkRo6d
WJ5+1IHnF2BS2/vdHotVLRcKJIozNLa4pqyvdCgvqKg74zBMMlffV+u4eNaHdVlA
lIaL5kIB0BZsY8hZ3FMEyamUAuhs3G4L4WVXnEN/ehdh2Q/fjF2PensmefwV6jTx
vI88pzTl4vQ8jcdLr7c5HSKmfAs2qem0ek/qnHElJqhkNJC8bXP2u3Q0BoPsEZf8
KZ1Nvzftf7R+FeGyfpIO2fZUjHTYEJ/JGPVufPO3W2XsBy/NRtNVv99GjNBxxStN
cqwSp5F6WBniUTtNIEtu4IbAf+Z27lqqYPqyDzfImjiIBA1opA8OlivmPO7JkUrJ
gSQOzNxUj5TqMM1Zy6kYmqkpt9Qhuf7mxmyqAtf7G4nOIbWhc5ypkYRHCW+OnnFt
HC3gAh+aYyIUkzx9X1klvgBBUAA02tyYXnM+TLzeK3LhP6/y5KMNKhARwoTfXUOM
MNTRFIrF2P1jXnccfpy68jEORUF2kpEXkSGQAtEwQxMfmMCJdtpIXwhldUWIDYq9
wtA22FfYQCJqbkWCc7gwL8NJe7RS98qcKhNKeGR39qYwCzwtWZjUnuwz0y0cDjjw
wvmtJxD9qWjZNSxfa2PWq8Oj0nSqx6x3eTbfUsAv/Z7pkofiU4+ErORYIUy4lqvB
zS57hhRRvkNKvjHgpwLzGCHL7ZgOb9zg6sjERIHTda6zBlB7J8lTrAJ09Sej8Cjd
9noowkYkpWD0Yovqvo29KkJ7LH9kDHdpapnLkCmPovGEi37931lcdE5Jldj9pd3R
B/liCsYM7l/rRlSeusg+ODRNB5wJoFZaXrzYaC6/JYptNEC0BEH7nOaanG9bmgS4
ZY8befqqK4bcSkANnLruhx1cUbx8lHIAbwKU6hAhcCH3SeVElfr4uWlslUTAcp5I
UI4Y4Y8PW6rUjDJxCU3q5rDag6mkHGzJa6A9zeX2sN6/MJ7rj2K2QgbwDK2n2Fh2
qZBM/XyuTwmZfKJ5pkIeXNYN95xle4WLq7woYLfEWVWLlv0yK6wvSDm43fZL5LWo
SsT/H1SSo8oSNURNkdz1OheCsyruFQgHCfoJNDWvW5rLsM+qeQYVFMucsmAsqmlE
SDCuAATPcAH0Q7FhZcgP9iQjwPN4w517+gcw5zwdkq7fCsAGs1zUWQdZKt/fLx5w
o5sOXgmdbG2V+Kn0l/IxFcoc9XKSMEQJ/wTpekLU7mP+43CYGa0+v/0pCu9Dkwnw
fjODqUHEufu6Bo4UBv206goMGsjNa9weqMvkKkzLU1k5wwQWR+EtdIKJPSZgLlu9
b3peFWuH6iidygs0ClwwmPVeVSzAraG2cR8BvLfhWkgjEOBjZlnmp0ZaoVPAMekZ
o4c/MnrYKgc2qTpIhp6j9JClPP5egOwS+El1mKBGqjP/HGPU7N8vKj32KZynQDpn
DIn/WmIyb0HnoGFFLopGLGybjagc6zc2bFA09k5blyya1W7JyCt5rG/O+a5hOIGS
Q870P+LfdBcFqpwBH4gNIEsGtC+uPSRALYd7ASneM0tQOiHw5tPBj3Qn6E3tIBjo
xzuzVlqMshyH48xC50XCc2+ZqPBGHndADUdrbG7uD3AYzw3XRKng43vEJlKcQloj
HiCS81lUGXHHi9W2qqEJpnUp5fRgoFm6uPp8NTH3hOPPNjnph80AGzBsDIxnoX91
Y9XMdUSgRELHzeZM03FwIL7p3lJCz1VRN8gKcO6qbM2ewsqchU9AyHwSGQUlbRqV
pf7FUkjSNE48eKHzEhcjxoZNWhFMPJwRLNTgUxhpg+HwgQdq51xEuEW5GBY1FG9N
5XbqZ4aFx8h7QjOdrdtSUNVe476cBlnSkrU9zcr62bPRbGjM0g7Qn+INGeHneFyd
8R7Ew5gvWD6HoanQvqGKFP/NbyRLBwFOlpjG6zNaT0x7nCWmm+fINsaHpETkFdHX
uh46kdVpV2LN5jfAifMswfA0OaLFGFfqQoohRo5JwUo2pIxhvIZB9ioYLb70siOL
XMa/OfaU6MVlfODuYz0hUo6ttMpHhCXCbZlDjMOnIlZy3xgX4TyCQ5OSgwWKYryP
xWLtmDu8STH/4t4Fgno5PWiOrCrd4Yq31d7VTI7Ezf96WIMkaCon19Ut489KOZwF
55BrDhQ2hetG8ESKc8NYdCGzWYrNjWWcGc6p45FLOKl4YHdT6+7LWlICa95JbNqv
j2YNFTWFoc2SwFGR6bmOAB+6wwK3WYsbrNsU7YbCGy/a6LHDL00u9T+mvMWfSZqx
+J3LDjDexTmOr4gIu7miaaYaLpv1pzM5vw741h6/HSFubuR6Jkhk/CAuTDNNQigD
G2Y83s/RUL9ubmeGCS3/27AcCIFTndkvRESQ0DDduiF4/3Bc1T3aU0UQ455Q7hKO
sBHGOCsHIfvct5evaMZZYo76G/c9gexVva9x3l9e1/XKCzG/qBdoKaYIkadkqz2U
R8sJfe69hpLZigtIM+U6OdUF3llCgtMDtZCyvKhAGfDQUNr2qmOHppkCAST226Iu
zgZTI6R/jJHxokbxX7YorPOomp5fH023o/BxlUBz7/4bYNW+STmVob4f0ulkoDwA
vhZ1aHhkZfjIZZt///Hjv4x9W/yf2V1iJZ4deKXwpCGlChzC+oywRyEYaRMEtFKi
dmXZFFHSDLX8DtG+aCzSDP1J/4AFrSlFQFdQXAWZXHcrkNlW6WKkZAe2dMUx1YtO
VfIug55HDsA8gh8MIbi2z+8thUQixKw/hBrjmusc19riayVLIWTFQ8lDNgLv0Xbz
qqAabyniGgF9y9XDeZrXxcmOQRrweLHXGhO5B31s0aiimbhCm+lC9BFjzTgX/J5j
JTC2cBr7yIh9UJ6yLdIPr+Huv7MYc450q7pj9d44NhQINWrHS0e+lXR5g+kqSbux
g/IgbFESYCUSrKrJvCxQVYb4a5qlursXrWJV9v5FOOIUIK8ueA7cuyBkLvImucdz
b8TFLQ4pu5Zc1/Lw6SqDJ+150Oh0+TSexHoEGl6cf8ymUfz9IbSDWtH0m3a8S999
sYWAMPd6gEfY1So4zVStGhfUmFMu5GAQ2To9NKmDng+tj7WyHhHcioc5h+2NYRHn
TMorqiatwwPZWxQ/9ATiLdXcueHT+5KB5aHEaGpm2jDxqlsIw2s95Aqjuy+F7ndm
tStp6mcpEuHvVOZPvRQ/Zxk6+vZH6S8xgMTNCWKE5+dh33PhQgzRkIfRuayvmBIp
QoisPS+EJ9aCApkFZCyjYoqpWBy4yJ4EW2kEZ/UIGlv/x6408bdw2AC9eIeh6H9G
JVvzl1P465YdAQOPJo9KuS/zgQ5Nq6f+nTqXo0c7iUaUIqbQA1JK8acWRuVwWUeC
yt7icdDjZxHPsotia85MGiwdAuMZ1ksTq6eOfN671oqk3/dtESzowehcSctdNZcS
SmFEsl3FjUa6pEUNSWav3CGih/i8H+bzneRs+djAPdV9bXJqxp8+pRurcyP7Lagy
h8CFBF6Kkg8XIRjWZDBi5pnvBCHFc3bpg7OUhVt/gQQbXLB3AnXwSWpbUVlxohu5
PWC9K57d8Q4Qzdk79X9PbQlIn1jknd6U0G1gW1SioQCyr8XDEa5S14c1UuKRZWlQ
/bvVs5/Mbo1wLzNHBc6cVtKdFMngJ/ah2ZjUYzuG5pSZ+GC7MuWFeZBntHB/4xwI
pr38GqIrD/ism8/1wUvYd5/+unXzXnz9dkXHXGdpm9XGEjF6mOkUMe472N9xyJjv
MKIg5Z0PKln8VX0oxkOfuZxUmYS2JW56B0iJC0tQvXBjnYIvuoK8kFppcLBxZ5Id
+N84FCdgIeKiJ8CTgwQzzxkQeOjqzCwRAjqetGuYiremUwLbXJvgCQyRnvFDIxJ0
qeLRrDWcWjnedgyQBo9f9/wIWVtFmZLJxxVO6zXuWR0LVzOtBR+Ti2Wnfd/5z9/R
yt4U5Sm985MN6kAzoWWwgRX8jhwJyje/7eMsbuJFYdYWBYukAfSLujwJMlfMgTg4
aovimu36aePn3jq5uJBxLLN1OhTvU9ameVA+URGCAyiPqUJAv1Nmhk0uMKB9BzC7
LgtFTAXpuHRFbR3cvj+6fobwhySq2g1GAxmkEs2eJxw4ExNQVKx0vflk23F7ddb6
flec+VN1SGB6xPX+6+B3vKOZIzE0k2oCEieP67bY/kNCk18jluoLWHJp6DOgm4JX
fJNeNInLLiTJ7zX65zNM9UVLnJdGw95kHx+LdAzVB4Qf6Rw3vgryWq5Ll9gqfDLV
Oo/xb+nAAKNawWVOkhxv1XiW3qUYXpRfM4xrHFgR+yJgIX20aNDFrOFFkIySv7dP
AkvXoMbBMfKT5qo6VCoYggrtVs2CB8mbaPAxTlES2Gv4WmROaQmcnKbnTwyXoN/0
UkeDKRhr/4KyfJj9xorZmJl6cjwfYdJfD2iY4T0yoiIiE7FS1bXKTGhvl6xM+/Ui
Rrm49o9vBD1+eUEpfkK67+fJhIprC6zr2OYKw6bLYGztdmH+eGEWywt7JQJ0fGLP
0DIhPBxhSMmktzMgH1Hdot45E50cq/DDg+e3/XQn8/JzkK05W24ogTsewvT+4s1k
s94yDpc7ENwDNLEuWxO0XDpJ/DQUkQkzDqY3M0O3dcRPfc1H4xIkEmDJGAC2jsgX
NaqNZDQJE5s4QVXMGWXPfVEV1ArDBqfBZJYbAhs1W1AlIGBzrlRzt/yYIltNKtC+
0temViUipbeRSOHfFgRSPu8I/Ks4V4xswyhF/ThW59mRyHVlXN1yjU3nBAqt9CyJ
DeWSqcvRJxR/QIXPcGoc9mfiEX9whj1SO6spYHVDpijbMs4F785VYEZY8rB1hib0
QpzdRG5UKNOkvTRqnjuRXrWozPLRUi2JYev5v/1djv31LCae50PrvOF5zU1iojZF
aE/Ku48v6ePwGtVYLwyRm0fnL/tTiHMUJUhUrpSCkXGBGtseZPk/8wuWt/zuhjpk
URoWyC+smf3YdN+1LVyKOpNyFReg4AYbjJupxe/6PR4emDFh6zf+8oGmhqn8pazJ
M027Vs4Kxh7HklbBfQf7BATxJTGAmwwUguRJ5If2L1TWDthzhTa30NWU/xU0qPIE
JPwHEdrtF/Iw4D52SZnCRBchnE2yqGBMJwlCi9uImU8X95MfEhtvkpBBTfBUiqxy
vuB2FByTXddWg6nFpotI8rHg/z17euBf4IEwWZFVZwlB9yTs01ibYEOTANGRthNi
RN3EoJKgnDrBN+8AK7T3EBxCQ2F8Jorg3hVSjdtgM4J2b65KyAE/uRcCx7por5O/
JJrv0usg5YB94VGq/LQZ5QF93kZM7RB5NBIFkxkJ83aV3iHr8OvQQWNDAJjua/su
FLe6hDPq5rIu44XN76qeV+0OA/M9fN1Q/snirtrc95xSDbmPIgnr98TVE2A4v+yW
z2Z4IKCMqOLtEj759V24+iEQ3l69NB+F0G4PzCFToDT1H8ww80Pqgtd8bL6pEGrC
33ZlcsFQh2T2f/Mk83sEVOmIxxwr/6nPqsyl9mLaMw7xGA0RXQCIDi9GA7iQS5Db
2XAPTREBIDKyaMon2JFcDWyhbIiBMN3Wmdvz5oo1gHi5vWJkrOgizd2WH5jAZyh5
gkfmBKN6vdOYwq7LUZG21th3NcbK3flz40H1dYVtb4JFkKBgIFQLdnp72WZd9QrE
s4PM4oJ88ZDKuURelyZgbD10wlYknHC9oWDzqmF3iMr1PjIsG1/jAnNmimOkOkNn
BiyazWMwQgkNbKf7P/wz6526pxGDfaWuvvQTqb9By3caE8nqGV/b9OU3Ct4RWh/e
3t8Ecw0OpjqOWG9CMLbz9ViyPkSYQ+GxRGGayUqhe/xKj5pJ1NfADhV4FgIgID30
GP42DGaBuJ8W3sAcN+hAT7mcADcJ2LfGw2bmJ2Ql4ESB5GhUo+hS/KgHzrT5tbvg
wYXOBXuWQB/6TNJx4EP+1n/WnLJAHo6NLxUqebpMhtRXxwQbX3YS9/4T3sAY9zg3
rfJUTVziW5V4gzdY4qkpvs5qwUfAAm/oM/V9JkhNx9Eqa3DBYyswdbhsoKcoP712
1Hmxb6/8mUzeceAg7AinsgAlRFXsEaYA57UxeYl5o7vcj0tkUMR7Lb/esKRvhzKU
AXOmDUHuNleN0KUJm4LHy0JGxiqGO8N50iSCEj/IlTOEjDuApsp28iFlFoCTmpVb
JKbe5JZVttViRHURtwLtSvWUum4/Nsxyd1sLGWyPGrOLnrmoGwQCH4/0aPd0/vP8
Ou2eLew07UgZwn1dFQ+eah8wIrK7/isX6G18hO+xkcPw6l4PvCFGn37qHg3JJSaT
0jtQ48JT6k6w+sBjEkAF84samEHws6774MBgtkVCk+PqHmMNhBMwm0mX/CnpLE5d
/bSdyNBl/umSEu84ZshcC6ig7r4KPnXkMcw+CJ5rXhMR2x4z1vahkTdlMdb2glim
Zmu/5IIdF8xl7xU472aoZXYV3iyNAARMETtrDwGDxN62K66J5m4TaD15rBuYFYOa
qD1AjHkEEo61iyP73QEVarFqH2VmpdaKqppmxjVSNfS4HrFppZCT/ilTvLoYJExi
743rwJxYAzdwduTA9ogP1SY+gYaMZxqdd+lllv044aTVydUfSLGJT7IKmjHwDp76
+Rr4K2DJk+quRH7Wmk6PEPDvm8mGEYmqWVEA/qKakX+Y0nH0ijz29joXsTMyqlQl
kufw6QfaSIXimc84m2Cwoa6u+u1vAm8W0zkbZgcYCBG60bY77MqrMbSZYNGuOb9O
fk1Zmj1I6p186hrP4eLGeQpQIEe++np9y9vk8x4lHiDwdvvT/Rvrrr+YZWp/D8wO
RMnN8Khj9FtEf6RgACqYsAOb6CyaOpIK31z7l5xqPDYcut74bDMMwBITAZgonugV
Ye5eI0cdFx62XSbZJX4ROG84hKFqsLxwWdlQjzYO3Y0hQloDl8rLI+ydotsqIRCP
nwTmkLtT/ftcfnMsmW1IPjyWrWiolOOCE7sc87M1C0FPqDjcNhv8jJnKSqIbqUYp
cFUWHgmPUngcfTP23DFSssq960FSxs7KYa0n+6lEquvkvuF+mRCptFHSR1ru5Mjw
xhaPC4GtoubcBg41g6qFXZO+Oh0FnTlZEo4OaBtE8jTKe/o54SgPlM7UNlyzWWLw
QY/Am8x4hypA12hoL8ps3gcr6uXusPsJjdn7V0p/YzhxDNyXOa0PCY83y/QMjoFG
XjfvYVvEFGtZPmQsMlmqn/Iv3WfiaskhTRBe2quVwJ/pkaYUsHoW5eowCVR4HGma
qpWNQqxlprN7kVc7dtiNtHPMq2iHAnOJn9MipgN/kWNQn5G3i4Q5pNqGmWopwIGf
zsnyK3JapFzeZy6aXBrA5I3LYWVAW6CPAvmdkQxdrQU=
`protect END_PROTECTED
