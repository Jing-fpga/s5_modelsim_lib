`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g5ruKwhh96Cjl3H3QcQVg0n2bIMkzZbFdcapSyhba5IBXO2ronIG2GknoVGut9nu
HTug1LyDi5stB3BvF597pzhLkAd7+PU7ehUi3X9xTSs1BHhaccRqdOfe5hnykehG
xdFTSbnohvVM7tmak3uyBAqhDC3r5XOpliVFnZ5kI/sbmuM31aj1sVvUBVCLE8Q/
pONzUuQd/bFjrtn0h2XBtqZ1ed0cJjvFxGmTJVIsw/ogt/3KIOISOYPn79Lj/zH3
jZ70PT4QcPaoF5MYhCweFffz/6t7/pVoVcqHB0KSeSuMtyfe67Fv1NJn35NFjKcW
fDEGroiBe5rEH/k7Npunhmu/w8T54I2ed5RpAELYYyHO3rxaZZWRf7deppiq4o4o
JxXIf33p9QejCyL7QBrfKeq/Vq8DRxjkh48KsBCrXFpJYR3CStZ0fIdH3AJ+/+jS
XfPNUIfztHYnHvRoTGizQrJ05UmxAMmc5O293qOydLtDQ3gUNMMSGoAcjyGnHj2n
WVwkNF7NPJxosU3iBnz3Y7ddWe3vWq++J4auIbRZmLO74Haj4VVm6NV+pF4XUsNI
etiYBIvNZ0bOqoGuX791JldwQDDqPr752ihOpoTZFmLsjx1Z2i1ybQf+W2oJQN7m
LiMQ/EHTBGWnFYfdMXRjyKbHE/5QwrMZD6zb2K9hph3kAlRaCoZv6iXkvHtkL9en
BDkFc792pTzvJX7xWz+n+g1kiCl6mldhvy7anPVWODKJdDjdfdPMX2opTIZADdnD
apAN97Pn4kj8MN8fQH7PUKj5N6lkoGs8wJtNVUeBb3h+uwnkdLKIueMiJkKTUMU7
dveEx/Yq9P99oH0rXNjjRNKyr0COqfRw0q0o8u2S2WihfU7sYxclcV5TE1SGERVP
jzHLdo1TLzx8wyT+d+y+WkTv4Vg1xggZMzauOkoFnTJHNKdhWWXmxsW2PeEpO6ny
`protect END_PROTECTED
