`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XD/jUAKV4oKbZ1SwRhPyrDR115cEkEXZTFTZGhKcYxIr58vKxlqrQRjLigqs+uOf
3HlsXL66uFjXKfo4oc3CqP1+bpfGWIs9YvCw5nsOpmVXBaA6TLGpqYXmPNzIt5rG
ZIsUurEEytcCNuLnUi03YApX1K3EhbfUuMVVtfZ3LWSbdzf7N8Zky/VJ1E4Khu0M
QRlwTNj62JLPLO1riaEFUenK01mWg0EMlQ7SIxVwalSs/lS9LofF2OZEl8BBShtQ
ydY+JDD75s+2R4a/z8XMy3H2DvKorT1RmH3pqjmTYmEMedfcBAuuG5y7HqFyLk0y
duNGi+Orc6tUriJJ2CuK4jbBbSR7S93cY/XPRINVSJEVZY6A3jH9N9AxW0tLmLRN
9PZOR4IjWNcXWnhWP7+8kba7taE+FcgjP7fRJcZYJ9jU3nRzR+8KlXhthnwt5aHO
9W3Tl6tTZoXD3rsQOd4Zkc3BX1coulrlFnj89xyYFeaw1q6jJT9rR8DFKxwiNa2f
e0lbebknrqoBfjmHrOIJkGV6U+Ya3NkQmMn5xJGijiwjgYUi6EhlB9N0fFTplPMe
t+ybadHYSwEk6o+NbBSXaRZh/1HeyuVmfRb9lXUjrjjUK0hRYVOOGJtO2UkpqoWf
p28KgAND0YWIj674pO4WkB5jYOQhVSKpdJLHCzsxj+5ZhpjSd0vW7Hp9PkR+jCrY
b6DXokKUS9aj2vS6kK2MRBGB0ZLMuj4pNb0vkGk2fvSAAKf5Rw90il47i4Fb4IMF
QCGfFlbR45GainWxAXjzi5DtjVg8CoCkifviEN1PSyOQoVoUCxTfH73YafQ+fE0Q
urZAtCxm3RGBoXINQNn9sIvQkNlTAj0R9c/hBNp/m8f8O+ADe6nPen07RGAwWexG
yj3jyMrForPVs2Q4znVtEpLns4y/GWmjNW2ogCZLjOhHC7lSE7x+1zlkj25pmyE7
j0ljwEjrM4BDrel2ozEwZj58dj5JpaCaGQ2HUu4eW0GG207N7Dw5Jd3f/Kbvodwj
MjGC7cJJxlzbSlVmagvXefmG5Q4KlQG7bZSwqFT1WPD9XHb2ETAO2iEHRYXfAq8S
T6691Ssp58EqEjYyh9n1hL5quuqu1NeaLWA47nJQapNff8RWFNn5wis4UbC7xcNZ
ukFx9McK5al1GESnkABq07+L5nvknLFEIs6nXB78lTYClvxtijhO6Ou5GjRYM2ZE
R5YG7YG/sssKgWly+Qbl5L1GE+nQuCokubvmRImQ2ZI7qqdsGWiVOTv7cKdjKjsx
IQ9Bww5KiP/os56eyd/QqUD8Xn93Ozo9GsewhMjGp1xaw6qiIIxDj+FOti4mmRIR
qvE3ZUnfIcuflyWgCwLg/PnOYBbxSsUVaEDFsSHsNbTByTSoOOPPVkQyCkejF6vj
/OpgGpAX1N7IWTuGZ7C5PGyjQSL12+CC1PbbuRl4al/z3RtNXM3FbcndNqDOMd70
5ebZ6in5cwgFYL2CG2MhFCuu9CFMvHSmKJy/JA5X9uZl3B6CC+5bigWpUmk92Z/v
f6xZyWQQHyjZvGhifnTrWMY78fkejfBjzbY7N9KfiSAijGXPoOpj/SATK4YGry7F
91bbEiXrWsy70YP+BTPxNNl/80mdrQUKBHksDET4jKOTJZ/ieDYa4sgqx235hAOw
Y5KGLvXfZEluVaz0K/vCFYQEUTUtn5fipPzZqgeZx1Cc23zZiYc4fx9m871fREB1
D1nrxsFiCii12B2p/h/mel4L6tuj43E5VZkZq8/TjoNnNudCivPLIV21yN+i1MKn
myIMAHvFnWv1BnKiEhOVa/iRM/o5c/X55uedumm5EbM+ZxPyepqVsU4ChVjyY4fg
gEa2wANtqk3xoYC666mrYL8HQHhRwGV9XW23kbm3pfzSJ+KO7XSJPpTnICa/Zj8c
glTo8y2f6jmk3ZRVnc9h5MvIUCMD0URhLQ4R6gWQOkTJuWAQXNh6R3HgaLsnvpER
1ItdHyHGaY03wKo3tENFPSZ/X0W+qZA0HOQf2acAZq5Y86UMJx9sbthLLDEmen89
x+80wc9EFNwlbkgB8aH/bS5lqt72D7QrGS2vwchD+mR3yDvy5z0GP4dTCIcSsRZp
Q4oqeW3RRgWPxxpWIR0K81JcLHHuK1FY1lYJWfq9t8vMZQriu7bRlYGdt3oU4Zsw
UOFy9zHj3iA0YshOkdb0Iq2cuSsktmDOX+n9JnTxT1vAAc3roVrUBFYhd1Z8G9ZH
ixdAouQhxGYhp+7Ml/e0pQ==
`protect END_PROTECTED
