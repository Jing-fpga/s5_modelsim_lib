`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bawhte8DiGJP03/PU5CSTmuPXl/CNnFde7vOdIOhLn7nSzDaS/1asZQbIuLfunOf
wUOfNfQo0kDOh+UqsFiKLFKH6e+J3f75NT1RPdFgu2ffz6bL/SPNNFYua7I4FIYX
j87O/I5pX1kvF3hK/B7poznbwU+waQtzMOKUlMXWjwUoClOM0fomgS1JPLD+DQ9j
Z+LycdAJhKF1FtV1gIrRQ14zwDiI6zxWNRU1UciZjSZRQwD7z10gPonjO37f5baP
XQlWV46tl5QvZUvfmV3lwicyj7LzLigVCY+YI5KNu17K2z6cZE+tUwpWGu/1l5u5
NpyyaXiTRlUSHRPVjNtAkaM8jviBYSJQgj4rm0//lsc3mUtsFYZYWPEKgmYhXaKd
R+Jn5dNDUe2pjoamLfmvqKi8sP1GWd01XGscCDBDNSv5fWGOdJd1/sgLb25x565l
RwMNY/YwT1xUsbZfCO+R0obLs7yKAiEduBy9w7fmU5D0uYyWRzp6bp8esexKoOoF
4illRIa/Mzm4tBkqR2WeB8JY0CnO8hVR3Gm8lpoBwC5Z2c/QM8dNtlteqX6Z2CqJ
jakcT/bvWBBHF9eSmZkbhzDNe6Pkaq0X6G58LUWFdncgQvp/wzoZ5Foth1F2W/C1
/6k24bQkqIzkGSKqxRyU4VjIubW8W84du6uGE4W7fY/vUIKAo2jXquwt9uJhU6/n
glB16w6H16AKvpFVTtlCMJM9E7VGfiaMYRTn7Fi954vSVqCPy5s2IRPOE15Vvblv
f0GI8mxDZ8ZjMv6wKVkiPYb3pLhPm9bzAqoToxtZfWvu2W9/TIhEwGf+5H+IQpKo
E0dG2DeOy0xuECPOQKnoUgdnrpLB+7dldSpzgDlEQZ3/5oFxfxTSJcPCUhZjoQwA
D5DT2JOlazrpB0FC9AmbfcmHVbzv+0YiMKYW6gXx2APV1ZcGecmYQuv11Pagq9NH
BnL5h5teDHGCh/ZRV2kKnPuuRx1wdYpHy/EX25IbsXbFMBq1grW/0OB0havQJbYu
ZIYEpZvN8ztTOAHhCrCklZJjxIr+tRcv9XNtR3vSLb5Cmx79VsBqs4mgkSgpLfp3
hu9Xw6dER5lten98q4GUkT8QH8pevf5VnWaRkUnmkpLI+5XnZdW8vPfrYN+EioDb
vbGfox1tokC8DFRECfWkbxQjeGHMAMlGr5x4fbVIedh1JyKMHe+pHmUcJ2uG5TDt
2oLhD3h4zvM/TAhAPBZE/hqys49oTu+3gRWYS6K6f/hRVlWV1DT8FwMeKKMX18+x
I5VA7XNoMl+52ix7lz9KaK7Wpo/JjNUFJ8njuf+coVbCXSsfjCbw2Icbb4RTNp40
xisMs2TBDYQtfWNlOgywgT7xFkiL+hEpzE5wFdz8kN7gOCKxF3rUnn1e16mW1tfF
x64TX5gQ0IVwNwbloJeZmnFu9eJ8Y9De9xs2ZuqjIm3j5v2QJl23cdPviw1WGw/4
jTehgThWrm0feUwGauNL3xKlDrmV3VkUYZpmJTGxcTut4FAeIP3mfBUuWt37ihHK
3Q55KA6FT8P4zeyQ6p0UeMvgbx9fOhqWmAZRTFK8iTNM2wQOK1PEZLofS2a2ANBI
NdPD6qYl4IvpUEghR02pvWU5khMLAAdasI9z6P5GmL/1iLNvogWUtlZFt2nJEi7e
ERA14K2wulXxz+rf+qPLWVNhvgbphdJektB2vgVe0aCIBnlFJurAtArthCX1UJtU
B+Wnho4/nYDvW82sM7cm4NOTMq99vdzU0q3ch6zaNkvFhEZ9xCoTHYtN6747fqwv
i6cnpduN/UCMRWsH00Qsr63uIKrDK17T7JY31Yf49QsbIqp2EkPlPATo6QvGFapV
xUP1RKYg1gbHI5K8J0RjwMOqUD4X0DHeEWFV3xrRiDAyDVFEzAkk78KwBAcO3W7A
bzmWJ73cil12OUzTEeRPwIFY4gndijyvz8ibOl4eXZKiN5vrStmKiiKjtN5oPF+S
3t3xmWNHPMA/xiVl603dg21dQo13D3sD6xpJnoLEZoef9IjPaOwvQChg9FYY6IqB
4/5pp8rtLn/NfFG+PowPxbiGRQlQqHdJr51lPtlwJH7rV6fGEyvnzfU2MwfitPV8
xR25Ibn2kccgMvIrmVPIVT9/Oskch1nQxCze+AZ8seYfk0VnjA7ui5Xzj5A8M6tR
T1UHB6KLwaSeJBZq9aKlkV+BG+DXI0wn/wil7fF69pUHdyMmCBK0ZVZZ4IEeXHwk
B9MJxKv8nk78fHvmrqCHSxBG7/jz6QHtk7s3o/k0vcRb+kw9Mq6KfY+zggcx1Zbx
9MCQXBdCd1QlV0nx8Yjj+jVgN9/EboK2uxHQg0Ip4afhk0pjASkSpkyGj6jfX/kx
M2Gk8L6xeMZy3U3zI2SNJM8RkedFq0SYVvD9LcS2XegLJ9hArURnEhEpZvZVw0hE
L4BzjhPD7vzEhA4IRvfCYgQagmSBxVt0mOM0jywAbC16bCPJCBFzVCEXMbcHNIeX
r66bbiFuzbLhui7vT9GAnhtQ3P0AkU+7c8A55QJRhJxkRY0/+7C0Oq7LZxHojg73
Rj92v0PNb3I6ZPpnkm6VG5cTi5+y61vZW7Z1SxzM5mIbLeA5Qfjkg1cT1zxRiIij
0R2QsKifdR729CT+NInyBu9OaIMcnIWDLc90X7XkNakWhKbPjVnePzuqrYpjQNp6
1QVoC8kMW1X20syLYvRWxVdz5nRluCcxEEmtNv26woUF6c2qZa41FA8Atwf/Q3ug
HrAkpmqDArkXvYdtercvBNR7vZ2IfoLLAiUnD27sVQqRteVukLLdo146utGCfyTN
7uq4wVOYRPXKZS/0vnHzjXMnpKBNibKXDSlD6qudzNw9jqM9/+zeulyc5G4OyZNe
DYlLi1wLkD2rerojSBMnATGTfV6H+Izbdx7cFuwBYbclchFPN9ojmUkkg/SuVhFH
PYwn9HdTWkBI8Ifn8n0xgyX351zQbc8YWNaTVM3G/Be7OUFzChKjoKuCNil89Gu7
lbxAZQfJ4h3xkZVZaU0eU6/BLD9a6Gvac+BT+yi/ievsXHfzBZGfLEu5rYoub4si
jcB0PwuZQLDiMNC7tUnF0FJtwMshwmVIKYuxgF6001IZDlZj4Hxm3alkRYfgb60I
fEkiCx1XnbUk17MDaRlIwtcqZcFZjpGZlrvjzrRylqQfT/Vo5CngrmFFsDDEDkJk
fs010VaGXzoOhNj4gApMMap7CTg7p4TaQKBNhkhF34Pslc/o9lfB1j24nvNw+djT
qEiKlBoIjFbZZysJf7XFoJexVDppHeFypXWinMSBnoFWA8m7y43vHjLqfGXa7hwV
x0t3JUq09z3AZCMmbCd87yGUneF/4swEzIJALtdE6vkd+E01N6eZZyZVumLMdx94
GXZBrMUGjENOfvD6RlgPfxUdlZH/oiE76U19YvHMGfaXKoAgu7qAP6zkftE0gsZG
Kw5HErfqCM7GtRe/AfE+6JT8kD4CL+T9j/BPCDAeiEpLKJ/RTjtJulw34lKRrdiZ
1NzHyCO4NE2G46B65kJca2ev5y2dscPFZfOGhtcmSALHKiG+UXo1pJ93Yk2oZqu7
QkKIZF1B5YN1QxfV34O3I3AerXlODmmtoENRfpLYX36lG+fldKBZ6Vd91zR2tDZO
hWYPV7Pz/c+CH+BOMMzt4ZuVaULwP91Mp9rrLmrGoeiAIqnPua2kc9owNUstTscx
FQ0mOtJsf/RFRTQZsLurzv6f2nFYb1xRHOq+5cc80iR3e9MSt6m5V3s2bY++NXvH
3tNSOmi0Tuis5q9qu/8m+MW6LUXcM08MJt25m6KU1D+Dq9aaj4SGeO25TNp/b8l0
v6Wm9YC1Fyg6hQIluRok05KKLtCfXOXdDs2Qt14O286rE0sx0FjWH8Vh2jkZDv3x
HdoT6/g5TolYxfxz78k/dBhRP+TmWTKLMeDLYNv5NZUyTFZzm11cZhSLePaHzrFr
TNgXQ5/2llCWxld0FQTTlIY3SuQAix/S60exoqZfhFRQLPQ3lD71x83fDAlvAHn9
bbmOhEo/AOFXjE54md4xP7iyOIw+YQ/B5r1ugNhtdEJTrQoptGvZbVv6eX1GKfzL
xWuXC9vGRSdN2fv0Vd6/vIE3rUNbKIs1t96/3423/5iSj7+gxH+CREKBZjS16xLw
s7jXMB8vJ066IuV7o5mSD2Wvr7C8mkhY+PgLmU5Oj2YLEBvo6MqSrf/ySMKCHX7O
8LVvlNXZf/obbt7e4H4z6FPbvegbnVGAtV6nW/UWW/zugMpwfYY3nT8XkmOGnnke
6BVJt3GeQJ5RuEOAjbjMx8QWoFa1fM45Gju7PSvQd4e7LWEaoXUw5KSGIBtyWB0v
hTWjAdvx3/NGg7VnUhGkWcnC4X2txlnWO1pCftOrel+GqvR06lkMssSkN4RsvW2s
8TG1rVn9AblCjehgf/pENKTtwm03JSV82RsZLtX637as8mJhAryh5xGXrEGll3GC
XVBtL4GI8ZDyC8Ou0efimQYeNDd7Mc+uuhK5lBpu5qmJ7mRrd1BrEv3ChFIT6813
OnjuTPPnWFbyI2KE2Wb4IDP/ld4w8TrjxftbMFp7mAfbCutA8E/aIpNfML0cthwU
c4beRlJAXDAnq/fI7r6xj0WlBebJJTSnS4qy7sHZp2+9y1K9B/tTYqLbjTQQFesV
wFH36rWJYBdEmr76dWvRnhZyuXdp8J1OpY8hGwD6iwV8CUfSgGZOf9TbLz2AhcCN
99V3gqYe3IYsmJcxX6ku4fPgXpAXVydBkqAXcwoEHPe1GjqvSRniOe6XTr0CV/oF
WcQthU5rY8qW4/rVW61q7O5uocmpFFiwqLCyurMf1XxHB2YuvKIpq/pigeTFUznv
zvIE7ioG20HrpMapDt9wnEoVeGn31B2/DsajticgVvCyGwA0m0KCcndvglduB6Eb
FOU3uGp1L7cTdEqFxiUYDe5RZlF07/adiTdGvxH80HPIkuJdYwWLwDceJ4z1AAOW
h6FvRco83k+hiMP4DFzFDSYAckF6g830PUDf7s0fJxOXgAi+ZYej/5yCBvCetVm9
26OUHMrqqRwwDryK9Ekg3C+2qtdGkO4rmw25SM1Y+eeyeJy3VsLTCG+YEnlJYkiO
4uq/h2kFKbk74d9xB0oMlCrwi7fY97UI+YN3JUYVOCjhDZa1UxGaTnPV2boKVo+u
XRrxU+eAOBR3hvivhG4ZtnT7qcBw0uvyIJebJ8xdGkamGwmBChJKaDVCvde1hRR8
GSC+RkcTJHr7QoZyYz/57LXTH2pZNb0vvxS9A9F6kHdLvAZhdYq5VJAgz0kbv8VT
sMIkA4hffMzpfe2Yl7DLkCx2a3zdAjLZXR4h7SdNuAUW6gXXxPtAMZNqL47clK8O
y4sZMyKIkNzIIBJr8czzA72Z8b3IMizgdKVO+4WQwjf0SeAGgWXfLjSXHJtj3BRG
azCTOPHDtVjh2duw1iXCmzZRLhbcIYNQzFi+tgIqmElWfjch0QOe8Ilt5IvZ11tW
IsTk+SD9cVjFRL2VOxTuFMrvOCftuNAGLSqpLFOtBvP16S1LewUNf6/7ehA7bLkj
tQ7UNERGoWyiY/yaprjzLW2HG1bRqeUnti4Y+UP9vfOHsMqCCR+cGj+ADtyVhbSN
cj607azp9RUsGS0N7NDlRn0sx5OUOMlVqSQFdJQH+ylE5MT5b6dAWLdNE2oNbrRa
mSD367o3Jdl4059m2UriNdaAOOJ7i2vLIn0acZSX6NXpXfEdeyPBHynxf/sKwPJG
QJfQAwvjqztgzz/p0wrDujDIPqaxNwaWe++mD3Q7z5S2ct5iffuHLHBObhiOxAq0
s8Yd/gPF9mN/Wpsf/MNskfMILUaye38+cgB+jOoxYqfyXfCbTtvP4Z3KptW7H0uP
/w2CAsw1N/KVxHnfu1Tqd9RO8gZF78sveYkganEZDd8=
`protect END_PROTECTED
