`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cBcF72Qz7bpCEOmlbt2bxvjFVjePur/51EkGbZhXcNfo9vOsRNXLL67hoNJUv0NS
wKoDhcCqRTx11gsvdvk1hTquxZsAPaDWdjjjNW5i6tAs8fVyirLNTimoOLfRYkGr
iTMr77ZwYYri2LWjqnzpZVRX1+3g8RaS6Ytox4206MD5DAhpxuXSAP/PtObKsgyN
xJ6tNOR+oTxR7gXMK2gwjOfafFV2anzVG29T8v1ahokTVA6ZYh4NjJLrYLHJuAAU
u/AXqTji0U4eYTHKlo6siChSVVl8MbbauOpjceVXyCZh2oR/yFce1Jsjgd5fvwhc
jJcHN7WOv8hT9cjtNTdeNHJGm5X+bEeBIOZ9fii4G8F2dfm5APQudd1kktls9oA8
30PtLmS0Mce5MuWJaqqn9WxNNdcOJrrgZJ5e82nkdDaVzqe4HEk0nI5NY341fleK
Ul3/pAfOePFRI/IX6w/nmjrb9nlLNTqvim9BveKhScUla0bViS01hVCyZY4xIDtr
boPyFiiZs0eSTOCc13rNQ3PIHWG7LzguJuSNSMZVkJUczFVHsCHtwFREDdaMFSwv
ObtIcpz7fyYIlXX04n1yBGmV/8PVZi47cFv2nzAqBnFoodfa8HCJgMN3ExwS+9U5
a+1vFzPqvdrAq7bpjfTdBvIuAsr+KnvJZgSKVgKbkvuwNlqE2Yg84unYE+MNz5l/
V1NX0TJ3gIWScSTk4c3HHrfTC5fQ9UhEHDSHKKTF/kEFq6eGEjCiA1+7/x62r8Tw
EQa7t/c+MhYLTmodYgJ5/o5vloeL37F0IygfRTTWkFK7a2IEXzKD02+78+MhTIkv
AyYl5RZelSXsmXN6lWqP/FlI7ZmAFkCf7VtJT+sp5hFJWJ5SwpVJJyDYlXHrmOxh
wmeS40bvdQMRi8dIyCJ9oHeLB7DTLs1Bfj1PDusC5g4K0MDlaMx06DqZEz62l93O
zjB1/EgJxLcvexpEswMwklo+I5Ze/0aVvE3vuQZQeS+CAH8M3M2H1jLNi4VzwztJ
edhcKbdWlPoAh+6egKbyohlob29a7BAzkwnyHW38O/XZWBhMTCSse/0P5KQlM6AL
eQ2Qd3gm22DrbQPxtTg7/jOVX3RARjqPMdHrWmbpaVl4DKgDCKh3D96sxpEgwcn0
zzKxS2G154gQfzL/F+hcn0GVUtGLytqC/a40zcksiAi2FBNAhTe68q4/4907dRVC
OUF8/F4j7uG38ak10kPRQcviO0qkEsrih9X17QJE9wDf/JGKBV97eBcSvWEIDtOb
7ubILgvxNGgwiHiNTFPxtNCPVujUAcUKa0dvt47I9+LpDa3FeNGGmbhGmqJgIZV2
wIk11aXu9I5zBcnDIsmGxP/Jyr6/tpQGCJD6r3rgv+Tm7bQPKop0PZOgrpb4+KWc
EPRDYxuo2h0nSTmhDFizFdNNcKmsDrZ3O0E6WNDR+zeCd6sOUo0xScPINvRiEUmS
/tGhI4hAnRlCCJzv4zzzAbPTMrbbLFH1mdwf8+lm00DB0dyONnXOzQX2iN6O+rKa
Ytmlv3YXK+6zQBZhZ7AiITN605yitcTkp5Q7p6RDaxDplstTvRlm2j3fkqSsznW6
HyYTJb47enWTRzbEsxXOp5nsKrMIo409dwxYKlM2bokqcYymJaxesTR9b7fgrFJM
4o0rzTncFxtY7G4CBNECW7hhh8nbCYAeVqKxWjKyIglL9H5cJWKmAnA1KjLGtXTP
ajtvz41ZCeOZ1B/k79wS7brT8TZno4A8Ts38ZlVtpZXAPZdk7rTU/TaaN9JbgQTh
gyW1saHFjv6+ekntD+dU/ynsRkD+SNbiMeQa+nL6IfWPQ6SWFVZ4tC08xdmAD/j5
XQS8cv3S8/4W5oKb71iH5q9ymGAv7OkuNkoXLj8x6JPVLW/eema5bafqvIUKDMAT
`protect END_PROTECTED
