`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zExdvv8wUPWsbprE771t2I+Ewa1qxCiRsz3rgcajnb9mlI9p/RAD+3kZP5brvh8q
BVV6HAETyiGcstMgVIZbQMgsfnTUWI9dshIQXUDGgZUlLjr6hZS+RxsTp5stMgKP
fPIr9g+LlPEjL6T1fsSAIrMNPvz7P6rkVMei8KIxctXmei4u8TSeWOWpMD9NmJaO
9qht9u6kqYmJJ5lGKoHxwXbx79zGpI0YatLODCsijw+1Hr+HMVc39KtDsrqwLLWw
DiUrwsnrrbjS98+JE8myBRp9X0StHCttJYW2Q1unz3KTzALJ/68GdgYlNE2weh9I
XWCcVm+V7+8nAbD8UYGFMz1/+1cXppUdQhwRY5Dst7GicDy2UInDkZHWSFOEDxtm
D57xAveqvs6/4fnDuws5SgecUmez4CccW3sgGKbgTaOgbWkO8miE3nAhB0xMne4O
gZ6fDPfslAIHDef3boKLILEEPnUaHShnTNop9hmGFTCHuRpsTRVcaBzqTb2r0/lt
9/Ek3KIJdq+WidcA4l25esR4+egT3brQj3zDuZoUyZ974Ov4VYuJEcU3qm3Zome7
hLhdb8ye6u0xZ5mlJmJVBMCcciQtPizeYQjKBSYkXXd5pf6yXXjdvHN5BSrVwdrq
hKG6KwKyohSPP1vye8tEU5F8vKt4ux3C+51tuY75RiSorv3a60o3J/u+cxg8x4Hq
71dIT8VF1b/jlk+fphKY4eKCYEGCCpdUfCF9i0q3D7EYXCTU8rYB++T0ymKphnUF
5pUoC5uXbB+U8oCncC6+lRqZWK5E+tK9nd9ClrNB8Ll3H2t/5zhzz5IoGyrhBXPO
WIFRVt5Inm/y7gxUfGF8SCJJyhAxfcUFC7EqZ78z4ht9nBraotx9tFMvKpeNMwu1
pBp7N4ONbC+yA+A12/YzC2067k8hlCV45WBaJdg2yGfQInDfYU4Dkih545O5ORZy
vO/bbsT/Nf2LdOPaH2r2S0Wus03Vj7Ioa+PdzIcsCcR4pdH/Y4RHRz7AGOdbpXw3
cy0hxKgGG7XftIbEnOZPqrs8CaGL1aifOiKPhWrwcy75KjOv86oYxeLV1hiOFulK
qkT8wIQD5xSoxQXsHWCH2X7mcc+kQwHejtTdrAvmNmJNzd5e3W+YV8SHVPP9ET/R
zZpbf5DAm7KZqOTXMkxbAFCvIyluT19dhz+WYx2NWOUrmeh6pExLnvNtXfrWIWfD
FrVDDlYI5UD0hJggFVzYAwIlqyT4LK23V8lfilwWjLYYffP8fynANJNZkwM9ouzG
Zac6/AFTXnDuTC6RwMLx2HnJFVB174qgJNPtjZGPXbuD40+x9ByBjiAcCWDsLTd+
PVfcjRtDWRBdqTc+APyZqxW7yj+A1Js2URim4fQzsfcddPeaPVRw283xkh3nfCwe
Czb12P8UTfGqhBnlqu+tcpzhEpw+iVXhy+CO2u5oj6u7dTRRylxPhb7KPRIyVUSD
vqjBUcbKcVkpM+F9Na/99ihMeBZO7qKYbRAi/19sJbdGxYfneGZeHpfKZWpUgW/E
k37R7Uy1WCCFeoApHeE8ocxvitK9JDfwht5+LgJabgGlw16YqUKQHlKWodnP76Gt
BbbXvTsF2fYkZw+bxHyj2OMwzsR4dYODil7HUmBosIoIja+bUq4cOPJHAL8wCmmU
QAkGcpxVg0YaS6Knw1v61HnsUqYU7RPOmJmdwA9MzJUkakBQVic/ZOfRJcD8ApiY
PuyEzc9HkUiE7Kzxvi+5mRIOn2ciURWq3Zw85ru/k41pxU/bwyEiFSWKLItGApRf
7s5Zp+Zc8oYdURIiI9j4n6bL+US0/XjxjZBsD0D2fOA0sNLC6bL7Lckdk9iSwvGM
q+cv3P9WuFtWtlTzKRwnK5llMH/cyO2eqCStXWOhYq4PjPj3ItH2er5u62ArT48c
UZMe9Jkbene7VeO6MVoT8Oa1IsQy9dMh3uwSDZbk/r0Yxt2Ocvo2ovqQEEaalFxn
ogTNZToheCZJr80J0ep5ZaNS8HKIzmx5FPKVpbZfq2Pr53VPPFg1eRKMH57g8UzW
4vr+kvQOk0JMvru0K5Umgw8JB0K5ytr6+8msb2RBh0LsVhRTh3K+t+3epvS39Ysk
MEsxOilP0pV+Fjm4Iz4/x1vOW5X7zpJS2cewLaeaX0pPNPQZSZ7hPjt4A2OiCH6z
HemTNuoteW1Wj7dOYj6mlzQfAqmTZwRo26ZvGMj6GrG1cA8tKEsPw7syZDM1pUeu
Od9B2vKqfXKaHBjWF6O/OY6aP802+T8drHtlmNuBptxfXtahvHZftfgPtpn3uqbe
FTE9rDC6V9t0YEfLBkSgDPNOSU7RY8knARBLpr/Pw7X/bKaXJwF605Y6HIH8Z7Zk
xksuOSVE4dU4s5N/9sUfcSThrcHByPer5444fCx9Ws5J2Y6VIt7bAKV9I7KyyXA4
hCGL8Ax5IAGkYIpbWzbKgU8ccAnebHV8NZ2IPEtcTHpwknpzW0LV+ysmUYEmxdAb
1ZZ6i/XOp7jVj8kApRwWDzrj9fZ2FhlNG8MaRucODj32sWngP4eanuYN0WdXHNP4
HMsIGvS6qXRXhdTIYvQgNN1QhJeNUlPnz6zxgQ4eJL8RDlguvJsyPhwX2CdAuSCG
I9QjZ4+z9ISnreH88vmSny2FQ1tO/s4SnvAOFP2NC3tS6rxoFW/6AWrS7xqHJUfy
bnH01MfO274u1096hOn7Af8tO14rRuEVeNpVEob2qMXbORcRHNSqwpSKr6iaYzCu
CZhutpFEGcbQZ/GIXpR6+A9KFrj4OrhkaM/hONoLufzwERZIR08mHhG0AP/BcHMm
NcIMHM0aQ2Z+oTkhWFfOR1J2j1DCgZ8s5VXskle6h+LJ60SITBQt7o6lfhmdtrtr
5TikWYLxtXuVajLeXoOf6wWjwU+32t109UmcCgXHKEmrmL1CkgU2Q9xLIeskMWdV
4fLTzQ5YvU0z+4IzN82CzloGxe6bbkn1p0tGLWY759qf37/lz5e7UeXMgA8g7C/8
5udenl31mzBMbXu4McHp3qe8gawmZqXiZo00Df2kqdP4F9yXZ51mF+TyaTSSvsmk
TUhreSWLUKg7rosu4AVDPWLCHY0ZvKK4dc625fvbowebZKpGsbBnIzEfna8DEgYK
Z0coterKmDKxp+BbbYnxiWtwUqcqQ7g/bdnYpBTIRB4LdzECXjGIhgCE5WLDZIST
SIb3vgVCo29N+8cq4vNjpe6TecnTn4+pTlmFhehMjCsKC2iNuiSuOB9omSZawRZM
99jZ4yqCsaixVv1Llen5Gk48AUNkvlFvUATGmLZJ/TNs1Jtc/jmn2lxuQGliJK+Z
cz6bg68keCHeiMcShlRiSr/VQwuMapIubwSiKPMqKPWiaIvweZ2sM3qVMvtGzfQb
jjAzBa25QFIQqklJesKHWGqwfpGbfabBXQJRmFzc7zpsVaLSDIsmHqT0MIs39lbC
BmkzBEIpRcinoioK00AhjAm6qBabgl/zmOxhYe73/duWHpPCz2KtUSsWE1xq+veP
59hfjogWMi25thiJShQV33Oi3RnocmORt6KtR/UzpNpOCGIme40qyoWqgzu5NcFH
1+Rr5unqgYFcoGMj2aS8bKix4FyfK+1Fb59B0qIHtQL2wZhThRzo8k7b7zdnjFZw
+4QqEpkoTB81mauIEUfaYHNYHP9J8/wSjHbwmr8FBwrE9ZHxUIr/688hycapL7Sl
AFKfwkReZyEJAX/0SxM8xcaNhb0bdAsMiHqBiDgOLPH0psg1uK4FxIgS3v9E7mEM
7CNWzBz0xGwE1T638m81boI8XaxgsCmPMXmR+pmu0nyAoJhlOj0i+t78o7pZCqoH
IzXzg3z2jQHvPLKBaGrw+SnwDGujMShi9fvTZAYO7pTzjXmMZPxu8+8F7NYUmg1Q
JgG33t2O6dEk+fgHZQu4/P2vBhuN0+FCq/q6LnIh+SKtesoBqw7Yys7JXPbQDjdp
4y/7vHSv5Lgli5Iz6Rs61IOW767sMXKec9Dwr7YSAA3w/v67xhL9lVGOykVm37lk
IBzOkIDrS6HQ2in0rWYi5sDxX0CbScd+MwyM7BOwroMcIsSULq5vfs7n/i4F9ZrC
m/rP66iC/aqjKRGN11bfbdXN181ORAnuEqOqPn0sQpwz+cfIq8IB52Jj1M8V5kdc
6dOnMjuuutI+SeBU/2TFGRBUDvs3lx89MakE1bHcmlmz75iJ42ayqktYSdVeG6nt
XUcFxSFAtSFb3g1y8ZYxn03b53aneMK39pWtcYa2l9Wpbqv7G4G5QhWWnLbp1uyK
lsPgkC6FBMLd57gfmXvf6TwME7Lvu4dodnxZliIlgx9tlbL0jTZbiOViLIeEzoKu
BH9qVKmFuwHI2koR4W+QdobolJpBg9O2hImT83l9Zoc=
`protect END_PROTECTED
