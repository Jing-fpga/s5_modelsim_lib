`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SSo6c5twKdGYoiAcxcrQTrfTE+v1bKGZYn058ePHNoxA0u5QLLtJzSxPfLB9fNoC
HLilCpVUuEIEcfCLk0OtEnGw2+zXYuy4NRDQezyW1tIQP5XIXMqRYLZypxni0Lct
G7GFTjeTMZvTgd6O1FARMuNaLL0YXXQTuxtmt0jOgKX5cXzYgBTSu0z4AZoE2jn8
acpVVvoB3P39L5zOuPOCLEMRHaTchbCQcpcA8S3boTuT3XmU4aPa47bRUEwxjWPv
VcvWTZa5Z2OAxSqyuHO7kD8BCBM1xrWpCwRNSLcYUq3sbNW8lLaOx4Gmo1g7LSiK
u6fkXnFs2qM6eSPSiP9BUq8iBJ9vDOnH9tAq2WyB4kYZiSdSpA9Ntgl4s+nm3GU2
q4AUSc9FkyTpPMgGb4W4heetBnzC3Gl2Dp7Ey9eA7eKHfw3N8ms2Bm5rp8dc49wE
cl8uv/69/zvGk0gUxtglR3debs9wJhxEDBq3Cgg71BgWJ9RQT/JBfSTbLszhwbds
Hxa90jIgDVNrglYQ08rwOWl7Sqj9CAd+HLpnoD80qvalanOj0oFtPXZ9uAGhoys/
YjFp+OsoH/wbibQ7Zxnh4tQDVni0+qBPADh0O4Xgt8se0zn/OXyGyRqK4/4pfWcx
4cTq74GlsLzB2cwVks0mg+7ojiDI960ztuauYt5MLa3kjkkoAI3Kd1vobckcDTPz
dN4mqUyYcJ2f5OLRHmEGyyOC/ovyrlpft3pF/olfsH0OhaNNf44IFAb/wqiAGCAf
ggnV3oqXKs2eHkDxxxkulhCsYleIaeBeB7INDpJqAfLMJ55HNzVysiedsskJ2Iae
c14txgC5B+Y1Y8d5UBhpTuZj8Gli0zgpk/qvtnImgqYIh8b+QS2yQTexciLrmmNM
VN+//mePyjiJihREso9Pon96a81bgePsQPae47TGHVuLGZ3GHfp7HvRR6HS141NN
ZrCwaNjJnOaTlzt7rNcSEI1/rZCkThfvLhEmea+6y+GpeFeW+Lc7c5NAjE3dJfSF
0jdyDCgFArmK7OrLZlBJcOW3Pv6QD9Bbq9QFCI0loAe6b5FBlthngfC0uO6ddxg1
kIoPx0brOQ5KL27iwxKAK8dpqWtkFjR0lWA/9bmW+MOi+HLHhsrd71/IB5T4zXpi
yIV1dpzVxLiY2mDwtW+HO7rvcYqfgtaFFg3osMFpeH8v4RdNx4Db/iUwGCLD8SEE
ljh7jlsL/y1G1U1gj988q3GcuWYPs7D6XmKj4VMXVkmVOXaT1aqxT5xSaIE7M1PM
7gnszhCgd7K4uKQ5mPIn/Z2mlBlnGb6Im+Ioo16rcQV1GXr76KIAPU8i5PItsIsT
Eo1AJoBxK3s/jzXJ/53QTPmzlZNxNJsC6YtXf1OkN/XvTr+UaFBGUHRo3n1BD4xA
ZO4cijh+QCN28Mh8UMzPXrLch20tURf9pPPlbPyxKFFBMYuGZ3SKAx4L5LqGKhqS
xdDAk/n7qwj9Ju4Onu9lUjmeVXTOmoi+w0O9UKQMH72zTTW5GTWPO75CXi3CgueY
3GS/wq9IjUSQ4FeUNG08SYoXNbysV/cAPAS4FImeKMSl4O+k0Go1T+gkf9I2L3kl
zzjLzJmOFf8sDa7hFzAp3l72oifvSiIG97iK3EFTdLVGcIfac22EQy+5LuY3uiMI
9WPkHb8zSuhnCekCLgtIzohC5+d/NVkLNe+MVFFkz8UQSz5OXQj20bpLEoxSwx2g
wuFYNKl6g9pRMVEAp8egLSNTMqRhIApMwumKP++pzwu+2iRNOoDi+iWnG6EzjNwu
jyQScg3Re3rXhighkO9jZOBNSPFpZX9+nR+Kg2phtDBUNnIVzEpctLEb0ZAgi/+Z
Yyouen2c2cPrRMSczUU215NgDC6duZWC3pxXP0GN6FgkD9yAtr+jmihfEvBUZHbW
EOXvGGKRIjYay6taiOsekxBmV/KTTcAMxjOQ0vkuCTzDpXda6SdavCYBtLipP9FY
fLri9aOw0kRpjI6FNt6atTK6ZTrpOiyy7oNHjTcfGyHnaZ3hPuTbh1mU0QUbp1WY
Hn8jJe9KczcygqvhispDIlA/c6WYdHArVDbV+Pq/LvmvSKPs0pPvJb7oG/wknUdJ
8n5RMR2EIPNSKBvr0Mb9NpR2Kx0vvKJN2q8F3k1Ky86rPxKxtNLKura3gPDQbVia
iW3TU2IcvQnxBTQ9usC1Xv4upwUQAa1IO78eC0hoR9tZj4BZbj8tKqx+bo+FUsDo
iGB8nBGHvpQEFVWOKvWaTsPsMGBIgLXDUdqrfUrkg7QDqWpzNWDPB6qO3bkOSfMd
sSu36jzCAJZ/Ua1+RSlTYHsmXAhlPiXzMC3nKu0L3Cn6oouubG2FGpseW/NZw05S
OL5W2VUaAORNi1M8N15fqvlbKzwU5mGz4wmYrO5NL4teLXm7ZFF92QKr5t2VcPOX
jL5DahaN0o1bJ+kcc2HbiLviBM5fBjiZ4Uglef7hD6r8g03XAFK9RVSoP2mBYtRO
PLdVUXVpJFzKUHj7nYRgtY5GF/A+z6Reu4hUdfQI3+QNWX8e+QWj4q40o6OttQY9
ULNRJOlao04P/vNucoUFcczfr/OkMrvTyL5kKsuk6HVmsC/RdmVCUbcLXK79mU6p
QpgpiVgChJWRHVTaPBBMcPByzPGpt6wEMCiQS/MlO+30yiYS0JVS9kXSr61/6vNz
BTzNeHze0o77m1fVnpE+l72RGfjOqePpdSalDlDR0RdepcICdA+nk+DnOI38Xhu/
BRpksobDkVvD1rIi47JJ0Ghcm6a+VbuWSrLNc7INRLnjuySSGpDWxFToJX3oK9kO
Fjcw247pct/0otvdzG11aXhpj4pummYlXBqcVIzTpvaOTkHfjvhSEWSWUs7V2Id6
3wbhPks5SzfPSkk49Rh3Gro6Hvp4/VPV+FXpsbYzwAFJ8ejl1GXAUz/xXJ/+NqVE
fOI0kLvOpYQe9JVHKBUQA+Ab0TjHF/KXBE67rH7pN/sjezk19z8ojpGkAbsB2JIv
4/fT8WgHxDnLq7dnu3E7TwEW1LQ76ClS93VF1vxeKL7bYc6Qd1zzPbIg6CEYRkg7
WppgWnH17ooYq/kr/GEdS2pg/F6uXKjrcEF20n6zZ5LUmKwDUUo1H29C4iqb6OJh
eCbvtr7qOd+AvXIjMBeY/HDkn19Nnn5h2yerF09qKqZ6SrlsNFQ2YNWlfLBSX0Zz
e3cKf6J5kFpuijcCZGWnS37hAQRUaQUatAkAeghHuWI76IzO1hKtzYO03WOAxAlg
CEIvTS0zs75z3bGAwOTcAD5lv618fiAp7tt40yZl7FspzmTnPzLinREHfve0myXb
B1Go99q5eL3rPRZAwN2eopwfMh5KJ80dZZFKUHLboZ9fLEHz0ygfe21ng8vMftaP
EoaulxgykYvxMkLhqstZkLv22j3SsL/QPOORc7BA3En6Q59qjII0Tc1hZRYuNHTF
ZAI7U/4zEnDgtZUQM9ZNstBGGB98ZDkIfZYkgV35AUkF5rxzp4VgWtp4BTVwSgBx
wBFQqj2zFaOjwYd/PH6yFFZHwtvhIhMtIU8QS8/aB8hVfWxqqN1CREP+xrKWyr6x
rxGT2JMw3V8Ux8jSb5UmkwxYZrk6Hrm00I3DEawTvu1Viv/eHCHjMCYPefpyhxRx
1tjwfeXv3RxATJjpafxYM5QFLVBczJhqN9nSx1NYTUA5iLyI4YjABg1gUfso3r4d
xpfsoxtluzPOiOXTSNgfeNQ+y14jSzJVOKhXtydH2AOZS10KzAPBQVlqH515DY3U
H8+p3b0us8sl+YpP3ZMbOgYs+aXKUjylSkWIJvmzSqY0xjH9vU3F1MWlofkl54EI
Brcr06fTmTAj3BzPmGGH/AYy4JCM2jkB/uXuYcR/gzO5Jq5t5xn8Q9CG4DJFdxDp
zZfxv4oi4NR4Aj74I25+fNnzAgovv2c3lHmCiKdD6L9lJtCJRCpSSxk8+o2/6v9m
C1kQ9oRjMpDKV3JYZUBj1G18elYHdKkxYql4uF5fvYCMZkbS7jnSVJiSqWoK0TOq
nYAsrZQk+gqjCmgwK92IAqpZVQk9SD9QrUVYCKsB4nm2USoywlCCyyUEgz6uGJhA
vPIGed6wUXA2Lsjeb01AJ4AcgZj6+SGgTDuuZXCUvRJnQp7l6v3NkgFk9iEqUTuO
OQzEhZj5/0rNzqTf8lHiy7FU7o5QDcr4WdmYa5Qhva1O/PtP7CHm91AGa9/jLpbq
CLiRNUWmUNq8nHBV+oXaesVQujGE06OyAKBsUU9d8jeakWsYADYMm6clZKZQ3wgo
KaYBw8SZl25XMR5i26e8CSy+82SC/hOreBv0Rkkbsa8emsJqRMEU/o+X1Jh2SuNA
Y8mE+2B3pPJVMa5dDdRp/2kWSS2Es7NACqq1tti11D+aYe8z4JFixdjz8hmyFLsv
FVTlHvpX3iHiFzraURJyhARCB620BKa+sRnHOapO68GbJA8CYSMVbUBTvh6du/bw
54cLiCnyrj/L8jHILgvuCMmXsDWSdDKoSDZ3+PiXkV1AZM+DyzHWN0IDRN423ZFG
lL0GS/PWQTVW5bB7yfg8AUAj5RpO9ROvvBzndkoZRI/lswzKvSCk5Xi2T8+p8Gt8
LsAbuuA3bab/NwPWZLoFRpN4elaxPVRtgoLdazJv4kZdSxwQHjJtQt4ATGyn/tJ9
Og5sYoq0XtJZCby+ZqfuhiMgOX5W74N+agGe7RtUZPOXuQWRxN+pBk/2JWD0ol39
Dht/BjZHBekvpUJovWu4DeJ1m17UGDb3EcjTSzkquBgBzwfvtwZMNvHEQ9KxWa+d
EzaV0HJN/LZ8HW4EXbjC60wQ/cFx9ILumeZLhPg07Fjll6gn/CaVrG4Jf5LO+pE2
TtVCn4pMIT/HuNxdk+AIGj1R1RFd4HlzFVgOwmAl1ynullzoGRsPzUXGpMH2/Y+g
FlJqiwwRCAOLFWuwy4g+sr+J+uVO0r7bWvripTLsI/a48sLQS94BSo4yerFoN2rX
3PgfANq+j0tgLO+LcXpw9nRKVJK1JFrkZLjH2KQpsCFNyUyPmGYrWFrGDezBDujW
Y8S1cvO7B7OTnXFaz5RcBzmPd6LKeTono7ewxptwRo5fYtcGJRn1/+pSeqwnEavD
Wj3Utuo5fkvgMBwV0CXwYxNHSb182xmeIVKUANetxrfJF0LE8a0B2/AzyZEkn4qm
+yF0UVLCCE55bEgaqgu2CVoqu2yMrC9Oz4eShLRsieGzAqr3Z5x9Ww0+zZ+XLM1V
vDDPelRVAxrfkgQYp/WR6baNK9QPVJ7P0lxwuW76t7w1gYvXs6UvI3QNTc3o0mET
w8c/kcf6273THOrJKWqTuMiwZQ9sXkqRIHGGnccErAY/X9IVDxxf08bXd4lwBZml
CLkp4vI+eo7DuDuGwe9lYlg9txTW80n0vVlIpfUfDfuTnvBvXGkKhtO5Tq7paP4s
I6QQo9U062GvntSvAIir2Ossn0ZuXPPzwuNrnSNkHP49fE904n4kMAEUHlGgLsli
38t3qLGr/eRrPz8uYbLq8ZFAjFeMRxrF/A6ievJIcDVtD9CazaSsP14uFYJoMDyT
pK5YkInC1iZjPGN2vJoa8egnbit9gQ8fHe2UvAUFJesOgIS98lP2BBSpYHevupQo
hrfswRsSH2rx6elEp3+CaDhTIZLVlORJwPhaVGZBN7akFxfOmguWzvRpl9Ze/IxA
0QdOB5a3VutKdxVbvZV2B/3LlL+Lw3IohXXdoiA2ZUoKH/kn2SfWUljJMzqoFNyC
FN5rOxphTFVRnluN/LXw2Co1ZC1Y7ub2dJnGVghb6a1IpQSX717z6QnD+cPuiAfJ
7kB17cFc/Xkt11iels/LBw/nv6F3yDVlHSoMDcvHZuqwvHZGQuaFzEDtQbAxgEAp
zNpPE5YCkpKs9I09gwFv0Y9gKqlE1RzzA6fBQeUgO9APQPu6VDMq4veTPUdu1Esf
ekpqdtN35OkwKL0/kcwPZFPO2xFfMhq4DgMFe6VJbA8Jw/qrMNOXKFh2oTYQZT5M
DY58ZPFQcLkxXws7M5OqE2KqEyS6mN5fhgm2ENOiYq80nMteabPt6C2WX+rvtD1G
znMC4sTZkpkG9e5QKLtA8AC3Zd+pKH0pEodStFxWU3KQWhS1s3b+XDBVchXs0Vs9
SZ8P45IDXyksiZQ2VP8PtjTuN4IwTpku+71t7XQQgpnD4/qeDftz2LzSe+isUQ6C
OGdgwizc0w8VyVKETCgejJp83v79lcs6YSZitB+S548wo0FRTln0Dyg2yVU9bS1r
X/LyP2y/PEqmVBHnoSyo2DZ011ek9nO7vwUR1+cPRm6U/wld6dQWWoU8xT3QIgWV
/nzW4fBXv7QNT/s+zLq+MOzmVhpWoDlwYwO3UikVLsyZEvvr6TSL+d3n4ohzZ6CV
Aaq1DXFEx88oJRKWLoWEY6XSq9o8wi3JduQ4tFfvTkP88z5VWFbtXIsjBUuGvKtY
j42xJAk6c8EK8f6g6CQVWC4igIlVa3Oz2J6g3ICuk4EcYos0AbFal14anaJWnal4
RKWDveufdkXizzojemouLZvKj3V2glwbF3I7+pMn6g62tcetKuYIPcYkmTheFkzI
NDBo2ywiUiORAVL0GzRSnFHG5lsaIYv7ezFPKy0sRcTIMrLUYkps0oW89fFW1dV7
8+y0VGtDZYRz5NSBLyD6C1KAJEPoClcNtzua0PapZn7jp+JxBhi/nmvFjUEnLl0g
tVtqh2PwoSzN3zTT64BDuVRYRVqsgw4fp2Rm01A7vESdeObtmS2xNVEzXRE21o7a
yFgQLSYeflq881ojysoEKBju/g7jJ3Fzr8fCbFJvrvI+xWCtZO42pL4ItJzrE35p
lYPh6RRJKzn+AejZQiD6cPyL7j9NelsIpnhk6UhS43m0HY3lJlhmAl6J+UjuxOfT
WIWGZRiZoX1IdUg68r4dybKkmXQlrcPz5KyAWZOlT9Cy300NZLB3icAI+kVI0SQq
pBHQbLdBdB4g0E7KUKNR8ruTFloMEPwa146Rqczqik8+8wErxZi/7F6Trs6UmxTn
uxLST9iyTtnQLf/0NGs1oUs+q61hTtFyLKt+Jw+/yyUhB85/p7Ff+gLfdkLvnUdd
CI2Sql3HRFOPGPfZlKfvmRNrdomMx0EkzwOtbZgJtq99+teb54RxxoCN/c1fapye
YCKj9ccDX/+WCW6Z+z/M4WbUT7jLXPPgGz3USuOJ1BnqweM7mLZgr2VYZhcuRjP0
t5s4fGD6A//CVfHUYpiLeSdBjp4Vq55qT42hPVr2dlihXJPCILnRRglvTv2coidN
UA0WcOVHH4Cl9aiSt1KB+Dq1Sd0pdjOAbB9aosaJdDPylpFpfqLmFIzLdiWgxCWm
hKwceViDZykGoGFOODPUWbvDezPUkIaHz/6L3bfDWUZgfFigFm3t3XlinexcI9CS
X5eI8tBqGcPpmZ5YbjF773OGy5sLVqDBsDHOoIgNONL61UzIav9RtYPlqDPREj3J
a8ss1oRc/EeKogTe326j1LE5NOfSbC0oMJLilI83GOpEz3V8yB0b2eb5Fqulcssy
GB2Y0qYENeuL3glM+ABHuFb09SM6AkZzfEc/KrA71FX6wS1iGzos1syCVibibKb2
o9ljxYj+DaBYhYAz1sxHnI5teTaWZwwiJUHIPQrTD1+xaLuz2h5T7ibRM9LllA8e
eqwWzK+bbkx7CBtkFt2V7XrgnN75+etufcfHrrqyfLFyHN5FSF1M/DNRHbNE/+nX
YV/Uns+doI8iKlZR4oZvzZe4U4PZECviahFZXvDYY/HAEUC04T84nV3+M+OgD4WQ
SYEbiUg4jnbMYfU0lz5Dxv6ACBqq1q0ev2668qic6eeJG2OGKv5X2u6aSRLvMt2I
/cfHyUEL3YSoVPOeND4/xZND7Y0xTW10ghzpN1csK4klDaEQyGLhe+Qb/0HLl4u4
7atoDcoJJ5Bwb4KltEPKR6l7OPU82yHtXY/EXXM4YeGZQj0H7BCoPQtTYL8il7Ch
lfglTzQjPGFMIhb6fBokYcLhSU9GRE59ObrB3ho/zwIZflKRtRn5MFxJCo7Q3sp7
xudW+A2jg1akUGssSPJFlwfvCFD3S5y+EDlc/Ka7Pe3+2e1oFuCD6BmvfYLcDc8P
D0JljJb5wkePsJfPmAUGu+g8g+WVAtRvZ5EW10eN0t7G83YDdwF9yLs2Iks76/WT
+DXKHjop+zAuCYamlYFeaSu7TPTA3NqotSH8Eq8WOAOyVI5FQkI2pU5ccp42qNVT
zkk2hne7Vz6ZdjFZ6YK0Txv9u4n65XvUGATQzja4q4hbFTGct0uDQUY3ft0S331x
v24DtC3hMaEfAZDJb8tCeDoO6Qg7i/O7G0bRk5He26YTi5/1BI4Uw6WEYfqKOY7Z
zl1bP0IP3ng2CQgPEJVEudBYOKR80fnaGZxKAAZIzFiEqZQ6oF2UzFLLPMKzsOSx
KJkklFSn/2HtSjwkGGNxslvq8LB05IUwEyuSZNT0Ud9GFOjatGzLPn5/yk9m60Vw
yFMAEYmdmAPS/eMKkr8Gs6QuIvIBq+epDpXFGmCsVwCNvuNKo3mpcO9pmPD1Xk1D
z0ha4WDJ/YZvIUbWWQKACi4/8/BSzDe2gteJ3o8YR9X6pA+Dl/Ha36BBSl43AVcr
7JAPWFNo/xrUil8hDJp6oC5G2xQpMJ0rDaKYUeV7glTxustfXBRGc8xuiGg/bPju
pAsDbyhwgyXJkQyXMCBaiNZIXXy5efXPY3E1TwAP1uYgNhZQo6GQYNuUqJl9B5vH
sheQsnA1IhJ8e14oB/FeHUaXOivQBu1v7nxE+auR9NdX3A3//FHJFZ5Y7eZ/uPSC
KlVbbwW3Inz/UeqYW3xmhvXn3RIKXMJhvwCa8XwZeX2+kVUvs1GZbA0iLsLCJken
mFB9qgoRf6zQU16v5CYcqB+ZSGmQNNxUkbQHJrKDgj+T6ULVEUYSekdsL+lzGJ52
T32TV9UInZfybzilCGrcVoeZHxX9s/pVJaVxWjphIfkniyl+iCR3lDEa3SdxGJjo
XzuppAB3w3CUFHS2AJpc+hvifvRdFHSwUHKVFz/3j2yUfve5LMDD5PILlqhCiXfM
qMt+57dR8RtOF9Ra82z8yFjlvwAz00/iIInYn4Xpr98RmR8Ft/DY45D6k4JAYHzI
ZP+Ay4T1P5BWlrcRbMdKpaIA53WK28SSy79pHSYLUut0C6RjwNGeHimRpb/I4GPb
rd/FATrsSdZ40u5Adh3TGeeF+eOsxX0FTC3RHZ9Hwe9FomcEbDQsaJJJYWouOrsq
VvHgSqR/66g8fydom0O7uZhzC+xJLsTFgvUJ8gwS94FxVho1VKSwEULNYAJoMzQH
M4znZ0ndkaYO/p+/egb00xj4odLdAyUwscRV6u8NqvzGOj5pBYQ7sIQ50gjYAKbn
0m94MC4or7O9V/BzEqqLdD5NcYUuVjqWu9NOWkFRRbH6+m15ByccKMd6hsqoEWJw
bEyTp1xjpTREdChY6985Y2KDu+xngoTRWtCr/Z+tvwKp4Rl4tjcUkrOBT17+Nhef
fzz4uram+ZMTxkTKiEO/MkQ3K1/WH6UhU89s2YB/8qto+Qddu2/4nqRZ21wlh7id
7rL/WZkc9pHK3MKp4YhzQUb0u2jgtlOV2m/sHindERs9rNX5JIjDkjA9y8Be51bD
rf7bolm54WBiwubV5/Z2+e66t71GrU48hsW+H8YORUHwi7ng3xuqfNnNA7P8RI5X
bY4FtsCQHAA0LUdrD6+h/ahudDdXWc1MVp62m+gboCjLheQBw9xIGp1mV2GxQ9+8
oLyzRjE8yya5qar+nXeNshGIAX8YLMv4MfsAei4IMvcOZYW+Sr+EpX05Nv0bBnXX
qwhZdsgq1D3RS2vq9LIKW0oXyw8RCj/fL+v2Lk1XXUk2e24guLvAn+pok9SDEP9s
eyw08k9Yxtn/m1M1CjN+SC5z/WSYN0jsrdpjENSHH3j6qwXmFB6vqjUrYuXU9kqJ
qzdrXSeJibe50K4QZwyKZvOWK7xWGCZbFnG9ZldOFA4FcwqETXvYdVXd7V2TQvwl
K48lemZQwe89Fz5+AwK5vHMkf8DFVCUqN8RELLB54xBdv6MGA7p65eJL6PC9Fmcf
gQbAwzTJr/i+l7wP6ma3EOncTVVYGcZtwHS+DpMZsTEr1VviNID8cHaXr17oBMzP
lzsJt8WEQYievwxiyUTk1XAr+lknmaFDyQ3AcshsJXaxBKEdfnzSduYgoCSTzn7r
9L4QvgZOPFwTgwjmuJbx0QcaP2rK3ExmhYeD/G4x/e1RJvJNLTobWhZ7iOZ+geym
w8elup2TgKFfqU+LYx3fxlGEv1Xw4NMyRucV+TsFcNC+hT0/wGwTtRRZSzvxu+yw
+awVuKnav0v1ws0eEVg0t5VCw2Suigan81wSiqGXTi8j4NXxDu4LxVSYnAxPGqiP
umfMMyq8cUbJqozbfDTm1TtPt7eO2Ba93JyKeCcg3rJaj4jiIvUkgEr9uWQ5Dah6
IAK2nG0YWw5fMTlPAUItugy7kKRx2O0RKi+jJGpuHSRpDeI6iPHNLGFhUDOfmnUN
LnBbeDO1ISNfaAYAJQTiOmixoCTuemmF2eDPCTPaQ/Wf8NJrxkAK22XZoR3OB594
oFd/ngkwGCZD9BuAcXRyDVig4WqI38kspM+JNL53MH3Afhk8owyzEHswk/j9E38w
NnTne4dgKklv7LrfBbs3UQ==
`protect END_PROTECTED
