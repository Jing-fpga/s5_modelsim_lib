`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IMnibCtb5cV+o1diXePvHp0zUrX1yH6pOJSxMOqRuCYE4f7q5PlvPkHVh0C5TcMf
2AjdG6VApqFWDQxvPMA6g84P+PIPGfdP6n2S+++h7+g5wI+r+qFIM5FnFn///w7x
0DgGKuHqEgtPKtObw+lmC1KYvL1XNtNzcZeenUMsDlSCE3G0woPvn7LnTubtcJ72
JLZV7mcOvT4A8dhwb50tHNkc5X+r1WpB393wnjvLP0IWNdwKlpJ7CyvwV4zK+aTX
qebRcFsEXHPCTtFOolTwt17Xoq3faw2xPAFy1zLPqvjRjYduIsxDGljKNvfpPPYX
aCtdtGzF03de1WcyGd+ha5R09hn22xAyO3BWByOhv2psjWdYdQNRlYLnvJSzLQTw
VZUvkT4IiE9T+0+WBm6YzCA1YrKebp7mZ3GkOU9D/w0eVws4ASEJ395ZWSvtlFMM
S8vQ6XYB+1pMusZXL/PFt8pwI6k/dOT3jfB6pk6m1KiLGU0B7y3ewncBdgpYcWY4
wGV3MyF/ZIBVmIPItWue2z/qk1Apl3Tz8bwngeH2BjnxusLNwuNd2lLQi1EMFX0m
wFw6t2QkECe5MPCtcVlHidFbqJgO20pe+O4Gymvt1psgFduqtpdCQqOC5wKT1XIh
XivaHewHaxye9u4/QW6A6F1FeleoxL685AmtGBWcq6zu/PCEQ2/dttz/ZW66z+hd
Q9Tq4AOQTvw/rlWGAmr6Yf60CdShbEBbY8WLDTpC9Z4iI8YESHz01rmH8BQHmlPy
GytLBFuNRunnYbcApEnIY00XqylqlkRVZJJue4BnkTzOtK9mtnJQJlelz6cGbpEm
94mvBC4Vs+sO4rN/lWvntyU2oVC91fV6i99LDSSwn6MkCXTFTt/JM3FmJI1s1jTO
VB2QG1iRvSKFSyZkADsiY1hwaHr9R8s7y5JqwEt4PWQ4AO4nAbn+rhjsS7NG2sk0
P4sGT96nDjzXFBW5Her8ez0J3RLxYP1qoMfHh02AbGbm+4KKYERhoNhY1PYohRUb
/h+Rg6VELwnkKyS4h8rt7XFfdNS5By3NmHyrUMn8NIxzOFfbED+9fCUkvboEt/Ba
w/NgVCztjIcKXnm6OtkHYgONqo7Llzl+mz3wvbMNdvZdVr+7VhCklP9vfEVAfPTL
FdTItBq9URHRhE6ykwCTdZi1pZ3JpLXPTBThl6mRVNjjJYg2P4i6b0tYv83JN16k
WUk9dLHHZ1oFEue7I2XOqUt9b71Cu7glqwrTq0cks/vrtZ0xS2ca0UlrZ7mJ9XeP
/3HKtke7Hxe2XZFXjtou44lqfUEws+YPxo5rVPGjtaFjuyg3hmkhMDIeXyaXlTc9
myicsRk53NkVuV2Qawk7/MA+VgHxex/SnBLgw3c3j5dsyEAhAMXz1K1E5TKuT1lg
VyRfQdb3xPJt3q3o6w8sSXv7Xfkv5wuav/VT8B4Dt2fgWd25fAArdwztdilKvxSv
h3pi6FKQuwrmZIKWlVcerkckqYGSnd7tGU73aHSwqbf4fP23zrQ2PKeha/xhFiVy
JEp7xkZa9cEUxREMx0BXXbNFPowFz4omIaEX9BV95dGbdCVQX9mj0PfUmRzO4YVw
oKxqoTMNDYElwrdkQGPbIV7Vk2jagILhoFLby/DtIaCRIUQL3v/mHJWB8yvK2QTY
CkuW1MyyQlUfm8I7A5j2l7Q2tY93IFfl3k328QTrNGwALO6tv+0F0yFkRtcg+BwN
kKsqbXX0R/IAEMXTCnkc7H//KWJun38Vu8EsD7zYuyATcRmduvq3Ml2aQHbWwI0l
WCnmfKE3cmmCQCKwq9ERzHgsO/KjBP+r785aKFDGd+cJcm8ZUBzcBTc7I7xR5v6g
qiYweAm2p+slTLGE3WcaQzmxgQc2AnwsxQ1SCrsGm+2xmoPe8Mg4YfNpM2yuxZrt
tEt/t/UqVl7ZBbKqwsUdy3l3uNMPFGSs5p4c1dUjoGpkUZ3hmJwNgqM6x+af8L72
H1RFDJcSSEreky/H8epkuOm/FK7j7gf6uqClsQIM03wqzA5PoMhItBtDpd0uG1ef
lZHTxMqCHl1vbcK0ePYzIsnuMwrJ0MDMoLfXUcrPr+p7DYp8iOua6LhbCAkvYWdS
YC0E/PIvZC7MIvPru/YcThg08e4LL12VqPpdgMZNlokS2Gv99ApP1LItyV1pjTDp
ly5FmVqu2J/AOpzIDw+QoIndfVO7cjzTHRRny8H9x5Sfsi9VLSxAovcEJdx/1kQx
VeCm9vNa10w4rChDj1zGKUfUQ8mAWd3rW4DewjWwn8dUcRxrNPskZYatmM7zwdyT
FagatvIov+I524W8QZMmfSTNUVpML9KeoMquG2/LxPfbheXWiPxzf++1chMo4xKE
5MpVoaBDuYIo1fvB8/vzYj4VNrKxWs+v3f+vcKJsk+fszoJv7XYY9K9tVEtgCjgM
1AixizGSIn+wpczhZc1KWCNtHMEjDgMxva1rAzSplUwC66ywkid1I2DvBZpYbVf7
eOpFadTT3IWxmXGeZWt6iLfCf67lVtynnGzCiiPxGuQ=
`protect END_PROTECTED
