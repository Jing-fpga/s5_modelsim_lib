`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N9EHXt0QZxVciKIOBXTxGoISCrqouLN+T7Wm4qs3JNndeXEtn/w59lilBA17IAUq
tkZYAl84M8DHY/HEZ93bJQPVA/0/uINpAnYjUVVBhIyD014w/di2fMW5wXPC1oK4
939dpRgAdFzcRe8/GRKXEXLc3DeGJrBmyn9ODrYbDD4ca0mNdvGyU25G9NshpBNk
l+tuLKJ5mioXckl5HGYtjd1dIQhP1zPDyma92p9pX0lUO/hmp7yLTUYhFFX2KCR4
xuJR1gy8IjleA+q0MQp/62vAr6ZwxKjBeiS3Ld2pNyPMKxE+y6pG4b0eVxFzLeZa
mIElonKyvbyKfto5322zAiWT/N9Ai2wyhLGFMveQUECoE9+BVZsa3hwUNjVNpDa5
j27GplnXNxPpbH1FRmkKSuTY22ED1rwNqH4fLGT29NyfnjSLz3oKvkIXczcwCv2+
rMXmo816WpYjFSJvIusqhkcrA8f92tO3FbnWX/ppPYvcv651lhbLRekBpZ2nFNjs
gHCwAZOzp+0R6vSFVwVnvFBX4BoKLN3DwdJf4rkdcwGkYtAXlemjAUAG0YQHO65d
PB11cWiO18z1wpw7Ml4ZBqQ9K5vUp8+verls8Lb2DyrSXAS4b8RE8Spz8yizg4gr
ti40rMhmOoluuIFpu9H7h2Ybbi389e41XfeZXMxuK/YnUSGfCaAxzdtuWTl2EedI
/3g0DgAmV614ANvnnTaTd6BZu6PSRerOFnlnZS/Vz8zrb/vgjC9QO6RVpJad1BFW
eQImjVdrdXJ3/YDwccv2KeUK+CZCHWo/0rP0c9skyKGWYpA4cTzik/RS4Rjco0zb
yyif97kDpnAPiCUPguP66T2ky4+fBEdDXPYZNZpZpTp395BOvU0KZKQZ5KqqiahP
tUPhnEuBobbbbsZGZqcHPHg3XMAItdWyxjIJOyrkUPLWChedrex7R41RvoRj1pxB
6din1TOXNlFrNVFI5GRPw+eebvyxp2FGmstzKMz1tWYgUhJ1ckTeKwprJ206kp3N
0WUJE6UOrQTUXCO6bHuLIYDS9bH71SCB13zfjBBtzelAkukdscexxOHCBYFnWoPI
JoJPVr39anRnWbNDt4AG9xhZZGE8UNX0Krr5C9hAXfCbgt2FcnQStGGgg6fD5HGC
575iXnE8oN0eXWI2zMYDqZiCGho4/nzj5YOJoBEtHQ92QFWSt5GoysgbjmOFwb6Q
4CdQII4zy542J+Da9jx87SnK5uj3sfkS7VqjrGUeQG+FmBdF+Nw0AK1LBZD9yrus
UNM4/GMp6p1Vux+XJmWE5XxyPoZSfRWPp9FcbRqaiC3LKWKohTvtNpmaMCtvsWL9
V/xLuBF+x7PZ7mKEJO9lH93LnD/QD5k2myMBi6HrEsTQRQKICF0Cr4DcMLeM24iS
+jUVXR+Pghz2shqjNuLZ7OTuX5/2J20vxxUTFmgBZh/YsYH7lBfH3y9evHJ/vbiV
DsYvvu25TSv69eN+vAvoeFlJXu1nCX6a++cMYVEXi9bp2DIdifSxLiU7Hly75B3c
No75nzmjt7XeOEW95zUIQhOBeF8PpWXxv+a0Hod2/zQlkFDxnNpI1XuLPuaX/+Eq
Zaqhwk7ezdIvRhQRQFglVmKlbI7hMrpgQWboeFMDpdujLernNVMyhSBjIjoTGeIY
fIt/gLFpW2xau39DiZywPy7a2SEo0ebzxUSs6w8sdfMHMk8MTf0S7X++PcQ9E/a8
/G1ySHIP6dYu4LZWqS0HQsLla7wHVqbtyuLGLo8YyWm3E7f0aBURnTPyGk58Els4
ZO6emhvYqTuzn5cL5/QOUQxUDBqLLHTJYKvJytHRCfe087loj6EQ+txPvr4coxrE
/k8C1gv9SasUG4Srdjzq91IbGu/M7xHpv6fTWlmUe9VSNUTJJS2vsSnzDAbqXdlA
AxhADmMj1XPNo1e4uJF4LSu9uDMFZ4c8Zdp/mIVRKazMxMhZj5CJhysdyPhAEFTm
ot6kkJaPb2oF/qsWHAM2YnS7Kq/x+AOGQjwXMao1utG7eJKzTI38tDZH93BwU+Yh
U5yirzp267sRU1YEw8iKPlasp6RRIeyZOeobl3tnPt1KLL8YpfKrnF00p686zXeO
Fiblf/8HNABf1ZbWpeyhwGSEgBSjmnwp9+AX+bys+TDq6zQlXeRA/HuG1NxjUv2L
xM2WI9n9aR/+f0VV+w3fBbp5MLCqrzfJAAHvAwZx7x9y7SzqE020d6uWQbKYdkn+
kM7PFq0pghYVCtWz1jmEO6PHgM7PIlXAicsMPKxKcWHFkdA6ZRd5LaUYH4DD7CfG
dNa6YAe+5j+I86M4PiyeJwCtdnQSi/W/PDfLZSzZgZwga8UMQXtSRZ8omF0ROSE9
gaEQw4H6q7shOctCr/eKrjoMnLM/+FgTjh0aEIZTdL9g1V+32ho9/8tNPrhGYqSx
YLqjgUQnDPiXb9ECgbNGVoV+nBG5STMB3mMBo4P9mPh/CJwZsR1yCeo9PZfru2zh
/6ti7wUFSAYX/oaxUf3cwMH6u4hSdoa0/TS48g/c6qm+zK1HDEI2094l6g9p2CcM
A4dlz1XWJm6hGgIqq7eZU7xqybUlo6aVBu6HmWZw1lIrBi7k/68sC7Jmwa7/6h2n
BnDgf2DhX+Fh5VGw5Y3qtWIN+qJLy1SdqI42DD2CFaLqWkbFBl5Gx5LyoJiw8WGz
uwL/WBlQkRMUaDKsa7VfC6qJ4ZoUS3NqQtOWACifvwHrXZaLZ72sRvA8IaPizn7M
VIqqJiOH+GWe/koj0OxFCOKWJtXukMqugFS/GrFMfes0J7eM0YQLahCZlSAWWjxy
omQe2MNiSdO92gPOwSlRq1GbmAmmMHnfi9hKs6cGLRy4q4NomDyCAbcCfPtatHMI
k/XSz6Jx2s179FrLZBYjPxocjXP5qsTPIr9VfqZk8TbCWHnzHAfDqrVCs2eFmUjl
h0QjpFVfqYP0/uZOd82GNRWE/0G2iTAetgaccpitHET75+jzFKO3l2tWWXQkE4qd
Lat5ecIcEgS4ROQrBZo1iJBIRff+C5xLKDFIH72m/kLG6sJ4riUbOo7ot7UCO/y/
IJdPMqUbJ9LxmqsPojdQ4vn7tyMNRTtFzOmqtixpm3GYJ3BJBmwTzLNdpX6Pk2wD
NHR2n++W/gbW+bPF9iuIC4Phq6EW6BY4dQlo+2GbN812kFA06pBhP0xUSrfJCKGH
/25MphjWzdLlPl9fzGq52jPHiLjMZwvkT2zTFmzRNz+WaCDhDWrOL17jtgmmJbhs
/BOaeYcyjVVgoFXvBR5/nJk0dTOUN/L3tzOEKQe1SlK2HTtYqZe13wz08u/oYwxx
QkHeQim4ithLNnJSVLAZOdxYfibECA+68XFl/h6Ir3cUVJ9YH+GammPm4rEU0M06
b/XXRjvUaF6mWfO8V1F0NrjeTo1Yq4OxVyZToJtnKBsiXARz1IhlOaChU07UGEaB
oxBxXdwZ9jxv9BMMQkAHgb26lntX/EL8CuYOeTvtr6Q5eJGOsrWCRKUy6eT4uEyN
hkjv4/kLCZc7xOD8XJgv8cE3aejsNs/YwdOCPI9PY2Y6GckoiAfxMiPsQ5bijEqw
fGWsVRJCTmcgbbpL4NipOHB9ObK9y2UEcN6xLzOOYlzUoZe/cfUcU1uR5bLePmjz
xc8wuJO8lncBZgwsNWmKgyGXkYwRFwkRL9BzHAU3Vl5tQFqAyql9+EpKSAbAzUE8
VCFPZc7tPk8ThgWDjCfHzB+nRkDOqS3DnVR4ufXC7cDcZvdNatXY+dOgVeywmUEH
Vw9GUZwT1PyvVYlOA82eZH5MxvnChECmmYmy5e1LqAaAKjc6TEGA3qDQIIIYZc4V
g7jnXKt1z3LzIKE/77uONmwo3vCHAzQ5ONCIq3nkp7wjo9tUZZFr6VeO+30hIlcU
9XMG2+JrumZuQ8EkFisPdd85/qc1LSiX7PYRrzFWCiq+LH9WvwASiQmaVwoQwQpQ
3lrrwhizz97BcxpubO7d3h+nNTB2juOh7pzMB58Y4NmJFdJK78nUpLIfYoPDPbnZ
kN92ZsbFI5mIFO22BPYt0Z/KPdplnjH96yU7WsrmbSajZ71UlNTnujUoQYhVAZUc
sIezqHQ1Q71udq+ndEnHdrxE0692oIXC6HM6diqdHEAG9pJK1jY6dBxzh15yUut3
mo+W00WYWnNZP0qUzAh7RfJvjJq0AmoyWIM0Sc9wCk77riW9Fb199vuEfT5B3v2g
ldtaOP/rSDrTY0JBVYtiWMsP76fVKaD2BUlfzvDToRIdQ+p6gsSiLtTvnK9rRDj7
eCQT0BxO4EVqn7LZ2DdyjA0w3/vQGD7nL70pVJKaWn2LKdoOJuadmjeTVjo19ya2
49S7KUv9Evqhb4UdulWjmBK6piU40SJhPnt0tF/8+iIbY6N076r5k4yBnLaHiXBk
7RJ9sWk8vpSOx2JxYEJQYcg81TYHAiP45g7l0uWxMdcJzw7N6Qit07YgySIn73ck
YGIw64fTrSIeqLpzHl08EjN6WbWobylrAf1UU1yBwB1t73Tce5eVqL7LjG3k7t5D
DjK6fYk31QxP3XnWJ6bfpGXIz4eoRl7yEg1J3fwX2FBGJxbbv94yS5QJ8XKESr4b
rLW+90Tz4Iae29WDvAcdDzGdFjKRn7kuXKD1dfOjpBavhZAxiU9/zpb8Iquv6cHp
xeNWWaCMNYUiUpuII+cagw88bqbaK8Ka88QnzSe4+WEiO53FIPX3StKm6q4oo0wd
Re5GX3z2rkcMxgDgKsCuC3vKv2Ocm7QXALK2qsgQrtQV8vFjBv+rZ52nN6yHzwGo
t+f5LngcAwBXsQkcqaEXC4JAJuOId2D2xhVdrGjTBxW72pgz13IquhZK9xKZBYbl
1/YRD/52ZY7pm77NhltFcm4k5JJrGDCwVyBOBJaYeVzd5SFieKEZl9MuvFUE7cKv
6f01fHylC5nTvnJO/DpwkmYLLUzxbU432YAWhAMS3eI=
`protect END_PROTECTED
