`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s4W+7eb8eXCNS3A4pjiwyHMXfVyGZmVF7Xfm3N5Ju/5ssysW7Mkr8QFdLqm6Qiy/
a3ElDRC2ydARqA3Bw3Rq4/2bdF5892eVjkxY+TNnj8op+rsL3rJ7lk423yrl+uXP
bvyg50kSe88zBd0K0SgSCTOWRTLhZlp4j+VGK6kWxBSGIG7cd3Wovxp/FWTZDkby
bZSBcCJsxlQhdW8JtJdS8txc3euxIee4UNhZryDBo6PtEVctSGvzPVtnOD3aMTbF
SND+nfYfr1i6JFpO9SpV7TiybrJenjReu9jIx0mMaseizct9MGSUoM0oh71C8gDK
AfwdxKHS7D0daaZrAV72ianJeFzzoom5TX4Qhtcc+LRnW5ryZOD0bbkeubrl/fsS
Hm7idVD3f1IhTWoqCbTU845FnmfsNKMj9RhJC9htWGuhsuN1uMvkK8Dv735Z+J1/
FLuyIx/r34xdP6CZXdPDZn6+MwVV9Kw5P+bka98W5n0NMjn5riWszY9demxlhOUj
v/RcMpoP/yRcMMz63+lqGLDb1DhGmKxoJLBQlArTHJhn/yan80whluHXI3f2clN3
GzgkQE+4Mu5qYgUPWWSPIEEpj9NuiPfFO5csmS85Aj/S5flY5naS9sh+Jaw9rcYQ
vqL+a5qe8FZ/Iz7LzMx/SHmW4jSfirvTDoIW9WoqLsYtiJoEIA/11p/uQXCON1zS
sp1Rrf60mNNwtDUNzDxAv15oxTTGkoCooo7KlOi4yWb5ktr6qS1fMwNUrng9NPV1
Wnw03kOztS+V6cjld539SiKlOvZ++B57C2Zo0xe58ReGqEaGjH1Cl959A5/GwNDz
fDSL3JRYDdTvsPWQrcnVMN/JhL2lTV7vW5CR9wr+ydtZZDJE5+paOjU08MOqOv3I
mr+3IhXHUqRRYCjqhfLazFjn6Zh6O+ZFeZpkLL8UI6dhfjM3IxKy9HZSzTdYvtGh
Lv6DhPnRKSkHrFV7V4AP4qhGtIJ7jLLZ4jZ6pwrm3bdk1A3xNpLTOLNNDjES9fLm
6RMZiJGHhK6m3b2HvI4K/TteAkiWLbpvFsarg0nA9SnIYpvkSt6j3Y5vc+4WWu6c
YT+45cnjaLc2eErCJYf1kLUCIxXwCyMs17ByzgOIXmaSnGvS9wgSwF6QX5yzqZGZ
yqu8bs1zdaDRKK1Z8C63qzKAD0HHPvvZeE7vqvXEVqqDsSzL1wDY44d64cl2enGp
ZIoLOCFX6ArmbB6/F+PMbX9CZPSpxJHvw7nhSGysm9IOOckUBB/jMZhLnZEwAJEL
yelV0rkkkqYlL8k0FOxzJxdHv8r2Mnzy7umK5vUDQ+wPLkDpZPas8HgKf1X/LgDp
088Chlq8h67y2y7c31D+T3A8WOXEmQw6CGlWrEfrWVMjhUTN9NjIhP/1bOqILuYU
K15XNLFS3EzMpXkkuIFJecKNjLM1IWGz8JJMIZl5uh/tG+ZGNMxmrWSapucJqN+F
6qv5F6rZ1R890SOigHcw2k5faYlKfXWOjpkzq3bv60WW7j81nS8fmz63ig7ccwON
X2lcXObfZFqMmBq4vkwIWVgzoApGACHmCHB8tLoO5Cpe/tPUb24WtFdqTUYK6sHD
jmRv2MhJ+xVIXE98sFMtx+g8rJ0U/gCnipT654g56OhKNZ6YyO9xvidVWlN9eWzw
`protect END_PROTECTED
