`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2MADceamQ2yaN5QKx3dN20vSqsoh8WNZBP7D5RFJOiHCqHHxFDuzQDpwGPNLhIc8
8xhy2mtYN+B43qyIgSWSgD0ers+XUwe+k1ZFInVu02DCJxOV7yOI/S2XTpf7fHDq
8xyCykMFjeJ8hiWj3qu7bh7ajhbte5G4Cvk/w5N5RFEGw8tIVCtIeLJWSecxNA8F
QI/YrnNxrRusBDyWLBsqWku5otz4EbsNU7dGYnv5BtdwUE+MCjBqPLugR9lCw1c8
H4UXn4R8kgzo9FuhleDGJw/S9KsFRLHbANOWtT9PbmRpeOs6RatOmd8ZoNc+PcpF
RCONcd386A2W1mOqo7zocWM+8dcPL9GgzIr1xonUR1IXLobLQCAw6ZJiwlwjhgOb
nETiv2cOHJEW9JAc5OP84HxVYk9OwYACoh89bOVZ3iLarqXuhdwSdOFNiHqUSFi8
uHQrDu43uRI4Ap3jDZgoiOLd7LgBkYspKDGwRFjTM7wp9o3UTboAUVJHfndtFcTY
bJ/XOs+y+67soiIq1z2RXZR6AMjDoK2Ibmkhxi6S3P7P0+04bdxYQamU8wFll3/h
1DAjFeMuG9qO1QZzsfjgRQKxqHmKPeaxPUt4DTyDsCoXp2p3r1m6fJDkp/WF5C6w
0xSqz0DDweGP1yW73ogj+Y27bz5p+52QO+wTXmbYCkhDxFcsQEPHsgjkO2OTaEjK
SXo4DoIT2JW4OBY5yZk7L/1V+gwrmPPI1AUSeehI3P2mdfRIq5zGv9+mVpIMcV+x
XRQcERf+Fw6ZKB2o0vC/4gwi87upedAcVpBkHEhreujk/6F7xVBQDHcN7A1Q6vDe
y7JhyRhpOkf/ec1E9tL30pwWwt4IOB0aax0dFZEddOKKZAn2hD7uJ8hu6JO9DLRQ
URJlK5HIZDYrNq5A2NQoHChKgvGk5cbn3QZv75hgtkwtQBrfnf58woqmbRzdTCX7
De/g5grQlTmrASyFrCnhhv4uhN3t9gu9MU2g7X3slNkw0B7I3sdTgWyaPz+oL0UX
CQ9tBjavQW4rwnnwdeO6gbjTQSTwXUzpbskdEsEel6xW4elPabzazNxcr/Kk1gu9
T6z2cKLKPctCvHCaCAsJM23TufqI60nl4RLkkLuL5IA2S8+K/ZGZWG/qU6Om4bZl
Nof492H62A61XF7AsWYLWd3OhSUHi4dJSnjMAVr8LT0x6Dm8A0O0r+O3bISkAl8A
YQX/1yV7//H7qA92mfV0Nl30Juql6/AgZ7VrmPYntIt2WfwMBdV7Kj0C9ZsEohWU
HsGjWyYWpJ+VzOGU2vh++3uYFqEvJwvnQG4DJgg5dPa7+uv+uozItbUh+ZT8Pf3F
WRVvC8sjSg62X4ZV96R4IQyIsovA6j8Gm6KZm/Wxd5O8jXg535m1Fg/XzzsvyPH0
cNrOFd54CrKoPBK2WfOONNWXbdTsxcEFvqHKPFF08gk9k8uKCmPtZrzaStyugZr9
DwlJIbbaKZM8qRstK09G/4DuzIXKvTMqdb6KjOt6WYs9pLt3L8Tf0jsOgdferRHY
h8O33KCnIhmNTN9OXkXDdNVIcmVPo53hj7nOP3ykd2UbUbBjya8ECTaYAYzJphKS
uga3Z2xUMyfdnlilDgdCmtIXNGaXaYNnDSqHQDsmkizMB1UARQScrRL09xNAimuL
gDbwb3NGWcpxiSgcFLtlk+AOOlReIaPB7t++Z3rjlgVSZ9RN5jQUDHQJypPgRLzi
mRlvhxw88dc+zOu0BMXCmdEmo5Q/CXlkWHnNTImru5hTj8ZqWl/JPs4F9hUOtPZC
cQXKBCQdBa9kxF/qM/Fhy5b54quzjb05iepe9ztv8oueOA9JRW5xRcc5Bd+gq2eY
DLFrgdxCts4jYk6mvVnCBvNDcEYMkmkwD9LR5qRzEIzQUQwdORu+I4sA81Y58jgx
6dtFcMFYLm/9ZUgpiRURpcsB7kPNVMliI5E18uHUcDeIj451UE7ktJTQDhOnFEIK
6TOhoi3ztgMS9901NZy16yka4bxIoSi2YQZocpLNCcktRCK4nNSfMvYFn/0R9QRX
UXQQjFhyS0bwDMXuImNcaETK8S1491+SydrrIlV+xAJl/EJGmymk3B2U9lDcJY+3
otrYIdLzeSUvaDFj8DfwdxYcMX+WA13EUd+rlC/VvgoRmzXMO/YOMLW6aq8pKI3w
YfkR+PA7gz72w+hdvI/FpwdnoBaG4NAFLDRER7PyRG2yGtoN6qpJCSh9vwpGbu6+
sWTelaGK/D6r/EB1kqPcvSe90f8aW89ZJSltQS3L75rOadU+5KrvZpRlTVm2fOGW
Xn0c3w318WSY69KT5IsPocZL689mF+ykXWu5Z97RBoQykWz4/ixuykcz3oREanGs
FCECInDsdPZ1oPDm8xHA1A024H0ryWx2S3EGHwFdsabG5Q8YSjOYmQ7xQjRArL2q
lrMJCiCaV7WAiLVSkhn3O5+roixjAlty1Lqo7saLXyr88F6bj9ZNICE3EbgdDbkD
5I/49u2xoSiOB19UaCyYrgCAaAt5YeIrwF1/R1wYVlo2+gIKo2M99k5tNM84lOya
s4Xc4cD1zEFb+KuWZV1fT3DxLIo31CdIuWTezymMIMxaoJSGAa1v5OFf21oUn7r7
Ls7gqQzX2yULZhEnZh84f5gQ8ASG6i7UTjtcC2IzXXVAgYPugK3y8LUIQuFo+G+B
Rm0u96znOA27KgLAuDO31+x+jJuabjUSWFh/rDLm421QKVQlMe0jJrmrt94wQA2x
2C0pw9QcGuoDQAcitolkS3lD2Jx7xdY0hHflB0LkIRXs4IYvysNOl4KvVm19ufVw
kTrHp7JoX/omFuUElCxdIjMZUGwunAPNF/mSaXYMavKbRp0eWxo3aKCY9oeRa3yN
+kxMkjzvt0PPD54E7BdeIT3u5f7ZV4UAib/AlQw9b+h+EgnRr4r/gGPdIO31rHmG
ByxPjxWgFacXXzCE9YH/fBV2Ax2Aru7DcCZgILGWdPHC9jhxq9MTiEU0W2fOd5cy
wwZ8eWBEo4ZXJ9yVQ04HjxrzLl6DqicNvT3szgUQJ0jERIQoTsFCCbIHTdSfUd5X
mFvXdzCSW8NraTO/jl5A0RYibXH7V/no3NCS0pqMmBZjPFPlxB4T6vZPqnnDFuFc
Fm8nyVCJHMzhVP72lRD5sZ/T5KCkliVY6mTd88e8G7k/3r6lM1DJpWFavt0jV9jT
lBvSjejwqp8rOrNFn54Ej7Ay7MJMC7/eEEq8RyQBYYhHfPtBsBWNYX5eZtS0yuXZ
VuK8RYCo27prFZChlB8s4fm2JTy22WhwVK0dzEUBOwVJxQI/6jmo9aLoNjqCs4TX
zVFLIuhZrX5m5h8C7Y7ky2cDjBsQO0Bfi8zxeAKfMZikZH2fQvolnNtUfr/z4+TX
A/O3jCl3oIgpmyljTWzCTL6JaTgzuWqjT6/qWVYpjtggw68M76ALlGpvWyIxgyW1
CdFHmaGLm9D0Ey6rPzDmNhGBz5XtJVC4MSLZDJkIaH4FrJEKJQA9suVBqK4lVRTl
CpMPTUzuFjBSyrbzs0UOC03LHa9vssC/l76ZGLlYrfhDWzZ+pjYNq+dQpPs+P5QK
8laC34vB9Aqyvf+gzZ8B+lV8ec4cCNHl+EYPkNMPtYXnSZwc8udh3ugRVjYEzjAw
udOOTC8h4NLdbKXF4/xf1zIYsXm8XAepkXthiXGTzzAYygBX8lRdQnmPgQT2NC3Z
6cYRTPptfdLI2dsZu819EotJ6R0rWEzuWCfE/bWzUITn9KVVv5hYK3S6ECVUmnEV
6HHXLLut97daNLUagf9v+4Z+/QWWTIdEPvu0Es1KWOaAdTAA8YttZ8A9Md0h9NU9
raxm5kH5wasMG2OqRsywbzOBybSojVf4NYZs47p3ViVMekbK7IOA4xch0ztzigyx
NML7Py2M2YgSqra9y1eofKetu1ckQgwdqwwXIepUIJXr/Cufhm4e62yq+2cECsbW
YXldsfrn5MHllL7HF2+6uI2EgLgT+S9lA/w7RAymN2aLyOGBKmMtLGGrPhq/vjes
CvuVT+ZxX7S8DHt24wR8srmuoTtvP3wx6gUPFk7XAyY5IKVaHn6qof0XBbk3WBdj
Hq9ev/DScEuA6+JPl6GVEgi57UBSVSDgiKyUynHnFtlRDJUBmFYVpub8LTZyC0lm
x7uMHKZfD0Gtp7rrkBKD1pvHa5vVbYWjemh5tRIeiLeXUaQhXZDOM3BnSKAZdg2Z
OgcXL0ndBkSIWPTTF6MYgQBfH9t/UV8Tqb1S9glTtJCtFrBcCggEpz41gOZHqOnh
oiGHq+bzpNAjxosHuNPiHg3UmPimTIFiUM61E2LC4d5Lw3ZjM/WBbTCsxZwUbwgz
glhy6oSaMXxClauET5hw3fEdWBhs02KcRAYh+pOa5wI7vKuoFSeX+bW39qH2ry2c
bm4o2bAgqx6eHRqb5+bok3ezJkJnr4ptYdJEZSrOw47AfoA7jqizhuXrTajDZBf0
DO1EJVJ69A2Q/7ry1OFQ2+xFLoZegYTJMNwM2x9/1236fthds0uRs08YwDJB2Hi8
vKEDK7JNbHa9Lra/nYxA7z0Ol47SynseeK82vvCqHik3Ml+DjWULqfC7qRNz/iJ9
bG38YsivKWWjyPJs4bmKhiaKTiPWx6Dp/gHJN3glHn7CSlR9wluYDVKmmZ/o6PoJ
43xn2/Z0Q0SUO7AAzWVMcTCfvD8LTlJabicvSGkHTqDDrf1MJo34bCQBtumEHMhp
WcmtKmZZoKXimSyHjO2GLTMe3d34Zlh06yfUKrEzv+5ek7skGp+BdaVA6YiUFzET
uGYGaS7JrIAkT5carOen9rwdSWlEL2F2jknkhjEWnYDUygq25Gybhf4uAWH9uxC7
xQQdT673rpGgEfF30S/RPQEIqFKIfvX5jD/jme3dOpx4FFvtH3r05BwTI59bARY0
VoVsuiqZjGOVKdo9kEreAbL19gndJ5NLwSGm3I7RX1e1Lfq5RowZRJ7tLkyrMLh7
sNR/WytDMeokzcgQIyRFYfweME6hzGWnGjAEgQGSi/QwRa4mVJMEzfR9PpcqoBHr
4r+fro81ehXrcXcnVRcOb+e9FrEq1hlD8vu6ia1TPIJMCdkopHNnA4TqIa9m7XJm
1nwlBWaRpRzdvbtvjkOPynsIfFdo3iQENpXYLIFjgavlpZCs12OEXY0gy8ke2XVh
Saf6099wkIR4iky3FyBe+KpPlcGQw48GsaGxGPzySKvSepMN/uOR4Z99vEcUL5ka
kSINyLqrPqV/5YEgprVZWOe6mKbMbJPjcASKf+PkthT994LDO+epsIH7CtJjNXYe
u9gShIBHexY8k6CYtZT5Cc6ny2e65jtXAAv2h1y8eBI67JoKt3JugvdFLZZsrVPt
jEi8fGxtPw869XXcsrn2mEW2xtpHFCOfaa6mhlU90HJK6YWi50423SlogSkRlSgm
pfbsjTMkxdU+32FKdFXVkLcOnEtFYEA83ahSrU0HJovpRxBQDznbbdayILdn9tpI
8MusO0tzof2wbi/tTKbqA87er4Z0tu9PMUxlAJwkWfv3fC9JJ3tRsnPEHrzzhNh5
yVZeCI+3UKyhsR6CCtGjiBrx3qkJMWobjELn9FtyVHYj6qrjluLsmtg3Qo77g0fo
OAw4nnUadVvMPCbeSMUR4bAme5acyOaHj0BB/CchB/uKo75oj26yZFI0rwve7FXW
1UzOpv/BACWodrQrdYm14We/DExDSa36uAHNMKxWlZVgXqeBlJkVgVz22ZjB2N+I
gPR8nkjxQppMBEUlLk4dPXq53NfJFoXeMpbJUbAbx36qGKtsxxEQo7/6hFZYgnlG
z3oQTbG9oH0tw62Z5+0nkGrik98Roe3/e1gWG+0mv3UdSxGklBAvhpYGJbJhYcdg
7bdtzMbGMx1I0dNWYuxhSbIUDidDuRYNg+EAR+s1MJal68K1DaJ9dA1r8ynLCqli
OEwcJHtzzfnNbe8rO3P10PYk/veUu4tL114nH/RVH0FqiJFHqDnl2Pnb9Jxo1uCe
2p5j4arZiEvmgxW0XtGLMtZ+TIY+5Y5TJ2E9nRVWzNUk1dGe1HqTMYCggWYMSBFd
L3Qy2KuN03g+JELYELKi+/LiqA20xi9OynYxF0MhqKsIw5uZr9+0JIAhWA8eBLKj
dnvbYp1fcdm7Qv99v8A/eqg2m8aJ0G0QKKZRbZuDkoQdt+0UeHIFHhYhYjpcidAg
k+x9KQ/4w+MKXVZrOyMNmysvVuDrmE9EFUBXNOIW5VQfOas5U1rKLmxhvCQ8WOKY
6crdtxaqSYE63X7gLRz0x7YlhZaC6Zmv9G5eI0jCyUPVAgWnJ6eU25vs31fsfRi1
WC9i4ubAAwETP5AcXBdB97Zv9/KWPtYqeiAP6p9Psb+6vX3WHefpbffYWurYRMKv
IxidGKiogWYTGj6Y7Lj935fXnwzLl7ThRXREN1vykD64h/hW9StVVVXb9SlAtDiD
P0a0hOwsDXQXkKRnACyKYhumVLepaoRFuhrneNyiTHdoMZcUwBURncbYFd/4K8yi
YEY+xIoJ9teLMH1j2Xlro4x9+tEQWU+rC08FexccyGXjEEFza9QCXzso9UfpQxql
4VhW/1k7ofOj53DA4vcaGlH1SPWQgLOz13aEfbdCesdNphdacXbk7QaoO/SAwl/B
C2gaIHHLqNzbpPOP2Be6m3GZ5IIQTP3laQrkNtdFNPXOpfnmsYEgU03MNuJoLKdu
P3TDJW4YzEdgwGljq7RELhte1/H9NoeESQajBkVHwyBB3AHowCrR335AMYrPEzlD
nV655qgrk8s21c+5NgJMMa9Tc103nzfXi6/nuGrO5ZjKXYYkJi4W9dbJJpM4UCSx
fHln7wyQlgXKOX14RfSwYJ5MFD49CqkXAGKbeaucDH6dLa8AouiBzQ02s2sTvOZG
fQtWmvwyYlzjR7qDQ4cC6WTDk/Ha1H7wKXf9WCqKLA14O4k4cVBeMsYYvSseET+C
tDAuCMj6d90ek+c6AjbjMcpvOMBZzQtprZEwyMMau4H/vNxkRkuUet9YAOA+S1MS
jAbL6LZa93k/UvweePULsNKtbRVWTFYPtKzCTTzXG9SV/gqCdTWNIMQT9m8i1oPy
YCUkHLRmcIiapndX5DYesAVn01igoj990DoBx9nzsrKIGpSO/V0msq7kxbo7gH1C
L6XLSw1LOZYlXPGHMcdeaszGytCMe0upA5htHLDPSqzII9iH6YVfET1J2tAHt+yc
`protect END_PROTECTED
