`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o253xMCU8sdA4xsU5i7PIIru6OX9XgDh5yWZJNGjokgqIpmTiEbHu5nwREc8uVK0
INIVoQo8CTzUxQof4F7R4YceVrCrJNJsYV6/TGxcSORfZ9Kjbz16RhKZmZORGin6
82YgDfWkYTkh8DktrdoCrr5WobNMDZZ1avDRdT5GSWPF8RnOVSj0JEK1TBMcB24X
B117h1NBzle8tqxtwco3xrbPOhYr18o5m5BDjQHscMLwxiNVVqJWvtIzO8IFz6Z8
QO9ZDk/zqY9CiVL0I90svNj78JEGcv1XpPJOh6GYKyr1SQrmd3sjCsSFoz0zUbI6
B2rqxWiKFFhMJVROZWH41H7pTy49W1cuSVt6WLOGGcwqZeODMFMriJrOFA4qvqzg
kNT4Cd1FQE5FU3WqNvRO5PgLlN895C8NLmxxZKGhsby7kpOqlkE/00e8MENDSo/f
81Bu+e66IXaVxi6DYEQXYDJfmXSe5bjVmsXOU+y29Cy9nNVz61nRE3/UU69i2rHY
oZBEpTzvMs2tu1TwslBx+CwHYQzQs9Gt0JcO7x+7MLr4h4tgFFlRcUzUfPrrt40H
y8uUqpSJRzIgfKjxa4vsgtQfxL/Qw8E+bEpiofdZ+9GGLLu9FH2CIOf2onXs6w1Y
GVn8dhEVY4t/+ff4EeuK6aKZTHUXHPo2glb6jAuL9GAdDdD6dIcjo83cQSheaZTk
vh/8ClNEG2NDipkSbVMPnGqXcLGPeIM9yabOVPh7cMukITQbTF6ovV/KgK3uY8BS
aQ7uXTae8ZUdvLu58RdWWZZvlRpXCS3wxcUMd7sYb8gvykJpguwL7EK06wKGIJ75
9w4Fw0yMRhUIw0Ejoz1JLRY6vm2Q8z7sfdqeSw0yyvGvvOff/q+EjDeNIoqNGcLR
iEOs9NVl5Nrj23EkltfaEKD1fEbq4Ela4c7MQDT0yhHUlPjdP7Hiu5AMD8Ndh2qk
EzGilwAhL6xt8x7+F52fTFYp5de1J+Z/Vprzf/CKiKjdXU2dqYGzyz8/Qi+Jo0Lj
xKxHsWAlXfvWRIQfwJXHiumpRMiMeup8h72KZFsZsGFfsyVCbTiKKoojIwkxNC/L
Sf/9Tiddtcqcr7XaXOBN8G5m7rPQ/zc0AEhyAomHcetCsoyvHKuJA/P0sl79ZsuU
rhjg4GB0PGc/yti3fxEAeUaxFNoiHSN8Ko/1mv4VOdsKBpTNc1JU0OWzyeoFqihi
0zGSvYWJX2Mzat/O8lincvhecLavBGZR9jsYNBXOjNuHPqqSyL4ymbop0AJ6ZAEJ
+snB9YEPeXyY+OQp+5zQfd7g4SKFH/vE4Uj/TJyuym2ikaqrg9SWMxYv8lBe1F0P
tNOb9e+VDwly7CTkITzfMlkPtfSIntl0rrnemebSMDUJsQJoVNhX0Be2DN/JUYDB
5r2uno8sUvr7LsgptV6iCZo4SrnOXfl5w6403omRVtDub6yFZvIOTh96DXOmbxqa
7G47Hoa6f9L+offcqd8QqKC8KQtqy7IFvo2bl1e4vkjhq4plLvnme0Ms86p7QbSy
UxDQ4FDiVUN0PWoVnZHDF1bAUxyVeTkAZ9leBSUJxPYLmdyg3LbgKA0Bc5QEha33
yqmnZ7S4R/srqNF2hPr/IL4x7BnacutA5DrSxYkPU1nJ1hLThGIdkcxFzptfNLDi
4OX7LaJAmqnGggi0OefHa8KCE/ErEB729cp+NA69IHqS+C5mtbUyrpAZLibwZJs0
MJqdVcGkaN3DDuKEqOjikgNaJ7/PKcB5t7xofMmRlffyMWfwwDMONGHhgGYLkg7L
+GWYTv5Dku+he3VQWDYFDDFYTkCAFyhC49+TumkBw6jHGw5CmDplWdSi3TvRyuH1
Xl6iSVqKxztPV9Wi4GaSQmHFUbIp3ldGnvUOzIwqMAewM8Vu/x/Hh7+JoeeDn8va
5UyRpwPtu34rjeM9ZaqanYCVKg1ccetwAwFp0GsmQTnzJneyMeGLxqJ/oUGWuBCU
Tz5XbFAI9VlQQTeHtN+a12OF0mYWpP3pMw5qP5onWYflMyedbFuEgli2XXxAQYnm
rNZyKqlygmf2RGIfB0eTgOlw9N7Uj4p1ATMe7TfDmFmJ7DOCJ3kSsU48atXfyica
mFwmtyL+Zh3fdxD6fyKV7NWLDYe3Z74fFYCgOTKy+gsnwHWNxVW+kH7CIzt+dC1H
y1Q5w8WC+qWG4qOHGPL1JP8BY6Ll7zkb4ohbAZxQD8gOz1mi+imIWgVvJRzVuElc
/6me8+XlpUjqiVNNOh+PCwv+dfo3nBKt4OoIQ8hDVekXShJ7XtMATSLEZy3mMn33
A2xSERFROsMXlSUYqcpVYF9AUnNFDJhoHwR8gxNrS9kI5NA2DjBXoycVHOz3R/oc
V0sh/osgg1zH9LQs/S/E3nqMKSlTHqNF+c90jebS2aB7w+b7LO/fZEGJcOERU+N3
JSVD/6PYfpLUj4LlsMjmBdbIFMlEOYsCfRog3fG+WsVFFDSAXhvHPlOeriNRmTKU
Zqg2tYvUhVix5VDx6praETkOTRr2/HPuLzwC1s1Esxu7ZAq3EvwvZkKyburwzjoz
585ydzBTrlH/FtY4SbdBJZXEbU9Zu0rPt3b0XYgukQ8BOErQz3JHYViWsCXZcv/B
K3i8cOPBYw8tW43rknVE08dolrXE7mP4gJ3DlVgWeW1J80E66nFoJDPwtv4qCRMv
vE7DcnZTxM3J/ShZVnv9KAw4gz8iLnFv8w7jFHXFugiYfk0rOzvqI4USoOtqgm17
DaFkKz1BDdsOD5kKixygbFuL1F+xoT/3uk+ITCxpqDlR5WqASXETI4GK1OSk2g3A
f0J7PVwgQQLoNm1QSdWWZsjdluRVQ2SrwfRaOJK/ea4qdI4rkXSAyyItC0GW4b0x
b+NEgJHJScmUfZRt6xtV43DbkSsC8Ym4kKGZ7Q+mQUi06fg2zNUZjlPcF1QA1slX
vjf9oiSr0UoLjBofsRqQ58iu1MXjoCfgQ4A+3N/7nNn46Mr9++bPlz5a3jJQf9fC
YOG7PbBGhvvZHve/OW6yedKatRlCQsUmvF/YGgUVbhYHGohqrZ804UMWVG0r3fNw
mu5BXYsavOvT9Z/+pFYLa4aOg4ubxfcpo7sFvYQFOafCS8WiPiM81+0K/70T4Arg
OsyqfR1rcECYqhlI7l9gSm0qQ4MhTcwaYoTbPwRb76pJB+KtSkeImHlWkXuWbNib
BeXqUG7W+ijWXmAh8yGytd7xVJPNq0cZTQ3T9ieAwTxmN+vssvWnE8LoBMIZjCCF
Sua2pEe5GQ6qXRrdjVzhdXFaGXM/3Be+xoanhMzwAVogZeX1GaA9gc6eCWBX/5dQ
HOpsnGiLB6oKeTJwlDQC5piqYgMsJ42UZi8PY9OsVKBVznKvXXAhi6mK1QbtFgu3
/wvlXYTq61+FlrjraUSRw2fvooZMUrg3/R1d2XqS2gnGWMj5S9Y6x5vQw6Hw5dFW
Tr55ydTKdh+9s+fYltcfJqBVZym8QOeaK3Z1ekeFU6Dv9W1yYGMZA5roSeoHEBAf
Fr/ns0Cpi9zRNSl/KHyA4zQ8gfeswHmVLTZVwBrONBvHkhO4yrXoOMqUqEk5Ob0q
VvfRttbSdLsoenveQJbV2kXQdgrG6RwJs7Currp9FGrdaQG6E7QqjdMASeFY/GIY
KiZtSAs7eLx+NkiwBgheoF6wyy5LaAonx4CsAY0q9X/iho/W19F6EdZqSQWZ3tpP
VdN8VQmc/ONGTGSuLX2y6a2zUfgIPs1z5RtNTZ/yraLXgKOzQcQ33rGAxN6WLste
GoHwQF/9i7WpNRhSuOWux5ylz5ZebpC3QEvgHhjyfEfUSu3BLGVjTTrWAVgKLAxh
DJgEshNSnLrugR4hq+x2HWi2TcWe68+nSfFLwNMZnKjH68z9fxOhOJuBvZ8jcx3B
XXstGlWdm/6cKbWB3SjA6CXdTwURPkUtrdNbADFrDBDn9QJD25rRbEu6gwhlyg61
nY8psvC/DfNlRCeIpQzlTcJkdlXOqM3HFNQFRGkoBt8SUc29T5MUDSbu76Y17pjb
jehFzWb68mDNbgsxXnbu0dcK1hbW5hRDMArLPJ4AT29NOZ/sd3KVH9b9i6oykMHF
g6b5jhr/93asATanAGWaHRO39HqXwQR0V3bBVDs7pMbisFGqN239BeUFRAcvHUfx
ZHIzZZ/b+cAoTAdKWh0BKrwZpE3iYMGuoHBG2BgsAnXOVoH/knzkaAdXia1C8bq2
Zg4k0TaqgSPq/UM9LIw2NWuhYe1IC6r9QpRoZHnd+zt3NM3QHhCNzG1HjHNReDj7
8nFxTE7J42c5/LoJtwqlSwjOgZUDcovehuTnrzp7jSOmwc7FpYEUlmaFaIJ2bP8X
N6TTIpuHcD497O8q3vzRS87KMUnqJS+OcKHMnQC7AHKMwP/WTCbA7ofikurZ1geh
2Qe+1x13zjLmr7OGEIaKxJtBqgYdvDPyhEk64bt13SKEuA1Xf5e+utWAcdIyn7lx
71BpmcqWGLhB5vRg29CXbcQ8vLgBpBmw1YpEpg2wgbJ/29PQXFfzdzq7u1bfuiHf
PTTQc+3OIf+Aek31x6GCyYfUslHThAkowQ8jQmm4ovfmq46u56zwbG9VhGKKk4yC
Vb70+3eLGQPrpgPWtX4RIU7l/UynpFVz1gLrPB8CwGyQ33cCAKx+ENokFrtLscQA
Rloi7bsDHCz6BwRiN4fy3FSxP/Q82Di9ejgX60OuHKbWnh2GYhjMiS5feiW+xYAe
IkykGDJjZ+sX2UcYX9a/wZwBTb9oogq3WJEVhRF0aVgwHXhKtGkGNjNvGFvhNgS3
3VropLJ86fQU4Liu25TsqH1yt6B6ionEpk0bOLCuYlCMnGEwmxo3j4eQ74IyFLbo
AlzqiZKvlxTZrzR9q20EhTaEkv7Wcw+abShnqWUw1sX5gqbk2F5k5uCVolXmBnWd
Ou6qCRZpFV7oV9enCFIoeQbPks7/xffzVM1reCSWIQbJqb1pWQ5kDMYbkzkKhoLk
RZUKmVmryXSC7ZnwXDAEHMXqfgkWLiJGB1k0d0u1/x+WHrESmm1vaDDl9bHnTQSI
FtwANDKRdgZd6cAF8KlsxRb4HH1MAXVhIUeoOEa09ixaUnledCD/h9yugAw9F9jQ
vhPLUmusGZQX2S2wkSkK6LrvM1NPh9maTXxVsXfaUpEvt8KjbP/VVUJ9shVszahx
KCSUv0mfo/KH/qIB4OHvAe+qEAVf7GUQ4KR6TCtmygPYJRvhFvGie1D0LCaRmusH
zTC9wb0UcKPBIy230xy1it5FFkzig99Ixwqqqa4Qc1EFMe5ey67fc6sWnf/pDF7h
zxBH3G6uFE3OXQrM3yXTq7g/j1o/c419cjUkHyVPUFLTowTrhL14bszRc46Rmdyl
FfOHh66qJRMNlSKejeTgqwsZyzLo/TILnig2iY5KjyqhNQdjb2lbouvihcv9hOUz
NIJi5RgsxTcdx3hziGKmrFJWIGdPcM9y/6e82R1FPH45T2lwyrYgDxj2U4Uq3Qjd
pNfUH79LHLPqnRlY3CJwkvWKb4O/g7KdMDrlz7LO97Wek7ah6ws3U0+wKqhucQkn
V5EHajngngbRmE5zfD03mzApUUzXfwaNsM/athZJ2VqiUYgRww+iZbdwjHor5QVr
Ou8DQraCvGFugRHuPjNGm6xWEDJZ2dEbGxmqZqUBcJh3KVqmmQOVxxhRGJuqc3up
ITF5bkLwU8mIHu3GA262Z2NzgsAtWEiSRZako9M/mHDZG31LjwziQUvlJnc29Eoh
NdR6dEgi91drAVGUUuYJ0Sna+fe2YHwL/BDsq0qWOpYMm+/LUpOw/sJNWA7mhdxQ
wEnBIj8GaNWGHnEk6nIlTdSxQYv63lWDRr2ylyaC/EtPZoDxYl1XA9IchhbFP555
btOJ9T8dOrmezROUOTq49uHfJWEIBXgS6sNCUlisf4ZtM9Fh8Vz/ByjRbFG0w5Z6
59pmRutoi6zSYVzYJXwkAItjFBJjbRTdA6hlINmm5TH/5WSYpr/5JL+jcGYSsHSF
9AZOdY1GB2fxiCUW4ChmRgnjI0thgtt37HCs6dymEOQqCdMqtEnHSuTQgytLXv1e
t0HpkeCQ4faGAUgEeA6dj6umIbBnt6R3VMV0py8HHH82xgL8sH9dC+oba+fL+Kcx
RqIW7ReknvtQC6FZTBfdnlX3aSuEeJLYGVp0epJoUjnndR1osizP1Ba9POvKm6JP
drEe+3Dy34mLHX2y+9Tnnm5WsSOWUKdp8xdOu91hlIANizfhTQOak5voLNc0wLhU
gLYqi6jdovsoZPjSHBsZ2SJkJsyVXIQhUeLe8FETbpqg54bQmupXSpRRU5R50spD
Nd9VnqQ1P7vYpI+aw92io1nt0F/JpZ5GUYm1XvfqMJXft+Cz7AoM3akr6PxAInU4
etW3960dP6Co1Eqj2xYD88skEBCud+zF3GdQkhGuIrrjx5Dy0FIO1Kv6FwftjgfU
87WhltDzPUNXD4zh6E29SkPZYYdsMW75mmlKucycdOChhjQ8BmWO3yKtxQos1S2Z
Cz0XnSCEX/JKAt4wZNOo4U2Bf6EhbaeBDI+iYpsw/+snKZS6G5vWhjM0KShRsu1u
0xF8jNNYGNGwCNSD6+0RBwJYXIw6cBxcSksOoGH+BToG2O4cEjGm3S6ciustA8si
xNBDJx7tf/KXb++IOeNxjUhsvWfctBuyUImGPLzm7QJkLyJVixLjEoC4tlN/NkSs
z8MUJo3FsLf9yydpDBUt7gOOVOvmXPFtLFsaRTilRa95sQE+2mLOxmbqHAjHzHW2
h9HcWjxG7VsKDNt458Pw8Dzt3cQEw9CGZGjO/H9fRlEVSWFAM312+FLrd99SdQ3k
serpA82bQZakEWm1+QT8XQt9hnbrv4Csl4vDolrl6lBw2gsnmL6WDmEPIcBS7ofD
I1RRg+PtaIbd4jlLWNDSj1Vp6DRaoq9HBAzQmhGZXxz0zMbeqzAVAszOXHiIWSZC
uOZtyCg13NoBKciqfLcsHosBQLvC2O7mLwGACzxfxPejp9TZCFuBJpVluERC90N2
2PRP4SO2t80S2Gqc2VuR739t+vsrIpKAJgJU03I0F/jbtruu+0V6AtI3jvVh7u2h
htGl0sEAZu+1VV9zadZ5Vab8zMu4XLb73YuqsPYN0RW9i3/zWgo+SS1YxYMdyZf7
L8h1wwn3BcLXNXrDSfOOmU0JbOkEsSlpuQ23jxHwWcBwt+5TxsxzUwFlJLuMtH4B
pn2OWMj2CvVUS3tvs1t1xFCY5r5rcXPe/SsYj+/4Z7dgZ2BCM86kOCtm7cMitDdh
zY+zVQ/UGD/z6TG3uQCBR5tTVqQv/4b1HZbo6APjx2UMQwT4tHj/YAPYbYNo1hUB
JJTMrhpWVqj2lxpoDdE9caBi8a7Z2jlj8DPdXWVrfmV+MAhsFbsDqJqoZEP4OTmk
vEAZ9OOrG9FdjOlpZUzLDCwj9ttGiclVSMDGXB/s8EZV6wbiSMhSvynvxqIyta8e
e8dLVF7uaB+89YuqIbo4JNb8YIX123ZdElg48bTZcXUscnmnOxObtq1gV+EiPxXV
Yjfeo1B6uYgxm2rCnC0s1vGbnsk23yGytXohPOB1OkQCYzXj7FpdU33SL/mNE3iL
szPTCiAD8LT+FL3q2Nwfces+K/NW9KQ6OLOSSZSQMIvbxPuy+Ioh/f7pYAU4slyF
bVpbDfTqWCLFhj78KRMWkFWFkoY/cnsadGfIJl+hoWtdj8/bS8yi+28bIlM9rLEf
B9NQfH50/uUAD1wqGvN3cFoGFCrXjjo/D7t585wzFJcehUB5aejgMot2Q00Psx5r
e4mFurOpwOlF3opiEr8UkoBQ1yiywUR9qI9au/utWK36YNVgaPJckhfjiWqaF5HV
PUPzunKp0SEbxZRoVtzbX9JYnWvwXY/dvl9P5I/+e2NHlZihCpZt/yvwY89hx+1E
jr5A0uTI3jZT3oqYCZT5WebPZivzyd3PGzZRLQZg4NCQsdb9Jl4Ru39Gxj04gRWO
VxVgagMB5j9MfRvC+A6VmdACX/dfPCGw8lPEuewH2eWLWrJ7DAd5xkEaLpZz/cso
Au0LGzvY98I3yx7R7J2HmcjdbmJjc7y+2+y27ucnRgwcjFnWik/CXlLd/zp7qvzA
Csd7oRQ/oHY34DMIJsZy6JPWzvDsddJItd8C5fGY+ZbxSMHtswFcrVVGpl6dnP5G
8EOUUu6QtQE5ElSOj0wzBg6LW/WJ7DgXbEOzqImjO9yuMz0/PVGrAuRkreXbRM9n
2eyG/n1ROXy8jk1Yh1rD0D4rm/YTaxkXca+XvhP+jT/pUiHjWmq88hxM/2+sxBo6
pYIxjoOA58MCvGITMRv9oBh1VHT8C5UQPy8yi03/OA4opyvVvrFF/bI/t4bCq48C
EhBSxHbCmvix5lzcv+Sr3TSl9PLp6MCcK6zsmbnOm/iL4vkbVWCoDR6Woi70Ru4p
t7LF6S1F+E+a1CqcDmmWqjEfbE/O9+D0wbg7fxDjUW0mNGo+zvrTPWWRCtcGIaMO
PBJbodHtN5l5H/wSzyKS3AcA1nRAyI827riAnKaPpCS4NwODFrszbpjMbf1hHMGC
barY3VClznW7+MLInvkXk7olsxvRQF9xKV963CBbxjuodRzmEldqkERGyl4esOc2
Wcz2zFMAKrdtfub8Bq8hscZMRVwrOIPikBJiY9sNkiA0gOIX8wAnNaK+vhdv4dEp
M4XXIKvXCu/wXPxNlXAC+sMcoJnutXnYvw9KKE1UJ39OhV4zupHHOnI2c0PxF6WM
FKjrrkklLXbgYKj19v5u+62zDkAsNrQ/l+/rrszlIkNETdPoTJt9fL+sK6RzQkel
dzvmrXV3ZuBCpZfGeQpr4uQnpUypdzaaHbFBOpl1aIjgVTp0NsrrsARCMhXAhU5w
9J+X5J8FSEnkX0tIgPopA4ByUbBEeWmHNBxh07a55Y+UJGfkWuyEanMP4VSK18y8
WVVFfek1tDAlZC3D3ULTcBpiebSXJd76rdYBpsvmG6hQEN+0ZuXfXNQjRAZC4sfL
jMbfMlbgPqGpillxCvoAJkM1Q9u8p8Be44lfFFB/+oTW2ODU3DUuMQJHivLfm9Ba
2OvTCzGkedvPmjw/Yn/YgHbV0CX0X9vEZ3GbyCz+l2gqcv71ZeTbkZS1m8/9gjHP
OxPJykc3NmB8CzSN8wR5uTkgedWq6wEcb6pVM2HW4XOoyF3h/EtaiPOrrx0+n6gY
hKb7AHTmoS5caAbzuOek5rah7cEgjHBTCGyXCMYD6si5KHxZZmnj25zBlo5RjlAF
NFRfMHnk46ssHQ3POyBypXvU2xSjRvP4CXgQ58Jr4n8CN+t/VHCgHLL3JBsdre8P
fQgWf6qu2MxKVClIH5k2RchRUDC81wxf3n1x8xQ0Q3gyhbBdaY9XhqXVQvaooGFy
0T39dMWBl8PJEuXy9l92MfnIwoxbxtsW6SOsveLkn8UJDRZnP8bxZiw17tj04XXm
FZ1VGpixfZa+wC0RcVm5DEXhCXm0PtoVG6O5ZsuRnhuGV70IvZYiRe5kDOCqy5Jg
tA9cp9Pw1jfFy/UkEdx7jMSviKpgs2DNHnmzMOTVo/qLsxYaxT8K6IQ3q/ur1edv
C0swIZHpkwhM1CEeJyEAfBKYDQO3MB3LSzPKAQpED4YY0mfS+wAAXaOfixQhbdo3
I58bgHuOnlysEDJiBLw9C3tIE/3mb9MdPy0IEiFyDDFU8LtjywYiBnvZN2zGIrJd
2Mo5Ke92Zei+XdZz0dj6u1A0AtHLgScDDyHM4IT9zYKnQZtA8m0FwDiXgJi1t0Yn
ohgAr9lp8y/DRQyPy6Ehu3zfb6nrzDS2O7bC7XSqjWWO1M/clZocseYMYcr/AV4O
TEs2PHVsIPsCP+rVfKHsPC38v2Av/8HgE42qe1DNurh3Le9eVMUj1HInNH7zkE6H
gIpkO+lPn6O+Fv9+T9mk/VyNcvPGpdoJ98Gp3/eJ5dsw2rZlo8VuRrzJe9dHgPyu
hPjDKR5PRQAfFYNmWrIqmxZIWxMpIFg3NW7I2cDLoZqG3yvuozhjrK2zzHt2McMi
/8DnG5Rn0D5vDXN9/U/y9ipUtyAKOBh/bYhModcHJ29gdw6Le2SNSrmtYcyqPfLy
ebdCNx8U/X/j2E2G78qj3mlLc3SEJSXR7ym9IQgnIXqLw/5QpNxQSF2l+9+4m+46
vykUtDaQPwffR1KCDG9e+SvctsYrjKxMOCMStncPex+ded+nBYqrw2Zhn2Rn65kt
QIYOUS7wNW/DSWMd+JqPPf6KBMR6XsrspiPbvjmIlu8DQ+rAMFA0maf2DdhI4opa
XSh0fz6haerxLXILWVq1Ujy2JwHP6okJ3pXGxkEVjJOALu0kIfSkQICwwF6iYH2B
KbMtrg2Mcb6LvnpLOHPqbvr4+iq30w/dfUbXJfzhcPsdee0sje++neltrEGF4ULb
R8/EfEFAf8HLhxfEAJkgg6J6bi0fI4e0CdFEb1J9grkRwu2/GnRqATYtkWf40mZ/
65W851s4qseuLoTSGu/N6hhpPmX0wLhMZM6ut3P1iBI4pMrb52Q/Guv0EcHISkSe
ohIDhXWqKfr9lCmgPtOEyQcxVnMfhpkCiFkCqzPPUFb/OmcaG1VT0I001S7fzOL1
BII41sruD8Cap2wbagRF6cuN40Z6Z2ty3O+cPtuSe7Tk/GPLfmm9bmcv42pMDvdM
PXPMCNVscJWbP0rIz2SrBeQHj6LGjcFvWU3bzwQ2weF9YmboMCLRFbybz9XQ2guH
N7LqDejhYhYBN3qESojEnv5uF120oiOzpKTk78mBie3U06f+ks58ivxl3eH1p6Jk
vCLyCyxmYgMks/yWVKhACbWuXm6uYbTtEXM8pq3bk3csSCl1dR1vlQF1BgfSerea
L3wT0JEnSBUNVjHYXlgppcmPqMj706uvcbyz1iXuyHJ2DV4mCTqnxguumb9x4Wms
yqbH036XnHWJ3nGIxXc8AKmj+v2WOVtjUyzjPkK4b6C+C2ctsV4J1i5qJz7THLPd
zy+WSdjH/qI+Q8W2VMvJtseFARhd2WJUzKd6ccEVY1V8Q6tiwba8LXi6OGcjybLP
Wnqgy6qfG9VVacqGbirtayqFh6o6xoOvNle8gcvcw+XZo5NUT1/eygaUjwZezBaK
3pKcPXSREP4knwUBuwaSp7iig45ciW20g6M5F4qQzsEM/ZmfyKMR9HNyy90ilr7+
HflzTDpmdPtB3Y+wy2dzHN+59tg7+DvHxnvGLdRzHxfpYj657xacv+oOJGITrEuw
kZy6z+Zp8mUkLIZdxTP0dAbXhuA1iaN5Tuwit6Vl70zYYtCDhyBboCtLpiSBexc5
WwYWEuDRBf+BySbFwjJEn1HgaVMBJ4G0H2lLWbcX3OwFfJab/7o20PxUoYcDLiBO
yIMjpco1pz1LB1vNmzN73A49oifEdFfIxas7WfzbrCjOMOTUux0jM1pEKFpQwd8S
oppV0l72vp/iGKtINTaYyEa2BDwiRZLuXTO25xv5Q9C7bEU/fsAZ1Dw+MevANAx7
a9oa2N9B01NnujVZyNqflGQt/4FtqBDu41VPfCAcSU91t6yEcSeVexO3IOzQf/W9
Wo6azKWxmxWMNPUt/h1uuz0OemSEROji8bJ7alwcCoiJgcKGp2dvFAWW12365plD
A3xCiOwNzyuGYZ4y7VSu0OcHdMlxqsOO0Duvv+Kxu+vdLJzviAbZFc1n8mE/hf5D
SP/MmmCRMfpBEojS0aW4AnDhpvdjlqFnZNNAP/OvJCkjySP5qT0axwJ8Dxy0+GXc
/NTghKrh8A/7vmQIU2Z30znXvCrR9eDQKV8f6EHQw/y4kST055zKMXqAlERpdOiQ
2N3Mn+7tz2MISJ2lcNJXkfaohlvUJROMa8FPRnrfKxbRWfixMDOxGFycgNrXbw7T
WiNqObb4ByWnbeFPGKU5siyURbUIbJorCEg+DoXGjqJzzO9wbA8qGx9d1mndtxsY
wh3uEBPeg6R/z3B4nf7L0WC/8VoEXU9tCiK0f8bZ5StUxvhILyoJb7bbLHqxCHgy
loR8p7wgT6s9+kfCo49tHqjiez7I464Rc5hYv/Q2wcVUEcj3KcxFn9H74H1Blrcd
0s4ya3eh1Wgr0BAZXsL/ZPCq9F3CGLlUYSOBh/6PJwY8gYdX5Zb6yWLCg8i1VxOd
m6sgxt/nhxSxbmzEsHMO9+V3FHPwRAo3W18mjP4Iij28JON5rYfpFgqL0NPKeEU9
6eUWly8QvskjAas/BLVDrY3eWq9FVYumj2H97F+C+3BFjbD13lVeflBJFtD8o3yi
8scp5HKyDLyJTOkLc7oC0LolyeIQMlMN0jRczaofR4qnVSKDybUgPwItfSLDSQ9g
hb8p7MOgHaYZrZrEvH+mg/DTkoyUiAZnfRwk1q0hWX1dW/COoMsaubr5Iz0xZZfT
CDExpWv+w8Ghgoh5bJYf1s6080BVdDz+BSrayjzx0vF2SkUAUCka3uW2fM+CQqbX
OUYx6ojeC7xJ9pMe5gRGsxJOXr0vbNL77Z8SvHQlYOWAKQRB3mgd1OlcaUSgY1AR
KrhB5I0arIxlcfFDeEarDnOKkCPQyX9/fISSeCIQeQZc6ValQDRIKSeGIUT6tjIe
0y9l5teb5GJSOyUk1A0SPsfDPf2HUrvxTbm4PQtDCMwAqanJtbqF5xwtlrxNXR37
wlDhUcZXtCyu1AlKK7XddiCdbYEutgBKdWeymidkTtmFRJK8z2AFpiX9Z5D3I5z8
pOJZ/JN1BUpN8cMW7MtNwGIc1FCg/EgIQ2PkiSm2P/0sqYS2ms2sgqxkcx1YmC6c
hHdd5ZlvctbrDZSgZwsgUvADCQKiIGzpNy+2Yx/BXpFa28jhYE3YRFS575ik9RDv
TETODNGJ/W+mkVge0Ld8UsJchm6MSkAY4OiMOWNBv7cY84gB+/YNLAVaV+7gGj7+
+iBDooWkDnY1Gs1jk7f5qj61ch3zu0fdR2C2kjdKaICaGkvnXv5MsW/t7pbHSwj/
BtIduMbFoohYfDLYYYJu5uuxGnO99KO7YKGnNfXoZpO9pvLLtD6smo1OBOmktxu2
rgv1x1bNiQf77FlT6iR7NMQAuPGVrMap7YeHTpYyhLbDaBIGHuFdtKB6FzKnzIwQ
Q3it0oCg2VJa/o0sL7q/W1YqNXj4dL+8QHjb1WMilUERzwiPGsvdoX5DIfO8/N5V
VKfhvzz2vfWG8ShowGeIesVrDRMWvc8n7/L2d34PXEmoVlVzBEWg2qx9iqJgKLVO
haGsWmXAZ/ppDguvMnjmFdVd9xtZMk79/WL9/9ljb++E3Fek8hMc4GlGFIGApx6h
RqDrBNr4g4vv5AeUOW0QWZDyh6kUC1JqBA24jMnawxcg/598y31+wZSnb2XkxPEW
+IwlQvHqGZLioFBrRbcIMuhbTDsBr1lsxFc8wBfNH4Zo4fUWVzfG/FMp8lJe7C/9
tXDmVeGcYuKTODvS7jaZ7ao515rPImmVoJMNO9QQc1v8zXqGtemmOEZIFA1vrOAY
ZBO9JAXfIofL5+n2mRBzKSlGUo6bjuzXWMQGTvKpm6rOJf91Hd6cvXqsUsVPYarW
61o+yK2dfp3ReU1CtIfgP7etFu2Rv+0wBSfrP4VGQU35gantKKISSm+uHzVqu40l
mkoTw59B74mLpP2W3shTBA+Ln6VF6KOXKJrgnWGKuNQ2gOZhDvu8f6DbSXWfulBE
SVTsVYunoWIuYNTZCvvu9sO8sIC+tBuD5N1x5DfmRkA5lwJx/RW2YEIGsv+b6EyS
xZJDftE1AO9JjXB/XfDcCnL6lpnUTnAH6wzhhOrgZPjBJX6pFq+46lViEkpB39hW
74lDJzGlTMUn7vdExZ/HzN9iXUGRM8ZVQqbEWSK95f/D6/gszvegysvSpZxcUC4t
gw5MwQBypAiEuvYtyQwNZp4CYxyJJByeoxRARmEyJ5+g0Q/FJXtVPae0u2KCKaHu
ZESKhQqT5Nk3d4KQ+voIL4kbBCfDCyNmimuWBXZ4ean0KI6uVbwkFkaa0QV9QVY6
8iDf+4TyTfJxqbjx3TcDxp+vdEEHQAQTjZl3yT6HtqPuyGi5XabT5V7qSXlnEd7T
FcUAt31GPAl3To5JiL9oXb6XmDHkaUjD6iYGfGLqt6R5BdqZvDY3Dkgz7k/QEUth
cxJLQ2viLY8U5B/TtrKJ4rT0SFNhJexfG4hBsJfPo7WeYeBJtEiNk+0fVGRkwLry
bGfCnQXTg2CrVa6yC4bbYzquHWMFOXmZkRlauWzvE/kAN3KDyCo/pkRnFdyrtLWz
RDpwCHI3xC8YOps3D+ZHpwVliJ3ifFjracGa2oDmgYPnXXMgetzaE9OAVe5qVAuV
ii5AM5J4eAng86rP2AsXUj6KCD1VPGQhwd40uvv+T1j9435VVeY0LglAbHsQZtwk
YxeJ7UTmAk4vGp9wKjN5UqG6X1NXw1bPKGBt1Qqz4nY1PYhKm7/iCwil0rodLMfA
qhUy05gQlBCmHSbE6tfIutv4Wp7bZ9tYM08sH99Cb5y0DQCYOvdeYnQutoDgJ4od
gH1if5eVOVtTXHoPlJ7Huuto9pWXxvQg05FrVHBYZJd1QFa+rkXlSDfWPE/5vAKs
eWx/x4d8PTY0LIbu2d2K2i4X6FCSaFnbfFnaXHHJsDWvGkbo2aMlmksefaiF/7Ka
2yxpwpQpywVVaZotRzCE6asUuPmh5DDX62fw5PkqA4VBYNYBSGcXYaTJzlfauLNL
uahs5tl0FWxqeEvHz7Op4WlEWU775if+e189BZFMV3tGz7XAOq5zSnI7e9PQmzWu
kG4DdOakuEFTCAyB87afZr+RA/eeKexZlO61oY5ETb5x6lhfiorbqTbqR8TS1FsH
1ut/bUfggfMUpXAf8cwNwKk/58fUgFh/BPaibFFeskIMmUqd+hT+BlJ2ZZsFU1Ug
GnlzZ5Ji1w13wqjfO33ugEIgnyIp6Dj/O4yJ8dWRZDTy3LY9gnrItUDsuNG9sGM5
lme+2GtV9cAY9utd+dCdiUxmX9919nxbc7XJMQQAmmjXGaqd43vCLjwsE9UecyDJ
0+QBYz3iztZ7x/UIJeUYZbbU7OM/qt+GnQuYyHv6vc2WexR1OVubXWdQgvr2n/2J
ELfZyXKV57e/ONuGpqX26e8PKT+2pOeZxbm/gWxGLppPnrvypmZ0DFAllvMN/QJy
ay3D67AHz92W4yXmni8Jfvyxb9KLUjwRcteJd9sRBX6c0IrPCYq//xfh7ysnOPjd
gLuWq0xLzBmEyQTN01pcnsTlfUVW2tTC3Q9jlAGnCnf0laZOjgU8wm/+zxGIdrR0
1DtALY/hrkmFItf51e2nK3p1yS4aZu0hoq/bEo4WxyqpU6hrIUiPeq+tWSYlxNq6
Q/VO//JK7DhbLofmfL1XfS7pdSdVyIfCsZz7rpn0V7F7DNE/MfQ/1qqkSpP36cJd
o1Kq1fMVcOrSZlQy4qECVvj0jN7TUtdDZBDjdM1z9uBIaUkYvDtpjgPw6cP1DNhx
olGRgcpKmpvGPwLq4IwFzelfwsyzyKBvu/WPLg7+ip3m4qfgmX7avj6JLAADPZgm
u6aVyL/JBJGvZz+hiQzph8QgVSeBtf0s3lCP9u365XuaXCA0QS5jhVDbjZRNAaNg
so10bbYlzukh5OpKgICfH9MKHMdrSw2Q7aseAM+Hq5QHfiXOON+J33WBXfxUR+0Q
LA6UhuhBKL+c5dUXCpGJH3CQujY6NmFaNJ0GoTrBEuVenGFL6nfTvrNo4bEw7ANb
bKMjgitxRousTptekShOdyGhjp23hswujQF19jPajWef2N68Pzo4a4HTZfnOCca7
bKVoX3LlFxdag2mYn22GNfLtOhCIpTanSIo9YMzyO/uUH+PzUksEbVVK5EKwP3Uy
9UcTEW1nAA7q7AhvTW0C7far2SSVzswy4nJRUEiTLS0f8oOcjXZ17FQxDClG+tTC
YzWHpCg7YTp4MkaOkBEQaMx38XBE94fIQCgTueQexNuVs6FsYDwNOtyGi9Espc67
2XbI/FmBczzPzQM56DOvW8eqHx7qHUbpIfOZ1JHSRdkmPBFBCDn8kmVAywkMQGCX
aVgCoOLb0qNqp4JCjVrqQY/Qf/E/R27JAt9xzUQ5jQOfv34M6eCObB5cvEK75wOo
qvVQIrwaBt0Cu2eCcnajfPaD4nYJbw9oEP309RM3ZNJxGBf9cgsl/f1/QC+PsDlT
6yJWbg0pGzGu2GYTU7L2UbsSlSkiRxuJqZYH6jr1MhNXkFwly3yzE3JqiYVPvzQ6
z8ZRO9t8Bv3ejxU0uxbg2PiIxg0WIfdgvDB+Fu+9Ty8dPRrTnvhOPhd4xXZ21yWH
g3cE5dA4aqbvlOkk+EXmlrywAWLvzOV+QFxGuPLzrCHg87demsROpYRPKS9sLbam
2BULW5TzRi0AChNNvr3EFMkisYCs4b/NVKGxFg60xTZvEPlpifLnBY/EXoPqNLwK
HrhOVlFymkhSF098Jx5VkySRh0tA+SwLgQNqb1EhMZGSQO5ARpeVMFJyzXwnK42Q
vpAyxY2s2YwYkIL9vFl0Ew4S0o75C0I0IbvTdDaHkF2QpZpXCUWr/DeSWHrop6bj
wEJuQ8sA8L7pLEdAr1VR2E4fr9cXQyPpx8IzIWruukPJQd80gY3Aw7gP3KUr/s1y
BEZEYvQJ9jQJwfueaQvvFQN3VegEW72ZfzSIxKM2rbg=
`protect END_PROTECTED
