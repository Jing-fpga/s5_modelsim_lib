`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
64OKsehc1ZAi4cDUy1Ewjec6cuqzSJ3pMw67XYbkkKVyuZbOl0SgY4LwyHkDVY0l
qcQ//KVWbvZIJPC8POGlwx5cqF/4pyJSGngJ/gKFsJqialjQUQnzvQ0/u4hQUvgU
RkHHFMqYyVe/2cXW9j5pNKdVPXga+Il9oL4M8w87oOT0z33yiTmCnHWwS35WIwYQ
`protect END_PROTECTED
