`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BSiEhGa+O4Ozh+gxuBy97yYdve3mJZIqdRmlstus2Lfj5Y3JBtLbhsG69MXk3lec
aMbncXNy/9O2+WXEMzzmPsGEQaYa1rbjEdMBIDtG7H4+6EjKGGW1G2mMryw4+dQe
tywy7QjIoqgpLWJ3/kzcqyP4iEjeWV2/9DNV/NG164zz2s9hK4Ds2ze//h0+TGkB
kd4Dj3AQ3fYeC1PmDFAK2/aFGoKgvEbDr/FvVZOJh/BczHB9kK8WcinkfMiaW+fS
Q0Y8J63nJzK8C+8OToYRNHoCh3yUeHe9jWKih6QQBYC7EHAJ+8mVJMZ+4aLr/Q3w
sMzMIFAjhsf/pg2B+ACewYmjE60EQ5PfHo78Le5vi4yZl7JKCRWQO/U6qEZyyjbh
b0rKPdYTH4F6W9IE1sOgscZG3nb/69X0zQ/MPvKnsJ646Kv/xErHHQPdlM11MRA4
ilOAyoPk2ckLGofz9kLiFGNjI1XGs5n9R/xkIUgz1WFsC+776dnRM1/o7+lbHJZi
gdI4OYYHJjePg3YhtGz+usGda0mflcJ7lIV5RlHvfpCKRXYw5FBbbdV2BljwhCiS
PF0YgyWbQdGzlbjUdQPZTvTwuIicOuPIXTYUBme8wKW7b+3JucOzOPlqKteY97R8
QWiL+Xjm2s3GmF01o5J1DCrAyUcz+Cx8F/0P4ynI7nZJGwrHhwZVv/5tUxw6RaWE
D6I9jRsEMpozAIyA+FlKxuaejwLyXdET/kzyVffv+udLvHaMWiCi6r7bgCFlHcDy
tygoZfd18bkVXOFBGBBMvs9fCrYSGdMnQknR+9ZaM3ztta2uGAmb8H/P0FNv/6qu
sbFIKw3qM7vrVlcd5eFHdUzPLGNnK0BTFHnS6pC+NMHKVvpciGK+jUXTHGwiIDX0
eA4xUVTxkiDY3CbZ4l0zJDADwJIwjFmCyNtQXwG/Nx7Ol6Ujm1sKxopFT2ICqb6D
+tb3xT2PYE9GaiptbIaMyuTgY2mGHAryg3N6PK0ZVwBHL2s2v/0P3Pkxv4/z7ddI
+VJg6Mspai4mBXaiMyeO2LCasT3ald6dVxr1kX9W6MAY285vJuPuGNbNEz2uEJvZ
L7cR462y7XYpPjbV2IyOGBnUB6WCge5sYCyj8XGzyECRJVTwLaYciEsSDRgGzDgu
dQv3AUsj52R5h3tNUi3fiQXDWF1Cpir98uOX4aJpvgA3xnxgyLIxtGvxUVcudhT7
VSQ6v6JF7ey06YCue7o4XKCZV7XLExCgDFKVcL01zvA9ns4IXXNE457U5HUk73pR
2hkmGK2df1YcLEvWpMVJzfShRmZ5P841q5z4eBMxCFIy7x0PdtoW8yvZaNARv2wK
q6kd7DiSjpycQntH0qQQElDFvJspd6rMRiKgfzYtHPFkTuWyBCpbVq1cCgUw2KsV
Oeew2QC+WbQ4zU2nXirMuUQWxDvI30dQYyaRELz36n1on8RScjHTjd1HKQlGHhE7
EEVCjTP1SK/rLDp1IXHMZhem40qkkw+dhk2kjwDIJreHCY4CNwuyoba0snQa1T2P
8pBwpsIoYZDi9ivLpJTAsqVQTS3o+cNXFxFfyCkrC6miWq8H1d/Sv9u/gdF9ObDK
mI8or67igfPokXviXp/LvS6HNJ6CyYW08hzyUAZG5kyOcE0MP8SUekSTRsKmHwve
upF30yJAyhE9YBWpIpxM5TX/xvwu5jE4yUXD/NhAzxb5N8QFsboyHV6ixhCId7jV
ed2PhzKn3NRNWfOx6q3f/hBDACN9c0gQ9wlup22LU2Inva87oLgNZlbVfmogO3EG
BCSSG349eko3VNNBx1yv4F0FsPcjbcuCKoOEt/arNXMUumaAmpSkOCqSF5ngZfga
ffRUN3RGlk2HMfdvtfqQsuiLP6DAqZh6B5CfWfdfkEnNsrFnSqBcP71ppftRZtwu
RtzP0UAY2FmSJJAZPin6YKoXylIEglC4vyktBIW9eYjiyY6Y374Brz4Aqci2DJO0
Vtvdu1gjeQ53MkCmS/zoofckNMArCAeEvBfWMGK392gZN6esXsnwXSXNzv/1CRLE
u+wq7LHI1qUgEerZEZbtbXegYnPXn9ZWQlKjlLbH0MAeAWojXiCmS/tkDN8Ya/Po
ngP9lKfBV62Fq7I2Hj0CG/HH2qNwynFhK2EjeHDOOJU=
`protect END_PROTECTED
