`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
359Ds9g6qw6atFr9N2Y0+eN3AVhqvVFzbxGKf+25LnTO+LaclV/r0amDfvAfOD6P
IPcG9IP4yPB3UhLysQtH5S2z2QrledAINyZ/f4UCdzhDrm1efF7NqUsqFAqf2CC2
GNbrRt106TCk6yIxMGE+u/3PFIt7MZhEk9VA7n7jSfBltgBm+5nbZ5x1ARm/pIsX
2nu/WLUFbXgAj5sJc7XSAasNddyB+6vbLp3U+PFTyM30YYzxBNoS4V+j7uhEcr5l
U/Ij81YYVGxWmoZs8SJ1wFqgdtW20BWbsleQpnyw8YBpTk4UX7xRw34ybgR/SV4u
F1PCbMYKHIwU2pMJadVVzu/CG0/udjYiw6AAbAWv+xtHjRtVbTBdIIzbOdNjsuF6
/VaTX7uvMHfq0/FI76oiTFNSagDKN3FJjxbqoV4FYf9BS1aCCrNvZ/zy+QH8F/GH
KPrLzz/k1AXmH2RjachAsYzEABWsl0iYTn8DvsoC6yVABPwGOdPVw6Fke9icbOQX
4vi47znOIUFD/0wVdfdfLclCgTnIdHrxOuOzIQyy8e1r74Lejt7aRceINVox0RfY
qwz7ieOa5VuwTfWej5c9MisX/5/nwD6oM9rMB9oDgD7ecQfxCuP/HDARLXa2J04o
0LBaG+hyc8qW9zWSEdk9qhQhmpRagLmuMHSk+r1PboRDTD5NeBz3App/NKgveq8E
3WaROYYEhKkuE+22zD5Ve2CmFRX9DdjdGsERLzJJDF3m4qx1d0wreN6Y42NjI3U4
G9OfwQCFC6EnIbYIuxzugKWqUHVr8XQyz47/kEptGdLb3stwGwRS2pZObQAgFyRJ
G/lAncnLVZudl5nB3d5EuiA2JeXjg1vLYWP+oDRTkLTMNY4QEPNK/HOj62WMvw9s
JhvnIK9LNuUf2LQ+1WXenJuXZOzlE4zJXCnkUlra3KCYcT2mpOL4J4pfVVfPaoH/
Y4jY5c1FubYAYIghspgrKdBqv9/uCszyuYX6ylPM4uY=
`protect END_PROTECTED
