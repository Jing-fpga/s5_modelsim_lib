`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KLgRXYvcXHQn+jrHLKxTF/wPu1pg2qW3b99mPGX6akpqH9kSpsVZ2Jc6yUDxQ6fF
YYUPd7bW70YMyPbmpua+ZZtlyJmkIJKT5zgHJl4tRnb05N5a9kHCKZuztRLQOCgd
fLlVWNZoYGxcEhzJTFpCmnwjsitamGLry4pN2inVpjX97LehIv3e+siAxJ5IcaUF
ZbjbU4brCf0qdKitVeB3xGpiiumVkDfbnCjty4aqOCXhlsyTJR8+8oENopJW9iQ1
IDjzygwtAdTIV76OWWhJMcv9CM2/ZnDmruCZ6yepdLvzeSVme3eYNln8UAWkNZXN
6R3+D5rrU6TR+/r2G5tVU25wRcxCl2RFrVMWQjKKZp6l8x+JzcpRDAtA4XuA8CEF
ff794B6PIPktZtXQE6GWmBh+A63CuI7hyPGf69eIBqRK5BoAY2pBp5cTF393aXIy
3NJ19JJRTall0t+qdNzuFynlRFVQjLhM/4eK5P9lBh3XfKO0ENkBPZVINh/vdxJS
YzT/b9Kiqu9nZ/gbCBh5nqUNzaovPaEcJM9Xw0ropW1+piUdJLiozinOvmA1uIj1
b+3UlVF9TXq96SSUEsxt9LUTxVwxoI8qaSmEWG0TtYHqzTt8ejmgG1OMAJOoF0pW
ViFjMeZOUWYBAOhHa0224icnXDs4DPjbbaPHi1vRHcRYxqsx4PiGaZ/jfgh4FEcd
meiPeze+VkjwtTA5mHZWdgXjLy7QeIuyZDZX5m1xEn0Ahjlo8BTXpoUNeV2ALMja
5l9Z/Aoyi6mwBYXQMxLcMipwbzQLWcDs4uVeVaIM1/oveIrR4Db+L9FJlzHR2oDO
VEAjlrkVAvpUO6n5OzQsvDI0kvIrGgxdZNdhVVj5jALOoHPwTOMd4kvLoJ85Svjm
dZf0B/j1KrnT7MGigFPzSZ+T7yNbEgu9eRr65aQZUd6wjLUR0tsWtcve0BLFMtph
efNod6+UaQz73QkzH8i9AQ==
`protect END_PROTECTED
