`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Td9RBdkLbH75bS8xsMVq4mMGFCW7WEb9YPQzZZZortoS0snPn4xUxq0yf7TYGak
35JibNHXnVJF6pOXQDUSxYGZmvyOYZl4Go1Q7Iy38me/GRqDBJkKFG28h+GeLkTi
v86kJvVA1VNpTxkcUeQE9PgaVmF8/DKOQOyeCCjDNAzl2Z4K55trMALLm18ogEq7
91EhbVoxSzwgQW6uowE5s5tIUF5VYgsg8Q1ossIcbcKQz+wnE0a4IgHo4XPmQULi
BDZl3WWgJEOtmvIUEwI6w8xHHj/0sI7RD19NrAZ7h8OmGnLgG94Z/t0ZT1D1qEkR
5Ifsw3fdXTX3TdEToYAOrIgBwE2VM6ZMip36Ilk2zQCgKXa/+PpFBPVN24c4FsLC
wBjv9Gw1fKnsjKmhf+rGZbU+1QGMq4ekql7jgWkLLc4qfkIOjHnsuHHtqVHk11wo
fN5M1AHm8Bq1MjQZD0Y4OS4kjGYX335XtbVmb6Ip5yyYVGRAJdi57Z211E+udFyo
muWf2LVzrqLL+uO8Jf9QvBT2WUoyvsKz7q5PwZ/srgDi1uovbH8jBDmnoQ0ovGtn
7YZnguv+3MO282YcLAKVvoqxUjanXetphyNzzgKqtazdAVbJ6FmOhz8PQY+fUGiA
Z3BZuuAwqccNShZ+Bklb4u/t6pQI6uSwPU5iPqK8C73382+u0YJYItDjK6CqMWTA
bWWb5coGCQE2XRAAX7KLZ70IbT92SQhoXYUIrqLrfAlZUxPaiYqd8RNMU0s0rIBJ
rTF/RSnePbZGn5hzC1I67PVauh3kh/S9jmcG6LnQ2gUAbUtO6NITfoIuiCiRIYL6
60lXAD0aD8tOGHopcrarP1UrLL5ijfFNiBwzh24UbClkbGKRWhQOumXia45M9+xr
tjJtUxy1S5keVPF7vxDz7Le4kYHJ7KVxzBZyk+fS+eqpzbKvh2o2jZWS3uc7h4eN
YvEhM6LNzK4Vkvgm5WT8Q0hPsQpFTKBw4n7s8Iv3KVJ06iNW/tvsleFMFTSM9U1S
cpJgKtgd09x7QV9SMpIyFOmAmvPGMqAQKqBgBmk/ecv2EE838mfTTQ+z+Wyh1g+K
qYHP5YrJM0987m3FlLAkGgHHCRAX80zy8pynO6BY++jye9v+lXICB/rMOuLbSQ1t
i/6lVI1PLAypHoPWS9Sh2Vg+E9V4oM9AdwVb2+XQ6DwdDMn1JmI0v1kb1qNDe6ID
e3NgXjY/NxY43uPXKvu1GFeDusUNaOyzvdSrNuIifDzb+OI3olmdFI+yj3C4IQBt
G0eRWgyai94s0nHRtstTIPDsiJxA8M+vmY0Nex9ErJ5MNJMS+1gMrcPLQfjjkqRO
41Uq9cyiSA9CHkEBE2kFxm0U5CTZYqLAmK2fAM6gYcdVnoIMPR89tR42CI9fONeU
OTrQfwp1Bdphmf39SqYl/IGCmVRNpk+kOzfboVUIs6biMmYAX5GQyWHzObtw7E7v
FPLc8t9CsT3jMTOqf2iJ5nQB3UeRfZmqQ+d2OsCGUTVzJwDEc7ricnPnOvuRmBoS
/q6YkJz9G8GfL7Dr47x4VWXHMXxgPhJz0tb9yhQUVyBfbmU+dHIrySK2jBIvipHg
l6R6ibIdvoIX7NAyWOLGbNJoAPqqvMYbRmd44rq3rZCNTMpkxFPtmH6+KdnM1wB1
qH7SM0sLsWRUTSgAD/5WhH2VvFF1wJmiZSYg+lv1zAN95unb13HBmWO4LqYNI17R
Ao3Su8TEXbbI8XaljVSSG1qdVTNHbdJPYjZ8geiiajuPlAlbdkkVcH/GYBquG47d
v5922GLfDpuI65ERFWzP+kf5+SwlJKxVXwTPM0p92uhy9GBLSia5HjQBSUlUE9s6
cF7qLLYZHpDIYcCmuOWwv9T0dZaGUidF+p/fnFIJylwMOPl+CeSjnnLaQmKGl4F2
tUJLGenox/ZmhlOW1bWsuqi2BhETYXtgxLCU9sZVYljx9LWYDeS1xwqU669jiEh0
yoO/5bYH/Xrcf3UjN/OJnOCsRpA2cjeWMSzdP3i0UoNQGSEuFgxtwjHQ2fp+oP0w
lmG+/OS++ND4ItjEaIR77BShDR21GUgMcHmGOUAHUTKuuq9gyjUspAYWJb4OB+Wo
9Faet81D6xLhSDVZh+p/uSYbrf/ebVlYCFoTB540dq28sq1PH8OrJ3Hktgs60gr4
NPvwsx/jqo6m0uDmyX1keLEts3IPiuxWk7nC29N7O+KdiK5x+mD+So6c6OJY6uAq
Eio2p6ai7LOEqsnH2DExeQ==
`protect END_PROTECTED
