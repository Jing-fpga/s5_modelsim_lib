`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
unmLjnmsauT1RrBb3h/QLQrXoSuvTAPOvs0/+GPjVy5kZ5Qb6dhP/tQOGpwMh/Zn
uA94Jx6yu2z53oqjzUjhNwbTwWDMJScppsyaGLKYMxesuGG73XYAN8TfZY21oC1c
hqXPLkaGD9jlkYyfX3ScREwRU+hPFIfLG3eGjhoqa9fR5kvqDQcbvLm9P450TX6m
N+MSd9FK7EB0DIdFx34V+UsyrpHoH1nrm2CSDBNxN+FOdPnokEPrn/EaQE5NIN+u
7bi+e5DjEll7jgFAtPbcOaiYnj6g2a6/pLvQCrlcfLgMWv0/kVOJ1ofMHL/iWD9E
gtHaB7IWu6gto26wlQbSMsgomtLHUEG4nb5410VjCHJvdUKz0RafnGYhZRSZEUK6
StTtDyR2uNVed5JuISs5vo1fqcMRPkkoef0HEAvuj+secqhmssHf29CpzqJK/MdX
oqKJYsIUkymLthop9MBjxxnuWgNoUBTfGahrkeaEMubOlwlpZ29aAIHNnfvRFybT
8PMGRx5aSSaXv0HHzNXayJlzbqagWmrVnLRFiXXb2ZQzu+J7tMfCcrFy+f5x+nmy
VtZRItLxN20oV4bHWjFrQCZHuRKyHFwlyomBEvWXBbBhVAdHpQg+R1eGjcrLr3K/
0/VHKkdpH0nQ4ZXA08Qrf7AuJgBn73V4OiP/etAfwP40bUDQUv+7MqImprxN8Ntd
VjtEaKESRgPfTyIasV2xn8kWvYSugsgyO2B6HXLsCicU4W+wVdxmWgh7SNBMelVY
O2RRyOhmevOMMVl/tOdJwvykYX6bEbQEAb73Ump/FbL2a/5mkLGddxrziKUQaRM4
d16f69SA1JrGyBtjL6vT5DCfYuvd74pCGcnvx0vFopB/HoWvigqKvIw3SKEI6Knw
yNkX7HAX4DUHGP7oTlKZE5shtBq2Q6weIUHKgg9zLFaRHSwXsP3IgmkVcKyqgKPJ
jWDrb4dehqzCpKCZKHVFbZ4KQ0/0bM2OPgSBB0iUvZKcEoS7XIinWeRLrKYoqeci
H0MYrNTTqGK+TLOscflRYkAjXzGNNKfRB7Xm/KPc/S27mP9On5pjnUhxJJDg3ZtH
Fh4u5CFN69kACpGXv3PEQ0ckxTLCtOeqLkRGH0MoIqDWEud9WGSew2eoEPTNCe6J
cC0t8LmGX/KE61IzrSA3sSPsrGrmd6kznI0eigJg5XbV1uLSEbtw/UlVKk4MJRCu
0PElXSMIKXKv1si7ZI34t5SX1IBiGGfG9MZVNOpnLcz9+kQQ1nj9Frz6+mqhV/L/
W/wuEPjIEg9Iqnpsgy/MIx1bNC2Yl5Dm1h1oXntMAsfOPo8HV3FVw+YVog2B9Xn9
AmHxxJtkhFcnOX8wUQnSW2px2AqeanXgqeauLPpOJm/8h7EqWhm2eU3vHUuvbJ8U
tKctEM0GYWAsH2NYJLdmvy+jf4diRmJqaXd52GpoXhL0SiY93AfuIxxgxTF0FgaP
VL5R2IMaEBelBM0DAlf119bbIy/4bXpORsbBp01X4egsgdMVghtghgzg6k91QLs1
lvoX/5aDnE1M1WwT0UelJA==
`protect END_PROTECTED
