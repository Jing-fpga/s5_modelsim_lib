`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ofrrDloPF0NS0+G+F6AR1uCaqTbMIqoMvTPpKpxNrqNujGG6gy2+BSR+6sFz8Bp+
ugSpByB37BTdXGDnn9UMS2hjCmuiHHQdFlmZaQ3BOcH+wgSNeUIn7y4BVsDchOGT
21Wfs2jKLJ8IcrqD574820YWX5Xha5PL8Mf5Zx5hxnKMSlNTYkYVC8jFVPyvDbcx
XmwfTi7CEhqnHbsaIloLQ2HjAcFsNDIhU9DaviOXiWlU0MHTkZtD6yyoxPqBRLBN
11+OdqKFkzWaB/Uy4YcXEsJe1FJSrG/qL7Nshl+/BQH6iJBas0V01+QS029b8xZl
Up441yRGtYHP4mUraZCMgpqPtDp1j/sDzFN1J6DrkSFAm8wieBHPdqRwpHZHgKWl
0UmUHMIeAG+hPodLRMD1J7pvDB4L/YyXkiJM77tRoYN6qZidUCm1wkSHIkcQ2P0h
ZZX75+mDxcpSQpNY/WCseWcgVhA7WOVd7vVFNMqO3O6uNjUkL5FeUANkxka3CsGf
I7NGB4LatrMSpQx+8Eb07tKzvbEHG3EPgSxRbzrJBoz1MwhK8R3yjWlbzpwb4j7f
DYHkwrS/+1Wna5pIUxtidNjXYHS1dzm62Jdx5F3fP//zMDmL2WVQXO7gII8kVimn
DyEbqZhFsns/jlt3Z3uWWBROqDhYKymk82D6a+149BNusezkVYb6A/yWxLJltx9u
PeNS9p8hOxVGIam8nHfGP+zE+FuNO+l+7ItTcIwlmqlswVFsO/f+8KpX7L6VLFFh
nKButGnvSp46t3Ab8oG9R8GuSxDfGqMTk+ELZaXyuJgdOrv7wld2V4reLVleEyNO
iTRe/xF9dXaR08m162MHKMJ2R5lQEYCtriVJLX6Cf0Vm+A+K1ZvUW5PU9swa4Gh8
vMZUVbcpmo42tEQo/jaAlM1+UMSIkWn8cg4KkiKCANi1XvzoZve0dQpV8uU1yYnY
fRVJNcuKmP72YDmaL5aUB0JHIB+C0zO93CpUIQ9C7N9aQmQFcLVhd8nLtJZk3H8H
/UOF8o/U7UC41eKk+9jAtmi16ZWhjCUWRFF7Eecd/JZ243umbIkj5mxNM86zY+K3
RUwabj0mizhoqggfVVEml8Yg3kWZNashnfMy20PSimHYVGnz5SGj80JXrlnXkgY/
WyeKbthXrjkwww3klpOyVa65gRr6BwH4KNKzyHvsy++dFAej3Vf7r4dgUaRd8iHY
NZBhpQshJW+/tgIEsa+jOPvemkEtYxkscg5Ld0PKdSKgNCKePC1py7PdinKEigvy
nQ06j2HHJeKVNxwz5g1CAcpfcqyBCT5vuUUgj6AVFySJQ+OypDPO7YpH4hRYyrK4
`protect END_PROTECTED
