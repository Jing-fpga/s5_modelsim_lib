`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Pn82sU1uHWjUEYzHQA7WfLG2m7IBtYEgPJeP1vH/FRfSZTch4GE1S3KL6XHolF3
bDq276NsVdr8ft5K38nQGnVxYU8IjdPjlAaBBAOKmfh36Ku7ucejlU3XcwSOB+iV
tWRl2LDNIoJbWVbYdR2BowAlXaEa5FRM46ypOUU0D/fq1yephUrWzFy1SYT8nw0p
yDvY3XzJpaBIStA1agNXtJIyTTkm81VuKIHSQt+X3Q0+HJtMQXzTpaO/5aweeG9B
tYSA4dageUsqreMaYRu4cjmFQDgoZdE2DqK3ZAJm67GSHVQWCWYz/rmhFkt+E7qn
chxu202qSXA6v6jrCw7smahhtqttU2PlBuPjfIpu7sbdmVAPHqm7u2lMDEex3edz
ClA1GhRxea06yuBcToQwhNBpysT0qN4yY1BsTSF0TMQpNKaHWACkt8HAiO5IkglJ
oOmGwseLTiFJdilakb+RtRMwO1r1klhF6wHHOD6wLa3c/eEOAMO1i1aOhHf1L8hS
ZMR1AOHM1RCe/uo88+iUyhcT0tEu0FXqITQoAoymrhXbgi6ytaV1M5Q8KXc92R1F
dqPWgDaM5NPfDCklaRzfec3elaxcHgZH/OuJAiYIomxWCPMYDxhZ0NaNcd0QGX9v
p9nzh/OiD9nWYXMqRI4g+YRuPO23xE5pY21hqaM0V4B70kGJ21DLXaCI8rUBie7C
Up34JdlZCw8kSJ1DTLvEWw==
`protect END_PROTECTED
