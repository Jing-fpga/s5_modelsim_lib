`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9ZDNtIczLr9Xisv6Ctkxh8jZQfaQIuk+AZ7oJnZ8JubUMuN1wPGyJw9NehIGG3G9
Cf4k00M7yA5mQvp3u2JRsQoJSxV+tMVvDVWnAWxcd3k/MN5rRGu7TarkXyLqncCG
fYvOqppRDQZhIoB4KfqLGJwAuvrPyOY7to7/65OcwEckhHVLB6Dp4uFCwX21+oX+
dguTcDOiHzaPh8H53zc61YiFRnldOwHbDXRURIHB8tFZhJWRpadZ4gzKwZQ46Ks4
UQWLCElOGUrCDSrhWvAZfR39a00GTYfYZST8rOvLHXQ0hKGzgUIbBk+3Yff4dGgy
fSGOO2T1X+8Brnq4Br9kYZL4Y6W/gruhw8HDw2qmQjiZQOg2D7LyoX3SdTyFx8DL
hp0zQVvVaZ19C7fLRbP0T6h2Hfh/8Yntx9F913z3bFJtVACmkXGn0G47JGjCmbzU
iYW/J9IdHBYc3AoioXl/+Mv198KSHxSDIEeWdLzMlsC6yHWm6YpoDW7KJzaA0xgP
uxe20wu6AQnTqjD7VWg3hhReBO0FMA12g7kF9Yv2nbRpGxzbvBoQKLXvE9kMSqsM
HUNwHM9WMdbRKG7EetDkVBSIfpkB3W0A4Yx32k18Av06m8RJT3m3dRBTWE9NH76b
WuJ2EcUY5bSrqaZ6t9QivBKa4sAYXF56aXck5uRxkXCqyguLLphqx9Kkm8ypVbIm
XFxioVPWuc1sR0HzKxXKGvbrESK6cbIV4rkU1badgKYsf8X7co/vRi2aD1dAkOmc
6Na0P73pqA9hRb50qKyA+PorCv2Fy0ZuZf/rwVC38xHw6Muy7zKA/eb99kDKwSOZ
lWrGAFA0dxlfGo32bUVRxImZWy7yxG3dQ23Vs37vHUQqWVwoMjX7dgE6ZMRCfGLL
f2iqbyI0Vxbj+IfYfgdr+rv2N7yIq+5fJziFKPiKLi91CQFZzaJF6NLJrY1FEONd
qApePSEfCKdTgQCMEESfIwDRmCUdEV+s6udP7cpy/+uKQ/WOfO8Sd9+L/aDHxtcm
rrWkC4KWcDj6lroEysuhsEi/UUMucubuSEtaYVKQk+Kb9CaIv5WMo6yAd1bROpee
PrRhUvaB9G1+FWhGJFsaZY/cVCLQHnNiWdwlOySfyK8pgQAshgEMxJ4KM8bcoCwa
FwBJ/aWx6BBc5zH8jJcY+E2tuD0sVHOzy5vBv5UcrC2AyNxke91KklLCJx0AZhYV
QqHYn/ub2RcaBPTDnbJc22eGsGoAIAQJGPwU8GiLl0+MqRGReDEFWJcGt0euhE0J
PgoNS3xj3u+5UBBuL38dd2U6p5cJkqSdQCWkQ3aSyRAV3JFUaWne4/uSDdCiJau8
OuIgTYjB9SfLRHrnKY4hGQNWXYijNzm+ikcfkHWYSbgl9C1Psq9PYv1BgV0hjGW5
r3BbclGgpbC2XE3bneeMG04a8daFLOx8CTbY3fiMNBRkyVnsXGN+ND+zpmlY3shO
`protect END_PROTECTED
