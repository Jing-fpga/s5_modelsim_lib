`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RYMw23l0WULpdkEQ51+4XZF/kwfDe1dQRhGp7/Ty9vjKJrOs2+RqvBsYfCjf//4W
43pyxklK7pqrAZo5wnwK9akpy92tsgOi+2cqAru8mcqDGQwkan36T+zPdKS/QmxZ
/rsBPeKf0ZZGtMY8ND4q7fgfJFh36wVYMOHlQJoQGnd8qBgQyXkuu9ktMq4XFl5i
EuKs9/Se6tCtGvrEo/CT0P1VZzVJfFoSehwFdAlcFWFp+MYSLvqegWFGLlKep9vy
RcaioMfCcEI3vymk+SUlaMPhuPCrv6YEXcajmZ+UrlOmwKdVvbIf5+FTHMMmQ1y2
IlzIHPjBwEvrGtQRKWgtPWVNIcSw33ZI5dkj8oKTvMLSzx0qkDibEI2w2ftpJVdF
qw82EhNAoSNkk1tI61/6kUCadzQAO4EsrNxicwcdieqYsILvvxoNtwVm45P+hNyP
uBFY96FcWUUJrO8FdR1Re2Uy96IcQr5ZHeQdbVwGqPz8FHp8m8WuupgsxsxsRczl
MkwdZzBYQgMMRT+IJwcErXVi/nIIp2dkhXP4O/YOXEsg0dNFY1d+4+gK/GKkA1gS
ThMgeSF/3BPbRU1nxMkNXpkIBxXaMSKCq5IzbXH+diIQ5rlh1LHDVtIGKlG/BWik
S1gAMKX8vFMZw1AitcMTyy9Yne+4CmtR04gECmJ+2COyChYT959jVcQNMQE3L+3H
QQGNbwfhwYWU1EuUQ6ut0538iOrBq57canbSmVEl2jsE7baTIkrZDRpQCcssX+DR
z+CnHT79+rparChrLatwQUtoT3Va2D7iMVE7dNGRR96LEb6nR28zYcpsJv/h+LVx
aARI0lS+OBkNQVzQXO4wvPRarXnqHhBoqIfmmeTwMPpkzFzprad1zU9bqNnkJBSh
k/lZQx6tbOkWaYCoBbXfiiRJG5wm+H4IqZn4Js/n02gMmqmeS7cErn+TdE3LRInf
baiR8el8Trtj/uPiwy5UyWe6hbX4DnjtVE1uEpt2njLUsy6zmuSVrWoso4nj9Q4j
yLe/6TQD/RKrNoRlV4PG6em5iGoe25D3nTEkesbP7c2LKG3lLaPGBKZ+J+w9Ga1c
sv/GpDLqI7IU0H/TuEajJ1Kg1xpTbxwGuc26nbaZexWarY0KYu+aXnob581xVcVa
BryXEgFV5xiSKFLr+mCHxTepekfNJzYfWN2VeEMJ8mbrBAPxkuJcj988WSino33s
EC67g82/koTYEC/FqjvMk/MW8xD7sTpswZATnFAK2xlBRquqAOewlnxhff/a9Ev5
`protect END_PROTECTED
