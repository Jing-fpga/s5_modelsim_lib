`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zk+X4N4IBmFQRbZV2uP0lxvQlU6T80Z5A1FGnMBYrmsS2UjfqQkAJF5DPFy5oPBy
KFUJlc4ZWJ/MWZmEC/tCCf0UcVq9h3HwEreZ4hzRXq9/9yYzTvPlHi6ooNq23rPz
djL2r0ny9E+gPGBL7QswbRcFM/FXvZMrvgW40AbYLrYjFbX0LtyDIfXsramIWMzM
pr9N+BB5Uw9Q/wPITcMrNBQ+h2f3SioF3RQHFowCOvuDggdabIcvqnSuIlSua0x6
Bzz0PAyyfdZwD3oGdawShdQnNh9e5E9CsP61Vn68hvPW/CqzKDfx4AvBJuTdji5v
+A4IsDDcrhV6Drh6ACVuJxPpk7jpccR8TufuzUaJ4YJBndFvlkcuVMZyT4XtnMaw
qDXv+j9sm6r/y70L5jaLGhkUq3Zr3wFxQscryLPfxlrdcxAFeV/8ZXhlq7aNbRhV
yjyGYrU81TccbaSTwtXkbnWWPx0tyt44A3np4rMPhIUmbn7DcWKPcFk5upBfj+PE
e/0+FaW8wMTojKTuKpR7/OBLH1k1ktSRbubbXyRuA9icgp7T7yBVGLL/KFuKYAqo
`protect END_PROTECTED
