`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kn/vSv9Rp7JiIFce8YNSUsxx54Ol1qpiOsyX6Z6mkleSILnV+sayqwMKtRqUGCNW
BbnGhJnysy08jrJwNjjqhNuRLt2Q5twAlflbR9C4f9jDPgj1Um/ph2RuOwMKe87n
2GDsZAndNXef0QFPIxgp0sDdRpVPyfO9Dwiult2Or2bL12et55FzzsZYL4f5sSQ9
9WMChP/3C2UKp9PDpU7YcogjmQtvCKh8LXGUta5h+B4H5tyQXoDX0tGdDP7SCGiG
ZTB9toGqONts73NRhlhitQk1sMQlxTlbJUGrF3bb0Ehl5L8gkgMnPa2C2iuNZ2ii
qB1igKs5BI/mgDF+1F6dQ2pV/NgzDx8cEmEkGlpNXxLz9G+w7dSbwWmNTRrroTbV
SHtFNy5bB6E6PMvj6ZwzTEAOP+V58vDc9+qLgj3vOjz1ZMXQWvtrtLtv3+gCEOK/
aYAt5893YAlBd0r1Om+NIN4+JYZzRILXEXqSRgctYpfIjGmmuhUFGVrvfoX0X2Ab
KsdDYih2tplXMcElykHTgVaMLSSY+bejS3Wp0lkzLW5ZOMBFJ1tgaZfM0Ehk+8nK
/8mhW3pVDozU6GqIhhjB09dXxPduQV1sDnycrZy7cKNI/j6s7EPrglFxpb5sBnuA
Xb9NeOOzFyx01fdmZiJe9vFEhSgsK1VY7gU86toedYAruFAx/e1bJwKCE0b4cVz5
ft2lRZGH+vC4mUDLaZtDt1aGTEKdkKoJLQu1D6C8oLf2oG7utYY98ufh95KvYydK
nB83c/ijWPeZn+AmmeK6WsMpmIuAu9E/Gl6DaA7vg8NPoYArUZV1qeyqThV3Geue
eQLEjG6eH4gO8y4fa7OKY+9v8eygCxrWtouVrcYshDs68x3Q9TWpoFSDOjXbkQn1
Lojk0teWd4P3Zr3acSic1Bt7MON8OfHiQR+GOhcfx2hpoxAELTlMX88SMZ2oi756
UkdfOxdrxydyRpPOdkUhLFlc0T9sy16dFysG1XtwqVYl+4dTyFiV93i8Gi17wPoC
eJpvpggKvh2W/VzQao7N2j1E37Rvrd5KOc62Ig+yVlQdnXhL4RUnGPfzCbaBSH9u
bfA8g6RYjPRBYNcqTg9HJXcMQVs82yyHo5E9sgePnAIw7fQEPTAWJ3bICxffPeu8
C4VKNkrdogP7C2E/BWQWVy8RINJko0Es4LLlDi6g031QWSZgN9EqR5huxZC525BW
ISIOFKtCNtjKv0p+SYKJ7AZ699jUZnaNXCFYz3XdHIORjfLKsJIFa+qjlQPWhOwu
MvpPkAht3nqdgOTXinmVyr/wVsplNPwa2AS4hZlbw+7vdG8H6CEu+3XlrhU9mcCh
DqOPw5IVJ+Zf3/e8acM8W5D5kpHB3lkQllPtxFBuuadCo2mbXlX0ddnasUeQNw8Q
VYr2qVBRjE63iAuNYanXE+7ntLs3iYl6cLaOMObQum7xjNnfYF7ZvvVum4XvZGr4
GLkk8tN8rKpbJ8PEt8bUZVsFdp3IapdxkH0l9a+NoROQIG6mOBzXcwzsc/Z+9gWE
UwjmWuijA0pg4lHHgrFgdStt9BncnIr0LSTCdKuDzad1eGTftkX+m4ngBynBpsLf
DOzGXkaE14qvGjtKtb9an/DzgXKwVNSiOqoPk3b6Ix+Z7uVK6TtYXnuJzaAS0QwW
IekJzwUmITEWD9EORMiYcJ03XFLP84gLQULUrMAFajI4YcXTRo3eNFfRnSoD0o0S
bcYEXafDfOQdSwJ1X4NKX+BvC8MYz56QXQOA0XaQLyxQ7TaAGYeEPEDHrOC191jc
pIDRR87cokO78nTyjoc4tyxD5KK6m2kl0NgstxHLDS0LBCtt8/EwCnya2SuUAPkO
C6LIxabjrr9KypS3wZb4tyAAeXXv4u74PtubKwHt8rPzZU2V6Uw++Fa2uYhVLPN4
/JZMRLYedBNmSsWN0D6jI/AQUi3IiFk9mU5lRtbpk0z6O4yYaRGMvAYut+D/dM9Z
c8yq50eGTPIC9DYDjUjsOjBPuNWb5txX9HF46dOJhreDbe2WZJnkwz3wBUlhQhT/
DLPr1Smvwo+UIxHVcodiawRbBjnftDXfB4TLQtRL+VuWZ8VW/rEOy0G88DpJQwQe
nGqVcnGOFUC5NXhtUt8y36VsOSG6FLbUssaxxZUHFGkW+PIrahxV/MeAe56TMAdZ
pEfHuZsetT2qV5/IBXBpSPdbWH1i/bUDxjmnKshkLcmKCcNio1i2IC42+jhTGe6d
jPIrTjE0UCTRJcMCF8GfpM7wRa2+pDY5DEhyKIs8/IvcNoILgu9T3o2EfsKE54n4
XMWlBLfL5LHNbdSN3cr61B1Qs+v+f4t9XQ7ENoX02bviZaMaWlKaXaEjaMO5Sp+P
B8kGg25mWd5VtC3VHA3u6WEnq3ZPf4jSL/BcmazHTYy/qP8VLUq8AicqqDNHKiEl
o4dEr7zuRhmRjHi0RoG//mET41XI0xWe7N2fVGLObz2v8Kxo6Cc5z71B4JgJBHZJ
RBdgM9LZy+Jix5J5dfuc9dcX8ix3Yq6upxVDdgTwE/utMCHz6HoiRkaOapjcf44S
WI9hUgzbGcydeZgQC5pMMhyhOCudXPTSgyRf1wmyEMOUvx571rRQjQYu9pMhyvaA
E1w0KA3V60WMppTqd9azcI4wMDM9ItQnsrZDzd2vTDtqvDLJ/x5NGO5ptroGnC6Z
uips4PJny5X1hEVdtb5nfO8MRb8kJfA8z42hlY7ojgs3MqQaLJcEjfaiUjkA/kqH
P9d0UAJqSMJ3zWFXQNNveLn9WxVb5fR1rzV3kClwqxcwCSOKdJ4UQTAoJnURS+7R
8pQ2uRbE6cMcE9XucThbkdiA7SZhJy9zfExCiS0hIsLKk2UoHsKcHa1aiXxFvB89
ZU5xvqE4RWRJQrDrX0QofgFqbZVx6TGGDMRw+q0Ygb7EgKTYolUKXUkYTyy5Q55T
1pqzBgchlblJwe1WXl1uXqsM/2fUAcb1bVGioIcWOoN93Ncm7m3lAgVtLmtbGNtE
+RFPyw1pqHFuxJfXmLW5CV4397FWeYEPxTPdh+WNGOKWs1jV1t+FG4b9+n7n7Ezp
BTsJfeWUIihNcwCou0U4FvHCtElMBSYoC4UpaT/PAGLTuQms9M6la6Q8lkwa1PdA
ygjPt15LVM/mFTjjJ3w7g+XbYkdELFEegdx0N/WIv2scNtDNmdJwep4MaJMlHfhH
piW90HmWRTCqsz4O7WQ53rasj3PwSAv1XSoJ9yFjZdOe6o3U1i/PLQuI28FV7vrL
wV47xL2ut5P5VqppyGhdEXo7frRIFN+9El5tq+muuGjh48ce977A4VJnqOmC/ii5
IkwcwNx6ixODYeElU44Ftt835etaX7Jkp0XPj3fapcgPUwXp7tVVzJG+E72qPDeX
/BLFiABAM5vAMb6f0cGn/prg1zp4OZVh6UbG0jokmycfFcfMr7PIpRklB1Jt4fd0
r1944bpXJSRnm+++efhqWIAtsOmPcm3vPzNbNpTF7z5KKBbv4ApI1WRua2ml4oAE
20F2MDl7m7K1gB99XGzstG7JSlg5EshUf+pFK3GAcPPuRPRGfhW3y6TNzh/fIK7y
8PqerQXk38Z+Ewr4ZUSpMYmNzcWTa06WBnvSAL3Q/WyY0W8U0+d3NhSDi511HUYH
vDJ1PfzMOnbt0pcX87FoIBC8XQCXAp4kDzOYxLzXCdWjy3ktZAv20V98+ykG7lPi
fY4nY1YpHEBIgEPNak3MJb3heWEEsP7tzGH+Dbvw22NZ96v1wf7WygDbw0AX7S8t
2uJfg0eKBJLKWTVvViEb/v68fAfVxPV9PHxsXk50su3rvdMryM+VRYYAMFylPrjK
uyYQFpKSbI6D0lC5xabDXEN3//dNYfc/RroqYjQGaPFb7nvTqBkpWt2yf+wRFgYy
wQxBylPymdEKizq99NDvkcoYOBxVEgVggu9hA2rLseZR2WX/GehFgg/biOiK2WTe
78qIEcBTq2mMRp/lxotnAighf69xyY6cNS313hSNnAEwTsIaCliQKICbw7SjeMfX
SlGbFU5y4ZZmFD6Qqv+DK8kWaeC6ou2lCpanFdWCk7T0WrW3jbo9rK24pPF8h5q/
gN07NDrm57x/2/h2dGICP9XholF7i2cSX2F7g5yzHNDA2JmxhUwkPeozKjL5vc0a
Fw1+8DH32HV58LTjZKk9xtYGoFmff190schgR1TmlDTrr0jaV8fWWxFmzM25/uuo
Bq0U9esyNGY2C9tztTupquLIxoA9i6vXS8GL8s+wTC+XsyguoUg9ORAugdN+KmMx
qdxP1bGbHaBoakJ2gM7CDIYHdb0jhdWksC85ZZ6Im5ocCIFRZfPqKpyEvp487hUi
8qeijTd9/kh2l1UgDEoLtuAQTgINrNCHnGC3+VkRwpVC+8a9nn3TEg7+2oKZfzzH
tZu/81FkJIztzijsXbhBauqy5Z8paswCkiZiECVqnPIaI81BzXl4lTd0w/ad8nNy
CqeeLCWJR5tyF/t6h9fnOEAfJ72vM2h3LiVoLXXACe+50BenL7Fpj7iz7olmQmUq
TOwKDncJ3Q9AZfYn643gLuOlRFKXRKG+KDFPTdNydXVNcD1vFwft1I7ncs6CcNRO
nBvmPf20RonITtqnhmHOF3x1CfVb6nMnVGXBj0iPhTIZ7pFZwT1j5yXZFJgzPZ8a
xSEoVoXd5h0o+HN7hZAumC2MnAjPvEEwIQ5BkupTpzsfrKxIvyDyLtowU1L5Qur1
7fz7+PpsvH7x8bIvrLARvl6eCvND1d+i8NyT7Uo8xP476T00p5cwcVClxvLiEZZZ
Mk77v0uEbIwQ0OJ6kC3bmqIV/CfzmPRVfiGilx46f9z7AY+Hcy3q0FNlKvBMGPfu
FZHstY3uLa7D5kTdclj4iqaS/Kgwk5j+MjK1nO5FAcaiqsioEW071shZ+fVBn9ZB
N9gQtmDFvvX8m+UpbsPKwW1Li4kZ/JAmS4X9NmGjnIXT4xhzbNKz39Dcgsgdhx0Z
t2PfzWgUxDA41i0CDv9OCK3Z1h9POT9FF6JSzGi+CVcdBUJ57G17H4PmVYCTAhen
OsgIpMb1SyurUZHg54JVfNRu8v0d+Kra2riW3Snxf1NmIniWCJE9UAW9x/Zi994X
uA+mCQ9xq6h18hlaNq3tkFCRMhWO79/GW3ajZADHMh/h8jeerXf1e7YXQsjNF6G4
J4ZIwMlQ/cNVl5HhYHKE9kFzo5ecJhZPWY+RHMwSbDVyavxai6lG5cj6zDG0+DBE
y+UzrBGEkQQFJa/oTl1WQJEKBnSyRvKgaW2ZHAFgUnm4rQmJjP+rVZaXdRp+2CxL
LL4HEr3PGwPo78pLxwwwIIQ1+dY5F0+Wutd3mpRomdX4zRmTzm7YOTwOtohf0G2Q
9nKQhMWhQIuJLa2rh+CDVnR73NYqcH174hJye8XmVAt2dc/2JHPhgoD6uSma1mrl
kgYdTJjnDDe+5K4A9dfIL2Ee4BK1YwfxLwdbnwNTV8jbQyKawIkEAILekAxW58+t
AiEZbu8vyER7OYOuV4KTW9yjp4irBp5mbUo5VeRSEC51bG3m5wVUAsUuYXohvHN0
6L04mxDPhbrpGuXsPL0HSPhQNx297HaE+sBgONknH48+7BzTfT2sHSDeA8BHp3Tv
7+eVw3zu+KBP8mXhDnTen62dL8MVEzizQhwR4nn/0heM/2Q2xSKQL4UurcKORExo
Q8mVdKHssRSyeQ32b1Tik+Opia4cQZ0+s96C9XDfla1m8/lLASpMl9LSARkO/66b
lK/Qsr8oZ7yQ28yV8SvH/x7P97PqQRT8Z4O3i0vZzN8FN4bN3Yco3iSgEPdztiDf
rOyELI0ybbknN0/0MbZVFmgCc11sm4U82tSKwo5RRENjT/I3UkMm6dRIODva4F7M
QJr0Sbd9+Wq9ik2WC0GmquC1u+1+gmt/uI3HMpxHFkmDAWdhe7Xs21u7GdrADarH
/eAReWl/awbu04FPKQry02c1jGEHdPj1srRBVYIRek4s9/rzz2VyATbX1cgzK2eP
FY9hg7oP0XzUvfdXFJ+iLgqcFl4bY+aIFHmdq+9M1AE2uRwu2DAVTOOEpG5TAlOC
xKP5wfpq8VUrqgRh8ivjtV2c9hpyBGoJKhJ54qHeMB92szxiYyRLGblTo9+N7KyQ
S4+hTsTTYTO+Kxky2Hz6UmqaIidbKU8ypkuCglDNBeGCfukB8xuVywJI/CJLxNWs
VyatgUGTXbZsMwUCSdKVVprBlvLfRtG+jwxv4db29xJKvS+/0Rf135wd1ug+FhDU
m7k5iFgQVmJgeuaAnYeorY49l5gj19CPsxiKl6+7fLGPxVwwJMKBtkfp41ia+Exj
7PNspX25NOEwhx3El41IdgP78fKqMi9XSpO3Bi9X8Lj8naZa/gYlEbe7AnIiferB
fQEL1YFhm3GjMHYNsAn5PKGG+OQv3et49LP5mH6J1FdGbuSglsF76eeJlpbGHZvW
XxOmuNRgyNyTlZUDimgjHtokTrwn0UuF9B8FFaQnUAos6cM+L4HDUev0yZXdamsx
HLHiEPBiqUF18dZVllb03pLJz19UCJHjQZSoDNFR5JdcB3HmRogxhd7exTQNLipC
F+3v7sTSbQutVpvQpLHFh5h0lDizqg11HDH5Ky1LEW804ggam1mU893lPKFTURPG
mRpkFxodu46sL76XkGrsTDABuLshd6/E16Hud/os43iVuKkihpL/z+eJCUgBYYgI
r4j/CWw41oRiXWQfQOUXT21MDknr3M+yyuHgKBPT0WB7AD6EKhnSxSBG8Tg2/z9T
Z7d9qc0sNBo9PtCYnQGhdU0H1CmQv+IY4tG0uc5PGm8ooxETTxEiPhta2yeZ9QSh
OoQHivSonmkk0xhqjeHEmawcIRO2f4kjz0TgtuLJoDYYcmHxfLvMFXefnAsXqQPk
Fn6AlgnNCOmDUd5GimHfk3H8KLCLKSV2DyRatLZ8ll8w+lrwrQDEZ92QZbFuIcWE
`protect END_PROTECTED
