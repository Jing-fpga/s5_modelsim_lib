`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3sQgR+e4D/fngb2S6ZdgQ8gia9bHKycEOzSCFCzgcWYYB8MRwpkGGWz1P8alcH8m
EsoFYVTVkd727/pooFGKlcGqtJXC3xdYswvIXBAkFM7rkCf2MA7cjEwUac2T9j+E
ZUJMHTWjde3Ypzl9A9LYKvWsRWzGtA1mABiD8fv+1FjCXfKfI8SVnbpI0Nc47cuw
K6geBKLhwZE3aRYNiSryRg==
`protect END_PROTECTED
