`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yBmutL+kXd1Ry/VWp9YMEouhtQ1vreY0tldSFE/Gu9hPFM4GUtGh796JvGxwAJip
kH3RFJxjG1UYoEiGzuk4Vn9XXv9zumRk1EVTAXkbjmgB9UfMIb2KrJ4oRaM2yMLb
UlLyZ9PvFRnBSGzNsJGE7oAJ8QToVeq3SkzaeODhSVdg043lKs448zFdGYk2NKtV
uZr0zhQOH84RRUiZpuwJiG574mpAIqcJTs4mMFb3FDhOInNLez6BHlZbWJxPQK3g
uwPYzSjQ5NULXHywm4qLcsAs/Bu/HN+GQ2ZOHScQYfAK0NUypegyJJiF452UXjFU
qRNZJxoPQ45NmeIoYV13tpcT2kLAPUMkX1II9aPeEc2UHHbw8fVtNAmGYMaS+x2H
pdlQRwsLrytBYGKfLNNYE57wTaFIav7MSItxQz6urqvh+CPvT/zDeiVQ8RGSemuF
+CUdgsuxl59JgeNrIPGrNixUFvSADEkzI3/091+lDFg=
`protect END_PROTECTED
