`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F206aXBejARftyy2On8cyC5dcANO/y+P341bewWEh/DpgfwWWBzW/dKIY8l0Z/KJ
uLFYytMQeIUdonNQtqkvpmdyipWziyDTPFuol/cnLqTqJOekYHq6tUMhr6DsGYmP
gMTVVBslPiVB6+gQMvNtV6EyC8BvygmduU8DV4+fk+atqG8/tB797H4vj+MArTL7
b/6yCRr9QEwrglcJ14rKlbD4NWbj70uDOf+PudosZVHwWMCvoew/TkMxXmvhs+cB
Ph5JmzKnhBDxe4DihnxMpNWhyAdvhZWia5FWVojFQLyYigoCOXY8U2Oon47oMn0B
1Qneg41HaQRoRD4X/GwmqjvxfKfGkT5yUTPEKcZnSNCHxT57Q11PJDN7FTyA8OJ+
ERwsSqwJVEmQSI9cynX3IO0+ZNi+YXg1j3UdFnVyMCqxYMQMVhF5R+qrVUZPlPDG
tArhe9WXm/PiJvfidMPnSkn6PrpiGeORgF42FnUyKqA8w0CGseWe3OehAZaS3UNp
5b7xbRYiET9hAOe4rZF2M+DJJrA88gws9qy83nIqFsw8S1/z1SBL61W/diVmwRN/
8Ka63ZboHyzMBO0UIXIokYS1emKsqXPBnFRc9HXNkFE0nY4gEnfQKPZQbyAFMK1J
rPbqGQ7PL+X9xvZQXiSXXQI4ZjYLN+RlfmOz4jqrip9aTvGQVvD/taiDTTgmiVBH
8DIT4Yd7QXXmUEA3FUfLpsF/nbZlduK7q2+09PnZd9zAIwN7PohO+ROsLHm8tEIT
/7uBDMPAJN5liNhKLJtO4SHFP9QlZSViVcp9j/UwNoxKbpzEilCarvzdgKFCkPIB
YL5BhbbvViI4eUmSDrzchadSPGBxTy2TJ4rrcIS65SfhZ7B3C3CGSne7VyllBFKT
j/T2pNZYiIb4YCQkeEG1OqThMMEBrIMe6kK29NVkgqIN+LYLbMJA2mcytBQJpdLV
r7WKGc4RQcgeyCTjffPcyNlodE2HZKvHrPEy9LEJDFSZOIDhjHDAXGUPKY7CmRH+
vu9QpUJhKy2xq3llikxSHtEm3ruatEzngBg9HEuNi+h4q9o1gjctvg0AAftcupAr
K0Jwq36tkHm0XUgi6ZWBCyiJJpEO7b4G57GL+mOgZbhBgFeJdnquwbv/9wJXkvR+
/fn+2+4ciqcNEMfaUB395VoeUgbMosAO6nnSO9CmxQrkcbRMychiWJdhlR6E2NCj
JbTzbxRJRZEQ+VTOAmMeJzaMOdU5EL25hv0qNZAEL3lOTvxPyWGfEg59ePb0Rox5
6hWoCJdfV7X7CdKIWvawFyB9LO1ZoECx35l5VcPZo/5ymQCzmqzYcyPFVD8rsznj
4tGONgVWqPnbsYOwPIt3NMGdeB6PM18NIDwCWbqUkA7Cug3fXUJvGYXmAvisOXRr
kuryOFgUu1AiWnBh+W/K2mEbTXlkbytkNCVUyqs8Cr59Aw5cMjTzKyL+qwJMredd
FbX4N9ed8C8nF87wB2sJo3mlCcAwMcHch2wqjyVmhIYk5NC0uqcuKgfkJ3LjWaHd
A4RY5HGChwhaHoZrwzo6CdjMQIeMPXLjtaVEMwgJQRx3UC4fTvKiwmOquCFciBEk
wbGNNBTiZx9H4Mx68Hst0U/mb/JMhIb2IKgyxjeDn+87P8g8CYc0wxBNhIlbAyPH
`protect END_PROTECTED
