`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9yWazqfYVH2RONHj7Qgl7EAgi5IEqgGCYFPBBoMFGAA1lk72OC9/WgXdRMZCua9f
QqudjekG4D/fHHfIbblnSNU9KEjuBkoDLeaHIB6xTQ93h5D3aGfcWQ/Mgw3GBaSR
qtlxyIOjMzfKoHI2jNMuLNuyTtR2hcu68MvkxC+fAe5R5YXR4Zdm5/RuAoPsJeyg
JSfqUb14fD4Dddja7nN4oSg5qJBZI1Jc9h8c7EPHhacob77waFL+bi1JdAQ8S7Ia
NCWZ84pO/BdfWTuHY+c4siEpxp36bpe6z7aUj798aXUXsP+umOQacJGfyojpurLg
voQBLPjFpnoJOunvILC3orec+iJUEaSW0egdN4kTOSye4fDRIRPhSauO/ORXN6as
U6BvsDy9aWo8O1q0wPF13dtuac+g30cjn6JDWkIAwSPYWu9DzUbXSuLpFXIDYo76
mIYkjJ8WJKVVCnSee/U8ehKY/R+EKyjQIt5dpxjA1+rIjMvMQxamF1RhtQ4pz5sp
BHQEgPsXnqn6gp3jydfEmOPSKdM5Xas+3pzwQjjbhUifSegnvoN/r7eByZNQpHmZ
MrFEHOTeFhjnklI92YI8B+K0e+jVLg0YfOXkV6YDERziQwsAus+M/tBgSGcklgOz
yj4VSRqr4fQhoAC++5TJayr31rn+VEzNUHjofsHjIxIUhKVV+YaDN8v+S+25dqC7
Wd+qqpOmvC1wA/Qdn0SPPw1I5HMlzZXNdgDjY4lY5F3FPt9I1/ZfIoYxv5jlot+S
acOV63TYBUVc3XD/dJdgi4UqbwJxxUX+CbmHfyEMwD03DTXlVXRFGjy25/PzfMY+
qAiJrJIbw+y23/4En1DO5dzMCEyQwGJ81EIRT05NttlSadpLLcLf6kr/n1zwPVFq
elEeiFCEEhKeZZF5yOIkoT1W0Efs0P778GPAxrZDGKtVGHtPpFMf2o2SnCz2/uET
eI4WGm/5ewxurhdl3qAHRi9NVlj4z4d9HgWEVxz4KfcdQkuvUzx9RE8ifc8ZIiKD
2mAkTdyqM07HjCYhQi4T4P0N2w06h6NKyYNhx8uG0906Gn7xV+dReBW/2KHnLsHd
cMeSMfLief7mmP3qZRtsWAPmvAlPxrIvDMec4M+CbZqy/0C38cbVicQGI7xhavwG
LEpN+uCsFjFo5u522Thv1UmifXcQHuuW0T+dHyQP0B9cRQjmmtaKrhnPFVS0F4W7
egRiLEnfS2vonTb4IIKJKBf2ehS5l0/7SJeMAyjuGicJukFqzYRF0SmIoIzmkfnu
+9oAfam/233plBqTQPl0Fla/DKcuR0xpk5LVVR4H6JdL4h6nW6GuMAyC3kPEVIXY
l0TvDsCAH+9cGVyUOtfuv9eQtIMHpOPEmlfpNBwSyCVBFoEUfPbw5qEBRRdabkDg
nS5S/OR14CqWUXMxhUYk+Ysz0+iLE7uZDb+sD3QpuUI/8UsQDMWfRo6pgSpm2n7B
xyvGBZ4nmqzn9NDK2Lzq8J2zTPBPV5BGk7LuTJ4UWw9cUL2ZwTznK10OQVoQDa9M
C2D26n7h8YDjeoYpEVeqJdSMJGaRwRnynwnL1ThLBJfKCWX6Yj12e6BxG0vZ25xN
8Ku6LxLWuuSGtvwlGr2kXP5QbpemERu9w04yWwyq2T2bam9QkqjbAYmkK4AegUDR
ekr7eatlQP2P9mbBjQ+lQ3O85Q7WT54MqmfKHJEbvt6WnB7+IucZnAGacyeAQDtP
upWG+6mohBD223Pj/GV4xjwCc0F4a5NrYP2YuXn4YxM/PC8976XP9vGAtkBnGY6G
7odkQCC7F3dTRCarFcQld9QZatHCjYWilFj4komfvJUmAKoK9Wuvi1n0eL0k5SII
ao2HNUgyCgMJn1Okb3svv9PXx3nuNU7LP5psDbueHUZKtmaoFDJNK8X4k23zzC2O
QDgqaRlqwUqcjkDvircpFcXhHoST9H2//zn3+mXsbdw=
`protect END_PROTECTED
