`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JlTLFym1vJgnhFtdtUHPIQR1zz8oRBUNoFbJRY0WaxHQWy2Kr8P+yvvT+sWXigkh
fVm5ove2IyIBPAZWVaaon9DkVCA5DbDAl0d8PYE1zDheWb3L5h9UgydilkNlOvct
z94eBAlYg5RBQXD87CuLO6DQ3ryuaf7qmbbzLURttJPgF8CMAd9kx00lHIS7gXI4
iUu+C+fECx1eUICO0SvlFNxtszVfA8AG6S4PlF30iVJ2Luzz8OHs0OQmlekW7D2P
hXU5eh+ZId2bsQLzaCf/w34gMlggHNbBYBHIH0AJvMt3ZHxUgv7SETuWzlFmZMZn
RQ9HaAi4zoSsyAVyZcCkIrT3OBR9at+04WpoeLH5ksylx8Kv3Y0htBBn59puw/bb
n2q1V8zBKs+yEJP+BOSG8RqlK+Kwf7uwyjMbN6gcOB3wJiQDWsJDRZtbEH2Gw+qJ
seiJej5cZW+CTp2AwdQ9/YjCXFAJrCeMfR6QQEtkplMzcteVrZqSC54CJ2Tk0lHK
eFWJYWwSu0RQfneyrclU81YDQoqVl2qo63dogdIHZ+d4yzELTyPNIFAeQNkbk8rZ
mfJwuFsiYDLRwVLEO01540uPGupyfHxM22LlB6zOb1WiCNkPWjvUeW/byj8CCC3U
T8FOcBbIbw8UcBcXsGPFV64OdLI7FInJUh0iRoODR5vQwi++9xAj1MmmCmNbwPdK
BPQ6zZy0ASlHnb1TV3U2ygzQFFVDYkRXfI2md11lvlPz/82lQkJJ9p7XsrBdgdOv
WAuLODNx0XjjjKGZU94Mjxh8lzmouBU96tJoEeNyeYw3aJ02xpZRvOTE08Mf9pwJ
YszC+px/NPk3iyUH2qWKGQbOPlHCHoxlA14RzHf75WyKTKJ4UkojrXy+BBNrULGf
V6j+K+xh54jxUq+h2alxh1cSPBWizvOg7cB/ZQ2BagMWKPl3y+WOoaLbEBy1+BG/
wAcg01aHPm8Ej5WzcQybaQOzQ/YTHa0cIr3T2iMJhKLCUfv1IwNk+js3PNQpDn1n
2Ktl4bNXej8HblPEjcmrv7zYNpVc62DA6twaruUMSfKWoGjvBUF1/6CAdAcsVyKr
i8f6wCOWV/S+9h7sNLCIHCE4mUEwd84MK4a54czB4Zw9kgPs6G+IWxNsRAZLoBV9
max4Zw+4OuwDVO+fGDpsgRxM/30ZSaD8hAKoPuMbnchryJ+Y9OE1YYcd+Nvwx+5j
HFTCIhxxkpQFngq+aANOFlbZx6RqveqGs9hzjF6bZC3DxhwYEATwm5Cp9exICMkK
rHjjhO6tCCwF+TgxC7qqQZF/A4JkdhXQQ8ToiRbMjOry93l/bfifQFzTusSW2Q3+
/4suHJKHjlKZdKCCVbgeab7lYDAZ/eDq/++g8LMuB9iWD4vXXh3KxsMWyxaRwY+R
nUQMET2RSXHU0UugrpQM8PFomLNTYv6av3p1zz+cusrFC7cR5KFXIHHEBfYCITqz
Uxr0odrNv+H4cLGY2EdVibj4AL9HAGI19HIoiJSuF5wNV38wESJv73goHPL7k/cc
AGO5m2y4DbUPoRtVd2muZw==
`protect END_PROTECTED
