`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RZyyauKHaPjaps+rJi+mFBk4vjgZE/7VJVmL+2hrBWKxqmBg06r5yz/mypJX9+Wn
VY/TebMSqfHkbCJOTtL0j5FHndcOA4CQdOzbi8Wsi/sHZ8E5pc/fkgvCewOYqntv
DaBheUHHbvvFe8sTe8ax2ix5F/RXKNH6SNcHmWEeCaqw3nmC7eQksywesWmDNsNO
N5UiZXuriDCqPSwoRIYlWVPeDrlxJFX+ylmcBOP0x11BQqKCGD9+hlc4IOemEVlJ
LC3xIINXgLPjrFjx1pXY944J0OOVIlOgGq3a/h0BQwsk12uqPLKqO1gJC1NSzqYB
VyNANMmSlFzvmNyLnguJ68bE05j1Rjz9wU++I3H2/TIMYSAz8V7ZXyefVTdFS2g0
Rzjtco84XrssbcTkKxSx70bzXrHP1LjXcoT+RTQtemJZSlBgnA0GcuT3P4Y770ei
4e9gef6yYsPXlPlhLIdQogBr52vmHQ4hfKN3/ocBwJD/1bFiwUTa8WJ1rLW/dRHL
H4w0ltLzVJ1l+LhrcZ+ppNFsbC/CS/BSwD6Cm3cvl+tY2Vysg2sKZW2W7UvIRVUt
byefIERhkDKB7EIO94rcCB03RVIZ+fSM1n7fsRGXe+IlSG0367G9VH9mSeePnoXu
2qM9dcmRt5B8lP/HdeE6UzJTXrMxX4Gd7rOPUy/9XjK0Hj+FcwkslRjjr43j1Zq7
`protect END_PROTECTED
