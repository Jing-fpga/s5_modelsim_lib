`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HjBI5Gretjdv/8DnSORaRh2x2cbcxPySLSvI6jmhceC+w66Y+gJEY86fEmO7HUt+
wrF6U35TPkBPmf1CDc+f4DR0fzxlaNvZfv2zwBOgjyvP8FSUzSh76YAbZyqrypnQ
XdoxTInaRKYTzdvcOa3sEXZhtdQlyyUfBqfTBjJzoBm9/BiB7QErHpazt+DQzNcG
mKTr4LhbSeDoXGjiOjkg6jtuNNlkA9SuFAbA8fmquWmF9hot/lbpPc638HGOMZI+
rmQorploBHYRR7Q6QthdDyX2vTnk88OFes/U36Kn4kG4ToAeID1YeW2e/csmeXjR
jk7VIF2prjEBNy7dtPWTsT5bq3cd/flm4pNYHIuQ8so4hVmNhurCx5h/IqQ3XWfr
VvEb0Khq88Vqge9wIQsJkdRCdrERmJCw3dwfaYWlw7rfIdw2GcKMoVLvDJ2etcXE
t6i2Itvji8LCGcsF9YTfhO4IbyJwDbIBuL+zc7C3Isap19cHEdUEd1aKCAOaCQgU
GQXMISwRlCJCg20LW5poAu3HZ0PJLMJRXYAKvbOAmDq1/r/3Sbee5pQI9wTijj7e
sh/l8RgjuYgCuWMyrP78kUNN/VwWQuhll171u4rW6em/MSPIk2zypF/ce4uynczP
1bxDHFdE/oBS3XerCj8CYxw+LmvVDX80J/p9rkUFuHrqVvOw+6xmOrUl8wI4VW/N
NeXbhZUSZ4J800vIqZFlQO2Gw9YY44Io1ZYRLpNgUAtK8B9cR+uOvC1II62ItHri
1OE1UZCjHIvQElYwOUQJH4OOEkp0dexcteIkEpqEk1Tg348C2A96iKzIbsFArkiz
D9XHA/VAsdihOU/onWTdgG0TL5MRNs8TSHMHoiCqjVbIotuPgSXWyFht5wzzE9OW
jE52s/qZd9sfEXA87wQ5cIxvirlR3LtANHZKb0P9ZD1UG70uqAzVR6dWFoVtn46D
qaK5+HXjN3N1j4rv3nWI3o/DVzDIQft+feKsyvZ9NczsTEe6eoVJGnvDDJMAUQ+a
Knbloge84INQHh/z7Km5uh5fBub8Zp8ATUvpsRXj9nUFrHV44LH1tV97T9QXqLfY
PThY6hWwc6AG3BNx3GhawwEEvgLp6dnDLkvf1QZAJIXCUIi5dff9zHqK77wVISCP
JtSAeETUhLU5mqDHIxp1+Qw7s0ByoZw8qn0Cuci4x3SX2YqpEzoSRPkJQfKzhPc3
W5mwvRZa3vaTE3vZMbfCSKNWJSFfFxZ5RR3c+2V08Tv4wuB01Nm3jt3JsOya0/Mo
8n/6+CHUv0vEtpjkZMOGjymV9FVyrYfI/s72WXgwKc0OzY/hEpNOLAyolHsCvqXd
2LAEOELwi46NrSrvSxJNkZVofgrFk7QB2EaE++8UtJIbUjwqpVncUj3ux+dwYimO
s3F6se2HS5D/MpbSqKNAVKVNXpE2tA6omFfFXWeWbBIg044Y0T94jSUU3O057TEI
/2chVMMcShWqhNT6DzRNKim+Bz1bk8xsktefgWiQlgSpr5zd/3dfAhGfxe3vyoiO
g282J/U+u1XNYyCdo7d47GWDsqgMfPgTulQzJxJhMltBx5IZuNXExvHAlghuOOVa
OELOohDwDw2R+ddUKUhmrMWR95aRECOaOWahh06/xNaj+mtQDdNNWQI32B8IfBpJ
dJqSuqtQPYJkQgxkdXEVbfJ8mfyFOMdUsVAqbLsixFk1utOjyPIrTfa/n4RMeAQH
DtXve3m9b/jeu3lyBVqaQ+RaaWVzEdVRZzfRu1vxpaRH6O4F56uAdkDFJ5U16/Pk
8Pv5fX8TWB/25H5FaMRibpPa+IO13bTBx10v73hVqjVbZsxMXo8yfHIxo4jEqtai
jJsqu2WI+xN3mohbXHtrlt8FhQsvt9H1xhscSRcTb4Qeb4SoWSsyZbO5o2Ijq7mN
OdFfk3II1DjHX1ev0AVTLXyfZ+ua+gwqghNcNfnhTpVVzHUj1s9cmwNrNuoJo066
kcbBcvz3BQMmgRlHfATyzU7sc04jhgNFOZwnojuSCv4PdwjMDCdcIvEYGL2pONgJ
pFve3FuWCLaVq7iyzR2SkH7rRZxldmr/EcRyAIRxbPjIClMUycREl2WCITekDPeu
KvzTxYHRFfPf9BZmdVwOPmHWAS/As3ECGdGTM5vzVgMd+bx4zkyAfO16cixiarAN
TVr3G4DmHupTAhpWmryjQBgYSmlxyOTf4balQtH4JgW4qXQ5rk16ewVF66Q5WzKF
xIi+9SvuAddQRQiTreDtqX8j3iOfXMJw9XK7KGVw/La26+PKS64Ey0Rfl7tCGdhU
jmWWdCQ4lnp8C0U1CE/4YlrQpxYM4JCM1KVyJr+PFZ3PNe9/b1nEx3zf7l82sNuE
POjTLspr8tdLGNnfcF0LvV6AUY3TYNY7yMPnlReVm/7E0UgmZt+A2fghPI4lFFAG
tNoJIzucL0W9NC43pvzK8saYCb//BJWcfIFmgzEd6bGXh7p4+JtDDzNHNvjHnS70
mf3VGL2NGRJoFp8k3V0pAocq1+PlIfO7olLjBX5zNc0t26PjxyML2wL9zigueIhA
FgjgxYj/UZMjjLDU6Nye5KCifD9PrKavHM2lr8Ic/KRWtKQQnIcuwvFkNydg+6xe
gsA13FPHjEwT9eSP6pB4nM42a2kAigIB5iU+WV8FqdRJp5Bw0PQG1mCbDw3kyrNF
HTQzW4ygfUXbvEgGnXY9wneFLpavaS7gd29miDpYWX1T12A1YR6knEaj51DsZy9M
IuQhxaZ6GYgbRS5Sf9Rgu6cpxg94765163Lq/hKfkMIpOSUv6FpYypiCd9BeQ95x
LzA6qOqx2eq2ueD0Zo/EhIQoFTqo3ChOUzoWOFC7VNkY8GPKExuF/BrRFjqXeU9v
xPrdfZRK6QAiQ7jgVG9OoWMfm03P88Pzdt8BLDBpiY4ZaFxwQ0rDfa3pBCg1358F
9+WtK/IkGeEDnSLTPVmBYtHwgPDzdc5pzSjMaH4v/UY6fOTmZELVUWDf7cufI6XR
2C33DX9Fa2z82SWoFAcph6507fmGGin2v/eJ9PNTdEt+58GQT6I2QERgSY8NNiOK
oqWWTnpfpd4HwmWvetLYlSz6icTn5yoz3vJ25ymEQVwg8gZhT6UrMeuTD4/e1inL
fggl/2ah64cG8jRPlxt2U+CTpoBPa8ANpKsQlIpe8HEfi1r0X6l5uAhNfjVfp8pA
tIaue3nDfIo3SGnrfNBCzYn0RIf0KrCmKz0OWR5w1uWPGGpbdXkRgS6dWXGJSPZB
QZcWUOaCjhpCthTDS8VMYZJZL19wesSuTZ8D4tqc1RKwd95IKBXzBX/KNkARzZs3
HEZ74kZqeE49do7OHqe1HVG0+wxF+6ad2DvjJiZJm0tWPqFQYDda+CGjLI37D/yl
EkaHDd5b3Xg2DMYNSYKrRtFnBfEgmQbm3ZHlBDlGTPJ9FYXSYAArrMEqsJ5MEilj
rf/eUu8WLM169aO0ourFgBiFhJiDjwfnISgBaLX77dBuIvG16i7ROBmXCQiJ+FYW
wWtdpkQr1IQVLNFAU7EMuvwMin6DSxZxajIxRz7qid+O9SzzEwT0U/6V1FUux/Mb
8GxSmQeEZ6JQNCo+4i0ezu/vBx67Ft3JPnS94b667VhUX0lv7Un9If/4LHoF9Nn+
+WIbpq45ftn4MBm8KoogCSzDJQMuhaGjNm2YOXsgq2rwQa53Qj9XDWBsJ/2h162y
rxDr8cC7EaIZQj4C9fhTmNiW/2uWOGOrjIIb+MsThdbYGCz2t+vrDzDuKbbskCls
O/bDzAHVfjbNvrJUyvPN+tSGs7zeNFEOG7zgVzt+1kKDMv2eg3uKNJCXKSU9FnBE
4tFjjdAAdFHnIj2LVGNW0rBi6rXi2R/ICvmla7GM1vNseCHOjUDSx0bvSMDAiFZx
8LDat7Tpj79y8ST6Ux1kZIHlPrx/XUeSf3EMTbbsRBSdmwJHL6wJfcVq8nXQSeFl
FCqmuwzsznbrXgitIEAgk1W+xE+bmgZu0WOPSxTbq0LdqZAvOi/Bc0BhTvKYsR/q
kwXOR+jEUj3L7+jOmR6q+3bXJrCwwcfsb7ejW3WGoXPv1Y6lC23WxZSkySfxktNI
by5mmyDvDdLU0ioJhXJKuZOpiZlFUW2AQvBZvQF7I39AOvGA8qYbCCfUj2SNkto5
Eo35ANC6m3eDio3yxTMcTNB3bPisj46zuF9mm7Ql+cL+8IDGyOIkaYXzt1CXVJtQ
z2vT6sSnB6z3sIda4fl+uJzI34eQLTa3SHTF5ufgGHVCcFzaWR9FaG1Lj5XC7yAt
DFta87wbtIvKaygSHga+J44e0rDDhEAhEjRq2HTqcbY0GOdVGN2Ra9JDkgk2i9X/
l5Im+QpX55qKUMtfe1pthrUdveLBXBHEl9h86sd7r2KnvA7q6+Zrw5UHkhkzzOOy
8bQOBDNnUPsB1yUtoMXQvPv6Y9qVeakQE4qs5YLXI6kSaeakyE2lSpddi8I2jhU4
V1x0Nb331kjS3tjqNMG+HzfLnhqpGGzCm1GmFQo7DyI0bsaiwraIFq/sAP3c/vcz
Hm0q4srRWm3TdsfDM9Qo3Fl+Q4s52n/Cnf31JXIIT/DX4CJgELwy+B0SCHTrJJYd
1gZfb/B66h5NCDccI5LCzp5xyzDd2KqqX/NINoLkKug9tGY/xAHuDwv0GwqfpZvY
dLzGNJUAaVZtnizfKKBjwe1hRjkNH3ZsEIE3+M9fLYd0xamkXo49+D/GBI9DIpYl
WsAIXd0SqzrYiD6o1B/tsPM2xZ9gkiiyDccA6jjHR77e+m8Qy39/RXjkGzdfX7bX
ySvM7raty8C126Atnf70FlIn7s/A5SjoxRaKv+CbPP3JPwXn7SPkWsYq8LB//rb2
4/zInTmXIU35AwHTCG6rCyeXdx3kZ0eue0qXF0h1sMKobcRcWyqWj0svJ66G4TgJ
beJdjIMxp8cudT8qFVzxQD61wyZAcIS+/rYc/gKcV2ryY1iI8C5qbPsnNiNUohYJ
+Thcc0Y+g0R8qYphwyXR2AtTLOKde1B6e9Qp3Rxy2QvZpMxfeG8+byr0XEtG9Vtf
U6mjtJBDlwgg5Ig+7QLSF08nZGXoDko4hiTDKqd9RQyE8PJpp3cz1Ets/uA+XgIw
HkoI6cMNjyVQ8llYl6XxNrGdm4kM/sMK2VpGaE7qyzn/c8hWUQV+jL/yDgjZYSNa
gFBlm9ZhBS3X+57kjEo49VmvHXEowVDwpvEezv3DBQm7lmUi7OzM3nl7ItD7zQ8o
vQClNvqWYJgdSOFX1IjpOvGIx5YZtDN/l73SgRzJjq9M7QK/iLzz5d1ZlmTMnfJt
e8GhCTV+xRXsPxvyLY9e1P+v9ai5Y2jx2c+Lvg4d/sbYahqDznBqNy//RkwrpiCG
AByi2PoWCPUPkZVJGKEKJ+Wrxq9ro+UTnxjguujIooKFuLh1/HZpbBKftBMbToxw
22M/zWWu9UeuuPkDi1dTmjVzbMJTsYCMpFDic6hUmYYqvg2QAD9JeyeWBwYzN1b0
imHdoJhhAn4qFtzRXEBuiHdsu0mPEIkf6xxgn9j5VmOHFqbKD9lqWGeM8yRscCvy
rKvBVq7cXdSr3CsSNnlcHSZjHJh68vfI0pYOOToonAyrjUjopqmd9lol/SaB0k26
nmohIEnMveKdaJ6H+rl0bUMNMArTtUmmgQZRvpPeZpgdetiUGCe6ub459EM8ahmM
7RLXlnknhQQY5a82rtXqLlnqFK6lQG23PNIw2SC+rZZklP6E8P4ki0ZcoLBgj8hR
u/YnCmtSA31iY4z5vRf3D+zY1a+oCzZ4YSFoCPDbf1P4Srry6AZG41Zk3adlZSwx
Uxzq5W+290eP1hBxWotobusz+wenurCyjM1ghpim9FHCz7FkLjTvrw0xcQPetgal
4ILrLs9NLV00eUN1PA/AkE/uyN4lHuOEdcHRdAE+UPgDL1jKiZnPZaHsda/y2ddr
OswImiwzSCkimGcHMKxTlcukyI68dd+S5Tb15Sv2AYfkYPOzHfkzqPK7Tu5Fi13w
rJMvmSkDR9KMkpFrOM83I3yEMDg6avjsUVyz69025EfHqvsCCbe5ncNX/kZQz0cP
dNXM5PSWw02uXiozzXAXIJltxzk9TA8d/RLEj/vITlmCOxHpaurUcmLW5Are/VhX
LlTPClufM4PvP6H72jddqMGfliwiSn99w3astFpQbI4z7XCBp6tNnoV5cQirDTae
NpsKviAeIVKdQ4tiWh7cozPWY9S7sNBM95GHnBKYiddnvooRBnnyvbyL2oNN7iKM
3wnnBAo71WTsH+U8uwaXrN8bj1GWkYZk1ISsjvMDcLRgCSgCU+urjKqb1zHhEMur
xAopGgwl684MyemntKojdU97Co0Q+Y1IAR8/Q9A0PKV7Skja9tmv1Aqq+rMGALmx
g5/ALINchLJIpbs0N9TBjQ08zzPcUHqoB/8Po59GuvGzDXRnE4d0pX9eV4sv7t4m
pRJsXSM+9Ezw1w9Ec1mjgld5b4U25LkuUeIEH/js5t+CyCG3JqavlpILfWav7I7T
g16Zf86LysUAvpcr8ftwDiVvw8Qc584Mr7sexCvf1k8k6g/VsUaYcv0mNuJO3wpR
WbD9u/z49/uYz8RiRUKprq/9Z8e6x2Gf5kg3FnuwgfnywLvZpBV7qU33lrLjBCOz
a/YhrG2pcI/nBP/5SiusCi+zEOFKVN/w14qirumJHfhKRyu1cFXnr5Z8jJsqIwSv
r6Il9XwTKj1n7ErMcwV93GGhD3p7gFg8RiD0CoAuGgV/yPdSGsFHbp9DNu4A/B1u
HPPxHSPJqr8U/bBsetwfE4if5aKTOJhH5/m2EdmhWP1kxZLZ8dx5/RiG/WROChP0
veGk4kV26rr+I8VP6c+MYQVdo1yvdHueCrkeK2faKpOb+K1R611MIiRrJ4/dR2CA
AuVOaFWiHuIApv9lVFcK6WA6zufScViXx83Zygjtc2YDZmXVgsXVA5O/NUgt5epm
PCgcbhr0WkMJauX5AudowMTF7MrBgGnnlSfLWg/RmJflKhJiWI0CmgeSJSL1rl4O
DmXJ1qVqLtYhkNsBmEXfs6LkdtRkkDowCzbMSTyy3ddK8AE330RKs2aiZyXYXEJw
ssaMRke2iExyor3hT8P/Slqc5WtVxU+Q755cHVLDvUWxFqxbzocEMntBAIEheJYX
1nTpn2us4OTSU79TrOV6at5eDKSZtyPPm5dOz3+6IT1QiIuN0Qe8pNDK2ffA7ULb
uoyodU4JnKyY3cXoxVNPJrO+Os55MRvjMRx+rIOVGq3IAtXnnqt4bsUpd1ZYRV5y
RlF7FwSWntAGbMb2JfdpnN8pQ2bvlBICx0rVv2B0QZ9Wo9/Vx4DUz+4c0ojg25pK
STZ17KTxpfXQ6umxu6ogAjc1W80R0P8ZdeygNgi5xBDx294PhsNNbsuzHCxPMTow
Kud6BHMHt5oQsUI1agZwbPdVha1KBLOsaVXC5UbMJlGkS5vqtb9vsUueSBfMF2AT
dqLw4vomtntv5kMZziNQEPL8mpbQ1Q4OiYGDj1Cda522lqT5u0eLYPNchHF4jZ3f
Ubq+B9qeygvyLPr78Tsw8Fmvaf42gsh22V/LzFm2LQSPIh9lWy7iJDA5xe1rPqhj
AUMCtimhpCV4RH7n3LO16249VZUnJbd7y3Gai6Etc3Xr6Zi9ZDz4Tgy9wItLBco7
L26WsJrnJggp6TZNKugdm1luoccrZ1BG1eC64+T7Td5vXc9cBWJkIP3oO0ZtfP5t
TmvIMER4Wv/coTV3/aKpeQto54ld3L4v2kEdjaa7iULvV+Cn3zMtOnOSSUBpxD+O
nQHdgUeyNLVnNev3g2Qg5KdYcbC3GawvVxonkKf1yMWIykKDwC/Gs/rf2Ye+H28k
z+eiKJebPMa2XRyd7WoHYWEVBuEW7gGIHl7xp35W3jMBFHAYCVJPqsVfhpVzaxsN
emFAI/EXLV4Yv3iEC66j1R+KGrswyctDmTyxGi9KvH0mi/L174/76+nZIn9K3PZ7
M8g1OY7Ga0thFg5Ha+qkyoTW+Gfw/Fu53XBv5r09BFi3WLrJbtyeJwoXFzKcNgLG
bhoqbGKe9bwgNm+LZSwAGnfHi73qHsAF++Jxq5NjOvH22YPts+xXFjsymALFVCob
HCFhFfEWeVxj0ZthElHslQAXKDE3x+H6QSS9mkS6sTn9iYvWLkbHucSCE0Qk8SJZ
hNxzllhy/t/6QPj1GwipnPlNZcyzNAU8q/duRQ7sZ4JjpVn4w5RJpfNKv9HcTwng
f+x6eaE0WQAYgru9LTHRB/v0dlByCE9CSlmxOqGnG/I2M865+B27ps7fo1jAhJEO
TYfo2zWAhZgKoQGlR955ZPaWksPfg8Z+AMDoSmVk0RN2liX9vu7sz5Zq2HX5jKUq
/hAKo0M+Z8Q0glycB00SfNMqt5K+wUEmzQywkIK5Rn7os0rI42OFsloTmPeYmhph
UdzpA4GSbCfv6qRhMCpcqoYPc4fZnU/jD7NpAbqkRtxtW9n0hU3YJ7gV5ygQYlCT
qcK6V68ayBoibNl8f0woGZ9S8V/96PeTKGPlFLg2kGLdi8AdgBT5Ap74D1+98YGj
HzN/Z0m8N0dgCK7XtVxbqbfqVlbRu68ykYKuk2HIMl1ZeNf3/D6y08VePeTRQotR
U9FSVleSI+YfLrUDh2avCTZWJJ4wusRVfCgjK76dEYaZQA435qCykpu35ErnnLAN
zKS+P23x8VrZgbeo20OsSLktUB94lKvy5eHAxs4og6AlHx/vl0JgUxTFYYNQOJnW
BzWPGFtAgGirnupR+7juux0CFr8DxAtwfBmnc/D3jDqhQIM45KK+04gktlWPwwKk
CMXIkufdOrr6X6+ONocorV2+V8LmQpmvOHhYTwJu0mVZL+RnuLNkyWH1gX+Ak+GA
SMKy/UZ/3HCwBHSPm7s7ZirVHm8oIknyQNqWKhi3OjkIsJRxFLsfqI6QZhWaqqlI
d5+yZfas4rFFKNlE5rt0J7M5ArFmWWqJZZ6f5SisfrsQM/tQNCLxnKjhelkfDtAM
BkifIa3GqJ8UzW+7Q0/warVSYOBBgPUViilX/0fLqnM/v6qqZOUr7PtH04EPp/Ct
qm80o1dTxKFlNg7wyQh5kMX0g8AgZy0G4/56FAnbJCrRzzmh7S+6oUJE2OSoJK10
+76JgkVd/r+0BIDWhJMytNarcwOdsbK0Gotuf2WAl22YgWjGudbVENjMYg6XLyfW
XYGFeC1JVDDHUp132STgqg2hooJxFrZZMDYhOBxYqrbFRM17mbzCTHncp82Bz0WO
45WX3GbccN/mhRNhZTMAIPnfX+AJTF5dbZKGXExFx+2gYL9vawjngx/PiqEkuZbY
YTtT+nyZTotuz+7FeUNddzsdp/ggEND1HzM+UzzUUqzjYO6npU9t4eTM1dG16bF9
qMAlQpHlsPsC0biLvVpRBEO4okaseyAOGUkJLBGaaZcax5BQkGT8cfpDQvlE5i/Z
OmGvVeIMjOwIQXxG8iCBoB3lyIOD8Y8bCrjM9oNMBrP03Q9JQi+qimgkyiwl6ZMt
cBaCig6v3jWFuofI8Nh5DtVgrU+HGxNg7QXkWZKNZkNMXfVTv6MiMUR0endgq3Ok
qvdr22U/F2XLQYgm0LPqbW8RhrN9grEmSFe8g+OI1vMHGJRPV7NtFgDJVVRILxRm
VfgGJSPCTDE+dDoIftDwBpGkYiS4OLOAP3xgogjC4XjccejJK8aIZ/PxXWimht6U
u4IgUTrAlFWFm96eAPvG280tFDPgnCY4keP3UVYMJHaFBUjyBkd3M5vBgwaDKRz9
lTdCHxdhJlpKSdpt4V0Z4CJBMPlpXPta+8wuUQ0JJy4c8atV9O9oexKG4r34ehB6
fYtiC932dGGGNCyf3H3YzZK687IV/dvMrSGBu3NCSc+oRBTCnPjHrzJ8TzCJWXeb
1icI3Kq+AaWeC7916PVSL+U/CefFa2I6WPGn0g1zWub/o9vOK9Tvgp8nLKvhhF6H
sX119jAjUUWs8go2JhHce3tw4BXU+bL0rVCG+RrfauOk1bkh4D0afxYkEzXwmtPG
+yRomJeUmD42t8TlkmD/DEANW0WcQj5OhFiMmYm9Oa+aA5nLm+tqZ5sywrmKJYjD
L+QLBReDanjOK0R6Jvu5KeTUi1oES6KCGbebZUGVj5xybVBuBhW/lf+Oh/MDoYYX
amxvvvgFNZuTW0WKlYpsy5QbDMJKJNITjf4PrllrcRzpQn5HDp530gP3LDfu2Mt+
BeGnbOC0dOrWdPIBLiMZQMaymmmVjlhzqdu+bOQzoqXZv/fAAGtziyiMWCLlf6Ta
y4E5hgz8Fk0eX7KvClsakkFWCRLdtcabQg+mIcWutTbqIAk8bOgAlV5c8AyRInU4
XbOd3SfzOpjCO46c1pVYCLVjSwJZfse8wJbJW5y1Q5A95jnbozv3pb6CN/05emeS
Yiydhl8JxhJVDQmhp5LlAS4w5qsniiOY8okwkQ8Kofn2+bChtJhDrZTdNRmFft/A
QWvpEX5rqs6/FWo3M7w/PQZKIhHYSvDAe4ipA21zH+BfL2XoUSnUVxOiBAbYoDXf
wxAroGtMvTBsD6B4pUl4l3uNiJxRDqMytj2rGgmxIutx/yMz7hoz1s3fNtmhTPLq
CEuUF+IMovhaQfjtqvb1zkjOkUg5++3Mwe8qtgvuwNok+e49O532PjjFjazWdLNs
TDBTRs7tzCMq427wPyQ1kspVqLfRvGhi93FfpwtgNPOejyxcpkDEIIJA1kPfN7in
TiplHp/PsIaqdRDlkyTjEpJT2fJRmdUc9ItSjUNvCWlwSbuFPAaMmVSnPT49uHcN
YiR7O8f0gzYpZxKa4Cc3fTYJ5uxu5W5S7Z8116QMJojRzVkzSHrwASU4gFIgfldf
y77l5IQS4emoJHIf/4adPJROAZWyURWo0vQpnMW5YBx5mAqFGs4N7FROV7UQxMlk
EVBZbhxK4U81pfrJs5bh38rxfBwL1rtAH6veDlFeMQGYfa8xuntY3/sL8OKIqH/T
uwR4AEAGqBzDdsL880RzFb2sXp2NP+ZnRJVKUen2E5XCB57Tno2D39cQtnz6EhCz
LBLeznZYeiIzACdiz7yC4SFHL8s0ekQxm6/L79oA6iyJf2uZe/SzZyl2fFk9iWUQ
0nGgawjFi6JLRWk9wo0u+rOzu2mTHRLNt37NU6y+0/i9cq6cAKgRsDEwTp9fgX8Y
/DXBum1ukziYIjArbc5sHLqczxUIgGoDICS/bq9h23vWnJufZrGcjjTY6xAlKrRv
92VbHSlidAA+XSiLxCCD1RLJ4De9MhinnVNYu4yf6VEL/uRWUpmSOCzO3PeU07bM
IUmdH1dvXaMP/Opi43PD4+EXZXATmNu9oFhiMhygEqXj4ZW+z5QEIO7DAta6QSTh
3GsjePQWPi8SID4+cZ/6H3WGnIQRXddYD8GmrazLa4qg6nvLWkxVqGfBF132UEKw
mXBtuSIhH49W7auwM6VentabqWR0n2wVW9i+1UhDPvgZ+WdO7SDF6eWIv2+pTHbA
Cz/cWhasz8tMQ9hbBAULk/+5/Kq5d++i9Yey/LQJcOjTfdL1WZH6z4QsB6JL29Ku
N9rTFW3fZLM9ilKZ/UsjMUW5l0D2PZ2P69e3cNR3AtIoWZZFUAWAH/hHBdqsbrFO
zuuvze1CF8JvqlYXnG8HaSm/9dS7lNpjpynBnsfBFBegr5H37o24n74nWKkfZwyk
I6k/RXO5yZ5XtNJ44X/hv63g6brWSGUHXM0UqMBv8vU1xo8O4lsCzckjHlKuH1Z1
UyCHJ9BQPF3a9bbbzRqdq2YMWkmbGu/OPQwV4WSNCls1BSI06Al1+uvXiUnhPYLV
9C6uDcJCEshQ0+26PS7xQluwzuIQ/15FhFHWKgei8iPSytYdjq7sLwMMVcy9K8sA
PKY+vdvlX4rU+ChdOeEAkVw1XsInTQ8s/0R+xKlTgQz7cH784ow/ZzEMeY4hKYX9
LZxm87+cec5JKKX5/gQtVQ3Ie4XcTmjMfPHbHFfmZiX3ao+FVrua0CG6QVWCz2wp
9hSpeYpTyKmMgk7mMr9UarVfeGltYO+ULxic/tBrmgukWNtfRRGTAMBPiXfTEo6m
QYXqzcHqBuJpKgh3qs3yngt7T3lY/09pQOe56u1XXij4hGZhYtJ6gbzRIJ1+xTTQ
WVvl5j8NWnYiPNQ3jG2HxK7OLfm5m4RReQ6ZmCNGAJeP5V1V4Kr52yNfduVcC+sL
vyT9fWwCWSQa4Pe5nhstboWqW9LlPuxC9nrrEhjDZsJ39xDxg6IYNU1G2I62rGb9
q/ZoquzAXp3EzwVa3a5ddrHEKl9vqfSiaBxnpt/+5/byEyFQRQhU91Lh6Z25SD4q
+ikOZWAjRweav9tA/2fHRwF2VZCzeYrbEYfy04mnYnRSa27cd5tb0VuXyCnX/pbc
+Pg074cEzXC+XzKFrV+6saCzIJVxN9G9Goq5qNe1J6AU8rqFZx2utCYtfd+a4qi/
ohxYHol0TyMUMRruiBPkrzYoVv9u6q1x7RW/Zbf/zawoYvpTvcqzDWOU5PWGx2hG
9Uw07ZPHDXwc9WOtKMSMHnGZ+Tt6VD0yNmn2meba5R6nDc+VBlGQnv+n4f497vv2
zRlcgdAuElYeRMwS0WaUqaiDCbnS1DbR0UNZojStpfKrOeAPJCK9711AlZdOgzwe
0kWi2kEoeq7KKeaLPTp6Vz5Cmq+ueXu3th/Nz+W6klH+MJVeNUJDZrBbI7Pb4GLJ
8W60crLE9e7YvcD28Vb6dKoSAYR7ZhfYEv6LKKci84VlFvIxu8/4Pd0ehJswdbXh
GO2eO8rSVMJQwBNfOiL2UhH/HAWw9vXtb6uvCa6+W7WKl+/nZRQbPePIY9gs27Ja
2enR8rHNX+A9brPDMMjaA23f9WLEy1Fd155jxG53IVLjc7GREVJLoSBI66UWWpRM
1zigaPIpbvUVUeotHS2U2+5TmF5o2lAtQzIpP33bYMqiD3BQpJIBHmwAb9n0aVdM
JgEGow3DBWOiD5FxZwOwi/N7k96c/Cd4bdUS1WgLmkspRbTnSKtoIUL+/LjaSfHp
tKxLAdqvLKlHLt3kdSW8eKIQF94VGwb+z71eHahhtOlODYp2oyDRrDgNHLYCYmES
+Ue9nuZOAfQgmC22zT6oqg3fwoIgzP0sbxT8xm9j/STSlbHd2+6LhXC6SKZMw4FE
/FF/61gj1D6p3g1+gBNtOPCU3kihLeWsX0Pya7UZWLSMXMbS7eQtMv3Lf8Tp0o8s
GrugRcd7D8TUzKosTFETT1JcWdpZeDrssEFo/mY1AZpziIckV3hgNsxnMtPj42pv
vO3UrLyeSRCbTPsLurYsnA==
`protect END_PROTECTED
