`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hBpmy/1imk/SDhxNUtujTQRuClZZ2lVdOhXNaP6nUKjuNaJf577Hhdx8hKIr5Kuc
kXC1TKNl3NzS+cnXYB4l1KzjTFmaTcia3Nbp/U2nlGRlBT6AUTvN9FrGKYLs215z
r/YlkhpzeEEPo/19WScH0H0QGmG6s8FE9VyNtfy/YYDXRRYpP+MO0XArXfKJLOEf
T5mhC4BD5yjbtDtlOA5sSAArxVvXeOgmspXVml1kylu7fKa3LnVQlN09n2pPdztT
zTQRbUleK0fWrsb8O6jfekzSkfuNeVCSq3OSMFkzo2uXgrh8mswqZPnHEWHew5f2
O2KZQdbT+2AZFQJiIIsexDia1UwUDpXziChx6bICKr+JolgptoqVjrL/asGqpeda
qX0HaVkJ7MA1zkE0NBpEIKckRShIkzEt4+bzBwXpFB0jf09uF8F86WYgxFn7D6O6
e/Chk356ylAAfvxe5CbwY2qHwMBvxguUDvHkRvZfDcaOQ2p/LWU0nqVAEc1NQSEK
TqOvjMQsRVYByQl+PzF4RF9+UwcFfDywNnhWBi748g7nUaa9Uhalgfh6wxKXqD13
+wOz59ahKJzIOwrj/fb0rEEkJlnVj0HpF4UI//9jhXhoCKWFGpKyyql53qqY1b2+
fgMg9v2P1Dt1SH5sjA7L9sE+3GuIpa4fJ1YtuznNAICHA/K2DnuoCUW0uheoAO5t
cMqevU1u/oh2wN3Hkm6mqf6Bv+qqJyHlFaRFJU/tkwV9E3tY6Bw8wlSudyaqbc6k
HkvJ/MlyooQkttkn/a4lI1MrLetnIoqZxq0yqvBcDG9klE969rZfSYVRooIZEj/f
SprFOtBE/xJEz0udcajbOx/PhBBRw75XyL4lzlmgPM05dEkL+X/vUzMztFej/Vbt
WDbhf/UJRjr1lH2m3xVq4wZ0ZoB0mfXwFEIXvg4DoD8WsRKM6OR37dwOPv7HxCHj
WjHX9w6S5J7/T19rX/tHcbvqIh2nxFWReF45/LK+3xrIKg2HiOh+z25+GKcRgXYZ
Qi+4Oc5K8eKic7IJC/fbK3RAuOGzqIvoJJALV6g3JI5vx25IAEKVRMzn+bhfw8pK
QYzig+QiO0PDH13wkx+ahLImCYI85GRbFykvnwtbWL46dzsQhHsuTOxgWONLHwWL
XgZ8ORGqGuesjVeObHZnCwOGfwwNVNRuOy/xYoZnGm5cdnD0sVXXfL9WSbw/Mr5s
ms5h0S618piMV4TfbQqH0CcyuxDX9FHCb+Iyk9eDqc/L0RDdWjEq5NhWzrBY6TUr
KypxyHQQO9gacmLQEiO04nV1EW6NBOiRz7K3AVplNGh2d/O0xE0ObeuGfn6xyvZ7
u5PgRk6xZLsREwVoNx9hkMlgtvfPok4ArvYXiFP/ksDnjwsWINQCV1NI10euq+L9
C1B4vI/wMerChlEfoOLoOJe1uFp2aRL1pyV1NEqCbo7hQTkRpBQBW/tYdD0GIPji
kIE7AuJ1Nc+3vcPWVh/vome7zUwtDiBeO2aT0Ar/WTg=
`protect END_PROTECTED
