`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q94uxIV2+OfsPyOxvy3QD05LGLQdYyPwvhUXvafT7yzq9WVfZXoYK0xB9G2OaVJx
azexySuxQKXB4v/qa1WHQbEZqRnOrvCIP6y4ViEUfUlvn/4qJr8Pb1JzG+CdikcO
dRc/WC6WeKukcOWftXKKt13UnxqRCPJRf27LQmNP6J7TFlmpNJqw3vhvYH9qjppc
dxeEySTYCqv5zRZz8zKR9D+6PeI9ivZPwJf0CgQZJwsku7QNyMxxjIoynQmd7lPK
4LMgT90R2zsdorQQhSakmZ7jS+ri2H0k5FsGEbwh3UUmQvGtxToJAhDvm1VAQy1T
9p2IevhrUKUffdIkhDpyCi5WuQUUafhKGiPGRb7SR7C8V5sWnzonM5pNkMXPPaWv
VM26qZcLPB5mAl2/NUDiE6GNohhvdfJwGLbh5LGPWQrbW7ELI2KA2Clm1U2t6MVW
TcMp0wT7fK/Zz/DG2SNHLwQ18eBcC58ZmTm9mlgh0w/nUw/F7K1Cg3rZ8ASroJdq
56QwwxOr67PTMKuVgmVU+yR4pllnFV1MCwWCbuGGBpIVNKK/l/42b/Lw6iR684e0
7xgZfCTZ5UbuxX1DpvKsAWWvLZ/1Fvo1sNnYTGNcFDbMshkC4uEVXe5SBQOJH+bs
VS9/WGNPS3mLRVOBagBvWaLpZ1cbuEgKI7eBe4EhARiMNo09MXcipsQ+p7hPOC7z
nU0lp+biwRfHSUYsRHy84XGaBufVGBym2fSTxeZZVUT95RytzCXvV8TsjE2dxDHu
2pkZnxzMlURCm4QFO5Yi0YcMiD1FWrO9hIQ45i2xrcOJwl2/9rceyKsgIVVQ871a
yhYhjSmCS/Tb3/uoNlKBIj7bCI1UxuUPO2p3MEgyCeuj3FDBeY9JvCyB28GCUypI
XS29EmKNMIV+kNprc121g6vbKJt69lIfXkjgTTWsyT5k+oV8ftk73j5wSZ4j/Kqu
cu9Eq8irKn3uMsYMwqQF8oRxMtl0BaYorqJldFZFlviTekDVDfFpqn2CyiTznjo8
f4D4Z1sNjaFUvEZOJYRPMtD8s80CPK8DbI+rjl+tb0ucAdHrc+yog/5HxitoY2Oh
ydiDTrgMqMJZVQHSmcu4GBn7Y5PuhZ//eDGpFmYh0kPo1EM3z75suySGU0Z4sEIL
/Zh8gz+mdKIpuycgUFWdMwU6W9c8AEUkVZOgRBshM/9Qrm6bV+GKZpCrx9/OjHoQ
rPsMIaJxM1l5anjm2wYAwfIxPgxdjEAulTtOvIqaw42ZD92AM2vBHejf5ISQspFc
bx/AYOsCXO5718MgaBsAmpitdfSOzuh3VtuWJVkVYPEt7o0OvQ/ixXs/pMRHUE5s
9A8DiAjDnJ2toJLoNBQywMwRhicWIxGP8NqH+cpGUmu3gI06sNOC1HX+3XhpgIdE
KvgDJN7BU/stSwLVpvuKN2Yed8xcESQ+4CswlmmyxddRkl00qhNvzghadT/1Kise
YfRn+OTrrthmusjctO0pW4Itq6KcRN4Cm4mex9AenRjiOJtJM1hQXdEPsswlg8sN
pDLqXdD8r4qFJR2gdcqwcR+tN450Ry1Jr/o9YUVYwDnNaMw4uVFyXkngDYdxk26o
KRpncOFfyFjO6HS63zaJmYyFx9xyxWFmHzF9cAVWi2uTJPszqjQtB1fa4sCysa3A
iUmkBR0z3Ap0WmPUkE42AvmI1utKeRjO33Gh3IIkqElLAuzTP1gqpxa0z2f1WvlJ
BTRMKzjqe3luCykHb0XR0w==
`protect END_PROTECTED
