`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2AbTymeK4DfTS1FI9KfMBZ1ujV25H3XTMQ47O5zHxqaQqaPeYbhjVxOm+kLnqu3t
bItSFlnJcAEMlcIoFzsfaotTNzdpi9n03gXulYu082J7gierBOJ/tXlEdkfDu8G4
0IuX9zRnpau4n+sZStXt9L4gko/yIOLkl1SMa7At46mS+00u8H0QPAWwImfxgiFR
8de3UEWcoAls9EhSbStZReFxU1I7C89V14VjpWnb8xiZZ3zJTSpke6YByIi3eNt4
t/nzTgmeRcntnbwrHR5HB8oSK3gGWJuXQnMaepZFmx7InTTexF+Q11FLsaoVMh1q
+sDxV0kT07UxTjATSiVGj9vy+Vqw0sQHFetjNtfOFZi5eRwYL17Rj4Io/8Wkz+4K
FvV8VHdg4YMBPF4DgFKL5BUP0NLz7igJfHFBV+djG/sy4qY0rdTUP6BRIRRQKpz3
LTxkjVXW4wDhTSKkFV8BSBMSzBwW2PJ21LDZfkIahpq5PqPZla6Hx0EAiHUUJtz0
uOUZhoBVYP5j2RqWfaun+5QqT7h0C+39UU4M2Erwcq35MKE4qbvCW4vppfid1ZNy
lIQIDtutUozFvU0KnsLxxOHMWGrdty21WLdNdvEw3Ow1+t3tKWHxG2xNOlpFUMnE
PRez87dTYqbgGjT9p1lq53P4MQ5fCwsJWcZUIaMW44wkpz1V7PHXouvzR4lOxqRf
zy7RIbgB2LOfedIAW+ae920e7ntnR6ztye7plvLwP9ebXiRpCw7XF4JiLo5VsFyP
TQM85mGRtkp5xI0+oCDzTkHQwg4tZwn6etp5XYr/zlhSqTeabKndC6N1tM/20uEF
zUX36rSbJiDJcBqREvO0s5ppYf8daveRoMdiRL3zOaEDB8CkJhTWDPoC38XA5G07
GvvXw+JKF/+VhblyXwVSkqnGs0UPsThh1zQ8IQVT42c8iqaHn82J3jxoJobZeJfL
oApf4Sm4fvYrCb1zXJ/E8FICTlWs30CCZI5KK8U6NvPwaio1igZ3p1QdbYB5Hr8j
cV4AL/1Vl6XlJDBAi0rGHUBT3aWuGCdjAg0vlgPYQhAw8e27hq7TzoiBjhn45DiN
yYG8dgrtvq/2K6j/kHbn6wdAZ3vFrem/v+tlBMAdN1+TfTv18E00LV4gOvj5jYNO
wBJwzV9nk85+iyct3GNQsPG6nH0DxO82N02Gyu2wwjRCp8k9rKuFVo+OjaoAgL9h
/Tp6kRXB+WBEqWKcQ9vGojoPp93KVyzQA3iA+D0Wo1mE2kxCc8N4AGGm6fEEN4KT
sB6AI0n5PWoAnE31LJyPft2HdY47GgP8i+akRS1phS//JSL6O9dQQgTwrj0cuzmP
m4NO7cVWuWYmT5SP+hadxlLKPm0dSXORj5kPK0t0vVtwevody4tWnMFov6p1nopB
k2rjLGpymFPUk4iz+IGbqAXQvwNHFguWl97ZmGVSyDh96Dp6I8C0zQqsmq6Mvwym
rEPwYALD4Axj7QksphvuUho9H/MGYnOermsZmksh2aP0WfLbXMBMY5Bk/i5Prq7h
8/gSMjM58EtoL7FK1kpYcL/8b8jEW7/mRA+79R68cxJpssv96/9K3UXyso00d1I1
CbF4ZrNCTghlt2wnycKpJkSb5nuS5rx0gQJZJbZClk5rtoMWGsePWk68c0vOA+wW
V2ZOkQC/Dwc9CoM0TJ+GgVzWDV9nD3QqAiMKx6CIWPnMOMftevrdTLNEOGa19EPN
NCiPkCzWyVMUEvjlUoGypjfRo/xU1tXn5i+kcJ4THSnSNnTMxrOmZ7liDVffnmRX
TlJnfIq6VCXbm/74P4OWGh8wOJLuyTmsVnR+m9aVNBjApzNbs3bhgLbiPqpj9ocL
ur1Mq6reieE/p/PI5inO9Koc927f2Z1sanEt8hX6+zjaqt8sU8pP9fmtb1tUAuGU
p/x+iKS8dXFdwXI+MmrxrwB7fhU5gazxd5GS6hcsazWk1LJiXBMb7ZlJiJr8lChl
kzXSjnIC+t/S3/K85jjCtiQjQB1wDn2VqmeU/8p2XpSk9VlPmPpPDHTNqUF+lBJz
fCVUMwnJW4hLI63kdVVkPb18WOnRWTV6ig2Nfsdo4upEpXroYKPmUbuO+8NkBW81
ZNbHCAR9sh5llOjvhk59h7yJTPQ68Bj8yXAgV2bfvMrFWSvEk5voj5gnORVCRLCV
sA8cKPXHBwrJYmGi4D+mNKyQGa99d6lyRcQt14KptiTEZQYakyi/u525cS7+FQTo
bBa5HdxNqv2oKfSrSBut+KdJSHooKTi/3YNy2+ic4wqBrWv1OesYt3KCoR6Slh23
qdG1tpI4AQfCltwUcxs4JpXtaaV5ruiW2LKc+vUoP7m4OGnRi1TD/4aA8U2xjFF7
ifB4jBku6VUefbCiErxp+PWwJ4Z1mRClLUo4wMP1C6TU2PNsA7F2fQZA9FPysOyr
Y+7GpLcLprFZV+trLrOsKlhDLAiW4o+PmLTSeFaHy7iUI3+LrdtBxfKuZQzTpn5I
06yR3tSxYUe+8eNVZ/mEdStgWdotAWf9HWkS4gKSbDQ6QKWlqs9c5l3Wo4py79if
kL9NgfYzlNmR53uQboXR+bnIipbeceoPUtPldIPUmkRdyXDa2BfIZKcYdvr3S4ZK
6a63YUhz12atrhIrjIfDAxjIWZRmtKMRzcQoKJrN8mpGleQlQBzlc2tg9KPvvdvV
Siw+hNsnCfR4uZrBHjO+KjAANHwoaMeKhrPaNgdKahyDISSLRrlkc5KSj8SZmD5I
CTmmRV4d2T0QlqoDsTM0UpLqaH0hWby3bLRcXZNNk6bwCPp8HQuzTz4+LgpjeLmK
Aqz7PI1/g/cnMWkG05mYSzkjImBRE770VVMvszXiN7VbUH21T4yYAZfGPvp1R19W
rvlk2HVdACJy+oXL1VufDLdTm63wYyAuo1B7UKmSpA2z9xdetDCVlqP3VuhJD/Xu
QrA2EFi9GhtvEYSVHcPUTn4ejHDeKnggV2R7AiiHqTsqzeDWIPL4MSQoXmH/PFHm
VqkITuzWP7kSDUfoqAsUzJuf94djT1UjXbd+f1QNn0cdefuwgSZeog0V0sMRi9OA
nGl+FYWP4Z+MhRqnCunq7TMb2xaE5tafBiNFTaeE7bNHMGVj40jbg8I4XrPdd46t
6SlZy23W9caJgGt3EkK/9OAUBQAHlK37b5YHS0zOipDNmOlU63r+vLoKBJmsfUSu
kfBFJYpKCF8mu11KixiFGsLYgQEprL1R+99aFol9tttXiXXdegbYK59lkBB7GVAs
bwnEWN10D5rwA08hSyo2inz6rcTsnmi28yMCbydxyqdKabQ4NcpLa5u4NOflQbjS
+bq+DJzCitrK/1gpEET45PYgT1a3Hpzy8v461T00xOkFr8/7Z3cBzBtIlZcElIE1
kO+6zVXqu/x0OBMhmRh3TI3PskEl2bgkPr5XDs/GgyWwBDKzQ4BJF65+zmTntHKc
fJsa2MrbWd8OVCku8UGKnMZhVQl5vswWEFQHnFA9A6InFjaZj1U98HB2y3TGjt3Q
BQq3++dsU2El/c/UDR7OUDyWBy2jteyxsYucZglkfy/ONfO8kpu+oWRIeQy6GXRy
31+TMjPPU1wvR6ZcplUcQTsgSAv7G5h1vMSVAIMT3hK0p2OWPGO/VGYoyyMl0+Lh
2KYPMZk77xg5/EQp8mGbQc+54xpiMmCwBPPp39DKMqpTi3C6lzwE/JnHlITLrcra
/aDpLG74PHZDiqVk0PT7q5EIXgSNBbQ6lxjZbvtyjPXT4AYJgivE8zMFzRjKDx24
E1TIr8XyHGTtw/Z1cqPpe4IbvYGytTE/4BIWfEGthl53Rn4c4KnXm3TR4PRA/29t
8U8AFyQaggcFFUv2gtE/IrUS61QiyoIL6+ICnb1mLNJj3sh4IO9+zWG0EAsVUvuj
AQTfzXCx6OOXNwWpBh9QqdJjvPG7JghYaCqrpodxs1fXRQXMQMq31dvqueNDu5qb
4NUuozKmSiypCSK3hEgecSsSTRPCrFztA5PIc3qA98YXRaOGNuChvtbhcx6xse0S
didYvd2NvcHUKw0DI/VMVw==
`protect END_PROTECTED
