`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QrJ1aYvmz7ctfOTKzMNM5YZj4uWm+P7+GGMPepmpDfubHabXauY7QGckMLauoD3s
6NPol1pHzOcHeGClTqKVsBUByKec+/60cITmiBAH3gaHAAdGxOyu2KnFlxAHllBC
qGJLLglYr75DUpbUxR0cJclQOF1+Ky44sDnCyjZasQJGzXiux0b3qRX/x9TwjyHj
3iWqkBbH+bF4VAeYAuG49NTNpaGqloKLDDQhEtinCICmFaeC8tQ7rcd+SIuEZ/Aa
3XeSWUQAx0O7G+EwX/dmVfZEKNmQzvWLjIHOVB4LcGggHyNKBoI+PAMZPPdbFw+W
GsWQId9A9VW+UnoIx1bda0r+pYU5lDhvkFfW9yq+MsrSUTgJAvMtoIYPb/360toI
4uDbMa0VVpb+zKFeR4gTgO59DTKdPl0Fvm4yOIWT6DzsyrnwuiuJVAz/ghLzCCWS
ZGAYm3GAFFdzAJyQ09yXT0hcbQSrbU4k5TnXR/CACkuxgy/Flwk+mFRdEbSRV8PU
hbtTVfsbm+AwKmajm54PpzIVrFhlaSdruF6GeYxklbJJxIhJdfjptW5TCnoMhrEh
qSQxaVe3CFF2yEzZOPaulTRZKghT6Ijv7DtZsH717+DXENXtoo6NrAQyf0+rpokx
g9ixZPnbrrV+3VFefVd2znTtw8uVW6MTvDfRBELuEwLP1UpRc+O95dJFCLM/bAZT
mlD4ccVgZfBhKw2nsFIA8PTI7Gd7lYNndC51676KugS4TNfP+rQ58MNxwQbBJZcL
smqgynTBMk0kjSuQ9P7qFQ==
`protect END_PROTECTED
