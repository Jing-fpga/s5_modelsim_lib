`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KK3Td1OH0Oozzq3rCeqR12ompbhPEbCY3Enfw9ehcQ5heboWI35A9Nf0vOjwZej4
r/7gsE73WqLj87sKUxa38GBuL6A/hmhaFdr6EGjISSzYyS+jMyWSoGdSA7kaVbpy
ofYda1yQSjJ3wjlbikwnX4eT90bQWgxRPTTf5cPbkxL2E434xytYP6Yq+b0xPLSq
210v7ydq5vpKm3aOtiP6qX03Eb7yhrZhKVz2THLiBkfj6YWIh6Wlj/EANWrlNobT
cVImqdk7N19MyvjlTsasNBj4xRKeLj3bY5UmyYVlIsMCu/qVar+L4JW/+LrkEgTh
WOLfW2pwunI4qGMw2E9yfd/8Nnzr4ocu5wtZuItpQm25l347rnDK2s/em98X0Yi6
AJ7CkPtOLTbHk4UG+3uglEylwZrESNnHS3fVLOVX3Ffjae7g1myzPiY/mJqjB0Td
cljDU3qlHXUzmojrQ/5LtkmIzCuRq0PhRhycl2DLRxQO9o4vaCmshL6a6+XTyloU
ccvXx7XvYil7UuM9+xjrL4ZIidozQCn7LjBct2IC2O1yEZh9mUWf8rsAdJ+X4O+x
WA+XA/DxFo9cO8w9SFj60QzUffGmm4dJciIxnPU7DZS8h/+1YYpvbOC09IJ8xBVr
H4LrBoJIvSRy2Be+9WUAS70IUzT8DK+18rLanLbpAItZi25dlxRsOEEH0XoefQe1
8/yM75ZcfDVCi2mhTdQNNxYsMiM1JDDpBXw2NQvZlAlRMdGuHZh4Gcya7tsp/DJu
pkWEhIQQuOlHJbdxeDXYO2Udhg0Czi15/QRl/F1M3wHy015PW4ItNubmw+7u5XY1
AjE3LlypTk9Ql0Q1KvAIrmi0jlvdcATlpcXWv+tdVUKlc24zZickmANL3B/05S5L
UD8ubeS4jmx9LGuay1a41slcbsg2rck6LSSz4r0Xhbmc0tMs+mHf0whmVmBJh1S8
f903v4yx52F5GQTlJqJ2GjcBeO8u+V6NN281DZU0AuuLg2eZIXdnLmXimXwNlSlv
qJ0KzBWo41ywBlDpNaJShPk0M/YDRady9SRAoMg66PSrS4C38+LCyzmJllJw31Uh
`protect END_PROTECTED
