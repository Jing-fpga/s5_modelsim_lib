`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lDDsr0u+dZcarJ+Fnbc4lC7Hw4GaPQqak4SwA96DUZ49ABrBWDxa/sQWoZmvw6K+
x8/SbDlHlBgwsMo+axSLh/HmL28yTKlnJINYJJKqUCG/4d/hMld2pgrSbBLIzyiy
fqKOKXM/URQV8peIyALxiSfar5WMvsb1yYHEcNAKz6kBAXaMgPIygds1pV/F8yuY
Pcaq0QWjFRl13Jm2YUyn4ui2p5G6ZFzfHBANhAWKiR9Mffr/Uz8oN6bZ3SCu0cj5
dEJBAawwNq4Ondtwm3T2dEgyHwleWGARwLQ4/eNLMcBxu2PhTmqyBb91I1lCLhGc
19iXy6h3tEqlM9vwYez86Jh/irJYVGyb0K2Vb9U9aDcNUPpYMzwKxoDpjhK3tbCZ
y/Eh1ZtuVFkhq8Wtqc4D58a3BrPvJISpbZhRnExEaW2biVWxwyS61DIvf2sC8fRX
9o/x83jsKJpsB4xSwkcyAQmj+VucO70Q8GEt1Kyh4s3CaILIsofwNQJf6iYiCLQt
yRKnWLK1F/55w8sCgQnlAiP7gdTf/taKLh9JruAMjk2e97htzat8sP9/QjLnlgEH
modyljUUCweMM22qrvd1owxJnKowsmjAlIErb0Rpo2MGjT6Q4tgb0r7LycjFVxhy
mx8YR9fPIBEOVfdMZNa9UfNerUETX5VCEfqvmKZkUsF3QxmvA3TdE1dDSd9yOd3N
+CIKh31HxS2E72wZnvnzjMBmkbyTfaP0Mkf9wlRRiDGasKMmjbk023vYfBdhOWlX
ueU72JPEKI5v/BzeSUedRRllpUlquBedWnUInuHJeDbMgXPYTO7C/GDjy6Ailqvz
DN4AwPz3SODwHsfPKBORYTVesdPG0mwJYM+yJAedtm+vKcvOAqe1PmVAwV1Z+SPg
GtbFnKJ8M1xjCK7k0afyUkrl9gIyRlO8a7/MTT41N1AARjT/HgT5rR9sRLc81ccV
Z01XhaC5FDW/bKck11J2roZR4tX1zJyMHYDoiMw0LT7UnZemrQEmMkDWZsn1JNsl
EeqykNYkkTD15dqZ6nkUeobJbca3fGoTYJPQ66kvWyI2T6b/mo2WdtgNnaubsei7
gQm1B9v7k1R2WcjGAQU/3ZW5FN7e0TnuhUVEtZYIzQ6uJZTigjc1SYsviolGmFG2
crYbzKABoaT3Qubybs4TLhBZm6Ur1kPX/bW+yZF+VML45BVBRCv2YVFQPj8SaZCI
O2AiSrZjTvKmgUnC2jV2knj7+ufHBOYOTnfOzOsIpiRrEXYp0+YdWLNWkmck0qPN
LJPB+oeLQrOQ0xQ41AeZqI7LcF4zj/0Byvq1cI9T/ajMZj1w5dAxX6Hz1lBv5ald
AcdKuCtS0KEjM057YWD2i4MqM34yR+w4UFjp9lZIPGFhBVxZO2PIBHK/gwgDU6ok
VNA8VN+Ny6IEe7jS8E6FitRNj2wfPeJgEWq1JoNWwpRYIfhrG8aKDfWE9n3RuRqP
rJoDkEWjr75E9btnzH2X8DC6CRVhQT5+B/8psl/a1tX0Qih4e1c+31azfg0f55Qp
MG3baavleE9vRybAyDGgCCAAVg9+oWggpneuAP7iJ/Y=
`protect END_PROTECTED
