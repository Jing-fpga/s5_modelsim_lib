`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vHSviGe598CKrfvFsgCXb83LhppbTn6d1/QH6vODlGF8lWcfG0DzlzO9/B9WMwr5
7D8ZCzED18BiX80TQ8ctogwi6axkYTRNInDhlrdbJMJ/X7y6rWc5g1/VtD4XyQRb
Ps4VSLet0BBxUiV6YFLKwVxskoZs0kDmzMLe4qkjRTG+zKFNzOs71IF7HTfB5PLl
BeiFC490tDlFoRmTVmNuX835NppeYKZHMr6yly7l8Wdq8A6lgnr7kRNcqP1zBdm1
MgEdVvyzz6r8s/CLToPtUW7d88fErxUooyC2NIGAHQ8sr6ElIpSXKMaetVfjUQed
C4LqB//sDicF4qZhVBa8xV5h07uQ0P3FmTlTafa6w3NvASS+idG033wT4S+CepVe
BQF9VAmFx/LZ+SEQJlXuu4Ww31pJDoSXwJEyI2IZzYQon3+8Sd3gDZlakYM9HkgW
`protect END_PROTECTED
