`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tC4LDyYgAVuDA41gd1otR95CE+UmrI/87XrOAYcYirNWEOgSKOP9ffWdLI3UQPRj
hUHUoW3UNdPMKYqIMFCG5BzEggaHlCMktpKNKVKgw2raxGRzJawryRmtM7PTdW+G
i3HDSrzzLxrfPcbvI4wCz/3nSK3C3+EGem2hdyf2tDW7uslDssJ593lzGVd7dy/f
UDgPqTqF3GvARaVFov4c4uWsvXrF84gQElVdb0z+DDBOsAXSyy66Y/dsBRtjtXX+
Nsvpzqjbgk1DpzK7Xu4QzAk9ZD2JuuLW7gK8NK5HPFZEz7xwxn9W6DJaico4eu8d
XD0sbQWGyhFLTQBwZXYGUgGjX6sMxZaimqwq4XqjVHE8zWnpQt5GdU9zN2y+h2dr
j92qlg3HQoWjxP74CkO/7UbCe3fpa8Qy1Jbym2skgPHhKOXrb0odxvZchAYr7fR8
UsW55xxdJHlkBO38yutihYo+8U8HkWdzJ1TP4qUnKmxY1k9EJEcStgYTynp39/TA
86XXIsSFKtw6fym6W9eYwsj8TnKYus++PDieqrNI+Dlz443LuLW7UktWW74/dxGP
qC+MhUUhQNT+7TJLwCp6esTBGWN16+s2VdQ0w4/piO25UyXRyWgVnGPwTzSxUK8m
knnQhbLXvybQhQN8fvzGQ4+fidDB0JmQ1uhljwVxxotn/6ykXeVcGazGKYNG7EAM
GYQrUeAc2VB0JrRFpSLBuzMhHuMVMZ2moND9gta6dtk5Vuv0QOb1GXqDS5KbHy24
J/E7VaK0S95eHAxtEOmLNSErsmcIWm81P5huOAPiPp9o2sqxkjTo0A/+Qaqyq4XO
01EsrCysPV8TqFSiOGvTJ3XyU9CADTyFkldXC1Ok10bzqgAn0A+B/CDW9MxfJLqW
buzPCGQAvZs4prAkm24Zwh4RKzWieLSXhiGoMBpjjwh7gFv5GPFv4nz5ElEQxoID
JerUYJIBXK0X0Ci97eILdFva8BYwsyiCEa/9xePQvQKipXQuyMfnEEIwheav+9Gt
jGXtsD7wu3Qzs1ZNAqhAouzyuYyAzeovDBAsXd1xwDCyrOMke8fBBII0GrU3nE2b
Ys9DkN57tg8jkZitLVVWVKoxsoiwxAA+egAuIt1HutvF2qKGeIARbzjl0CvfU9C6
mAvvJc9Y6yC6/EiHJemnobpiOWGcxHZt4iQ80h/BNb9boSkxwVnsUHWWRCXdESsw
ujz+DCNaZIIW3HCme3i1lIbHPEoto501Eg5QJHERXa/9FrHH1QUfBYPnL8zIPw+x
VF2QNCwRthtTshjsYdeR8YkQTvnFKMaBTToSH1/4Qj9I8d2GcvgOElgWSCKZn5n9
XavkMdcDigF7aalEpKzea9eRlG+cbaCFFO1+wKJtrBYkY0hmUQmy/daPI07per05
UDkf0UV3p/LaCDY3TB5hDR7g2dv4BrudNp66wH+nBCfi/O3kklldefnzQqPfRsHF
rS1UpXjeAMrDZcg5zEhthRZp8kuOrx53WzyZvyoNEAp5wjDYuBIAiuh6m8VuBcCr
ce1695M/lYPGAVx9+Tn1A6CrU02jKXrOZwMF5up4hAf/CnQ6DW012RLOV7JT7pjI
NvpAl+XRFjI9b4qRIVUsRfPJUENRIqNcbeCnWgcIFjBvvMbe4S2QKh9f1/k4ZgUV
jcCm6PT03biwguVHfcUnvhsfPm6DrIiRMIeu+ztRLfdvDTVSkO9ZzahPcthZMlud
3pFR0w6RgiOqf3KksRDqVW8VhVLWIfUU8FuuS6qXlzMAiz9Ucon+Yq8vvMf/TR13
aLEpVpXIiDjt5ovVJQx9P1CFXo+YbaJHe71+nmxNCC34nPW6WGPgAppJRA+gdDpK
IcE0ZJtIFxSYj1QqTvBRrcIRylIIOAXGwMZUIy6rSo021F/gCYoI1rJDlnS9/OBE
rGsLBI9OtNd49hn0ppWWh+uLYUAKUvDtL5rQCpP7fElMnv+UZ4kmttO7wGeZ9XMs
1kKVEvxehRMM5VC9oiwUgNVXyaMTJosWOggIXYgE/CltS/FEVNP9SFSUDx3m4U2u
Blm0ame91epO5vS4p2QG+xa1HZS1wa0thI+NwRiwfp76vfgdqoIxtdUkPavSnSEY
dg8DLElv7pYlDemenQ9f2IT9Xnjoy2O+p8Rje3Gp6did1wmRxBgJdMF0wzz9w0zO
xK74W50uUEo4GJqQ2E5+RQsseSgQjvLIcsEEsd2r8VCNDwULgUYWplyyS7mdEBas
lyCSbUgykK7aCrbgXGPBUh/2fc3Y2T4YeFV7pQpP4V/CvZ4i9xzrW5pSg3n4qDUr
TN1CsGEI9cN76CIR6LCBR6U0YQgd0wBWq3HSxK7fYDqWrbXzMvYd1pdwJ63I4fok
eoqHE4oLmKX90ifaHBXq3JL1GyF6U9kUg0XxLpKZ8s2qZcf0OF6EzljIcGRZX87w
LgnBRaey27Fr9FlnkZ13JB0F8C8cIrV51G7VCsYvlRh11cV7vShIYXjZ4RWay4s2
/v+QE2JcRkzzaH8xiyENnXsIQps86YZovTj2N5BBTy/J8PlbAyQyEfZ0prsZMYeD
FPrtJpDhxeLhlAFfGBc62CRs53wGFYWUKb/9I16ZVAQciRcFnW/PVEuBD2zsiwQ2
86rxd8HJz2HnV1wQ4TRWXZHpTSwzJ25QGtghcJ05RID6DU4R6YcFQJacPUkKtC2L
K6OVZa9xiwXAvuXcuFIuTcxuR3ZKMsxcn7YStK0+yq40RbAnoccauAbkpulmhRJ0
AyPfz2KQnPAWkMn/BewY9U//XGS6/UM1ktX5wUwlKlcEO9CDQnGDsaHw4vv14xCs
77lq60DbirONW8faTd4SoETx4XF44d6bkYaKkjW+WitSdetDI/2Yl7DrIXcN80Q3
AoUz+d/WoN+KboNxqHhSKz2xPZx76rwtrVHxk2Kh3a5shG0PsBHQqt5bxfGtA3v8
L3hMaS9/pI0ADx2jw5R2zXux7FWDXGhzG6F1doF40fbwghwA0QVDHo5LibWyVVtS
TwE5KTWGkgi6CF/QHmvCAk53X7bGj4eTtGwCKXoTsUYCKLCQc3Kzl9p4z4S4CP83
Btwaw23GB0C9Nm0RoPZriSPGZH4PDOyii4f6TMLb0dY9j3++Hv9kMloiOvnMY2PA
V5U6Il64+wGvHyzS7Y7tpIyMCING9sa3HOv7ws6rqQgg9mbbSJ/vhfSsBbqA34gE
aMpwAiYLj+NUG0zRj+dTgWcYpqEBWrqNhcn9gSrV4q3skxGhXp4mNLUrzOuuSl3K
XCJWRo5TR3dPqL6KF/MwsOp+M8b2WMn4/mcmp6RRmW9/FxSkMEThmkrRvC2q12Xy
IsPKCAMM/bp9YTCC5OWEsIzS8RZ86ZGrOgXK12rmNBJLbUqdStXAb/SgVRN2HctP
x2yZN0hRiQrThfn+ZW2knwrSZbR3FKBaRPjn5F1IJO6xaHeJrswzlW4ujldeq9g7
2mVxPYUJfI7ow54Xp3bMCRWDS7frZELJI4hlP365O1SIdnTJ8mY+iOF3BHW4xeaV
otIuWo5hzicMapNcjYM8+l+eL1K/NkBmjhGdCSYb3r7euYf0lLSHkPZl3ka6Nr0U
x28cfbzgMp0UI0pEYV/dsxrXnPRuadbK2RiLc9PHW5V02zU/w+Y/l8YBRcItrh7Q
pE9NtGqc2hcVU/YeHjQpc4tw6bTH0WpnDPx9yoyWDvSk6/ISSZHmu7zhuONhtSpY
UOiwkXQ5mbyYJU4lPTS3eSBcaGO++2Mt4GXdUCmT4xv7JAbrw9YYh77NG5QmtmOi
HXaFY+Xi32XDR+Ym6AztIS6GUzIZCNX5vNbSSHBQhKQzLNIWBPSYHhfrIkWZWuYE
HRdsBfW/jZtPWXgg2jZkr+jnrAz2UUjns0Ia6H9LR0f75Enx/v7nXqlCVxShHWoL
kFZoXYLRwZqEkAyhsEEnqFtFUbJLo3zyQCXRhe/OsgFrncnvCyOWQM5P7MWpIeud
P3zloCUF8M6hdP2QadXgFSAPdqyLhMvYJcUxyiesBFJDmWZ9/9gTjeuTOKskpSBD
pyyEhBBFfagyth6I6cH5Mc8MVw+3VIPlZFQpwAxYYxOLtc6Wi8tglsVtb6ErKw00
dtrfV/cR6XhQDXHMwyb1RkWZunClhV82nFI6Y2FxdLbQQEbJG21g0ljsc+2FVCez
w2ZTS530jIHKS101fcJaYV6Tk0OeShqxFEH84YjhSoQeqFipRB65y+OMptMrekad
z8JXL+XOI3UY+Dx/NRBWBAW8T1VA79LRzFKOw1ph4s0s8u2GB3i/M1LFKFZ4SkWO
hqFTIsX1/F0MOP5qJjsnVS/oWVf6mQ3i5ZaabYqSdJ990lPIGMbHQcrIx9AQg2Jq
qZufKWbRfVSeuyIzRfli2BelRS3NNutT4Pux1iC5/KkQEJENs96YvpmXlEd7IngA
JeDBGEluW2WkdX8sLD8cbmf7Ovd9kUJtJ0+g/M8jJFp0TjKKIumPV5w1Nhpkl52i
pAZIYH/MxE5X9uYLG9hf2pL5PUauYvOVYqk8pQy1R8O1qiCRz5/WJlNIBk1PaEWi
gMLZFbme/RE8ZJt7xJMeoVUQCbXpxJGoDQriFB1RV1hOfUzmSx8Swb9h7JF3q/jj
4Q/SOEIui9oS4I1R1kd0l5jc01yc7xsNSnX9hQdUZgJjOPM1ohbpJP6JhmQnXveq
BJbJZB774QpbjIhMQ42TrVND0bY7BAwLlx9T/NVsvwSfQkMdr43ThtrqqRY0oTIc
UJCdAWWQMxrdiJ1Est5rFCpmMh0zy7v3/Row3GQN/GhPTLnyRArsE+LBRgUjpsnD
g7fOQIpgX53GbdHZOjX6/ljlVFdZ8KLAjKcYDWZ6v9LAAGzHHSCnWezov3HX9wPn
eacSlEuQK55Qi9PkBiAF9ousua/OuMbMkSrU9qWE+mazTDzELPVj+XIsYjQ5L28q
rJ9XfdtL4W9vSfCkrz2sYDef19ynuUKz8Uay26E6q2JNAA6tBGbgJ+NVIgcF2Dzy
Th/1p1uCN3eqjYa4is3WED4aCSQuRC11KLkR+HznA4pKFo+AFWDFdR2G4JS9vdEM
69omNrH4IWG5T1/IpOYpTnailrm2VimbepgejwnqMHqNsUfTXgPv23Y9rc9u8yju
36C8DlQtwezFVB74lnBhNthZqS8OCad7oFvfhpAkE5kHDXoW5ruF1bpy+w0qz8kZ
kgpUnOM42nYSMMcmj6aFrdY/swnuRSvvvLToQVzNEA6EG71q4YbqiCBhsnwa6FG3
MsgtSShX0vtj6bffsSUuEzaDlvSJ0B2nbapbuh2Ij3Q4cSIjRUCgmlAcYTXybkYA
lIPnPTx4IOXdkhKSMzY8JoFdBCWAzcq5DJo1WQ9pnXEHZuWm49pICGllBqqBpPn+
mN2P2LN5qiIZe2YM/7Y8AyUykp/sYdCNZ5yFb9DL0YDwy+mIG4jiJEMogIk1sFAH
OSV7gqhlURlANs1SQwFSY3t2gRiE2yBT1sGcyTw25/ySr2/7yX+Oip0GQYPbiRKU
5+cpA1d8BgLPOzq/75lvA5FQIu6t9wTUZslZTEAXRaF77nthX8L/1CZ+U/dLMch5
pLtT1vR5byP1fj9FoP6bsJXkz/REPEitXODPTFNg8whejyq4vGv8kLV0OMtNbjc+
0BgTvphC5TfoKyju0m6EIOFuByNQv3jD5paDtBZDKUphvXBpsqlOL/KQW7POyNXk
X71zqF0vQl5R2ff5aLvjnTduSMW3ElpPXuzg6C6kA23eBoTlMYevPtZAZ3ysLwAA
6vBSxp2zyvOaVCERm7HG/YpLL1myby8QLZu9Ql8FBkdOWYpMvEvLZhoe1A9pEGKe
LpsMeJs65i1kHtbrAr7Ve1Z1W2Nj9ayO5bRjE6voNVgF7uTjfaq92ANQyvD+hcxy
drIHIUOj8JnO8z6sYcy+/2rywRY5osqtxcFGKO9xw8esxDCIU0rDpztA3ojHNqOs
heHzF/AlwEXwD6zmKduSaNXhmrejs1SmpY32sK/6JpAt7M7w7aUsWCfmUVEQbhit
5IP2HLsUlmndJR2YU5L35VCfrq7DWEhZMgTcIbWcvtslbnfRCTkV/+s7yi2w0O6v
ulrWxy8UgkPco3QF4pCxlksQS5/N0QVU59TlPCDT8WxcgcbgO3RqanNUtOnuujIG
3tqYLnwawISu774jl3Qjk4U4cG7N4gPJwJ9WwDq3psSI5pHfzjQLHKhyw8it2tLK
n6iWGXELCLi83llx6H6DFF9XBeOFNvMdQdJhrC5OgaRL5P/uxOyyp/0oDu/Wivqp
QAoUfIFDaXxB3bT2TzJYkT48UWaETRo8fK6FwPAKU9qHAFjZscNGXAUqhm/95iJP
gPIA80e1YD0YWedQ9KQ4CBgLufMt7IOx4pXL5YJW5FuM/IczaNL9DGX5wIzakwXi
buBC5CgGpsVSNVxWmUavoVe9HXVEzSOUPMOJ01amn5CfvbFtcOVLK5565B1MpnqE
F23qN2xifRy2SGLLh20g/eEqMccehljEtewADU/ms++OA13lXqhsq3p+AFtU0JuY
xUKCNmT62XzVj084pynVKwd7EkHYdXZxn+q4w0RknyCtDwI04w9THwDQ2/bzeAW+
h9sRnFBpCeOs90R2ZRg/sknvQb52R/41K0Bzux4ZYuKNdJR7dHeI1k+k5VE/jHvQ
kmDOmZZKrWGEDaqj5GNguyIszJItNLCpil91BGdqSy8ne89RahJbpWr7URExUe/r
mDH5JyxWte/dBIJYgXqTsJM3j40OH5TRK9V9qgK5taq+O4WS9UOAA4Nj1UFbN5iU
9623AICtbcei7F2GDYLoRh3Myab6nIYR1Fe15LFosE1NZjEI0Gvkoz6M0Dq5ZOtv
Cs0hq20OEuDaHchGNkPk3VgICtWAEjJD9kdJgNES3gLI1DxIiabFKriyd5vpp3xS
AJPVAusiW29uQpha4KQvMs4XK/w8anmVXkOQojJ4a8Q6EJWK8WWi5TbzlBKvBNgw
CY2Vug58bcc0hmMZcF5ubyrqJMN1rLFi+BILy2Ndnco7gOt7jlwESvdOOVf1qnmK
KKeaA6YW54wSl+7yS93EGGi9T4QqNirDjXZ8cs7dmEZNuzycD4VgI4G75c2HxSHX
VL3K5/fxbFMx16VdX4eKVXmGqWCZSoQiD0Mp9ZiLyJPQ0R9jc0VnEtmJ8XOLhvKJ
Cl+Ea23OsKtJu9THl+NkLvHRov96o8+CklLhE6hH372TzYeHoPiV49RwmP4vToUS
Ti6T5Tw1avi6fkzRa+PC0qm+NmdZcBXVKqE5kwxOou5LEW1IfQ5e8QDAO7471IX6
siHojZz5f4KBOuoNdyKkJE9m1zGntuXF0pUETVCYTWKDc/9y7WzqDac7qfTEG6Sk
9D4/RXPaoVUTRHkA6tfOcAsSmCBFuIdeK17uiRChiJPMUNLHVn9Dw3LUimbdB6lF
jIT/pgyKUxW2WTZiopFKntrhkgOi8JsSU7rdsK9QyEcMd8cZHlT8yu9b3A4Q1SkW
R8dAGnoL/kuGeqhLzbVe+5wazwhMZv7KRnyGo5UInEY/S0j0wsz9JtuxTM1H5V0a
jjfsTjGw59R2SQu4NUZAUh7KaQNtbp9XJusZWttrGKcND3xRI4PHZpff1KSGfdpQ
+jvazv5BpuvX2eFWsNmJ8OnoPpv/aC/BDbGK9qojmyN4bXuCMpg78043Cjo8jdQE
J4QgtCSprCqZrh3UiZRclBg8ubeXSZdBv642YjlhK8aAbGS3fzJY6yvNP00BeRYG
YmAELwYEPpuTOVt4LeV2G9gKYzWgfqUwvJR3d4Lz6tb/ewySqXeWurP1lb0k4p8w
lIBkAiJosvrcvtoqZKkQbHU/E6k6qWoxqLtOOaaV2buzkTnDMrBi2BgJPjCqs+cD
A+l8TavkB6PIiomHUYohbUnPgq4TLCnEqUd5ANEgwtqarNQRvRS5QPmRNWFmxXSP
9mWYk6vjYW6a0XaPBNFCeyU+ZBKlAYVyP6oiGWplUZQKrfnDO/Gzih7DhTDAZ97N
pBQHmLAy5JGI38Py0hQeV3DUvUrQ+zcVjaWATUYk4jZKMthWc7/D4OBhte3F5bvu
EdWwXv368eQM/V6rxEWFyCwn8LHnhP4QQqX99U14y3QfWZNkyXtl1x2/7YQ1sDjd
chz0KQYD0CEwDuVBx/E2eTYNl8RnlBGrJDKSSIE4pAZvpTY7iMOBMYv5IHYAsxE/
7d4n4zdO49+KPZ1jieGvdwPpd8RwW0pwTmDOwon/L9YoCabIpdsfrO0vnotMITIU
3z1u4e/4nZRE+KHDurXl2ukr47mXRSn/OsZ7/0RrdaV6o0CAShGbcQ8WBZam40DL
YstzTJcHkpOXh228CXea13hwnfwZ+t+OwrbZCNl0p1EGNT3qmvtSgl0mPCJj6rDV
h0HFCrUXCQGT/WFHA/wrTvc2CAZ5CHD1yGR8FA080XCyt88DJkTR7ZgM/PrHc2oP
bRq+0abshy1BwwOFvTtZ3FNf/1yZnkgbAuj8gtHrH+/eI5sl5kjFUQnmH2VNhjH4
7XF7e5cn+u2z7VM7Gcm6dLvRPiurp33ex9a7oU9rEWccnzeGuTWhBUATp+wM4Ky4
ZC5dS7flHY33q5KgCQgjZInMkAyt4509KYN7gjjD20iNL+PNyZFPkh2be117yzpC
cH0vvlBnXlUrWZxcXI2X4fQ4nJ/8nC/6YKu8kwq2zoUOw3bARBwWYPq/v9PgdLuG
tnP6tehf+mFylw7aA6YAlYegUk+4DUTw2v3ErhDnsdwSdB+h2LYBq7rNJno653za
PnvAXPk1uYeGTX1qMGUStJRMgzBGBblNehgwDl0hf2Pjl50X5XS5SivY3xdUBlsV
sYNwtlmwLFGEmJeRWf4Fk54Z5xDhjp/LEyS8zEIEv1+LYQ7LkdOO3DGPGWWyXa1a
6CoRR+CK0qgYSMiV56mZozO1gk4+ysRvjyE3UpL2wzwJ7jEetTl8HOTChUpp0QP8
vOE3zUINOKy42b0TDi3j8zjJo00hZr0KfXaOBlS/18xkgpqZlywpR3kFDunp3MPd
7yJgQV89e3QzukZO+3W2F2XT7nGGHVupQVtS56D/Ebi9XNrpHj4cJMLEf9Jzo9Tf
s6LWg3Zr37Q6vRJ0+ShKkIyp2eKUgKvCaKc8cvrBvZ35lCk8I9IQxZDlkNyq0RWv
7XzsvFrun5P1I9KLFHvkAphXoYL5UpJetTbbIqYdNU1+OQGYOpgiagrmpnuVT8sX
VCpqUUBczOItWJUsI7ZaAbzGRaYXGqx3YCG0P95RhNeA/zXU6tQ6tYrCvDUFrBjb
3ffpLgDERPGELVnZ4OEE7oYdsnV9dZ/DbNATzoo9d2X/PRjc7MW4UKA+IxOaeNDz
A/L8a+KUkM7WlDdga2Fx8tvVi1su1yY7IPjOjuB0DbF8fuMiLIzpfdilG/sCrE/E
uE4IEFtY6OSMIgqhHjqHXheVCgAv2a6QlvhoBJ7M8i0pVzh5FI7yTW+S8XhL7IME
zOBZH3tq2u8kXnHSMZOYqsMQB2OZGNIFFlfkFgkKa2qWo3ZzBn/FXNJ9pXJi700e
7yuTl9wdti27+SoinYaQ9mlcTnA1a8dA8iYk82P93rXEYD1y5/3NkJPOo/1kXxwQ
INJYOhjc4T6AK4FpwRo3rTYpG++GiFxuOmAcFeFQcFmY0g6HsI0QyKYhPCaWgSCR
VggbcD9C79GxgeClw565MPONl+JU1lod7QwVmG5shZpJqyTi0CO18yyhZMO20n1J
op1ptASw1ga0ohMbpOVEvYWGOFCUhkCQmDjDdrUDkZ0w/IvJ1E0DcZ5BekciRAaj
56s0X+38RJjN0VROX42GXJDATaeFR05tlT6EG/tKyTjzIJ9HyDKLkIZC6/QJsfxf
qyYIYTFmzKctVNyVwMrXgtDjDInno0662p4rMGKIYB77cAIA8IwIuqNGJ+XaPU2w
lJO3vZQILK1zuzH9rgTnt2SCKGTuXNgdqc+Jj49mMd1u36hz+od4lpEJ9USoOKK0
0hJGF/beBXgzy62CCF85Pc+egeRm8u9AG6lIPCT7/Lmi9JT5szNZOvE2HbFUy0ud
Y4JJzTi6eDGLtBrqSX2nMafBYtHt5z8KAzSCur4aJp9Zm/uOHVJ+a+av9+FlM3yo
qnrSzMkVn7HVPFZHSjsoliJoyQWyPQcVqk618dexWWftz50yWKbobpAlTMEMr58R
vROwZD8Mlpskj+v+tS2ANzP5Y0DZWMed1GYGQ6T20FReSGv9stq3dL+XBU2sIk5L
jgEXd61tIvGeD+hTwLgb2l/mBwGaCJvVJBLzXikP19oPtlBLBG8InuOFzU9nE3Uz
ByekrM29FKDuS6jOhsMToU0PvHAILSGs3rEOj+TQZgPnlLLEvvYND1GQaXATVcNJ
NeA4jPeYUPM9Awg7zy2MitQ58vQXGHpgZStiE6PuFHUBMNkdNXMb0PP2EG1Z8pTW
i5bG6QWRwTUCzfEm0BMyyVkDjc/Uj65Kw9f4JqdeQAk9upKhJfYyW99sUQorggmp
zfsFen6s7nywQWqA1JlILTo1DDEUknibRw6UlMBBvwwG5prVz5YLqKySlsOYUEU+
ppQXZAQKfORPwbnMl11lk2FqYEyi8edRKRoWXn90SsM7xCv/gkBQxqp/Ehk4/bk0
aTwyVcO3VnMh0hVhubxERPSCPi9PjxNufif+NQUhAxvDLg8YiVn3tDTFDM0Nz/xQ
IWDb424vxOYEVE8vZfXYRtcVZF5qmg4g0cGsxfJn028dClbKubetittFrmJ/tJGg
y8AC2i8gYup24YV5HHUxP9A/aX4/+3kN0aTsLoh9pYbjEYWCh8U8AQKefW/SHuXY
EazAhEf58p7Iz6GQT1PY9fGUn3Oy7S6KNlU4wb5MevrctFOaPvIAy4WmmGR/N5L+
P6l328p+OqJiRIPfXcPuyF8PgleCHJ4xJuEFaV2Toz3tr975DJuUAwUiyawk5Dbg
TouK+ZHmP2DcuzHCmV3AhJiQCc5B8ciwZpWmhu6a2LMFRpFYSRjYZxxYfOzcF58w
3v3RPZPbT55q33KKGTsVHdvmnQ2l/QXxC2msfMtVvaBz8aRpH0aGbQWBfNHH7u18
KLg1CWeZnP9217xGSfm4PfOoKDmkBY8bmdY9Kn4+WPTW7x90SYIixnNPfoqpVDbF
8bp5PgbKiNR0Ex3c01CieOa2NPJBkFrD0s26BoGE5bX3ZMBMw1mLSoRW38seRiBC
5n6zYKqm/rSupEk8vfJkk7V9v8bTJOXsbA7kJh+fymx6NksEKGqy8QPr9bQNBGlD
ghVwEJxPQYHNeaGxxZoWcR7/4kzLv6IGjkPTnXElKZYcqfa3JHzHhSs20zLT6NvX
pyKq2HysWRKFKvde7BPTv+y8/Cy4l2PmAyAmE25z9k2hJkv4KMTayaCZ4efK+QWl
JJZPIT83E5mXlTEm4z6CyjhVoaR5FweeciGOK9Y6hqSBlycKn1ir2jCpLfszp1QG
9KR34eVqMzb3SFotxtu5pXmBwZuX+JmgxMo6bNAndwqQWdNteXMgruB8Sf8A1py2
QJh/chfZknOX5oE8uWzCM3E0YnRq0M04nqTP7g2HVa3W87n9Zb8kqrZTkCDYQ2Kd
cylWc8TAs91oxAGDHcOIDqWOus9+vVsG1EE49br/G9sPvlzjcJugAMhFZ6jWz9oK
4gNSYOWGtbsyh3tO/tJbXUvCIviRiUqnxWePtXDlqHLMupDWKbJAGpvBHvjM+kFf
WdRUKtcKycI2w6lS+tFysilgNqMTSz3UdmKSNaOOaeG6yC02QGtkKE0+elOzmddK
Z9gsAASk21dw778Gi8u2HAzS2bXzaM4v5pKzeVoqVmpg0NzcQZujlMPLX6f39glS
AIUBYRw5a0s25/dS6IpDA0ouDf845usPl+qKN+XVQFeNL+R53RkquUnvN37qmTd8
23j4ydlRqeioDvHRWhBvk51c+A1+qwspmJukmJMJbOEkVPk4V8+L5KO/hadZ6Arb
6oXLbUA591yqk64I9gnl3u55xNKiE6R1OfRRJ2ueYRnJbOvI+ju7C6TaIHYaDrvs
ZQp48VNB0jyjr5nzVQa1fTQd9GiviJIgkZxGQ26hD9uAXEKbzgprjvOb7wv3EGmJ
/+OONFEfpIgJDjeUIeV2+K1lTWdzYI1I/veJ9wly7TXc0amG70CjuNaOTuGx1PFL
NKGZ8lXPnk1BPdc9MbO6D/4Tgk8zxXGRgngwizruLftnh/MUubU3U+oaQDWa+plz
UGTcI7jASxFUFVWnNuEIIlQd4At84scXKrGJ45X6IjuRXb/wuUzdeirHQOv3bN9n
QYeqSh3FAHloZPAG+jvlzeKRYyqa2G11l7pdigOzflU4VfmYJWk/JzmgqTO6eNye
OXib+jo6J/9VCRlM7p8gfIJQOr0eBhwR9pNeq4MQVO/48VZRHVVj+56xPHMsqof2
g1Y+usCGkfuRtp0qOxtn3j0dsFn/79FXJceP5gSrGMqIdoApV79yCutpdwNh8Gnr
SU5bPmYERicgyRRASnEWNXN8/eLvbsqqRKaFT6st1eAloEXx44sFrNLeSiXalRZp
hieqGJjwS3W4UMoyXhXETwJftipIwJjhFRLtmF/Lm8hQYi2C227R9jf41bgFsig9
/p+skWZLY73FWJESCE7MKgDFXXBheVALqsX/UXQRzAV69YNje624kZFPRqOTNWgx
tNcRO3xZJYknN/Hb6J9+o23HwU9pvueTKaceQzMsq7gjE05jlucRIvao1DjnmAn/
wFceRwZxk9bOUfvwsjeklgP4jXzGNwuLDNVL8dlGqhFSDkJRg4Ih7CthshEGICZO
SpUxKyCU3vjvxqHzGxkZc1VIMiasq1G3LxNJEWWHT6lIhtDJKS/ZP2u5eGHYnIXG
KK9qqQtNvlNrU1WMrdPbQIOeKUATp92dpSD/nB9qYKabUapfZnVPCxyjOOvocvJL
xHHT4KMugDurOqfsHIZdjP7HWjED4QaLp1cMMMroThPdOETl+01od5ruYsqEY72J
Ww9sXK//jWjWF6cmSTtlRFXTxvxrCGGRYjhbgUZlERR7WHvdmXhnw5Qs8e5kvqrf
YnIAUxkAXI3fgYfklpZfpm8T2xh+UeayoWmmvIR1w+YwNIUbX+eUSA69PhgnyARV
mVAe9wxZ5pPYMVrGtkr8M4hLVL9a3ar/gisYIs0cYW27r3Fl/+DjxKy/2bZ6FLob
xNirJtNA4ETnaOOHvteymDeYsZhleIbxNBYo8gzUHOXaTvoo+Kr9R2NulpPMbWaN
jITNGTwoHmI7K8GNyD0c6MFI0v/MjUqWZmO/waNQZJKxIXj/q5OBVX+C7TkKA0ZL
RtolmerrcONPv845bWObf1h5EUPxK1l+FsguSGU7IJecTtgQZYs0emzKQPJBjuVm
Hkw5j4oOIgepKUPyrj4KXisKs5j90BVEwsUvLENrpXzyN/MmHrMvwJAjXUDlHxt1
OhXA6JIJVuPN/PQyVJVAgS5g6Dm7FRx424LVQc0AsuJpwBHUHlYNWor2JCQfjHsj
EVP5/CZ+UdhFFgJVRllOaG7k5Zqh6lOLoWJCDCR3gKH/R/LFr9HwWD37t/BkMtTk
DyzgZ/+gpSy0dzNP46rawkN4H7bPuOzxwP2cUz+ojqRVoBW33izrctpZczS+vaoM
p6RiRA57St0U9cQc+TvamuR/90tpOAUBxwo2scIxmQgSVz3Y/5n1XE0tXJ5FicN8
S1UrOlLn46nWxEwSGx2pFLg2W3FV5/eExAgoGBvm4TOaR3H8sDtcrd4BlbrpTp8p
b+V5ThDNJ6stm3Bg780B4NMvbHaI9o/9G5mgpfmVr1C6vxhDUzIayg2ftw+vA5l/
M3XYZOD2JMJnxsBNyvlkg24zuHkCpBaAVzrk/ATkxRTaZa2Fw0cHn/a3lag7aec8
btyt7EcOV8QtLstit7v6MvmZkqxiPX9LGX+8BfgFCHs3fAcLLv0vC3Iq0IPQcTa0
6aV+GN1+V6gBpXyNxbs/2g1C+7dAfGroT6asI05itXeqTSufZfuEWFiVNMAVnqiM
rpaK5/HOrRZUUmUC/R9eQ/xY+4vkvDcho8fGm99cLyGOC2WHze11TVscuq8V8Zxk
tNp/vKZyKEJ/ZuxW/6d2ovrgMZpn3abU+agcfHzrTyHjd/BKf3EXiu7D3kXaBKCf
ID/zNmlxuyrQ0AAkRBzBkWbwLmrhfVrHqtxi8J4sLFwxyZPFQCp1/DifDc9H5f28
Gvjo8kNZkmFIjWGMXqjWpLPESD7VuT8Sjgz+iliqB7Z2GxOF4WxIhDt2ew5pPinq
me5OMMH+YllAOQXyLEpq/6oInjp71BfnIoKssmGAYLgs5L7rbcbJUyfNpdFZDIU/
Rw3VRTJubjDlgX9Q/ElW0ZVC9q5RscUXFrgz78McDGVUOxWwhPcuGCXjZLZg3Tsn
7ohJjYgzcYuDCXUxlL2dWMskwSwyoe36S58hU1fRscbWiHHSW5pbw6mYulCsZeJZ
u5Zus8+0pV6H7pTyeIGhgZvH2DfVqjxFWmSOdxVvRdYZRLYBhXnpaTgUaGya8/ek
6BGGRNnJJ0bD7FXwFrGe+80NTR2km5B2ROsVI0QY4WMlaGD5OymJfsfVWsNf6k5n
+bgemeQ7i8ArmSrt5YKelebpWWPUVqDHMNA6S348VCAMwxTeoUxOofAAyKuUJySD
00sni9lGUsNpZeofYaxpaf+O/xRFTEA/+3OsNqvyrk7+FRQNRNGqgaoUpMWXX2DA
lEeL1Kpj+7zgiFOrd8i0jdEqJlzEj4LrFuFdjLHrDDm4gHWAN1zCFN0djfdIS57V
8FqKMQnMw1ja8zMMIThwry7ycuQ0X0ySPtrPmestSozrWMZRBqqhEvBPWP+FNKq7
Dji8MMl2Vi1E+kT1TrUpRF70FITRKxtqXk8VAlP4jWuD9p21UqfcX72UMKueY5jZ
siFrepU7IjzpY9WsJsVOluYV6QhkspcKMFrYqoI5JXhgUBI27kTx1l2dbT5LFBo9
XGBrRlV/7j/JNAv/KEkJaLI0r9rQpuLsSY+2SueBYP8lACGDXULPjqG3534h/U1X
60tc/de/gyET34XuKr+HjfEHmREXY2xSXcAEF08tJDG5LnIZlgSQ9dvWeRb521C5
B6r5EP1tc3OOdGRjMVMcHrH2UWP+fcWUlamnnqBxdmFs/a4mmWYlUSOAbWgDNIVY
rKjsVpNiLtXcAydwDUH5mYMKYkOrh8CScYtHt3ExY+Rgc1h7ZipZK3McKGslmQhN
prnqVouH2HSW3hCOQOzOKrXzWB+RlrKeZ4kSFY1aIHQoLth4pFS8yNBG/XKCrwL5
PIR9cjnL83DAAevwgFLEGgwqV2M8cIx16ZvWO7T/NhTckm4ZYrpUeT7142JwMGuN
S+X4cjZ4V9CvKI9yeC5Nx82g8hoWYkNu6x8TxKg5vUI5MRSgx9SC6FUEi+K41iGx
nKyuCbHUz7s5qZfFnG61rl6kCdg5kPv01IZfvAlD8xlpy1jt2YZwpuW/Z/3wb1T3
pBOa9UNHqFJUi9SFUE+U9BpiGsFesuUHveTIkPBoBZbAkp5uO7vllnqV3zCaMs2y
BcnMJEhwRwTygdktOlBicpBfD8hIJmvNL304bfr0zkVYx2oui/VWbT0ffKpvIogh
zLOrIfrOE+TbglS48T1xm0zFsKsIhcccbc1e3FBSCuv16TzePyf5CF1aNGvhn9pZ
S/fqqIZ5YTrhedXiQiheaP7OxA79rWPJNMilu2sbYTXBDMqA4va8C0LFEXk1Idd3
CS7W6qxSMJubV/XWm4hfWcQoSK8gWETtQNAaOVC1HgPt7Apd6xNx7haBYbf+PBUP
tsHWF5FLB8enf8UWwCY0cJm1QkQjaMckXlj8zXNFgUAnk7a971o0JYpzDxP9ww9q
RO/7p50c5SPxfC+L09pQeLzt4cZ9VFwncKSe0NrPySxK4jII4eE6rb2OCKhVJyJF
l/WsuKTmzM8KgGTqzssYeXlstttNqK21DZQaLqlyCLOeskJpN9ZsNs5I/le/J9W4
p80bkwo/qeqdDYBeiVvrjW28ko4M9IYazOvpDGc5EfUdtQ6GrY4CCEnd7T0nsmeU
/D61Z3SKarHRGw84Pold+4o6rTpZG2M9jH0hZv+OD6zn/CG56yCqZ5Bq77D57BKV
RnS+HOoLZz1o8MYZ6bUJqc1AneTsYDdLc1wVFIDk0f1Zi2nqk/yWYVwKVuST0Yxx
Yr94I81otk01S8iBRMgVN3dEAuMjyY8XOrbcx99bkk3HELzQbHGowU8PWm4tha2J
GJ+3hZPsE30Um1ZHSWCU7hqESLSV5nrB3yLbDPCwuIOpXwfRqys34ubhNV9iHgns
TLCBNEwMec6qpadfLnx6ySwodw/jcJaVIgZWJdS0R/yCaENf06gBhftZ/Gd94Kdj
p5A9H8TtKexc6SBStNRRhEPt+Z2aRSaHyA0CfezrkDOT0RqNAnoZFk0DgE9U5g85
B3tHFrXlE3dvIuQvm+ikVHUAiqFfddA6NVB1jTq2pfel1cPAlUIIgzJ7+BPL8oPb
w4ab0ww+CW8R/4srwtO8Pb9kjs+B3k0tk/PdKJegYpfQUMb/UMv7ygIagzgg9F+c
yf/apv2FgOSWq7MTGOOnpP4s48upKpyciQu8L9vrNv9aC8sdBh2x42XP79hqroDb
mEZppq7GAje6wEY3dDOW7GATuxTVX9VEs2osf+33duZ6Ko4VEgZ+txTMpch3raX6
fxC2whNSZ83QFQ7FHJu6pfYc9VUeX8gox3sEmpjsBI3qHFIq0p3IZcxYFU4Oc/OL
ZkCv8trEbDol3bxQ6R9qC1mcvCheYRPfCBM9LcfeUDQZB0oDyb+IrlVnJobYMfkV
U9eeqO2qiSAlUb/tUHW/2kxDs/L1eXYuPArPIMTLFqv01dN3K4BZ8vR6SRWBCVr7
V3zOFxx/M+Q91RTpyTNZ4s/RRvtGCDW9/zxJkeLSBhG1gjPrFecU0FJZBsJRo5Xq
jue2wZcUsXGp7uRmM73ISnmFRtNkZ97WvztfFbmZIgf/diyOsK6R8MuIRb+TldkJ
uYsSTRTkChPIHaQyZSv7eHytsjkIk4i5YYezqqG4av4kE9vnTNQ0KvSeIKWlMMhM
46OBi5vjADjABWWk5+/GQ5uAsgNqlrtYoKIccZMXdBPPO02CDRqxvGPaTredpoIo
pNrxqJYC65OQX5qDO2M2HKaauWZJ3fWV6oUZRYT3HFhKxZ5s6WESkWSOpV0s9FMS
SNxwsjBNjKRNQWYzVyNe1eAIcMGbKv4i9j2LzOAJ+TA6aa3TJTIe+JW0u8myGo6s
t62z7N59Cz3zgBbtDzR3GTkh8HctoaDBwWXySrqUtK3quLv1nX0y5FDizhJcMHN0
LJY2PHq3JlJrDwWOQsDZ672SoVUQ7/rzw4w/tg8bbefGbC7GP9P6ANi46tONFwVF
WrnrNR4uBq8XFidVyIHvuAhN+hDS4f8xMJ+Wnew8dWtVN4FFaCVOX7+907asVo0C
2utJZM7pGx9/pf0pOY7B32ed/3Ly7WC0+KHUASMDyc9O2yfEyzk2+CgAQkK14W1P
04PjCahB3nEs6FT7piNF8qq7hPKYkg9x+01MFda3VycDjd45+w+UgCE6e4NmOWCN
lELqyvlOSAm255QIeK55udaWmWPgKazSJSo7ytu+Tf//NWmuIX5eE8zFLwhv7Pak
FUR69s8RfM2cuHOKjWtDhM+AlFVtQnPHeypaMXhiz7NZed6WsDjyn9IQLaxyXQ9v
Iiy5hBKDQLUuj5XY5QNTMkYvHyHZr3zjO/hQ+yeg30Xft8EOk2OORPg58oxqceqR
d/b9BbgZvJhocbTf+7sfUBokD2eaN3KyDd9FnTR9W/s1eVqQRM3p/lZZWHiOyBqt
cErOWXzOCE3fxSUz8xgNLaYJvr+ZcSM6sj4Fp9hqYQ4Fh1Rusv3DDlhrki8KIu/m
2A1UgPFMEJ/nQhxdZcQukDsBEVg8xiIjnaP+L8y7WKMU5e0xk48Ws9vaxWPvrFsr
oY+W7VMwhwdLqEpCb2lrwng2KBS1KVOghSDA0OcbUal/ck1RDT9t8NaxOonSOciu
aGuWFKnx67jm+ksqb723YGszQT2erQBZt79YZXIt1cxfcWE4lSARTtS9v/gn8Gw+
8OSoOskmSXt0/T+kHmhf5+T+79gafbgSGCkMhB7XosD5JtdxemNOABEcx4amEIT5
uKliXiuRdnZfpLJntCypoZgfUPjEmetv+JnEE9QRIMRTGT7/GREQ25enyf894gPq
DCeBf4jQXbdGQTUtlIED159TTGSbWHbWSw95gl3opXM9Ng+dO7+wL2bIRRLgh/yw
rXLy5TosG/nXCfmr+G/M1iVAkMCV21OhvjZ+MWgZQir7ye30ZvHRutJAEkBqynsg
SxaFvdCe2S3joRxsz2Mo2xql2wq5Mtjz7YPp1r+f+aFF5duNuWOtpJnk4HibpyC3
oZMMs7SkLdSkDePKXXhPQuFyLGdPMosPRDpUppS4vL37rbFfuC376ZdZhq6VYor0
HbgptOLWfNc2fdxwlVFJCLvSOYFKor5AJ7YfXvRibF3JNqyqZlg4S6UYwyZm+T6q
7q3SRP1zFpywY8WDGNsO6ngTnS204+FvHqwRVdafmXLuQjTbs+r48L6jbLOrfSCx
2dTxco6UQ6gb2nijHoWNA8VgUOD48eLS6060ZO54iX8JsQUPXQ587gw/yGnby0Rc
pq++PoABFmkc5SKk+mazW8mGccsoHvIqJ0fMJ+Fb5dqtVpN2MZnAc6zqPQSGE91Y
1cgBnyrrWLH9wL1cyMtHjprDArAKkJiNj5ts13Ea3YAOzeFrwYkfzDcADgJlvzg9
/219TKIRqieRVuXUyxJqMaM9cB5alpIO4x41YjmbxnkVsRJoaqNI3IRPTNmSlSKa
InBj0OYwJbINU+MPfB/Sb7GjQ1zuV+p7p6cEA/gfQQQ1FSBSrkLa2IKuIKZnbivw
awzsekTTnhL/Qfc30urucWNBr9aQx5zUmSf5z6GnndmFSX+QY3OeVq1FXHihAkUH
W9iKPsbpIk+ZSGrJTJQJOYMuJcnN7A/0aW5ZbW/EhE2vkk+mg4UWb51j9EvaBxSS
7XWG59Tmyd0XQ29C+lyiXFIZRIScOJ4tA2Qh3RIqyqkJh7ZVm3LUtuxxol7Xn53L
jnSDyZuivP7MU4aoFep6dR9XuxgjSzpAMZQ203kXw13hqmBqk0Hj9XD2l77Hv2BT
7fG2anNdTDtwB3lh1SYHStthp8WIRcc2f5mimVIUh61Ds+HK/w+oUjGmqLjfHs8n
jb8IebXq9CNTfsXytTellGGBLI+rqWsDXruCmsxEhyQKDBrBgiSlSUAna6f4w4tC
nACJyai3/qvpWj33jLVb6Kl4kEZjLcOHBSPFEZbEVg7bVwzjJknE7FWPIhxoel7M
oTf9GEyVy7xKCPksbLCUPEjBkMXyGt4bjP7zib2/SM8fslvJ5vk/PVlfYtPpQOYM
dGg4zhhQskloZBBMtjAwQcKBoyes4WvsP08zynb0OLBDfkHE9sgY7XHJApsPsXec
eqFzosrOQnEoVdAuVd7SVx+BUPn3BK2ypJ6KMpN0C99qseMnfmXsKtYOkEDTOrhO
l/19w1yyklugVzUutZqkWlNUpTc2Rwa5ZmgLGr7QUQqAct9rC2htQta5WTNzQkm5
K1ac7ei0lDBhEFj+xvj6SkKHwO3zdHXCwB2UyHEpH/HoUYinSWcYYgR9ecTMhPap
lhjr7Z3JcAO8MXhQuLkakSAS+MgRazKN5f/vxN8ruKFv71HzbGwgOFU6DNqHfLyM
3ht4AVBpfClcrJ3JhhO5lsqiXnYwv5i7yHiVK/Wpl8B+pUjVNHhVZjkIGJLYEqPO
P84rfW3iMrx0Pfh1afWRboA+Dwb5WP9HX0n3LDhiVdy0YCxZDKYVbGmWHkHhAXNY
b2airNTaSQ73iKzrzg9+z4JwvpLq64QZ0R2QjmxzZmi9/7tHErn3dK/430nTd/yR
Dnddvei0xByCucOPfWetPNqPDN22lMlae6A2VJAN95jtMZyIHDhcgWXF7bZ95iQN
Lrjbvuj3t5e6MMLXM7Gy9gZbC0+zyJGsnt7kJ0TncTZWdHcV1LZLJCU1Aa7AmaMt
H43yAu2lJMj1zupbMPwbXJiUFq7SzBFQt3EL5fpklV5spLN8tZFLqEDUvNErdCjT
pozReNDfEgc+x7AFyLsF1dfAohdIPU3vZvQa7aT21UcIxBocEagN482rTQks2xSJ
Sk+n0f4Sg5/+3KTmViyQpO+lhPKuUKB4WhSYsd6XddgeMw6JpcApkUe3ZrrHCaTT
vjmzo/joPhIyRpIflHGU1FkqC8Od09khxzHC8882zaQQ7+vSoIFKsalqxU/otU85
zpXE5Leq2qeop8MQ4V4YyUD29vFnt3mCeXuqwiDkec01YJlArWtZkCeMAOogidRM
vRD4wLnRLskRcyqMqjDI42Qqjbnwo9oGTB0jJG03elDLx62YFE3TYTp+Oy+40g3w
DfiSR1Se6v+CtY9i5soITJ13ym3zRyC2Y8jVuAC42cir/8Q12oGGqjj22A8FCTp6
KcNsaYT9NVQ32cQWqKGmNXax7wfe4XVSQEJ6GsVweyyZILX54Wt0xaW4Wh09C9oq
6081h5KiT7x3+jqyw5YsJZWNb4AJYJxm5YHhRVByLXRNDIg2YzYHoFKRFpgaRa4W
ddvjmv1duBtGuV1eXtn2at7GlEPwErI0Vmp4sbFuWuDW37gZ0BFGIVIjFU6XavKp
HQEpDE8iO0HubWb9qX/J6h1mg8MXdEHLwXPDdFNb2E9XVxSmzcpru718OC+Don6h
SC9Vstx3hqGUXlz6aUjdxaIFlnEu6sphHCeWlP1ZjuPnqsLajEly3LeLQRP7DaO4
BxEFfppbcyF4kD8DKpnTN02U8rAVLEVevxsOWd4jr/C4ZfyZI2UEfS8qekVNAk48
uguNgHtHSyCYYKwt6BY2GCuyNOjopFuTZ3e990zuruDQ5AWGaYMiPTh9l+2wiqyl
mQ2sw9vVZCJPBkoYUgFQQ1/5GlWf2AeB+p73ZiK+cO0zp8749JdFGMpDjdu0EC4d
9jxFfE6FgCPzhQrkxM1CkWNO+0Be0cPKUWm5Rq1A5fvlXvQatU1qVf9XznxfJrp8
u4AUhPihGdCIx+aBAMdBIwpCUZIp/CoIxV2ibDQk+XrqlZOeleEgjh2wAF8MgDbP
Hh7O3vRSYGRdaR7CcKDCKe5o3RP9i5Sid2yAIcIMRq1DCHoZoYfxfN9WEWLb4z0g
sMvrQKJrM9LEhHa9GDPlboGx9zSjzjoPPeFXQlwnQmBhUuloxncufiiuhehmqjnR
BZy8VTZNGuFbQIV54NUpPJeybWr3+sexoU7qdzWahnMZWByYXKW3wkWc8GOJpAkG
R/eChLFYxzOqBgqsPN9SUfSMpr75UqWzVah2zEYpp+xF7T27WrvseU/vL35J2/1s
otDEMCvAtAfbyVYGrYkp+ihwmOF4mKWIqP6lPuea3r9yZgA9VIaCMJAdj6Gc5FG7
EjfN8s0ocQo1BH39WvE68QaXXCRI5FF5nJ48wZhTZmFpSpXBTFxRZibz/OmhTJMn
Pgfg//i2gwPjCmivHGvxhhw9iur64sA9U6uJmhxj7X4+cGXulPe32J2zjq3SbfcL
P/amij3sEfQ9TS/8d4mDDT2tyl1DdG6OK+n9lTDU567jqDysE0ZzeuWbT0txT1Kp
Z15+vB7JxMSTArnhF++m/rIMrWn7pF11KE88bMVSwRVUjPxWxfJYOT6yhvzrsIh/
nI8YwdWajIIVQgJvRYqJ88pACytdJ6/EjlggtH6i661i23ZH8nnI9D12CYhxC0Q9
oTwusn2yowKQgMAFSq+vVk2p/WnHQ4DzRf+GF7v7hHUbMZkUZGDj8Aq7gRNw91Yf
xEsAdcfN4VoWsqJvzYvpP0riiar80TaYGMhknGXByVbuu0e2P82pZNpOMiiMNYbg
n40fOmSneb4MXcqXxliubQFouRP9AQI6Fr0uYsVJa1kMe4PDNV3d8L9rIlNN2R4m
QJO4HPGGy63hHe9vCIaGtzJ5nhnJnsELoKiKsz6hSrWxDfuEpVxJu0In9SVEnJke
urJ2Omq8RohPwhAvGEh7nP2cO4E/WJ9wys/BuRu6DL+JyXPB0RRhbXCVfaCcsV85
UH0s3vhgUug6hBBk+DP4nnk/LXf38PGbTY9nJQVEAIfTOOJ330mCRFgV63SX7j0X
ysKxEb8ljf2G4SEh2najEoXfwIIzZ6Po+AK8r6VHOg8D3Tl+fnkJOjytgCSqA2xV
up8/vbweRjeBvTmbdp5Ti/XieLXE0Vly7jpjpreFT0zxz1hfuWwGFTSmnrPKRgYr
uLc36i7v6XayNve6uEDWHecaE2BgRoVKb2zrNoso+MSFwLXu1IrLlqOwk1h8S7Ik
9rHIFF7051NlN4XWF/CzZ/wTBUMEm0IsBjoUe5NXpvTeOXXJet+Eerp4UYq5dpEO
Nq3G9w3MMs7SIbtFYNAf9FWp1gOxKzouAF5FoxorgX2aDFDGM8IxtxdfUaLhajaW
O18Q3utPuJDlJiBJGJz6ciD/XrlZMJ2F5JtVRDyq4/+gbxVvF8tgeMxVincAWANF
j5AFFFxARavRHqdwyLr2WDlDyjSJIT4ljEY2NIDf6Gm1BArUAMJeGSi504Y2QPXz
5Vn/x6mlnS0wwtg16rf4ZEje+1YIcaFjS4n6UCdeiNwG/EzH52HYFYBrdQjLXb75
p/1oOrKUGXdyGH4p4gnsab3uN9LnZPrVUKgX6AOT4pbacP7jMHyhZgJ0etrzzGo4
c4iA2n5a9nO+xJzzTxaBFSo+eOKfnVP4syYhNGKPwdnI+tsrfL7Vw4+T8gOEJ5yA
8W+l9IJaBes9cFLcg9RV19CwhjcDiCgfwjJfVbv3YEKPGWpEAdaJuCeCY16CmEEd
PjOIxjOb8+Bec8QAK++kUIFluxF0kmHjrONMAXmDxPERte2qZz+gefkOe8Nz1tL6
4CcyZOH7QaQTA1RVAuFNWqfIlR19JNcTAJPancww7xTk1miVbZFxkMOEK/sBb/UL
359MOnHDOCY3Tec7zlRVzzB0JZDbvmeSmYST0DnBj+6wEQXX8p+thx8zXNojSaed
4VQ39MzIZ0SZpcQreIlreGTWi7vBWa4Q3Ndgzo7YigWH2HqOtGNl0l3QpZ3kxVe/
VuJixJxbypHvINXu90M2k9dwibd9Dsnxqj5mJWJRfg1bsfOxI8JP4HyHLshi0RiK
CHKYEDoTP0/pITIy50cK+c5D/O9iM8ndTllz6NeDYW/b5jkec+G/CJsGjW0rOOZG
wajIZGsMhlixmQnp5U8pSWjeHeGTQ0WsDG0bkzWkdSKbXXE9BhnqqqpyUOrFkASQ
HNrFWTdpE/ABwvwwd3/iSpY651L4cgdRtXwrmNnmDpcwi2SBXHtNuSEi+2eNNNMA
UP9rfzyxpOWbbom5m5q9lM/22xuJBpkSDtVMhsWroRXouV8w/CDBKZamJRoZLj/m
jLUe+1CLr6Igwi4F1wqq0OKUhddvagy0cvJ1HLVl0hganYn6pl2GghW52bLg0Z6X
X13RluGEOkAiKh7/Gu18gENLLJejM76NWa39vZbTBbjhObjLhl3oJXs3zwzasRjG
0hcnXsqRUUa2xGVR4UHVs2nmbHWP1ko4RQUcfO3PF09MQtWKLra1iPnl5yD87wVc
0PP5FUDrdruKq/XuQoZeyxQieMQ42+tT1uWxP87cocy4Lmi4slDspIv5kKIF2mTi
EuG5+1rDiTD6TKgFMvuESmWxIkSTsk1PVdvnQuLm2i1GdZPU+4Oxuy7BKlGj/EQt
1kmq2j1VJSEriCo7YuDlHxrnrChO+pD6fBpM3hNZGp+XMCUmbSplp5Shpjf14qBW
iiUlu0W8eBdlysSNi5t3vSzOFBvuIm95Iz1ef6cRMI2LrYSFo3xuh6MlkpZKTJgT
vpyp/ZuhR7r0YmTkhO51jbrbd6JCTwYlEfRAqIFHhvI/CoGdEIxoHXMf9g19a5QA
8/Kz1Kymu9ZoT2BMGjsbvsX1btdWRFV+vFtaPQ9aa1O8//Ucpkm92UUeNJIhrGar
E6tlSO8w14p7gbHUopPx/DaqMt+jl4zwTv+ThLKErfyL1aZ5CKEmlQOEiRm8/nxG
U5qv4UODksBtJVDrLhE7khrGfvIzwvVv3Vq2z8NcTN9tBRH/sVHVHnfHUDA76OxK
7Ehll5n9lWOBkYs+KhSdnSdOipCg4dmL1v+gpXbj39jDQYsobmDTFVk59bZLD+qu
8GFBMLbkCeUA0Y7v8CWSqPDrRw7G6YGbTWQPA9W7O1tPR43Cy3FKp0Qa+xN/02QR
NZmkOVjd6uw1hKuCxJN9j3FKgJgSNTuNuVJc9FLNpdhZhKbZ2LgJTF3ojAUpFJqP
416u6UqOcQ06CGYHazzzzfgCjp7ZyeAl6l8z9jKcPLtmofRpOmQ+UAOdMZJYm556
epbtc1rXF3GEJX7cdE6D8pj3usmpXfSOd4pmdqj6UI0ZqOu3uMZwIaOh/ht/MCLH
4AFcVnq7D/jqphzywI2Vi7OtGLBbmwjOALtL8oP+d1q1JBHqtXp+y6qDel7kl1s9
H1MO44vFWMvYDSLQFI5LQTJLC1TCoNEm7d3vdbTPKLpZsAwlhLbty7C46mmUjBQA
vhwPwNC6X0S6kkFnUYnnyem3VfpvdO8kPCd9rHg10JVhFtDYvSGEKAy7H7RoBxme
9FoFkQoWORhhfIPYvVr0PQfCvWtBeKzDka54KJV0+P0q6REAkqspgyG6tqQTPjqw
3LakpaUi4mWYx9eYa0yoT8Z3p9X2qiq+fjbBV/pK3gdJGZ7XqcaCr1hBfdWGt08k
Qy9G3kEs8JVw27N9EM7m2Ccx0i6twzGf5auaw84fZLH4zTfTS9z/AEULrTTxa7QI
+1hMrZKB9ntefXoJDKwR4C64+Esftyd8laSW4Ygxox9zOpNzaX4rRRiUeHszGkGU
cN9Znk6D73Ourl/GszSSNKqKSCgJzrT5+WfyvXdzc/9gFhiKyrptKhp1qhUcKGCR
308nARURgWCLDq1Chad0TWuOGXSzw4nrb9UeVjNbS+hqVAddfMMAwOa5t4y1SWGU
X2Tz0IwsEIUMqBmRWohKEHebAWmYWJI6fgJjIEAfAmFwtmeSkbBrUYavgrDtBuOl
4sYdVkY0wlBKOKavCZFNMl0VHEtQ6JyTOvOO/24b7YT8lSCN1e6YKX0E8VmzrP8K
gu9knOFJn+BVSB0Usa91Wdk25tXp7WjTkFlvknXSIzEcPjL7My6QMIB44kM9HDwf
njLyTkO6lNYJtS3AllBKCZfkwcKVPxxFRWVrtwunJNyXqhn2GYGkdQF/ldFpZ6vK
NZSnnpLhjmy82nPcM44g621yKeCPvNuM94WTqatUs2MuQumX+boEB6AhDhB5LfBa
VZ/e/zlZRZ2bpLonHmOKLnHUlK4OH/8rVNZCWk6QLliWtZVtp7Rv6wb4yLFCMsCk
+B9ZV8+TQsIQfbPg+Q+meLRTGZjdg2K8kM96LBOLtIGwOkSIflONwtQfHMKyr1Zo
cxpaZBtYRCA0YBpQCTdVL+pVCkjzZmoY+Rbp2Ogdsqw+QVCR5eFmZ4v46V8myzIQ
WlxwxRcQCB/qQr36gQF+OPYraDsy1WI7wmR2I1U40pcqtHVpHBU/s92J7LqrM+Bp
ctxuhfvFJCmOzEJ1gc7Fu/GKbYGV6s8riyPIq/a3xBwIlPD5gJxYl/1wD9LDlXin
RJtaSTMsgaUz/Wd4zJOXhnzORqw+AX3ws1Um0HrFwvbdJtQen4ZcRTz8kcsPd2zV
hFNQqFuXU4Wu/B0cHa1ki3whybmOgeVGceMccMdiw56WBMoZ0uMWB+26KL+YKyRv
Rey27x2FPjypUSBj75EDMAxkpzCVn6CDnZ3/fHC+Zi11t7uhDjPoB9lgHRXmuS2k
KCCQNbIqsyK7azygde0H3bl9+/g0ICuTsGstncsoGoKuAh8cokatrpcvZ8KIMtoE
c5NsGNXDodhLIvV6AnaETHeuqDqmbNEz4UhKON+UfvvLZTNLd6NErjefT+qHDrez
m3i1iwQ5rxPJFxwxROpqvVa40zJ7eTGjuGcBbqhjSVL8tqhA652KJ36GYOG93fyN
g/OgN1RJmOYUJp+J5SIQ8EMKOeMQve/Koqsoc19yp678+/RmnTzhQIcyazOl4d5u
+CGOS/mB2sRXY/Wgh5wrC7gN5k0mCiiU5SDBlmgFMgAmLwb/QQQXhgcrIXswoxzr
LD8s1LZD0hhWMbefPRiD++eEs8wvRjFgeW8z0cCUkhKPFp2TVyMfjpko4262bnxm
/9Vpy//7P0PqsbUaQrmhvdxLw5IXdO389vGEft1IqmU7bOzvVIld2YU//mp6Eh30
qtEOlb4Dt26EphdVDpZqrA==
`protect END_PROTECTED
