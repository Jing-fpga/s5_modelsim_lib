`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J0OifKAoK1/lICmCKsUMFiOTcL0iDr29bd3heE6xxTnEP6ionT+OWTqH8x7Ll0vI
9ChQ4nTEJHGAUTlaZYyGqka2xphQc02MkeHPW/TtGzOV2uY79AxFaafHysddl1j/
PU9HFSon1g+8TpCgq/XbtVlFuCVE/Adx2bbp89hBOLGf78WnfyOo4eDLQfxVx0OM
DmpvHse3Mzi6SOuhkEiZQiw0E4v4BfAE48gkKZw+YahRZM250xnHLDede7JvqCiG
kbvvb2rjm/1C0ZSUalyaD5aS3jqEMaTJ5O2mj9VweqUudofVfO0Xj992BQRZdnVO
7b1D9ni9fwDW6WTIzPCaRTO3jtvRBINrNbzCjcKCs/+XfMB+a31eS+GCrXMmQ8TP
9uXdXdry1NMJHhSrv9KY+aM71XxKShIbjXbaNOmygF2CKTL61eG7DXMk0L6Y0ogf
B4dF4ypK0cjm9BgDR3I+XXWrm76xRU86ptSi3uLn08ymrB4QqNfmMmttZ6IAMl2F
rqXqdOtunxj28bQSoIG1szJoBuMsHjVHQVjK+SfJjdE+vRTUqFUGPYIB5LLQaMNk
fEy3R7HHzcWX55zd7dteyd+dTwBHDX5CjzLmqlGubiPMcGhzuPe2dEdBOlt0afa9
RVAcpiq4KDX52eubXShECKMQ8WQ8NQuDrzfltrATctH+HslC9VjH6jParNC2EM+k
QnML+88JrUwtL/OKDTyB60UUO+TFtnHo+TjjP+4ZtImR70jcuC7smYzhnkFN1wOy
f+0RbDpbNQcaino44Txn9i7vjR13k3jG9SijqrCI6Xkgs+xT1bcpiqrly21B4EJu
4bzb7QnX/rV9NGaVA9YWcui8ySk5zbD52qV2whGMKZaOrlaABcn1Rk9QifQftvc5
HWrG+xceOz+pkw9jSd6zSpTZBR6SV0K+DfUohnaI+wZwcaCAJYl6/9ZhDpF5BN33
cH1RCVwsakGsvJZKFGTfIksiGmvRHLfkSITe6i0hz+3qgq9twWmtukqbz7Y1KMkC
`protect END_PROTECTED
