`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QB5rvLyUma088wvpmX2o6SDSS0iACJN2RX1Rs3aZy5hsHhqrpADy1VwkvvbJSXNA
xSd7TXmo9oYPAk3ZeOQQXcClD78sgscQ7kPslVbFLdUEg/opXlGeE8plYAbr3SOF
MznMC7wwl0uPiXg2eSHFG6P4XIjWlC6INyq0CJhUcIMLKmQwk36WyuB2kUe2KAdj
M9nL+ow57l+VEI0FIsGE1CMnNcQTwZOoFGkLTSBIOurWgaSRGjyZ01sqtK4JBCDF
9dvRHQXA+r3kPAROAtv19FIzx6sgjyRYvenvKf33ymkkI+ImvMz3/rpiuEC8POW+
sPs+WHo2ROuM29g6c6XNJf8Dq5IfeP01jxYNnx4+uuKr7meOKmkb9r86vJvKq+SK
hlMH126WUddNbmcLk0ZK2JKGdRENBc6raxHeu+iDa1H9H6tdTd/Yo5otZ/wyZ5ws
1s3FI6J+h339ac/T4F5bQZtpjh0CPU8cyKKyT8kgCqVJh1/fig69g9aieETzxVjl
vPd0PIjwfKlX9bn5drz8a+5WWaEpTYaKC/xYr/5kYF+VdXLpjI0pgzWNVR/0IuM2
e5dXqgwt8QbF+qsYm5LYRXUlXDPQHtOVdwQ5K3uHQwg=
`protect END_PROTECTED
