`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BGg7UAcj1gy40WgK2NVgHg/NC4I11bXS6KWiihAD/87imzGtOet+52dJoXRKhMPo
PRb+Jn0HBEP0LU1S/FTiWW5m/7YgqrJRIba7AFcPbCynmaet9MObqEInmLxiXTj3
BI6KGjsazfoGhY3qw5rTsWzZFIJ42g2bVeLiWkvDpkifuBmxa0GZoPfltldh8a5I
hKPVhc43HbDSW7lmBdgb+rtpgF5Nd4SejKEyP851lonLXdNwzuPq8wpCzWIIXAd2
/iL9jYITEpsNqBHXe3UXoU4t08eXg7yOeNVh8mMq8Yen9oQ0gO8sHJXZ2O4S8uSO
jvPGuhEGxJWJxbi9yfBGWNe2g+KNTPxXzCsa9jQdxmfdZ3MZ8yDYLUKLRAIN3dTX
E3/eBBh3bxUhJ4fMt1X8fKwVyavNTMft96AhB7hN43sN2FT1o+KvnAd/d078y1VN
mi2J4fob+r8JnNi8/vkA4WHdJ48Xs1nDJrEFFYn1lao954yWeqtiogZEwZ7RT6mP
lugBbWEc9YDE/qsjF7r3N4eLA2O64wcDu9ArAN04kFu16yeg03aKK2QOpmRKlfJk
2qc+4uYtLxbgFaGl2U1sPbtjSy+gLML2j7kGgU3mWQS5fEU2H5zYroeQQhB5tPOn
mkJeIYXjrJyyGE8RbZCcJJZRCy5zPnVmklyODKDGmkEII4RftjrDRM/aq6rxx1ZT
CKPYA7JK55+6HVEyP4L12wwT5CIDJaa6R5r+MTmsUf1QlBKiJ4HWNGHIxNnSnqsL
svq5g/rQntiYBLxt8N4t9djF/T5c+o9NculThog3xFOrVAsQii81N+2RL163MGXO
TyaeivxHvuK67uoF1ja5wvr0qq3p4Ak1JpI2qRo3Okbjw8CAaJ6JhrIRTp1gyedm
LsFZIzDjzeknTM700AukjxX2tPoWnDuh58fA3qxj3SjtxMnh03yLSmQuNVUDgZPa
QfGxzN80T3bD9o8ePWrPkFhpMJ/umGUaGo7Wd4U+gSowVnnmqrl1xq95Wd8jYyZj
Bi3QnEfWEe1oJ8ecrDp8djWCUV5gwN3yoIxBQGILNEXMOxR1F1ndf7XXMC4NUYKc
HnjyPaXSg05rsoMjZPQLMnmFdvzByrsPqhWE03todoK4QYqN2B7We3ewPIgOkNB/
rjHlp109A746h43n1yQwPnhcRfUGW+08X8F5ZJ5IaUdGI+KzasUKfRP2Qg5AUaJr
bqT9NJXciHwlPzHB/Y18th7/+t51mg9Yt8Z0BTcdCuzNqJJLBr3U54aY5oANRgmq
IwVr+0F93PxsOLHFObH9K4B3YR+4IHiXqd4VbQVzysCXOmV690hCsDHG/hAnsN3K
6+/vNC8dvGDGUjG3T/vWbY/LAursXDisehhY2aYAnkKwt+qczlowfO2zjFJOsPMs
J5uXrf9TGSw1S9CXn1O8C1ihHBuZeKKkjsgLbngYwpacxAfhthyw5rgwSmn0BDC5
vCuetzC0HNESa8KgvpNa+Gi05a0mLvnVNgJcCWNua+ZCfzRNdSAWVqKNE6XwvtGf
tjDEg6MuvigbKLjUnYtf2KrmbKdGbzNuB0TROSVRqJVbJGCDmWDpI88tQvi94Tw9
gOvGFK4wvXj0HKJZdBsT7qu7eB5V/enki558w7K6AZs4FHmbxBzJbc1zCcyqKfLO
MPv4vquq3GwuHGOiV5Ix5Vocx4v3zFyLd8kwacra4zSUx8FXGKhbEuo0bcELnGO0
x+mbqto1jrbDnEMLG+YD/ky5p6ddT/fxWFBQgpPZNDnBv5ufrZ3JZZWAvYr7wTBv
kADHef6NmThRJESfHavd+6+YvUEIWHeZpBp2s9uyCaVJ9lD4qMF2m/jZL2FX++R5
75HdsXpw2bWvlJadDp/qnDib6UeqcsCYzt0dhAOpJrAB21s1K981dcVPHXEHK9i7
+ggKiVf6wxejZbOcDp3lFZ+0/uP9xF7vdpDxxwdv0+LyvUOxWrpsRz/OniEbP5Rm
mnaHyWznMNAIZBTavZ6YhV3+yonf410cfcEC5E+gRWQUprb2xzEJxlLhJrJN/RiR
8zfDjV++RDBVnLmYVciZ1b73cl+e5Pw9fSoCIHmIB1smFk26YmHvXXKqm08WFa5p
eqAVEZ0pnqDkcyZ0BbgCQ35rBl7OubsRQX6QfVRzoOi3BhIAuzhJGsRhCRFhsApQ
wNpzG8FdRF/S2jcZSgQRdBwy2tVUESJaWlqublV0QR6a0Z+HYRsfhZjBQXT5A4mi
aQGyIiokWKE7kpyfHTLeabRWD6p2TFBuc9oTicXWkIntg29hS8rClRBtyO7GSz0b
2STU8CTuQVkBVuDX4NMby7T4p0y8BTMXXyFI+5UjIFAZFMo4FjxvYovN72KnucfX
DLS4zm+WN9i4wgyqh8PwJzGFmELIT3aBksOqeYW25PQ4Gfo/C7/WkporAXc3HUoa
qqQJVbAKZGENF/aB8Yv+rFWa8Tqs0mtOrqBSu4wLTx5qe6U6uFPjjnl40wO8WR4C
ui2w7XFLEEx3yQVArDekoh3ylvYuX7sxYVs/auIn4RYej5mDLdpKU1De/+E3kzk6
rJbuK90iOJa6mXwntUOfQ2nkJNLwigJUdp44LgJcWKix3mhd9laC242JjJ90zbDp
mRPyOhvMFPL7UMx+GC+a9TsxEENHiapkM4djBPBgYrzupoNyXJTMSFk+wcvAnLES
yuIlEb5/CU7O01NlAkodBQ==
`protect END_PROTECTED
