`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OpxwIfWxXks/Xd22EVAYVotNlluSntCYKMTghlBi1FQrueg56NUeyLeiJa/RDKxU
HMXl84w3ECeNxEVggI1ihewqzB6FBJmsO5OHVs8i1ojTM1RSZrxKS51Th5VvgUpt
wlnTFmt0gFfg0whqNw2uZuNwTC7dVPRarUbZH5lGE7T2bL77gq7rhktNowUnQAD1
44WyArhVCvJWmFzmuxPPd8FWnKMHZgYchlpuHrjwqQvmyYzX0iarnD2hydicSZCF
e2UzrqCjgd5FAbCs8yloX0cJppSgjNbvhPDMnkLk/PXiZlhSieiSQ/gMtjzkJcGe
g1BspoIZGrHidwN0SVezN9BL3iquHZe6TzG+ktGVfPa7FKCDHl006pdR4EiKuOuS
Yu1omHZ8LGzSWCnDLWkuYjs+Cq8Qs55O8uVGAY95fZxoQMcmwhIPdszl+TLxKdz/
kPAiXv5hxZfWDEfJJl6qEKf9MOKuswSA1M+fSiA2PiGG3ZQEoAHe0dUlmKHMXXco
dWvlRvLM67QePjVOX6ET5w68wuJ1KALxhm4cgdWsO7Futg+zNG/eaU6GzOTQmTzu
696E5pdo/IER57vdiywnYx1spgD5X/xbZPGw8p9BOjIhKDdOXKpzyiIdTK3lyG9T
BjZK7PxCmb2+1nt+fqcBmg==
`protect END_PROTECTED
