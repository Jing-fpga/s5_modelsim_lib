`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cpULIKxXf4d3mmLFe7KPQq3oUCSHfwl/cmfxQ9NHxxf5YurNlxe9ZtCpzyB+C9rS
ljBdLRoU9I/BilrHX8cebRLTkFQ3QwGpPK7jvHP6MkqyNqDs8gvnQtp+dymuLtb2
D8Ptzj5dwi3Jj10Ir3D406CKLCTz+U1kxMiz85B7p7PARuR1nbctMeayy3jr2cee
piT1+/Zu2J/qrhBnaWUFIp0LRf79TfhgAfudAhI2oXD85rvexINANf291NQW/SLf
7OYJxwNV0mM3uAliETUYdjpsx5HBhR/UxaOOubMWF+n44kAA+MSjmyV8vsgpR3mS
cvnLxcb14R4vn406WRx4Sdz4sXRBRKY/Nby2CXTtrz1pPYJHfIPyTPu/jNJolPFb
vmvXifHVE5qmpKb76CYMC0sKguBnRHT0V7PTdjuIKTBYiqW2mYtVgbkikWe57/wx
bfADTmiwEVURpCRrVTGnjWIg/t48+sxjv+QpPbYhMDQIR8MflxJYyiY+yIGX/fNw
gT3vJwIymBOoma5+UzxHxS+Dn0XxnCnkpg0fksoej5XLQiRGD3mUxvkEa/i1LT9G
++qT/KwTRfihhEr1hElI+a6YB9geG1AsGFbHPt5L5txVjgH3H3T39e1BF7UTe0A9
kSMtBmYGLoXrRjPifeq8gG45Fio7ZawbWTYyOag9R6SfasWXF05R/HVsrMvnaYFX
Hb33OefHSeY+XLlFgq+3/POuG00XgZafZAREpVNPM+BPTap3LJbSSUnLGmmyQhq7
53p0s/Z7dTxqmNonTERAxJguH3PFKJo/Y7ftibZ0qYcF5C65FDM6SIkBI0sLgg/H
oDpSVIyDAStyFpmfsa5JUKjg+Pzcf5RoyvAH6r8uB8u5WwLzNw8YKSZme+W8Lwc1
La9aQz3jJOcdFXXkLcqiD/x3er6R337O4AqoqU4MnPTPAYK7bq4l3I3pDjkARUyk
SiuHXItT3vkw5IG0tduxLjQzFDf14t4K77oDkIDS5pqKdgwWRIRYp/ETdiPvmnfk
OemSLzkxcSUCywbb4JzID7N+NEogKQxwU7Gx2yBoMD4ScYmCsXF+9o7nr7AQr+QA
x0WQOIKtSbGphFaXzm7Jy0MryRyAsmD58gRtQQclMOITIPoa6jr4PmD8Ywi69wXS
maKhYkmWJkZYyLuEpTuzUWTQoWHdVkTK4cAxHRMiUZzjgGCb4rv8MtO7xVZ2gbv2
Vc0U9ISb9puhoQ2kLZtLDbA13gWBl92EQlFKWOil9vflan7Dyh7eariAKX1JpPvf
NQ1DOJ5txrWqF7N9qY0jgNiLJhgCPPzz10fG0+KRQp8rUoGGZyAlFI+xzJ/vH6bk
zoD0jCSYTNVG0qF4K779q+NTmFuAZ93JeKqayalkaCqYL8V3sE2cb5WUz9hZWQUP
uEetXuB74990RCywICzoZ0p1E4W807c0SI8w2bDxaBXWXKaWIBnDSDlWCgdepg2r
3FR9IdFwrk2PeL7wwQtYqilBgoM7+4dAFSADHZX+dTzZZImb1LuJHn8eqorphZvw
f+DfzaAVd23hjuyJMj7J5oujjxBAfqHKNTtMFKWQGJDZrr9YXeFwIarL9RRICLef
W1sRfOtPDZYJ0W4nGw3vojAya4c4KQb7UrHRHviQIqXRYT6hplnQHU0XPKJMWL/L
IQdz8VWf38HNS8dhKbwlEHIsA1GLHrvJxc/DMO4zQHUVmpoJVQDN3fKCdzVJNI1l
j6q+xaJmDjvmL+vOPnp4UfMpC+LJIj0JCoXm2bLlTV3jRaJVUvkJUX1g+JWvwhnM
7P0nqrUdyXvcyUEXTEape6jftTGOL2RdtLFLs9Ddstt+DBGRZYZqc9GYkLUojaHe
xVSM6XwgLYOtbc257FsMNtCfW6GA/momVMupcyF+QlogexyAJxw62ytOPVWOjWnI
GOV0xSSXpeD/I4oDtyHJ7HLEM62Z4sspPyD12jzVNobwfvSBiryH16Gv9sJ9j9T0
GiiNlLDgQkL937QuLSIWOPTzy9zUw3hP45l6LQ3p8sv7wrazWY+JC74uVBBK4atS
cabNVYBU+/bksUcTspJHLV9Y1MOj98WHhO+87DqvGfK7woFb728qZvyPxf/N205F
BNmTNgtElO+6I9gGyLsOUA2TpVRTrnnckseQagZ91M6o38oAo0q44pFUJoFN31U0
kEpYg1BsQwGfwoDNd8Tq2AmdLDv1WgKtWnlcsuEQXY+7rvVcytuEvIfCf7uLGojX
0ZrpAq00x/DjoamIAeVBAVuBcKc2lcnYtPIRsNS7u1dsU5e2frNRViegTfjJG1Uh
HiUjR47hiv12eEl1AU4O6vRYZiKb/oH2LxEn+YG/4ktoZAi6mROTDGw3ygQmgh05
oPe2hA9Lr2hBcPzWi/malpydORSqhZ+Zl2V43jd+gwuYxC0NbVFlWnEL5cySV1kn
EnpIRPiEjpk6sPbZLyUzS9+NxFfdcIb8yTcsAE6vpiHWEDT+f+Kbz8cRVc0EiRoR
lz8GQsT+yHusPnqDozV9PyDgaLdYDuw7EphtDbOTFeQONMdtWI6wypf0B08IaSha
5ci3LnsxDmmIbMOkoGA4JmBb6LgT4YvzLwd/f4O0XT7cyyUOeXUy2U3m37x4p1KV
7vJ/eAEPtVDjrpwHiNr+fNh0G5t+GL9D7moRonwLVwoHXZFfhnuyWtY7vpmq5jI8
1qj5SLpfk6XOZS5IljYopSWFbWKDwWoqFEjWYMtROg58HRIO7KaJbdH+XoJSQNqh
JErUsfpIFbKy1i810wmbMaU1LIwwsaxrmMZvThTJJcSX7gGNG7v/ZqOilLAgVvVY
OhTSJrJjf2VV7ErLRolEWr3Sq3c5nwqirigDGqgjOP23+iJ0SpqpCJEmJEGET69I
49bap7Hn6CeCEO5ZPm1wwFg9mIuPhUb9QMsE7bCHLequwK6tqhEQX2yc/Mc8etD/
RfnUJy8VyRDMjmZabybzJzVgciyAj/2IxKn/Vw77KhXtOZ1ZOnsZU2dFVa+lzCUU
9bAe4wnGUQWKZG6yYflrFk5YyllYxneaaZkJ83lXORvlhEUsmHlsS5H2GHye3qIX
0kY5YRgKWbwmFPRQP7seFBe64j6BsY8G6l7GpOlBc20nsISPOTvIAHYRVlSjEnQ2
E84mr6GVFWXPCZOR9qhdTdv1AVFSUUpvjrjN7k2HZt6jhJdVMp1mjNRy2NERy5aJ
Hfj63OaLYSIT+X+Y6MGhisP1mNx6TVGl2Xoz5fVhzBYp9XX4qmSFKOI0la8BCgz0
rZqWv3DtYX0KmKjwjQJxUl2SHWbGy9UsZfcHSDMprKpRbt2AmGgwX6y8yMMGL5WZ
POjyL6AS1HHBkvPAyAwY6JzAio57aDeY8ebJm5fIY7G+2BmBYstkH2i92IjlTuSK
x4IpgU2Qdx5dg7DffS25dZzKNHKUphtg5eGElyUjQW+bFCu6fVISwcuM3+x1vv7f
388fVO/PJw4p7rxy7+l4QPDKZOMdJVjqw2Qtd57ZBVMqVGWibEKZQXIttGp02Qzl
D5DXzfPK1vgiLglRn0FdZo+Czni8Gdm00miG/3G658EvxareTQu9As2h3VJ3+sww
MqRG2HrEue11e53rAnB+LW1LU0A+TyM0q16e5EJbarDGQx15YQvpoT9RclrKJ4lI
21dGasR5cqHlhmod4kIqwm4MUSk0eC0Kugq2fKx5G0c0fMgDmkuhnKePbdHcdvLZ
DVtx+1gEoMLY9fxb3hoELRf0Yn7kuEC7o/kK+AAJIjyIYTEtPi9889TGVB+FgAPx
BRTJq3Z3rNaHyzGCYAbaBxScYY7uwmVgagpfbA33fLXNbY00BPXcOOZYWGAabS6w
6a+8Sx6u7Ejj/rH+BDVd6CRPf23+6IbeIVW/5mg+tsWQwJzqquhsQCLo9bE63Lsr
dvZZRkd8SuUbQ4KlO3dRth3F/1pj9Hn1HcZRBTnf8Ncp+pYcqFbFMPnlGyzfFKKl
Pn1hajf5WiPGttaB+HuAXcxXY3LUkjCMw4l1AMa1mQP0lOnrFIbJ0G5SP8ggee3x
gwSuNrJKYzTNBr3Xtx7TKlO7bnZVsubjf8HHQNq7BkKK+zhgP8v/Ery4YmUYpbH4
eq+TWWOwB0LAS69EtC3cuwuhbykhFU72fVms7BjS0uonZL9jJ71UhcisSotQ2aoF
kTLbB1t+T/8P4qYNp18a32HNBpZE/19CgY+STzMapz6paQDC2GITElhOauPFI18b
16g+RWnE2MfOvMWq+bl2Rh4W8pVbOTKvSMB9mbTsbOCqxvnFaqzghij4CtJP1p0N
ey8X9sJVY+QRd+OPfTNfCafzuyyTt0n+v1fvq8tvCp24eCte4Gz61GZbkkaXw3gI
BMQjLznfK4vq8Uyppg94DUnpdBQbuSfJ+zOBMRVg/WblmoFb0Y1489Jh5u3zX/4w
LVYfuOzmc2XbjgLN13Rm1v4ty1O4wPIQZh6HI9tOu1FbM4eC750eXVF7Kh2RauSx
tughsBRn5x3zD9lYiGrQuU0YC1WN/MKylKTXwMlZqGYC1bgsVfjAZacKXdli2pR1
k07DoXn9sJLwH653DZr03Slmikl7k7LyIjgdC6DK1+GgghzdFLFvuIikuDLRh1He
IOxUBQ9If96mwxO4JWl+jRY1CzZDkkCWMebxy9yc2q7TRO0DRxCEKC+j5PwvubJf
vBQS3Yj5whkN/4gSzLaQzKLf+sdXI4sc49AdG2+ODHA8HJbhrKLWN/LNJ3wHLoam
nuji4z/h2Z03g/e37RNASgqI+5yadgyn2Ahu7VGmz8AQa2itMMwdnKiqKRCi+tlM
qBfIx6wpwMChYpLz/dJukO0rkmGi+S7Zb6BKSOPVu8RhbqFOQRHocIfOBi0PVY9k
Ko30UF1Kmt5FoylNoz2oy1uo60UGTqN7cqX7TnpBAJxYfEFxL8EHCbTAI5uwAnr4
vKq4vA6hKHsy28r8Zxb0d376lMTHVj+JlAWH870v1D4E5ak+Or+OLtzIkh+oaQqj
t2nSGDHagntLfCJwgd3BcaMyeb8u9C4kkMOWFYiSJF7uK0zj7lDCtg3m7SQIst/n
4080xqfKsx5ak1mbwjQRzX43zL/WDdH+hw9mbVzUnvHSv39dMZio1aEYTA8f+oW+
wwm5bROo9/rAyKK/9PXMX5uwi6/UClCfFJnDJS1mIk98nRUeUP+Rhdk4ihmIoWme
vS7gdnMGY0ccXks8uroc9njhTCjGSWrAMqGnsLEEJ+s6LLXpkdXNzLOJvdRGF02D
zo5haQoS+dMhTzV4V3/NdbAD1SxOqtY9+lM7FB7z6ckmDL6Z8tnJsNZUK/4R96w5
+q6POMo+PvEitTqYGsvlgXYyXSJrPWbXA2l4zkYKWWvdPlM9rbL3fF3ngKYI0ERP
T3jmEBYx12rDkfGqzbioeyXr3zKDEP5OFDvoU9mb1ISY69neSe8rvli4+iJBv4n0
cxR42VMwie/aRMrlwc0tRkiSlQ+m42Vq4wC8yJ22eZv0EF+Sp2kzYQODMsxIoh4w
OnZGPbuyxy9X8CLc1rNWrUBQcvBLSb9vYGU+6tFRATdDRryl2S0Czvvk4SoFl7P4
xtMj29Uk41GJtZq4HNz5T4LwALpYEPxgMGz8bvgrD+vws6DQIhVpeA0MPyWNgIRG
lD9DpqCh6mDGuIQ5/kmsFtSfakH1uBZiOQ4N+Pk6oSo/bxUHVJTFECh8uOupgYuU
6GNYppLloSEvy3A0Wc+fwPoyGCNWT4X7kU1GYzWkBsBxxIuZXJP0Hz0RACJK7oSN
fEK4nkcNSikHzZ1VfvDGmaLxgQJmo9rZbR7fGl2GXSDkAU7+oq4ln5t0YjASr693
m2SVWngIGsA3C4yziHxbEYUjqwHGcMNMLG+jfd80epWBGd8ONnupbWpr5xTY+Bvv
clXjMeYn5cxmDQ0Pp2CF8C+MNVp0KF9fees/cLjYpwtb6iDVdEFW7XBoLnl+2w8I
VonjE0Rrhg4d8BcLEHJx6Dwp/PSt3DYlF+zwEKy3IHO7SSFVVMalf12pbtEwBM4q
b3h2/Q+N1hQoenFqaZytjthwVQ/3baeBzs7BZJw9k8W8X9qsAKyo62upWBxbtVY2
kaPvlhFskcLmlHwh/tiQinYg0xPLhtyCimMDOailS5L5j3TiNPL28Jq8SEHELRmO
RgdyzHsCXOFlYxhS0Cf4BWF7n0yYha9ebOT6dcSH0L6E4NjtcXGXdFK32YSmmO6Y
LssgXWByRUw8q2azXJ7bZsHK4L173aCSP5RhKcQxR9d2kWBtW0HB4PJrU0xHZ3iv
kcyS95BGWQieCmt9sSql/LuIbU6CekYnlfkjg6UnfuoyV63NAoFgO0I9rR+SIdXO
y+iKJleNUYIr5oRYdzaA6fCg23kjaGyJf+tvF+hZBJzP7QW4Xj01dD3s6x9n9Swh
b0utLcmLObBnr0KvKshfnSY24LOgxsRLpYpsdjnGkoKzxxfamDQuwbJ/Dm50LDJ5
XbsrilYCHEoyCQZFP7T78ImzpFplC7LgveXHkmGr5lC9r8WORnC40HoJB2szc6ka
JfXkZwt5S9otBu0wLgzL0iewDuuGi93yAiPXGW4t1HRJfVnmuJ9MlJecNygTGDYa
4g60WjVC5xoqCPODOsBAHkM4L5WlVm9Ovty9d9vHHGkpc1r/TbIBKmssHNx65iZi
zWTnhCSC4ekvsj2mHpy3SmJ2Yy5/TdxXs/BXJHTpxFL/Ark8lKAOwILpybQvRuhj
JjW073zojYBO3zENElNHu3TdTdj4wCp6mHL5WUq/M8T2qQiEmkQelPnHxWQv8j+X
f6e0dBuh0O2l9lU/julXLilWBz+BB3v+leU8ijXSgMIupzdoywM9tcsn1SYbNwwy
9lIBtEoTDeMzutPLlKvetoXUIbu+BS8TlNa0Z/dflmKyHUWhzrsy12eL/z+PRA6s
oS9Kzc/SeG87nYnZD55SYsM60XVpU5PMy6EXXeAuTqOl88boMLx1euagy5hf6pBP
FsI5mbKhD0VMCxhX5Fz04XzKwsGRuaIGtDqRDUp0iIWLsIJ7ItDo7+G5igiJ5kYw
pmJDq4UuKADMn7qMMTY90d1Jmq/DK364eqOXsGXQREcZetphUkgsuKWx2muKmKnu
QOsWd8B1HUaEhxpqa0l0J6uxJ5/kStf8krIiLG6NlJBax6aDMQkoEVHaEz4mk2ih
/OBagafkGksnPov7TLurKMmufAf1+Mw2m85WfxBAXsMPrm6YsyL7f4u+U0MkHqYR
yyjI1GhYwSzX2zU0ugVXV3g6pKw4ClIPoQBoGPAk9nPQYkq0ZHvECfaSSbxJkjAS
0xO2MTuWc2KEaBbyPyvJEIDlEHxfEYby4r1gYlLAc6La/wYEA6AUS8MyVYaWzB3X
bS9WAhCrL5IE8MkRyP4/cPmS6/aYM/fwL+emER2SY6TiJCh1meR7tkzzp36XNUdR
hJGqw1dAIRUnBJ/27Jvqelu9dO18UQ3rmxjV4s0vQaYxchDizYQn+EDuE/FJhVuF
5Hmbvq70XPNWY1OJ/vtwsVmqxKtILfwlEL+nNvWx5Vm4OxFHkl1538Rc9MXietux
/GzKRzeIdKuI5+jRecmIdClhP6B0UNDALE6y26l7XVrwIJbV8NUMTDxW3J3S+58e
AWNWylJw7AYv+OxbTQ9NQwNhiA2VQPr5BT3yY+LQVqtAMc+WUq42qP7PfXkWCS4t
jK+QPZEuw3+TqsL686db5kUN7iOMey3tWZfVqW0oOfsq/VYW4QnX6fj5zD6yqwrl
tBu1n+boPNarfa3cXAExd3orP2o5qvijZANVk2mj2tNRfjbHO+xnVt5eJtfjCdfF
w3/9RISNwo9qfYG1atdWfaUPJHrKUPpCUwVnGqIK0jGQIgtJLU1YpOI1Jq6N8t3d
iiximHL64+pndNYgjS35bOXesyPt68DeX3CPTGtjWXIdGif+Q1lFf4SQXT7P/hyf
rGSKXCE0h84yZMcAuat/npShJQ2knOZij9/TYo3HIlrROo2wm+onV8VeEYw41rc4
AymoRUoIYRBWBpPVZZQPAWYkdBbViwqOPg8a7MfvsnM6DlFl9/pAEl8dZ8JTQAJ9
EApKaIEfdCHH3n4W7MlhmNnSQyFXHgaOA1/DxWK5AWXraZPD/sehF9tpa/Vw7NAh
Yd6PKhDfgJtbXWawop3z29R9VcDVSt0i/IGofAq8E5JmEqc9XxxljkiOernZ7mOd
9gdYheRmH99tRT4UpAvyX/NMmysHSHQn9OynI8MoXeVzq70PkWPgp9XtZTFsb7r2
rAY/YGUYs3etyrcbW2RpRrgt6aaRTOak/xH9anrTaUUwBkQnd8XwFhS/qQ8dymFE
YyvbQYBMbdMEyB4hUCt6pFKE4nm8FuoZv4uqdULVEoRykfYDdXeGM+PwCg38NLxr
pYxIwdCUdImW/OqGRHeQwTw0iKkSOgc8wSluW+Qady6p/YZa/Cbwq330lQJLkYVA
5XAKKo9PtfH+o0khv1zee8Lhn3rbH6qOJ7DRFTiBJqyYJKXVu95xp3ERxrFyRTVI
t2L2LF1WLGNH12/R64pzxWEqaVSb+P2nCNErz11AeRt67y4tRv4DLCm11iraN7Fk
L5aDCQAjhxuHNH5urLWhBIykaGGkp/x618qPPMzm5f9hsdEGY7Oww9nf2++0hfNn
mw531I6geA9TFFgbYZr4gKeenOBA/FczG5ef0Nb8Y4E7IUwSQFEWiq/QQzODlQ1Q
D2P22EmKLEh2AgebrlMXQ16J8T2JwZxV9bU2OiZPcg6d9Rexq44pGh/GSO0Tkb4o
UpshlI1bbT76Sk2cgXR2y+ny63YxWYUjW1G8tN7dvqI221UPOUQ4OxJf0S40t0BU
ZNAExVnYpmuvLHisVYfi+qpJQSFDPGIh1sZc726LTevz4FvUZTl18kKBhTa8TFSw
CK1uRYX8t1lwPKKxHZBE2dNhGsbVBb+bARYX1n45QJ/iMPzmJXnZb1WJmzkaqb2G
sS5OdwqMZ60locLsqNcSLtfSyG2IOOAROZiOt2/GAvtwdIS/G42aesMAgOUqzLS9
uCFMPG5JvuRrvp9jqU7JPUXDaPLmrpYrbS0caBduCRg8BIMEfTu63AQ6t6dqX6l0
N0HxXaGFEI/W7KNbqp1dpWqWtreFxa8meocW+IeKUjNf6tz0F/q2JGrfprJLKb9d
Pzfoc6AiVxoCBXtc8AdU7DXcN1MMXRog6KDwhCJCElJR+euaaj4AIkV2VyuPNU4r
acX1N5g6hV3/CgW+zOz5sN1NJ57ZlvJpc4AnKsIn2L8+3tPvgjTna+fzogl3g9s5
jaXLvIrAoB+lUB19bltgWMLWEwiz4pl6u1aI49dggMClLNnYQSFmSQekwCZfFzZF
qF4Zu6oVf/y7FbztLQayxJ9iEbMs43MRuEyLWLg2fvIa0dGx1vPcEECqmgHU3/9R
qlYZsmmax/5plVk6CjvTxOS3rRcmn9T4Z1k9bmSN0eHIRjk69IgS3Ec9Cq04lpzf
xYJtQLHPAMSPoTp58aW2oxXUQ/liWH+9DDwByAHNS/zU1VOcgDmOpCJp8SYWd09W
7rILCcIOzadP82GTur58+ufaxdjZfpOsIpYTs3yyN4lkoBYP1Vs/uisrbhrFNEJu
9odOBhXQkWe5YBa6eWfP3jZaOAZpM7tbcy/EA0MqjXYDT05YPvK0YruoaDySZTsi
pcdQznsQhFAfKs/QpHAaZn25om6I/CmNRzpicPK5M+6aUsXmK/SuwsxwrsnCFAld
FPHl5cI6WRJTLu5tJV4gW3ZwTLZHnNY+m2/fczYY2jY/aSlm46iopVZabUPaDhI+
EMaUiE71lIebIwJlAxl73XZzp/AJ07vayGfxTfT+oC6YjJpF9V9zjLhutu4MQTh8
P7i5EsQ65SkPkSh1lhBV9twhSdBTtuAyfYyW7HuFG8RSuFhON/Set/T886vI0Fl5
pfo9MAjowUnYtkpJpUHFR8F7rQ1LJ+hJlJ78LNVzW38/Qi6vz7wrKaLf/ganlVhZ
eCKp/bxTYyXh+YmnZy9bSTXPm6WEE73XA6bX+K90bZM57Nfq1zjNq45pf0yPHu8e
4TPU/bulv9rJ+4XstTxN50P/JiHi0ZXmgjZXKA5pI9zYEbiXdemXN6c6qPcURrwz
lD/JoW4voyQBp+zKDo6hwHqaGJSgG4NL+pdLELv4ATr6Ow0U/T1pDSm/LnV3Wi9K
DZIBjeBXQlklCzg+Bsf6a4TQ5i/alfw+DxcABnC0eQWUiVEph46SGomcgoUbZjtl
/g0weoA9XwWBn8R9XUTKUGjjBVzDkp3sUhttlM+gTc91ziuVkjV2FiLishvDVRqw
3d7YxHqMj+Qo3GGfzwfOh7RA7XgWS8nNbTbh23D8UiMQQQqf80BhQihv6blv3JXd
WhWeIex4vQqk7fvxYFESy7M61aGPZFZpw/sfLJjm/F0=
`protect END_PROTECTED
