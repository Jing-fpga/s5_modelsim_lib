`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6GylbVvfNx3jUyqxBRl2xc3gx0QnWC564oi/hacXiFrGfoBHI09G1b1fMego5edu
YfMRmw033juZSKAWSWeIJK6riHxNH0qVje4C6MzjkJIX851UcEUHHJ1bu2moggkf
gfhqcXlcT1pRSA7WFQUd4SegEsUYxSYDG6erQ+meb9iqepHvWwz3oGkLWdPcVJXi
g9X1SI23yQuuxk2goHh4P6N/zsmHG6KeRyN+7DJQq+LHBoddxgRi1KoNNdH0HSNa
IfEN5Yop/Y6H0dPI5Mr83C+PyndPRqV9BZHJJafx7xp5Br9p9/TGkyq67tXG2fmJ
y/8UZFTqrF3FnLz6UzcUdJWaQOiWFaGj9NoHMzBwc1y1YOWugr2bBpxNsHn7Tzc/
/K5zafFwRAeM1ehHL2b3NojvkCXlR95tlYT/UcPHMz7NeYFsJkvGwAFKNsctIqtY
B6U1jkmX9IJsIkYqosK5EqcYVqz8NsBiQpblA9UPN0KebG9cFOG1fL9fQ1oTNgIt
TCTQZ3pKS9F3HP9BPu3FxxynNyNq5CcCxIP4/NDuF8g5ADaOapZifq23M71+QHCX
RE3eioHDKrhDsfGsSIev5ZvffA8hZoYpxY71duOOiRZcAH1T9ioX5O6b0aMkcYrd
G6HsT2EYcN+s6xtBLWfm8zltmLyJq3Qu9YOZXFx8ZfAqTHNa73vr7FGayr+tr99n
kkpoiBwJ/qYvOjcCDuZfu0Hx4LQL21/p1w+UwHCxePKZiWuRnxA9XBE0Diwtn418
z2pt4vqoXWZteYUrSrrHyaMWSO3VM0YrTG8gCoZgxrMPhn8anQWARDQyi3dEFq1b
n/bCkuq2pCjXyNTb1KROXpWWwO6FfOwD00+6+NdDPm0X1lzmE9rVbMjTETdgFy2b
1fwm67JHrrdr9m2CxVi79Eilz+vZ5b5Rx9mpDkHheinjUNTqXH6tl9IJ2Pr+JzG8
uiXEaHU588uw8WW6lzYaAxaWoX3ll0xGxDCMHR9KPil7z+eQqfBWlGmqTXXxU/Co
2wHJWNFfTCAZzqiG1ShRdIy3sMMVKV8siVRW/QBp3cm0CQx2Jx2Y4bb/GaUmKrZn
jV0PPVYYSTzKgFJmfg1C1tZoCcK84V6R1zfZu2k0eTRcMKknF36rCemFN4BmRer3
SZZbcImo/Vd2XbHyEK+bQne/4UvR579B+8rrI67sblVILb+fpI/NbFjxx6fbYR5N
a6w7/oMws1o7DhvBNUgiA2e4CrsF0shGbcVjnO930bKpj9N8zFinH+jmXeqPBbEm
o+SckDz150igtJ6eIsK/2rcQA3d/lyHA7e8xUvp6iCNoryrdtGnC2h4lIbtBqPwu
I9nFYvCG36xLd8BB6werff2hRoTbdSpwy66s616a7UAZ9JxcaVtWRpvXA0ZRc0ZH
NEc+R9VyfVqLvogzhng+iKLUs2ZWjdObAc5/C9B76IAFSbetWcR5vlNKg3VoYU95
Bp1k6ihN8HiDimUUafUg9EZd0PlSMOXnnScrplr7nVe6xxyyJO6dsL8cwntxVugu
ToCL6ViuzX4LPrvCKVSD5hF5yf6TMpQY3lWVrpFMPO2nRMnuXKl63l6FykxmlPe8
fXfXsPjtl4DaaL6/kBYpAqwAMlIsyJ2BIdcGfoc0l5UTh2UKcA5c3ZDeO1ILQJ2i
np5/cgRCD+GaoqmCz53nxDpSrpQhFoaF8Op4npK/TXQD2m5RuvcXYPNJshbWJY+X
5wSKGX9qf2NrBqKE9/taZgvD23EZDFnavNUbM6rschgtZ7ZAe/OByUAhP1xSUI5V
o/1WkK/eYruamjpPSLRlQD931CNi73xnAL9sSgtsd6VtHfeSNHoCXGf/bFuRpoDS
fwpfed+UWoLjstTovBqN9U3wnAaQZSNZiqGWjbqSAAeeyNCMeuD7RcROFTK03FHj
d/IrKrDXWSfrFg0e49Nyf0q9gf3B5hURcylrEdfPBCUSt8rQIPp0duWbpuKMbM5W
GuRKERRSBzMVHmW+BXWAF97oPg0XLTyPFCWfdYNbVHMJCJxDQTBevQSa3TcLWMnP
CmhPVxdYLsb4dTS3dZOixGd+vEhsLDkvh9uWWpcOoqfJKDs5P1CK6EmzvoGZjQhL
CqK/lopUpL6EpfeAGmJBRx0V0cM0TWszHmhkKb51Ggagsvk4XwTb7oJxGakOnBTc
tKzf6ju7bl/tuldoC7hEP0wTC9u4qd5YOdPe3O8pXwFRptPkrcR3LmS8Embbc3TQ
1dj3t78SylY96At9JITu4ApkoplbAsORMjRbAkhXLQgJF1v8YYnk7FeuY1JXu1e3
d0XVfAZ96+w2Y68nhh3iFqrBKTgda6Hfy2jknBEsST6n9u2Qe3B8mJlosGvZMb1j
uJogfz4WvxkZC/GerWvINZTKH6pQdbDl+qQUdPP39eXlCaFZmZIAIDEOGP6wziUg
w/n/YDWmy4wvnQXt49c6rKxb34SduvxPwMdXPQ8FpdLCgKXFuDUCubqhWtsU3d8U
KUVP6EZd21wyQmzxdeERYjJaEUWvJv/6sbbv4KGxCPAKtGFNO+buIZAsmUtKJrhj
eaC/4tgAoaOggla1lv5oS+pY8mEm/J1HZO05Mfg/GqNm6hTh0jNu8mlkknUpaIPM
ffd2507S+SzvTuYUg2R2AsnONuQmsEe9DI4PW8nVKWWI1pV7tJ38lYVYnZzB2g/s
Q+6B9NFzuYIJH/gaKb2xh/oQ3M+LO2+aIGLL61zPEsg62kyc+FueRNMf63RkZP0G
RdU1AEkLI7GQz2tY/4QvbxVgatuVpzN2hScvP/W/AhH4S0IMLhsEczaOmig4FP+q
5dFFdKVt33REo2tv69ZsHP3chjEIFQ9cB3oEe2Llj+pTCehbDK0qNlOTn5dEHnbA
1KiBaHPRUKYVFherKrGO4wtQwcHq4LaufNEs6ZNSvPNpLG5U5NZd5gk1eHtoUhBD
fARE2OqLVY1VKaZcHJNgjV7kXjgHXfyrGzcdGVbiyuU+yJOoJ1ZtRcSYNespuE+z
sY0tw+etWEsVLsWw9J8ft8BdqB+xiR3AwgFaEGjD9a1uYgiKA4oxdqnUswThpBC6
Z66v4/vJA0vNOVc/WEaU0ELofIZdg1M1oJXJeoSueBHDVZru+pNrqug7asna80tf
ZYGZJSbGzaNambLlQMObQztCiGRzRGKlaIBDvE8odFCI47hOWWK8mPz1LmFsHcLE
S7pI8CGUnyzqZ8/0L2q32w4/cypwaM1b2Hx7PCq2bXFFId77fLT3/rVmksyE9mkc
o84UcIjEyi5G9qeehklRc9+WJuT0im/84OfqB2kih7vP6kDvGkZMYdiAj0DeN6ld
1DUYbzCklw/nKqCMNfSAYbxExFlu/sydCS6yuomzm3/lS9FzOQlv6cd00+Moqj3D
jS8hQyXMcbd8LUqfhsXMU7Gw7KdkqR1OgLYx6M+a5a/oxHMo/jmL5sJGRXgYUijA
+6fiy82TzeAKi61wRBxIaigW89UbsWQDLMsI3IatxmvB6QyPXL442F8hMbmYTG/H
+C6IdipiW2Jp6bqCuonl1cWS4OlMBgsh53gqwbSvWXQf/e8kQW0TG4oeED6hQZ6G
LOEGqgOlUuz6Ye7fqbjYejhemC1oG4QaaIe1AeTJERP5S7z7ugBgJa2rhGyUCJQW
x8AHLxZeLVAcx4+pHzBX/oZN6e/vpANVboEtMFfAPVNsJkawK0/zcmJ65KUrlynx
/wDTU93kNF5ufUv6JcBy2a0sjp9p07aPITAep7u1JjSsULwJsQlk8PFe0+c21xZR
BjtpsWLfLnZJTMeY5cLSU46ECULwO3+0iS8UDpHSAx9L4HzsCLdYtVCaUxEyjUA6
t4n7/CIJbovqvU5ZhV8MfA==
`protect END_PROTECTED
