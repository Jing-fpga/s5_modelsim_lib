`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gOVh1bu7j8uJE7KRBA0aZ48iqyGqfver1jQhyMkf5M4vIUQwd9lx/8j6gwk5wJha
qKx2D+69O3tHJfdqHcsXXWce4OggcoPVL/HtBRjlI5fM5IYmBn6miv08fdpCUfwB
CiWgEF75FRq/xDDbXPiZwY/5DxTdZdXv9F1dr+XCsHP6y47YXm8pVjzUnihP0mRV
OaLNnldL2G+n/CFKmPmr8jOXtLp48xsNNiYMq4Ha9i1AKTLe99sz5npndX2cKt4G
GQvfhI0N69UmxK8t0Gj5tdzTjlaPYkEQRa53hg98COa43gAXcYhArVSwHGGNFm8h
4VX0d0XDje1aAZhw8MaARM5srU45LVT78HW37XSH47gs2QFC5nHPA/DVxsAPAjKM
fb3YnOy8yoc4hYRAU9MPQgbYo8Vf4c601VoEa8LBheYl3EtGHuQNY6wOYe2SVtTi
4aEKepqBriHy2p2hmhUC97/pp7J89SYH1d2iTPAhS9XCEzYlOeweKmNtOkfX+Zh7
w6wRTyPgexSgqRfe342QJaJX01Mqs2aU1GLvDFgpwmWqXZinkjAQrgFrb5GI0XZh
5cpVCj0KQBwGFYLbAgXrCUGmcQvkPY5jEcnxV+Z71EZqOUR0tPzjc/3r9YJiIQ2I
rzn5+7rMCgYIEGC40yfqwdphyrP11ngziSt14X+s17UAP/NjjrWzeyUNHvP+W/NF
N81nCHfMEMAIScdJRa4hipMkPUq2nhyF0u3xHyxww2DHg4TnImKctvwtEmo2BzoC
KwPk5noh6Yq/tPNsOfe0NkBpEx1xunXv7r7YyswaIaOACMlLL0cABPdY4KnWB5VU
WmcEpy+P8MzT28WtCOuSGY/tjVNCRxwGnpPtHB6iWXgrU4MdgHR/abgrXD4N1W7l
f6wuj3QlfFdCxptSN6hnFYRUX88Ekq27GQVptiZHjAJ137OVVOg99n/VyrYjd7h/
7Y0hSsZMxqQS2zY3FbRwZKoux1dIbCT/U770EZ0kTJIT9zQlfnYvaao1ITw77fEE
TaQYjzIoZGoBXZVi4T+VKyhH8DOUHmtZ9h6dPErSdfzBIJvrX3E5RjDUBn0xXqVG
/KE0c0c/P3NXBn1TMqByUGHO0xHq4qZXs5PwelNNzjLQ71+nXumqMjZyIrpAaXfY
534NzeyzHm++kSYnagf7pSi/imZlhnjTX+A2zO9jSLxTuBYdr1GFKYVRTQoV/Fsz
gchIi9dPlkzcyTSnzFkyvDR0YKjrcMKuAf6upYm8/Y/x9NRZJHr73pI37wBzbYcZ
hH6XCrzDGKreOfSes0s0+sXroAi8BrlOfAIybk16d+kn0Vq0oIjsT2Ra8Kb1/yIv
XsF+pAQIZuGH1AVddOZ7oWyqzHPXTIaJa8viq8iUOmIX3/nKsgOEGqvhNJWwjroA
++ugCuEFE5l+0nIKwHju0E4b47T8v+Rxpctgy4C5hGjdTr47jqdGnMfiGzWBbIQm
b43eb8CrhK4e6rmmJHWgoH9JHTJD3hyXHAo0e2o+itLCYa6rYy8ksRENjIRfjbvP
fBH1p8bztOMyfO19e4SJgWIDe01FIobKUAiYESBv17KXO618egGbiQs0YQpghBOy
eCcdiLlBDB9Q6biqqf2uofa8qcBGeTDRmpxXMCasW0PuhzyBbaVZ9P1P9uPRVq66
EM2EeNxFQ/CBtu/TLjuzm9wpmdqh7WyrbMsEFCxAnxtkj35pFv1tIVbtr5cY7H3Y
LV3p9Tvy0C1ATIdupbE5CJOBKq4RcGW24fhWnO9D6BDKK0ZAbktfAmTEEAdZia80
lkupobFVTvddUOoTv74wASpLtwuo0XcA0I8vbJ+A1GdQbqMBY2YLfNar4A8PyE65
30meYl9BC4lHAwzBuOdTPG6bEL0mnqVbbYAj5jvJGcn/uh2ZsrWyoVlu9F3CGnSC
c21TBRTMI5xVnIhhPYfypSQxW3h5bOM22Hm2VlnFoPf43gEUs3ufnqBfDehK6E+9
9p4jZ/G8Plxv00x15Oe8sAcRwCBIWP0ommfgxKz1W8rRZeBKfD4ubYOYQhSkcbl9
h34waxA1ftDn9fVgIvJH3UUn/KAMLUM5Oi78RABX0JyUzQgln+hYCyHjjVYBmoam
ZKakA/tccywP171MqhHB4x9p6lHSmDa+FbhMv7qZRVQayozxIZIqmR7xXYUhvrkE
f6Tsiw0nektggPg6esK32bDqLWYg6ZVXSCuVyYa3qASGYadQOQHmvgoCiHxBC7kX
ldAkJii7PpnmRI24/BcTYppUwIi9FehpkDq8w6CriW/PdJPF9o+1AMCx+WWsaUaN
78TSxp4wN8eS/K676qn3xAen04nfR0A8Pv+kjr3J2vow2ZCnUjChbJJ/qLGjP9N/
po2VW7836nrjeD8XqVRtxI1a6j+fVPMJRjsgp5fHb4YaX1JK7d8vnSD/JzGq5p9T
oYYYa8V60B3PNkEUGc3/rmwuALxTdHuKGQbeEDRsadhhsL8SOGA5emXKXRm5kikW
ANpEBRV5GQQJq8glLgSUPKiBlagWV1RP4lNOQB/zW/YlKv36VENTXs//1LB+n6sj
vfZarD1i/6zkz3gvd6HmuwLC2C2vi/wryf8NlfgI+tegxZ8OvCxAC85AzMdkvKm8
acNS6KkKUZPCP1yvorPB0+QG6CYOjmNeiYl0jM3ynvSzKOZo7aYxPn3h65q5Sv3X
lVU+ywljD3+tXMo0f7NuUxJSSTc6g1M/TIzRv2ZppYMaLh0zKriDK/9wfFLwz2UO
1EMqUXaVLEcLa26mIC6A11sPgulhZrrpWy72jBD+cDMnB+2xPkq/xEqPCdX4r3cn
VO6AbUxvzsqYohbnr9FVID1vTAR1CdVfzgdQX1F0+ldoGFpWO8bCpoKPrftrpopT
dwWP9MrwE6qmAh6O5rQsA24LzLOHeFlkD0uMJ1c2CqZ9jGofy8RU/4c3NZGAYqh8
AdK0uC68Kp+fr46qtCb235nsObgM11oFbmBocRVb/1v/73/6OrAasCi9KCCQwlPP
vs4uD4vy1I5an+iZlmKZvleMN9AY98Hkt+l97q9Yai6/uxCEw6oF3yc9/GLrHvW3
bW7PW0IcRZKhKwU9edXs3cQcy7/vM+K5UUO40lFWgJjJnrjQWt9moI5jNnQOXIOF
bo60wH7Ak72GNL1zlYf9OdbV6B/pIcgeThlX+0JGSABqnbRX9rV8EtHa6sdeNWRM
2o02fLXEpylbAPlySF3Z4Nx20lVSJngYtWc8Gt3sIsYmUop8MujJJEVjzVOzTTrb
0GEHzljO153eQmdV1ZdCr+V+rHwGfBFxeZTIzkrBYS7bt29eR+5Qz50sL6efS8DD
LDkfIJTFN0lARRvHcp8SVKJtvgvRTrD0ZZChWVP6F0i4j3MfkWE3Vd63DETUpZ9v
6cOZOzCDIehT0JcQ3IsvthXJzI27dUBIAKl7j7VEV7+qStlmMZl5LdkO44KwLYrl
PhhuaM5pYf0ZdhdeUHNArCfQv4nJYxh8aoYCb0ay0iHoehqJLq4z2LJUICA013Oi
vYBQBGVxM85Ofz1weSbPhWDe8jMmzdpxRqsIpLxO3jeVVbmz0gF1ok7kiW36k8qD
78e5utR3pSPKH3dPlR1gdCdwznszICu26KO9q39mWWfMOa9pOP9Wha4FXwy3RHVQ
Bp+HAWEnygmmAmpMLIrtTKCnb5TWh75dgoDmV2HbRCFYxwzOC4caS4F/LQmApx0k
t0KSLR8+SxJgvIJtk1rGq7iAcv6xtYM+NwqWvECjScCbhHm6JPeYjSkXu+6lfEbC
MlpdLPHdEWHpzyclIcdWrFx4x43cON6B0is7svIwXYJYtdkHbUamWpmTKNYvZ9J0
0Z627aJRk0s8TTfqecCmaFZXJ3pjAEB70joALm4VZW2a2wlA9vBaHhwwKFH16ab5
IkcYOHLBFobYTxWAZl9nj+McBOffJzNkIhWKIdsy6VKhz8lN1jpBhd3FLj4Giltj
iEhq0zO7Um3znDGrRlSH1qQfj5mn+E/Fgkoj4Ok6fRzCSGKAB3VuNhvCyK4/ftYC
BPZYfLUyUfcJQyo7jpiPSqYQRKoJaWjaFqNsenOvUYjzCGskLpf0sHVXz618nCU1
Jl+7WI6Si4E5brQtLALgi7HoNVgoYwI+V18CvnhlDvr8p1Pk3LcOz/lOsa1CwFJt
aADAiSCdY2SQEre9CJKyXzsJWSfpXZLjDngkkndwIi7zWfVhXEcib5x5M1tLFAMI
L37mRiohiJ8iNt9jNbNdIJtFMyNpbh9blws674rOzWmSm+AZpXbZPOx9+rRU1MqL
joTsfDl2G2jSB+k3we/YpDiSvZhYgmgUBTtUyqQH1B8rrBvuF3SE6+dqMVakg2ad
/8RMfr6iggwevctw2bQbYar4Tes5TH8Bk3jCEDXvslrp/oS1mDohaL4ue81YqE+I
BH1tsFmRu5rV44xg/tNiUu2iR/ngp8qNYAA361Gm/kZBqTgObfKywK014q1PZMYb
BbRA66ysCwzC7oMeWkeObWIpbMAa6ZWH10UnsgujnVUwYtuaEgoM6ThFToOk3HgJ
M3OmpWyLOtt2/kfOBrZAYAhTumktXxYwuI0ACYCC/4yHYAhC8tJk04eSk/KhwuiE
3/mmwCmbQT1U6YXkhho3IHGuwmJ4Sds4aUFpRqwArAPMg02Hm+chD817YDLbCkyi
96LTByRHWoAB1QuBsT7jqsihdh9r3bmlsolVPIWXVWpF5RfUrRPzS6WYhoBdyDmF
7kHFmlb21iI7nET3wCX/QPDkei7DolAp+oukm8UftllHRtA+Rkr9Rh7Tkza2jKPh
7mzXcLGIqjdeE6/Gusc970eNKwUEy70+E9eJuHDH4uQbZwQKBj1sOEhLFT/fGTQc
oSBPOeyxV69Rz4Glcvpc/3ozfNBjaIqypkiQlhbyf2SIHE2K9kv3hvM//ntRLSE+
BEHgW7iq4KMOwjSjXdV38eGl/culmIiUaBtysqGzlYj7JSYrIXFjPai5DPkqlAQW
jfRK6PpE6YFsGEjCDtBGIEJi31+7qhdscWzw8Na+7pH1707GQZf27i1j1OmU4BDR
P7x2VGROhal19L4sXGdLtozXMuwOhbWcM4PXcYLPK0NUCg5wf2Wg5TWPjlrhsLNq
1fqv/yOVMy0vaR7Ig4vcCLdTfUkAXBKSPApxHs4U3g5YcJ/SjuDyow1rdz6N/sPB
TgB03m8ddziqY2zufDI3w6jgSKamsMW/kwD7joua2ZgLNIDgPB8BR+9ImeWskjC7
Q43myWEotcJeNmSAKedXtfyrnZBiBaz8F9aMpZ5yCpaHPoqRDcUv3yKE8Hx0LfM2
pRJ/xMlEKySaAH6Iq/zM1EkUO6VlATQuq2vKl9lgKFFSt7Zs/HpAk/SwBfHEzWpR
6MO56E/it1z6p30nNYIzqrp9h3Rh/dpzZ/QWn79un0mY+DHnbFxW+54yaQmI3iM1
aUcCaO3KBRWaY9JJQz4mXXKXx/JZrJ/8MCJHJ56k9ULp85skSOSFugQ4/VMYX6zL
Fb52BnzspPUn4an8Q4dVzeWwtV2CpXLPJyks+xGvzyGv/VQDfayn3EOpWZZffR9w
mz6ryDfDOwCDvY9Iud75FDOGmMg5Of+H4jHrj/zdKt0msVcNZLRRuQyxYETNDplt
VqKutrtKTAu/NGzIXH9F1vV/obikRFEV2kt8+MHI1u0Z8Tw+S2XFARCdvwpc6zei
zHPLZkfdu+nEYf9WpE1zgfCa8z/+GmR4sr2B4zklYno3qvhtxQCBrMwsfU0Ui2Nk
WMQYJM5wvhNNmUFsYPW81dfj86WU40eqzUo1K6V3tlsy3nr7aPioMG9s8GQjgMw3
lQgpAnbNvNFn9Oty5rWDNc8D470N34Oly+svpQlOvrBi8ToEBkm5AWmrQqjruqJt
UpoCFXCtBT0htqWPMhOtAFy5Lkxy7j+fIREIwlqZTt3H1mUBmqg27ugQfVUqCO2Q
uyKrxgvYvUNby9Mb92KRY8zo4qHdurbXOlJO8FPVKnRG89VpmAHDP0K83cjOWnNL
x57zr1RcZxSmGMTkAfu3m+SjBdWZSN0vQEXHALwj27jWaX1EYqUOnIkH5cQfc5Il
D1cMxnTO2yZsoexWV5XCE3663hu5YVKRUlFQSSXaOJaj7nXHtliBk4TlSRgsKBpV
9MphlgTR9T6W99unCwP7quctseQ83RuHX0aTsv5QMolf1L+sBSkONcqto/rCDQ2E
PirmTQ9mG8LJYJpTXgf2LQ2ImVjhi5JZaHa/ecJoqVkyrimMuh4EOx9G/MtiFl2f
7YcCNCbzlbAaChwr1/0PL7eZC7CT/Kxnfhak0LfryVPqXRCjoypUnzO1Z9Cp6NoK
XRou7RpEL3bIodsIPZ3FO5d3+DitAtuots0/hqRm62R7cO37INwtSmey9ohAxQnl
pzVVU8FufTfyqjVBrEgUIMOvPX8MfGnK1sC7O27xQaFEVjHVm2FQU7SQZ/T2oPDY
n/iDKXNstp7brS8a4jgn2iNSK1JoSaioKRHRMBO4r48DVPVXDWGqLb90brHNQKru
6b9Ui9HellZLwmgSm74DoJXH2eqM24REeZy2P3sO7m3vKc+ha/mujwRSaGo3Pc8i
zfI+J62dPyrMxuv5KOoAP6tQC+56dnzUdT92vW8amwX2o0GvlKQCLSM9j4lDXN4w
0OTMK9805J1MrD73HIk/ALieUtoiYujSlwA6kx7eiq+mZHsNXGlOspYa59ymiiCw
LrFk4SgjjfPCeUV7wBID/DgGGNdaI/CZsGkN5VQgDx9WqidH7KyQpTOx/BJtIMF2
D1x80Aj2l5WHQla0b4t9zeSp+0cMsI7zZnG8ayyYJ3BAkCczAs9UNxZBXHlgCeSy
4sSxmhvOWVl0bk9NKRs2VsOn7q8Ex37Czw0LbtSePCm/C7dZvhaUcWaKhzYmnhXv
abTyS+Xc+8Eo7H2uK0fl/9uyvzI7nPbTbzeMITD2+L0OSnU+leKOdKbykbGlK2/z
t5u94PHtBtjmk7doGRgOcrzDZpDHoMrUo57+b11r7OIKQh1CTcpCg5JryIKw6kWE
lQsK43zvEAjEOXs99iNnN2cAuBtaaVUOPS0mFqsfmOfRven/EfRRzR20FlH7Gh15
pSGV+WYbgovJRdQcGqpIc1bO/HcLaiDVHCIZKUCQogH7mbdcQkxHR2EzIY1Q4zdY
t1ZHSHVppuxVSp65ugfoms7edUQQiGRo325pLy58PKHnBHTWARTw/VagypiPaq3B
hvCV0/Xr9pih5LjLnQPtRdlI8k/pVfJ8FTRSG944rKkdPhIAwW7RPLRy+fJvLApe
vAUiALCtrpZK5MsEKcUUtbMKbwycT1gykqR+If6TJ/AVfFeZCYeOJ9QUM+ubOWjV
uA3mSJAg8XTsKh2ya66wWDbUiQAR+QBEWW71TRhM5X2dV5QPEPxSlC1wk7Dbhlb1
9J3XAxw96ftH0aMdLdLxHQqQV0ovllYEwPgiI6JPov+xM+U9xa9y83k86M94AkB8
he0WcgDaOb+6zvw1cELhMaJBus/d/Mq74wYrJxqI8Xhddt6baav8h3z62QfSH+UU
nzdjiLdeZ+fVwZ6neqmdu9jNUvlvZz02nFSFvnXOQ8GNo9ZpFb9jJCURBMCof8Ce
3oBk3Pb8yyDw3IYW3erOjRR0bpQEEy174GS+PgtqPl+Bt0D99bfUBWDiCQdZlHzd
w7gmf5mSyiXYwMTHkNIbh8jIkZQRM730Lkkkp829p3zcb7KXEDUhRar26YT4D62Z
opf7W927j+326Tg/7qzkKqclZGvIt7SY3o5g86EW5BNbcnxH5HOdcqYDM3tTc4L3
+xvxZWxFPdq2/D0/oZ7Zq06OYcgo2nKHY/D+hJNXHb7ae9IaRGPWKuEvXMoJX44L
pwsAxTVNNmibV5Y0yun20MZf7S5wMRmUZhpWp5oFb4VNMaNM/UR9SmBDyQaCewJ5
3210895+Cs1zWeutGYyCDUqIYXsE9Q49v/38hukw+fMYm03kZyMFI5GArpzhcsxr
`protect END_PROTECTED
