`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3vrYYuiqJMQXL6FJ82cU1pIVBTDoR5SUDApSIHHHzYttm4J2nl1avwDGB2/s0onn
Bx1WSMNZj2nFNRf+vTOAasiAHmEUBEOOZFyycYz1ol03NozAHN3nvfIyvc0zM69m
ccM4r9rlQrGQXo51YCk5FWGfyHoqo47vEMb0E77OPnALME4gU7LUhVvcJaws1msE
1j5x+LJQuYl6fmOheX7tLialDGmZAcSpEiuYhHQhN6Xhvg7cIEIjyPv58z5CXN2T
bL/M6zTkrnzB9c/xXu02A9EuPNGVbBLrQaYwyUExaOBtaxIA5Yj3dPK/R6t4KsgV
LOwkBZRx21JcwsPHMADqIIftvpdvx/3KnP2yT/oYS+7CclTizaEt7YZnsxd7NIpn
jMAFQlWNm2Hhcef+6LQeX0PatBp0+goq/34+8jNwwlFp9wM5ePHwJGbDEf7J2R1R
uqHOBu6n2c/mldD1od/havcxIjrXun5Gx2jXv4ckpe5qwDvzcN5ZDz29RkeBgmhP
HPFl1jRkx8CncIrwr29sETdHaqT5xHdJhVEhUdRetqrj2xMZVlL8ESlW4Cn1Yv6S
rgROgX0ivLkZqgRzIcp59A==
`protect END_PROTECTED
