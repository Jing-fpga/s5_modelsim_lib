`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HRx97zA+CQDVaVo+NT3pLOdI4cAwCarzWZg0y+1ZrAbWwroPD8xcoQIrw2m9CHH9
mTQkhhQhliVee+jQ0/sRmWBqUiXaBCqgtVD+ZobLhzYRwc89CU1jNmuc8KmAUahX
ADqyVRWBaQtMADOJCXEAIydt5GvGdLjlrDk+04KxNI2auAdFfAfA15xRjThiSykK
rQ/zWtKwCThpBJqZNlM4N4N2wDr9Bki+i3iMq5UgNd5mbi00HcCuKCbsQQPCwayT
qsXoQ8xvrRgAn6bdvpg5uZBtmmE/kOVXnySGkAW7ooABAOLr3Wr4mPdC6vPlwHfD
jYZqd/Wegt/T66eOvX1qUv6WHv4m0VdjnZp+Ks0DiQuf6e15ZTyIl9alnS78biCk
q5UQrRBKP2lEza67P3h8nQJZ8fYv5iyeUbupoCrUzesJsA0sC5mE7U8KhJQn0aff
4p8rTA039dkdlXlAsGGOu5uHotnv+SKTgifsvi19QfvjqwMpr9GkbwLcq1ROPqDk
OGUjxOM/TKycZeoMmyzPoYP3gd/gL3Okk4PWyEw7Yt0Skj/qOTHdK6PZKfx1wcf8
wfoGSF3zkVotSZl5Y986bPGi7w/V5WcmugO8E3ffhRgbG33KlG0aWAsiZjBFYkIV
Luodaj2Nip2zvuSkA5hAsUoBNXY2ITIqo0CPvepiDC5V7T0BkEWxlgb8rVeJi4Vl
IGeeY+cL+2Yk1VPZaX4vxyh01dCqias1G5q9JBEpxAetJufROGBwJk+YHOF9cQrE
DvGVAnpLl9cVTurknmv1mYxWLPCeRbd6XHPXZWDYD14PYXNu8L5PC7nXJfK124q0
wFAc8IrY/Nqrn/FXj6oy7ZjfcY1CNEKSkFW2RJnVbkWSOFx2DNUecpyQpWLssA1B
bDQoFEZVQtFXAVIHvAPQb5zbHaGQyT3OGeQj2NKSUhQM2Lm9zXSEmYthZngHK9et
5xSSNFX40tQd5usfqWR6++AS+787LMmRIZunMXLJq0k+1uBLGhTHWBTKSqVp/U30
evuKVVw6/ugsh+AVlNMH7STZZawJe0Ldqec6OwPGvGP1si6vRyvhek7Vn31NUAOX
4QvatvWP1zGT31lKpbAEd/6XcUi/o5Hm1X8aFNPXGFhhpJ52SS9djS2S9h3Qyr+N
nVG4Oyh3SwLk1AK/f+jrkRUR6qix6mU1ypUjkB3VaN66KAbXxPJ40yTW84SY+F1p
dAgit/S3np8SeBpsrJhL7HQ4reD0IkgurK1pSPEeGRc/AdXCu+5p/XzbCLSQk+4a
wBQLxPPV9aloFZhMpA22PINBxgx/QQ9qcrZrM3p5j7SdA8TcwdRI9XBf8Fv3ui2d
bgAVPuTE7l7MbAJFFZHGvQAEz09rhWmSaUfTA9axQ16HkW7j/7G81dqLrjdb3xLw
VcdvFnAE0wC6b2KlyTe5C/H/dalW7pJyNF91dlYawwHNjHGrURYcupZpz5+2B/ro
Uay7jI75uSbXnMkro1nP9TP+AoI9H7xVa9Yc++yB3NDKyqE0nblolhMiQf6g2DpR
Zx8CvYWuLs+QGYGi9AAIAx2+GcU4GASJaUgTj3yHlAPfzmGcDapTeT8POatLHT/5
kxSJfkIjiLUyjPEuahNOTuDcqmRbQNBvVpSs5QfNr2N5AUOvpNtiGwdb91Hggqag
eryJO+FMQc331ibvqK6w66ckWu+lcDAtfk+xztgNXLy3CweOcmyaNhQoM+uvqT5u
41WdqM+dRc9KUOccwM9sgLuZHb1iL5xvb7lR6HJLmU6NDA7fkbJHu6xzvcw2FOvc
yRbSEj2HNevISXZys5dEXUfuQpPYsiyBJhJGm6gtwgCqLaroQPmvbB7T22fBG+sI
p08DpK8nKyDI4luCGz3dmfwigEleEhjJSBSKiwWPMySw8zniTMsmwoGjNZuDuZxt
IyM8Roi+zhHalJXMY535t8cun5Ot/+YcVOeCyTUFid2nC+VvBJQXjoLS8Z/07Auf
cydQ4uWNQLE8VksYdYJE9mLm+cePOwaxGVxyzbSgRA/ITdctJeDLePaEicSu5Lja
aytsNU5DWISCXkAIDYiaytY5d8bKMPAs09J7Ihmz4eXAZDyfxPMWxyw9KI27bGyH
BBICT3SACAcEsowh4ex3nfbbrJUwLbA+TWmtcPA8MCBsycTCwGRoMrGXd4txRmF7
8TfJ+djrvezUAASLxBaWo4lzpTLE+T9Z48s1q50X/Q5ATLTpD/wa+OOj7R3qQJ6v
bcQCAKn8w0ZHyeIAIx/mwv678N7YQz4GEkOgrEOeCQd6xPUkxe4VX5TxIxfpmAEW
6whDQewKE5Rs6JeLiklDJ8RJPrVl2/kniNJH9qtuoDRaX6BFhqOBrjUsz7x0IToK
ZgMLX3vlLPHtf+peW/+vSwGV+IdFGJzrR7j1Hs2bhLIJqiHtMCM4bav0otHdP347
W0crpRSNFYfgCqPn2Ypn/H8nvjQXOXqusahA2AQSbUCCof4IXy3b+peIUhRVEfGX
JB8Lvz7Ulf3yV+MpgA/TNSBCA7ArS2VOUfYvFhzAaKf4v8Omtf39YqDEn8S5lvP0
8IGt/jwvisEvIVGSa9NINYkqUDbJzS/qkFv+fMG2Vkj5Iq6J2/agFP1GHl25eMMP
EigYKwB54h+IrM8nDXVDhGpEeiqQ93juI8kdtN/uF1KFoB2No8CxmelO836n0Dt/
WasXsNq5zEiF79L7NUhfBZTKHLw4SXVOMSdzK3DQy6DwojJIXFVQKhWqYnjFfygI
OuTmAAJtu6QbQ0g5faWNlOSijLGknV/F461hp6Ekz4HG6IV7mZqOyp/s4iFjQ559
s5x3xgKSFa8ECWOLNltxPNLrAoPV41eXAor/TrOLpNYA7ekf8AmKVVJDWrzeCuEm
gBm894pr6jdtJgyg5dqxzlqAO8w0b0UU3uPdnE60aXQYRJadegh6JPONevrItljd
KFtK0yRhPY22yRk0dkxk7tu7BmP7oGJhHGMKm3WYj8YGD1V8qu8ToQVE7iSXPTU6
LHaho3cipjryWIUCphkV0XO3qXrs8Wj9iXvl1zPs2EmveKbmxT7wbrjDH26fwNB1
sz/e4tAKuYes1YiLXRxLNcafTciPnqD9S+wIvUZIyWt6cDaOwqdTPaZnrJCA0/qI
BDHN/qAcl8QflIJT80iOYQTXeKyEtwBd35HwpJdyQXlAHVnuHinJ+OL7BdoOCT9H
k5eesMio4l8SHDrRORejLfWdW4DitYDGl9FG9mQqW8En2mOBzOJWwP1tJQlE7BHY
GAlbT3m8m8tANuuPOre7hdh1ACWXKJyI0U7Dsra95/Dhqa1ZTXjw/LQ8+U8RXf0M
kneXXh6zLpoNAywCYRaHLDuwWipYG8Ee844MMG1+4kFT1npDVoykd93fU3QEgTFh
wq93V50JqnKFPJ4YidUpy65ongKwGQ49kpTPALBp5dhdzifNBK1wgB8GvZ4fRkUB
v9gXotrwljdOwwc2TfMObPE9WYlOF8qXMpNiSh64sTM2Kxo2MR4QkjEWaNxCz5n1
VMgwaRB+3oznwbgYQKhriVWZ6OVx9hwAogoHgst9gV0iDPxd6T6AhMogwuuP7pzG
cEAyB2P/CTvbDS5tNCQbTOQVIhhW6bvNL8wzNcvlRIxXz+yUAu7UIigOn9eLQhru
HNhZWvkGCTXOkOQ+2lmOohny8LJYrTwDT67t0/7vKANBeLwth/0THbq8nEL4cAGQ
iJ1BcwwrQETppdvdzpXYFwWhes58TT8MCexwzofmPzyLof+9AU2w3YNuzG6Dj8yy
KGmSvibYOOS83LX/eGEsZfSMI78VfxHJn8B2FKsi8XSHbmPOj6tpMdIVN36Q2MFw
aFn8jNUiEl36/4kRyKpDSTpKG44rAv0FuhoSbK43D3wMZzCN08Dlx3oSev3ZHn/L
MoV7GJB0rtptTRspeMDJS6TTbvyS2RQS5ppKke4Pl54vDNVhV3blRXyHNB/Wkpz4
hj1UWPOwn/5N7PrgharPPiYs3ffCTrfTqs8fP3GB0eFegI+2UNMav0HeZZ1Qf+iy
uVOqOQjgSpHgA3ykLOU7O0grwgC48mZrcLUu9/4Kwqo6kFkfF6MiFwuHuc5V9aiI
psRax4FawvxPbJesx+z7LTha7YC7E9TzrKVl4FigqkIxCmfLTUzNQkH5ayQ1ys9P
2Piw9zLgk5CVMZjLyDdUcje5EV9OL4I7sSP82bxj1aEL4uqUEYponaQNQxZZSb/7
zmJRw+s2e6Q58FNf3BJY4poFaqV2jxClbYgISGBluK726nl3H0sevGI+Wl2aioFF
RDngwXG1mrzAOY30+6qDTUDEh7tuRsbevBO3pL/uyJIB+EA8ZBIXUmBWsVeXvBc+
438UaeIF7sfhxuxDKrnhzPHLmwHZf4jYwECRSxxnEmo9nGRQkPViQEP5T/p0BVn+
zH6lNkyZzT6GhXOnIg1W/295k7XwmUD3T5vs1YxLA+YwkbIAunLylRDfszCeU9ts
c9+PNk/ranb/puJd1L3bJ064WKM75yd8LMm8S6B45effaCcPgCy4HeF5wPAGBVTy
6WFeJH1ffgj3Z5x6xY1voL93i/VCf/DY6nSDuHKMHFLQqQ8gCMJYWeSPtzEvjFAh
U+HuarG4pNvgLomo8WAk+bDuGENRobBXYfFu8a4wXxWc+DP9KXtZAVLsEu8sdu4t
OTfXPWzOn6kbXAPlg7UdeJL6ktjIqVKT5o4j959cxZvBIJYGxfNmFN888WzI0Reh
MfNyaHVAUW8Y/2toB8Ouyn7m9QszM8z9wUhbPsHgpBlt4g2PCfzlJkTsDbyD2L5j
OvSWti+cU4nmySiLCk55oywWMp5JyaI9tMQwveBzh68+lIQJlwkgdIjV+cbk2mCp
qWdb18zGaSieiHkWZMkCz15Zy4ybym0p9kakrACB7cyJSj8NGataVM9NvCpr0xDp
IW6YIyanc+Hn5Pbhkelzb8109hyv7jzP7EpWFoKH2ZYCcrm6PlLDgAf899fmFojX
iWZ1mjypZUGn/J2gyhS7oyKvvG9Z8tU77SEwyWut/5pPW/vw4IKuXCaeusUqtx79
CvnaWT10d8mn2yvaMi8s6SRdDrfaJHNXbSeOSUzhboUuIxupi4AdrlYYE6Hawd5o
vHW6EOIv+HARz7VS71jvQQ/sNX8vI7MLdewhjbu1PT4V066gUWQXlRR/oY4erArT
Bg8QDibHUsCOl8jeVUAl/hCJbMrFvBBeTNs6pB7krLg0fBRLQ8FGUDZiv10VSh7R
KsxOQQRJ5Ho/Otnk9VqO1NTq8uHiffa64YkV3GIi870Iw5o4EfNjq0Mi1NQCQKId
RDlhZJYQBMbFbFOb+hgztMGNTvXfFv/J8OxUkyRXabNalT/sb1ztq0PSHaJiOxZi
N3LC0OyWa9U+pEOlFjDeL7cHIfuApiIg0PkuuXMAJ+swAx/jX045t3SGgkaD3UMH
vOJHPKZqqc3D2EMb7hzcq6oHeLpWU8ImOqLPRF+4/Xyo3Er458VZNWOYzTMJ43De
A9JkyDA3Ek7/lH5wlVfSoAqXev5GvrbiUXe7xSavMPPnN4d9ef9cpw9Gy+xUo8jM
MMpFW1EouruJJt60nwN8kjH/XeZu9FY1zwvvqa/p1C5UNmRxZOgTB+729/z08/Mt
33iAaMyTuPcz+WSWDuJR0eeO8u9bJBArv1xtB5zDMjZIW9RJDVD2P7uHSmw9ia6A
mr15lHLJXWWdgV/NcSXqatGPUSFKySBn9v8Z93TGBDAu+JGuDURY0IUCkcsPGZ7p
NT3pATSzbN4wdI81gDPJKsM5N0hM+t9cvddW6Kd1Ohitb8Ti1GD0UZYmM6ZexkZH
zyegzNRVSAc9jaiRmMzLmc8epVQ1a8gaaEE+5wO3HPWLmd7E9q1T5bkKPcMtLcN8
zZksK/7f29jxgGSa/hhN/HoNCVs6Xg4sTghzXpXRy45ON+YXqDT12SJe7C3UIqrI
AqqVEBPFxaHC/vL9MEXaHb1F5K6IyHjkC2TIqxL/XqLvunrY0azbFTBZQBPNZ4Rt
`protect END_PROTECTED
