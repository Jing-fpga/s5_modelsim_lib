`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/X1qT7J/4rTTIwvUPLpL75fDy1WRrnLuSAJxTlVBF5183M970vLplV9tQfa06tE8
Ce3usBIZvuz9dDOjnBK4S4evymNopMCYxARRhS/8AyWoiuFsrXw8PfQiOMHbkwvQ
JQ7MhRfDJTAlCpeWsf/pgLXPM6I9N/wZCuqCOCEjHrcTumjd/bdaSHYr6wCx1pXy
41R9BoVFdDblEqanhu5mLnVjJXfIK0+8dV4fQC+9CxPQIMPaC8KmtyKPQTLYFNVy
XNwLRWc11X8c00mzFYToMqaPGuTwZMYoaAoRXkFxIX3brZnZzPVd/VT7uyGSFkv6
JSMNMld5uLSefQV6/sZcO+KMy6CxJAV7ktbYRzDF48S+L39PbbJTE6jXdKzAvqzl
6R3kaXMzHZRPupyoyGTq5C7y2rENrU8OBelKAeX65WPN3iLehd4jmUUAnjxQJeoz
3Wlu58rwJ3YOj7ehOVsU8IGdxBrxNLVGHFYcmGQVKmre5jz8YujV0gTY3fGHksV4
wUSMfC9UH+hAT6S5GkXzF4/iQ+eOHZX9fNp9Dh2Ci10OTmSYDleHAEmMCMPH3/FX
gJLPiU21Y2MWd4G9Ub+eVLaqPys0PRsPPZOcXVvUWHyo5d3DTcCP7ZvgzWsBcEGL
FJ4Tiqc0hsr1n0+59hqK2COXW+TuXe8Me+/mdWUZBcv5y9vDP6mFkuAbFocSPtYo
akTF9ObHO9jvlwvh2STSzRzJOFb358aUWnO+AhElOTONsbGyM691XPRPm6MbC/ui
YEG+VO1Piwov7My1JFB0r6e/57OX+1oPnm9CzorQak9fZYzFov8qDes63KB6pDnU
RxiazT9DhQvccLL3i8cbF0p6JnaOBa8HGcL82+HYyu+aJTIeY1q5AOFngrggH57W
QuD1Zxi4PzyKKXPTaKIs4IzRjDvQLXk6mpMfBkwt8vK10zja9PXbLDgIu1cJBw0b
QcoPTenGOpPpo02U6MdnPLw7lYykshCrShuMeqydpR9Yub/PdHXYiT350CSzEWzI
eFuIWJIn6sPRwCjdVNUPz5jkLTSf7GGvGEIq5hX73ODBajdVLA8UPS1NKlVbt6/7
+BuxqlSeB0RuLAOgbtGTy+x7XtEuSdkym9jJnqj/EODAmBr/mWxHaAbMy5zyIp79
SxxFhHV5JSZv5++x/0Lu+wXYXE4hBFjjEJMlMe59tao2JkMUbmNg8IJvi6GgYTgX
JrkkgOjSws+JO1OJq3PWZJMFw571lv0bDnNcnl0GrrQjmyJh0UF3iq4+Rc4v16XS
1e7yNriwAQfI3NwmW2IMzw1RTBCwAfqWUUyFEqSAE4bktchr5rfYoXPIeoCExHFV
NCeKUqdTvLzLi6c+uakF2cvxRY4QGrxtJABYOnI0qq2pEPFxdzE/azXAMz1N2ZS8
BT+Ivi8pEnGDqR6FtKMRJIgrojfBQiWGqRykPuj9CzYTcghP1DG2v3uD1wsv/Yxk
DocqQfbyLLux4IDd+Vk0lSkkL2LdsaiArgcK+0bd8F6+0FZu5msmdoONXeAWw5Q5
hdI9wMwMYq7K9sJ0LBmeI6WLOdjfCIJqIi4hZj5WfnVGCDjAP0kLjNC7g8/caXvM
vIlVxYEUE6rI3J/iDezyKftx+5bG3dKK2f0Jr9rN0A0CatHOP1Xw7tDjoU4J84wZ
CwJmL3ntoSS8J5nXZ3yVfSM2E175xbGkZoEfrTIDS0VxJC56kC20PN/XN4UNR2vR
jJLDVSZQtBA1xYghnXwK8+vJqObPD67eBBNHGCjcq0WL5y0l/O2y23TanmPHckAJ
+rfL4GhH702iMuxog7yY8BGlaqVQEI93Kg8wxZd0oBxWhFxnShQM2kZphU2etoKp
rmrkD6l7ZY82qt+gH7BueqMEp6K0vpZH9vqtT3wXF++wwSLEtTJfEKu6/4cUndcD
`protect END_PROTECTED
