`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7yJ+nqTWrMpNLP6OzYpqfxJa7XlQjNxTwpexDDtSb06pn6CkF4YfuTYk/bUuxwUy
6S5rBYxTGFd7+UXejXnCfSfdkn7TU7HQXXooHoak8ajbMX7i6m50hEb4VDspv5cc
DNhcNeoe434Qt/RbAYaulDzefiPBLpspMTrGFFOGMlr0tYOqFs42bQyp09sI9IMw
eQ39P08KWF99gGXRRACaVIR6iG2MNktjTsNlaiim5LlukyJOEzlS162lcO7lkNQX
cg1mD6s3xijT08/3Riz1LygOIjJV+kkCJXwPJVI7m1I0MHPWIgAO5+AY2T07Kyc6
gPFDjOWYbRNGEKKzW3UMBrHGJ/Ji/Ky+SfjpwGLqSNv4k/ejEKdrzBTcQ5KgNxye
3xwdy4bJG3cHH0mV/yn/4F44Gz+D3iuwo4pnprB8HFmEtHC5jTtRG4z1Ogtq9J4f
zvOibWzoxkphrpFgttaIru5NEAPZcvFPISXwDRFJ6IIeW4WVawl9eNfnn8kjaC3P
4+PYrJdA9P9dBsRCh/Rk2rCiGYej6gBV90uYRur4awN+vvEtIDdKfkn5fQ5BWmY4
UAigZYn84ljN6b31kZ0q77qO96ZcUdkmGBZww2AC8LafMzLZv/EB7IjJSxCJ4kDa
fnh7xD3Bwyxv15B6+TwXxQwgNshDXZ01twpdsDyvTzs2+/CCpD//Rz1IwiLO29mM
FWa0nHvkGNkOpRT4ZagweNFDPeZfBIzTWOwrdv9yN3WCcgQHSoan/ZQs2eqrPAHH
mqvuGOB3mQW0wtjFrLnou/RENsH/uFzN4l9Cqx0lGT4XqyDYjOO+BmzjeOwg8atw
B9P2jy3rPrcOLM+bgXILXJMx32ucHVXjyYD91TYWOZLCoFRMyLue5b2zwLnP3GIa
i0LfJGgXzLIKSaJjUY+4sONknI6nY1b5oHX/iUnqFJ8Jq6G2cfYbZkZBHJsNUj2i
0z4SGpsKX/KJpu/kSJbpn2WtmQHyOi7I0evIW09yU/JqGHoYX3J0aMgtdtKQMsAL
B7rk/J9Qem4iCsojPwYEKBCYi9rLxeDbiqHovm4DKTRkJw3Fq7zo9xID0n6Ylgvo
//KeC8m8MgZUjpHrTLj8dUv0p8Ga6ZIrMVjlsARVNG3t0evqAWiltwqqZXB65GSZ
npHHDA8xmStiX0jUgiRfB6IbUT3nP7YSNwIfsrDTaCKl8GDUUeaO3x6YIZqXdBMf
reJOYu84H06s4vODNezHsH5JmK6HBBjLpXDDbcU2RCOV6s2sQTah8P3yONnRGa3r
LJw+ZovC15OvEiQw4Y6mhcLi3A8AhesIlYXOsl1BW8Sgi18afVgq9zJBT3THSdYS
WVTCwZKE/35GesWFJDBHbpeO79dfpr3xuegdx7IpHPDOC1sOpyYnsQvxLbdnnRf2
v9Vi2YU56QGUTdoCswR8Snq9ul/ezAPs7b1Tutw0RLeljSSQnAq05J9m6UozQ0/l
EyU2UNLUH+E4oLoEnpGH/z2izICnG4RxTtMVyXrZrwqD2bE/q30JACJLBztmD0KJ
iE+V9QQoTRcT3yhi1VdOJp4OUYCnD0nGxAp+ONDOhiTH4LiX/1ne+s6kPjXXsF8z
pOJQBpoS6+VqxcIRLsQoAEM0uYS1WJSqKB72/1teYRVqI96OxAZRL6boTEDn0Yu0
wPF2G6ngTCuGQUQeIIPBGBsWkzq97USkMgo4tI4ilYpjGg4yUsWKD1cULfEjLLrW
DWYOIs4ZODJvztTrK2/01EX4ebKHfy0ahSltQQmkZP55jqX2S6jvJxLDjb7h/MjQ
C1TFT7hk9vcOsSYk8Qm9xHn19srJu4ghjTQnrv1uPvbrwekqN8Z0qHIgt4tfk9Jx
Wp1E8y/KXubOrxXchx0+4rBaHCEhefZBTvwX6gUIJ0St6JamkZWq4D8JI+nhPzLP
oY2+qfdA2v9NuR0VzzZERiY9JAWcG/2boj+taR/PgTlsZy4hZfpagHrDY0YNK/bX
qfJmctfbrInoNryH3HumK7pgJ8Yrnn2QIgVGtl+oCfsIE8hMt67RNQW6cuPEr17Q
ZSLkO5C5wn8xZPepe+50GUlA5Yu2ZsP/JLWSP2tB6rhTsUg4Mur5wHdUf1g04wpQ
q1Nlv2OYgDdhLEPnz+lX74q6y1KYDur/Glz3M0DMDa8=
`protect END_PROTECTED
