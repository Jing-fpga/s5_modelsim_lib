`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ks0OB0oQtI7hq+F82G/U8lE2PIDRPrlevu7RyJ4q6ihjC4TwzAvKE3vx1nB8JRmR
J9JXOMbm3pmVik5HGmVMLQ88WhNS1bY7fUxj6s5ZYLdJmIyb3LIM0HZd+w6zdJlj
KisfqPV8lYmXn2Rf8KrRiFz9imNxu4YFOvQinA2evnuC6EyvxejNjtKtE8vDUfMu
qKlHVF8sxEciiDNGQ0JYY2zX6BRj0ND6ykxZI92HlGqGKTN08PCMYFlEJtzlpUJq
afSPmYIUJ6gCHMirDgYYuMZI2y7NQrgSEt/59NPu4+wlFNL2Br6pPLiqDtSTv7sO
/3pDc0cgZOROKtSwcazro4f9OYq7Sou4MXzUI7dHLeWIFOzBcuZfWKcFcqfxDOnW
Rb7zMIATNH/8Jc6U4i+72EYgrj8gYdFzko1RDiFipcXmso3f1/+U5bi3jvkjO1fM
D96NJ+2j2AS50LluExSDQqnu+pj4hE1NZYvqfSaax6wa+hiXliIHcj9MvhshOpK3
K/e8u7Z+jualdGlLwG4Zc4iV+OybCCufm1Moy6xGahAjFaRBdxnlgFEIEEXL3vef
13nTtbzNCGGX0Z75rkClQqgx/fjlKQy/MwHOY9JAWS0F74O3Wv9jGNWgsHb/A+qk
xaN4X6ljVYoFyfZ+MdIz/i5c72JVAzng5i/MMfGLM/37WWbqdOrE6i53XTFgJDxO
rdiSw3vs7B6FWzP9M1G5BmuudGyIe2Muy22LiaYYY+WRls1h0gfkLM3tlmQEzwZw
TbbfWdg4k79RgJvdn1AAVYvxL7zb1HhvJSvuUSz6rZ//HymUOvN/mjZ2D6DWI6Y+
YU5cgkcZTu0O1EDR9VjOl0qC9mWJvOdZGb/997i12RR+KLw5u4TiGWLjKd/zfIpt
jOpJ3DO1DNXULNDVsz7qPERWeRkgMI9x/qchtNZp5k8RhdoDXy1A6S2V+h44yJw9
ysIjEpAksJLmSY6HQVcCdX0tPVJiIjeIhHcZCXO7i465biJMDCK3YQlTZ/FLRxY1
m7C6mbb9MSAOytjIQ0900uD13CLK4/L7uWF7yqakFw8RNYwoFBvy2tEFj9bKCua5
WRuScdGW0fIIafR6i9kmQTJHKU1SrK9w5l6GruLStkgqbGpdfQwsAf0Yx7Eo1pSl
yxpMYMxNdI9yE2aqX3WhOhf797NsbHfzdfaqtlOVaTp3djV84vHJ6fpXaVou1t6j
FVso8o7OtSswxL+rMj0QYg592hALQHCqNw1mj7RpYTbECKXfyE6BqwaYqm7+1KmX
7XpJYF5rY04NPd+dCa0DG3FIC0o8ulG8x3aU6uU7ReE5F8hSGWclN+sNB5+o6rRf
Pn+DOt6J1pTsrhdlfnh6x+246XRdJB6/BNiju4+incKoTV4SuxEauV6Q6euM2A97
P5S/2jg9P3obaUSwtSrERc76KwtCrs4kD64Cc0Qj9taWb1j0eHIg9m0ozxWzZOnV
aYCwbsccMwuNFCBQeyolHdbBCyQgzhqmFvCcH9hHrPBH1LcDKs1Xm71/7Z0nujBH
zmEGQJopKfrDtjQz0+9BvpSOt0ntBJSdxlzgUCTL0aUbbqpdkFICKPpb2qXu0pZy
FpmY+q9jJ1PDw/tpsUY82AKh8EeISgMEHlaK/pNuhCBO+AvCFPBEEkblrMkawIlh
ziwJ2gGZ7BjgvxvtSX6OU3vS05jjcDT4wDxtWZrPFxgdMnJsxJkGYFXqBgtotQU5
QEVmQiupLKkABggrkY4CP0VPLeZtgqMwdukY/HXhidhZJ7iJQhn/9WTxUKHh33rP
yxHbUcitrUuTFTQ5qOA3D8NdEk2IU0AvAGNNivnCOhPci6Eiypaw59z60tDaSVys
4I2vocyUwiTa8iC4wINLIoCBaH2boIluiwF4FeII3T6mnjfm4xXrctd9s7sTtQ9C
e/AFPCdPtv1ft7/a88E9BUsPqH2TK9iFqiO9jSDXCgCe5lAPl93zwmGB2nGrFVhV
n8Xel7S+krnMFSODoutvdD6d3/vyO8eluS7b3PJY97hmse+mSwmw4RxCohzMnEhp
ikqFD/wpQ5OVTpMy436BgVpBx+RQQG/mnUHOSqebZrlLWh03rdGn696Lg1/FRrtp
usQ38FOEa+mF5PeevgP67zFgTKi33xtQkWUTOYJFxeR9ZefVeIFcuZDzSElylXY1
A1Jqsqh5r8nOGndOUXuH77OI/tYsmKLPM+q2z2ete4XuoAcDJ/dgRSN6GbdYGHCJ
iraAVmnkWDK6LEqLwNT9lWP52LS8kiR2Gl/v8rMkfHQ8v6SLQWZdYZx1xWpQzcxL
2stJeZpTq5ulTLCOFZCTpT8USZhBMDJQPMgXPZwhKtNN/vnDE78H8HeQM+UsgwGK
KzpOCQyg0d2Q+Oz/ziHubQ/wRbzblAxnKqZVGHxvLgfM7G7B/v7gQ8ApVorAE/iz
GrJh9qtds10u8P89NX6oyrNiCu3qNpaVoL+UF+6BEX8nyzqh27MA53+IlOUZTyNJ
NO1/yqJig/3FQBPtXMLNj5pKIsk6Abf7Udym1SzUEyFmpfs50aoYdJA2uFOLdZ+b
28WKfuEbb+LupE9aO2NTlgRQrFA54yRzaQz0iwLespW259kiSgn8zRTnejBtqTNm
EbxBxHecnEnWxSVsJSYXXwbwZpgesL+Ie+diYM6J/H5GL2Y7DrIQwol6Es4Tj3kH
43pn6oo90vSRFOY1/N0gWq6WSUS7nTW6SvFQWuOJhbiS6Fs+dyD24WKGGBSvLhc3
bCL19Q37jgGiXNa4+6pWbeRlcAOTZNBc13RKNbghHTmlYX6aWd44apIIWQWXqjpH
rtO1vKHVaxaKCsanWmMjerx1EaQJhtozC/6GEqYg93sIeMOKjsGUb7bmLxiYFNxP
EgkGCrizIrIStLMMu4cWf1lOw3CdX69576xsro825t2WtWijoLF4yKRM1ArbbKzv
a96XYhk1CccfBL23uIzWfAk1Z1NwJKNluEla7pFpfnWYZ9m0Kcdaj/N1YIVNEaPv
Rtl30HvvpY40bEB5+JEv6Nsfju6hqFb4NaQFmbtrnUdKjcli86mdd44Xz8g/vM8i
BmyC3PS6NOnnWB4GPnUkKuXCzDLJ6NGARaME+dZu1bqRBy+SUwdjqRu0sN/bBmlh
ASzxEza1NR2FuhzqF8Bpklj5ROGDZstBJiYdcuAAYRpMhDVhVs1PsTZA3z8t0DJi
j6nhUKzvdLTjLXNgA1z9CW0j29RNZCaPxVhjJ6X98gXAk2/uKVZZPTpmmNtesY1Z
GbiMldrBHzRL0RxPb371Ev9XXozTNBZ6y6t1aAOIFaXkBiQDTj4E4TM/Sl7nYLa2
3N9zOiAS3FfFf6awbMK7DPJiguEqoScq6DLkNRWrcPpdCGqLVeJdK5VKThPav9jK
rK1mhWeyoqThh1Bwgb+22nNR9hcDyARihMhSS7/ZXx992v6XK363Mbhgs8J4+vet
wSkt+nwiTdmtg+JXCsMJOCvrK/xdIu6h/jl6Ga7W9r8FFMkEX79uuL56F2BPmoeE
t8PL/grLytLuo2PDEzZsZWX1XzqjlEBw0dEyJObdkcVNjkBImykjX8pCmwVgOAMH
J21gd8lLJAkjbSPw4YPHV7cDv8QfRsk4GyE3ILUKDonLzNBNrOFUQjaDbaHpeuL6
6QRIuneazeGMVzJniEm/cGicY2pK3v7tD1RfcPS3bNYkoBCr8KUC3Fs3kpO/toQx
xXAii5R0h9qI27PL8UmHVRci18w7S+1X4fs+iu1EiBOFAdzafGJCwXB92mz4UzOL
ONurwyJbc0EHk7LbzRqTOZ9Ki5m3Nt2pVPYXXMeApP/ORoeVi3CNPQWhJGdkWaay
7GkppB2kKU7oWGcaztaeEetRfhpYCjgIvnBYZH3lW+ym/eqd53z9ijoboc9D1iSu
O1zrafqdnkjpIqmmv60ZBTuYtAGxS5RSvjOpsXfLgOaK+PiFLOyOMFqKd/ad8wkE
kmjJz736e20FKMdzPbIY3JKgMQjmeuYRe6E9tfyi6ulNSeCA4TQfxScEktarQrfl
YELbJ9esYUwyorSq8fhZnBQkU3zveOygDMbLRmKQVt/9SAfoffRuBslpezf91el4
aJXmNqbXbQmVFqMsexwJ3Twe+hr56uiBN//JVx5bXAv4xu/ZmAOjVs0Cpiv3xU6R
avNwE7LN7t7gv0Frx2FpgGdsGJ04nlRjy2/Lonh09Le6nxKA0b+MOldOXrlxL6sm
80SDsHfKsX/IrNHzBH3LroOrpOjrJEdIdYZijC1r6hFl8PF/kdgA8t6rxtzBlFpI
DxgUVMlCBINHx8N6Vjmuiyup6rKa3eaqtyV/nnrxgnhu4Ufx73DCgkZd/BNhucLi
YSw+cv7a5ichosMXu2BJmySd9PhAfLGZKNz6tuxXUV5Ywr6FB/l7r70V9k8WBtJR
8buqBueD3fEb62FaXB5BspGMz02lgjb4pWZBnohZN8x07z4wsOTcPpPPXP08lGKP
dDgAVFLIoQx67cOrIpsuL57l/+W+f0vV0FapuQqI1A3ZV7cWBH861w6s9qfGGH8j
13ulOKT8wwSqOUq92SMO2WpBnmvRVZBw41yk6w5SpDGILfhBCcmsBQY1N3CfqgE3
UPzhoESbWBILgT8T1VjpGDUTRzzahqyeovOgBOKZ0b2D0wS4BDrt7VRrm7CL58Ak
SjlG5344rvei2+8nLm5vA5+7rnZ/6HzXd+raEI7fQWysNmyDIPd7Z/7ZcHpJlY2s
Wsx108heWPnDzZd1nUqN4ro7MNmYXqvaWSy8Ms5eZlykUHacHKp+825OILdhYK18
W2hCEt7IIXrJVjdU9ERF+kRqbyzKT7PPcOgX6J4TjMGj1ifsFbLTVs77PpaZrzxz
wGtkPeMIBaS2mW1Jkyq089gqqpKsNXU5fGXBKLuKBbtntS12J2Z37L/FuqPI1MdT
FCl5aP7Eh78LJT+uvTW3pmMqP8ajyL2YBmbH+0nMc0DeeHEPlRV9s6VXS10w+QZL
RSN4YF9U8OX+a7tqbIQaz3haLgpD1AWpXkMadYyzRsZiHDjzuyMFHD3O7lA/SPWs
6yg+MLBvhR/8y5hnnq/3KR6Zi2v26Qdwdf9mIjjsT07M/trHKDYTM5b+U73jqhzr
N74Ul9AshKbQyZeYjxJf3L1APH9XgTo36c0NOo+SQRKMEPPM6O1gWa2WTUStfZ+Q
TiCKZW20A2tSBAuwXWAxMsw7rjB8ZS22uv0ejEG1tfIcWO5ZGtc0dnMAvZVHKF4P
2w/AWOEeMD57XvBCmInQ/k1z8gM+1260gltdljtGgmAOwpsNauCekmgYByjODmnx
N4ZIX7iz3W0AbgZwYqvuos8apdlFR8EvKuTxh3A2hAl2o6/mUzYPq5R9llLD0MqV
PtVpLDDR8gz7RgtdcQXzJE9pO1uLoozEMrzHsKMcVdb7lMazZW7WJnljct75gGt2
wRed5PY4XVqjrtMZPhafa0wbifETZ6uefFC1f/vK38oTO2KFnTUnNHF0XJdX+gKL
I7wTItBO8aeKSCMWJgCWa/uWArwF8DR529gaFTybddlsI7yVNjdPE8ytu6JLEHpQ
Q29aTWsEBNAQ1yRCXGBg6rgwteMtM6ACeR2hC71RBgGRvMGNFsIVQ+GTBGwCfamw
Tb2okcIE6ioGoYZXj5ra2T+dhHUHQE51fI1o8pYXdFq30I/+1c1JRAkrWLE5M6dV
el7sux5uqH0YWM4Mf/ff/1R3A8VRnO85TFWw8A2jE0986/A4rHFvOhQnY2TAScMp
oBF7cVOmCE9W0mRbiJdBiZMqPNIwlRIaABxrqAQavJxih0IxkxXWEtvSwsIsawvo
QRQ/AizOXMjRgg88I/lJf7BboJyOeyOOsBJCt1Mt/fNDQmOsFSfBuUczuX2+NKuV
fhisFWnXbNghQUFQ+R1PktaL3aoooRPi085M0Au44FpsWzJJy/HquzYZlF0F28rW
9ZlrleIjub6Xk97mrqCUKdM8OBFm21Xl36EZJsz3RNT8IaGPbS79udH0BwvNC91M
wjhsQIXRIEHpC1BkNaR1K8wHLFtnXNtHuP+fhT/jl5gxWJfXKBFwXImLyrymJxBG
Ado0riXbZ6eUH9J3AnFadmg26mrqT7h/sT9+E+B2vE0NqMtDJmxs9jfYM/32TTj3
/h8Lckf0SzVkj+AHtJCbYP6SdDJxyCi/lodR8jwpBVH99EJ0JzCq7pJe/CJUCpZt
a+odip6ep+u/0EOZjQduCsS+wbNO9TMNt1ZNjja/Wq5Et4LKhSwUwgfWtS6MqEob
QPa5lts4kEg1OfMfvLO4cUf1UAkQYVP079zptBPAiF3qQujA3fUibg3U6rJ6EzXw
i/qgczzQRWDqh+a3NvketIl2ZJF7KpIGWSgd/soFuaVrfR6cvDFCyQU66ee9fVL7
P0L3at/e3JFB9wOAgbLbutMpmhcwmZnnYJk497s9icJzxEhnR2wh27TEDOHu4Tuo
mY2dIgbdB16bIV/W9An24Vqn0jDnaz/59WdZlH+rsLXF5zO19rBZNfVXthVBCAcm
YCUxG/keVUrbsSFw9S7iZo1AAeVTr36tbwxc5lRgCCYMN0s1Tb53rMgw3LzeO/p/
Jg7C/d3QtapaEz9R894BvZdocwAtOLxzgJORzxRjB+friDn8rm4aj+aOW/miUbXR
mZ33ablMJWfPbKOSp+4HjuIMsyzoohojMsrDXT3FGhOG3iRiz4VzghETDoQAUF83
V9DpsZ3Tb18nGXXhnDBAc50qYe3UhyJXLtfAuj33o2m4Y8IKcA3ohTi5WqSvz4B8
vT6i3HtC++h0FXUIWO88c7fWvDnEiB3nfPWGUZnWHfP1f201u0mdo0A4xyaVSJlp
3yGJz2cB7ijc+9MgZHV1VobRiI7Mp58UcMasAsmAQZOKZy6fwT1UDvI4hXjPMtkX
UjQgURgSAXAMegOjK3os1LlAt1+HieWIH46gLa9+Sr9q5hJoJraZxXILF6kqFK5J
2Kh+Vg/kvUpa5e7h60m7betJqPxPZ6ZkQfFjVCZgMR4hcJJ04mCsA1aiNDLzvzQY
mNsRAJqeilCFry4B8lPodL/6XgeqW3UaMsA11aTWzr4okc0pY022ytQg2OCXgZMI
8bIz8ECZ6OQl4xuvt69rb5CJrR0eGWgmn57ves8PWL2T4lH+dEwQHPtyEAPPr1W9
0FAErPge0AkeX7ZzKWxmk+vRrsskb4fnLf8mFOdk04OAEIYsGd6fmC+Cpp00VQea
53n5rj1bFDv7+mKsTuDTr8iSRWHnXigrPWWCUvuvOCzSSzskdF6T0JRVDNCKlkTq
tkSIx81tavUqGj0kNBZn2PYSA8li15AD49U/qrmJsOYkUsmRr5mhad+VHSOYIhQW
uZO9XSJJ8eDoDFXocT/kqHIPM7ZE1qNI+X6z5H6MQNTYba6Cpl7ZdpL98J57yxii
jnfenre5D0l3d9wUCSF8f3O9Mq6wo503mAvRJ8B2VNxGbiDpBL9lAhsU6u/BnRlJ
WWRBAwUPhHAE2CMf0oVStD7uWoahwUNFQYSCacOdmFJtSvywP5XdmruJ35JZRGqf
dqybWYK2MAaQVAvZy3l0EEry6Zc+QqxtPjkZAoLR3GDWI+CJd0HXVhmrinI5qLYJ
CVn2Ix68ZxVTY/tEzq5vb0nn+FLJC5pdSDIW6Vapwl0wbDtPfuI5/9dQMEIt+QCU
TqwXtGdbijw0P1d4dPeJzzzAMzpUf+JqWlhpF2PXJmYKxiGnBtzMWkN4gWm+PP1f
p1T8dVhVNBCZj97awYbaEuPuKgIlmJq5q3S7mOFQpS4FwdaNGUhRJdzKWjEbJyIv
Ayho8WHajDk+6r11ZxmHO9uJGnlbP3TETtgQ68/7T5ojnlgxLlJiR7ea+lph4kJI
7ltButsJRGL+g9gGbGHNNczRjVvpDuaXGB+pLUbC8qu4q0eBLmUaN+yHhm0Pw2zu
4fffreERoIt9hrNpBrxFWl0fsc8vEDWUx4c7O0Qf45hM7K/CIFaJKxsFGbZDOwze
IdHspQqvi1wMK/ZazEqCgmsQQfh1Se4YZdY3MKDj1VimRW1WEQFqA6wbmhR8LLTo
ne5i0HYYk0b47A1ipsq7E+yqRf5UyhSXDdTHxSxLEi+M9iX2sHTHF0/k34N0yDi0
1xE2h1ScE5nES/qHZtmowQGe1qBovQAL4rgAS4DwKwQj5YNeiEd5jk3d//Vsr/2O
1aFLUfxJO3f91gyvILKEnpn4zOa2zhyfhSiYaLtyWWs7LNdWuXjFK1H9Js2J6BuB
vhQAyWhj+c/KmLwBhgBttXShwWrrC8IBx9mGQMsOQfV0ujhOv+ki9LqlctqvZnfZ
mBJiowUM2iLDb04ffaJPm+Xtoj1A9D7Wmvr2TM/UI3PtCvEegxQb5WiGc0eQ+Lcl
wMyd0j1JAtVQl4p6vrODlTNpcBD9ZYaiy+hNlLhhPe0nHTSw46+TpTgA5rURYTb6
cPztOF7X8SWX9gu5tx69o/Np0cVQbJyE/OqgTWbD54hq7LiCJ43P0S/oWPxnQ8rw
F7glpkXCZHtNoTJYjCvX54TZ3DDNyhBS/e2UKqzu6Q7v/qEnvrHZNWpfSmKZU0gZ
gEPJIIAc14OxNvke+S/OgrtNsNuQmJ0lyRioCJKBJb5SyCsqN8jFv1oQ3azf4rwn
3B/oTXsNTGuBGwNYvGVqB3fssOLNd3hbGzaI+wqp9wyEuV1JP8jo3o/hKVLiDq+u
XUBJnnwBPR2cBbwW2GV1cxP9ulrU4oYHs/SEvRevjSuJuKjQuo7pg7ou8BDJaxoN
gdzUO0JjjEsoDuE8KICVLyREWjXJXo7lbmR6LcNYPPXYkK0nxbR7IQVH7CvtuZcM
ef1fxkAlC+bkoIOeaVKPn1jlXpmSRnVrzlMjMhevsOwwmB7Wt/k1gRjTG9e0zfyN
HMz1TDRNIM8COx6AWVAvLWkaJ6yCth3wGfXcgnUYcDyt/iDD9I3ly0LMETUyawfA
D/peMpAquRpOb7kb920+jXNkuBFEi1P23KtmHUz9rfA1ck14PjUnmafvnI+8NCxv
kCT0pDr0m5q16CDhUOf8DIaVCIKRIFiZKiyEQHRKdSLMQt5mfSfJUc1bqCsK4hxF
jWcVny00GQJxCdHlKTgOgZ5200lCoBRE4xI4bOIJNWfKxhMNovSolpzRsHNN4yzG
MbvCBtO3vgee1T9DAIBBx0lvDWY/0WLSHXiofnoIEZUDjMgBztlTuYyjqrBDie8H
qk7PQ6RFcWCQBYjMW96rQ73xiuDFK6lS3QGlxpOQlEbZETLHxtGB0s7ZW3slzNuC
T1Sq2N/K3aYWMX5X9b5p30WA4Vx458UAXW6vRFmulob9khhbLTlPmbhABp4/Y2ZE
donEfoJlW3O82yTu8aj5822QJ0a0E+heUJNuP/27Haz1jb2t1thom44xIeh1Edqb
w2tuJGmCBNg6bLBWAgR8Kme8a89JgTg+dqHD9cgygIprhu+62evjMokmsZThXy4b
LDbommYLL4lP1a/+yCuRYSVCbNHo1BJSw3Wt4QeiP6F5+FWgBF+U3kanXbxJdBIV
BfDG8f6Z2o9KoO0Ubw6PR8J2nhZy7rjnROy5rL/Ed5a0Ai0TWoRUQ+d0o/1WiC/F
qZci1wIYd4fuFoM3l3j5rhSKEOqa9S28JHSqrbto2IMBCDkbnHB4zTozN0plBjaR
cicBsC6yeLq7QTKEazB4ijmwSTBn4teuE4TofBvsjG0ifatNx3KMnuPxm+SmaMAO
XOmu5u0QfeNEysdtFL6wAqnukww/51xB8hLQsXF3b/FLoXqncyT29qkmqKqVlEn/
AQ7YlAfXal8I+LDfMkdYZg/i+6A0iHYtJ4R0uyLRbJZ18Kps7yM+0k+aJWhgJnZ8
Kb2XPZyaQSpWdH58QXfqunYeXguRVG8wL6xWcM6z0Wh7cqyE/GRvGkAAtmBA0eys
yLAJdhrK2ThKC9C9F2siq1L6mw9BGNyFRwOqV83TxCx06x92TkYUfsoiUzh7pHyz
6RosNK35ikcSwL6Zpl+ewspFm/yPygEuzeF89tZny/Moa0sHChPVByc/obk9NBKI
bXC7qS2+YKRe1GMWz6J0LG5otgRbonTAJPD9FUJxjqu56jL8Dq/xYRiwr60alzve
BwxNNVz3fQ/rd/pyc5FFmcGX36zP1+bo9GBQXgijlyRKmXWQwZYrbWmikbt6oYwN
KfeJnTguPOraN7BviLf8nc90d52UqtD2TPYV4edH0R3DPQ52puZP/68S06CBbt+N
7QiP7JafaaTQylK+jAKNr5Js/ZQTlEHi52P4kUq2qSkAS0Zs3yPcL8jIazk73FEd
5KYBPo2fdZ2LIeawDFVCQxHMWPWkkMm/neCI1wuZ91HT3apKpuv6VU7a4T6vFMkk
Kw21tGj0oLfN9J+3S3FaNrtkQOsHSAfeXINagOn5IZdfK2K51iLQnCztyuAjm6u8
7cuyCVSoZLxSinOIlbW4t16tD83yQzNwbmDd3hxmFxJ+3U/l8gjwcKUHHSUoWc12
nBon6RRkfBuaaBOcuxGr1MFUAZZctkKgHUOJXZO7Ze9ef9IdDDKCvNKnqFt/xUBD
vvfrSw1dB3lRL7B32ytYcJHjwm5jfA+OXL2BCQewhcXdBbi1eIBvY37Fi3IXmFlr
XEa9VlMJYCpTaKR9kY6Jdcgrf0Pz3S9I6BsxgXrAHJ0Oper0pDG8TqRsyjNUmWzB
b1zM8Uk01UJrUD62qfpmbZzcVE7X2tCLIRWi+I/rJjog90Jw+fSYllvaKWHBu2mq
FJnzgDmma/RIJzif09vjnebiBM/Tk1rkYYiIzY0FiJ45BHw7+Sjy+qUN5WoCZwvC
YPJcbQoAdeOqzOjtH6HNrFBzUZdNVFI5zM1lytNn1oASXXc12Q519HXvw0VyQx1p
nLBLQ7FTgrYQlBpL/epNXU3QLDoEtkCLVKbf9F7rpMz3VGd19lXxUAuJr9oU9NSG
Mip/ObLaLRo734AFWBV37LCfBVLZpbPu4Qke/yRbvD8R6J0dCnm/bt9CuUqQXSon
I0EjT+wgC1lDMDsaLFjIAgHhk7S4/EidzKozim6CBBBIS5W1oVTojsBi0ldHiOJz
AASyUw/A1uy+CYgkMJ3tprHdRJ+ogNCnY4bGWixk2lr/o3C2bvkM2/sRpEnUbBel
tzRfidMKv208bOH266O79qiEI7VtXJE1MEHLyisJhyUEu/jRW1QJRy3Uxq6CGMjJ
9CgDqrpxbJH2grXlh8AHrjeKSsZ72IawoHN6SCt45RimVOipka5W2/aDuw90rYh6
ba26shLwcmX0y6Y7Y1vq3FJJbG0s9aOG45C1OK50VdxYIBXoKEdnEmiLynLaM5Q6
JaPPDJS3kiYiOHp6F8SUXPD9inq1M4xdoHsEbbOU9iFJ5MA6coES874SSeNLTQIK
RAZ/gu0Aan31Oan9XXDURzrB1xOFbBNvkeaBE0F9rk1cxkX1/0bExK4cKUknMrtz
X5AzX9JiSBmiL2XdkSwNvvmv+j6z36tUHmmchPEhpqjmPsv5ZJ7qJ1ByCZ1kM0AI
EA63ygxvTTWx/s0AGoKpBoRAmHoKt2CKYoRbG/sarWVq7NRAjg9g84it8+BX3mXU
0HCsyMbZ1kNcPtpHGBWco91gVaPcpNXKxbyq1qMpbx0sypZbJ+aQzQObbJQCkKHw
qJJqr+sXR4rkw7C6tgFZrMwPhClwL4G9U57Sdtx9rA7SBxxx0ZdBsLEmmp2ZvDso
i8w5etAq+THw3O8n2bxgo4+FOkI/teGzzPF20J1KyNG4fcWTEei7SE1vGMYAtJ3J
t//1h+yJePZJVGoPgNg3UFBszIckfexhKUUoYmm+q76Mxk/9m4i+xUD1rnqPxSrU
ZYMtG8IMIFQOvH0fzuHcli4FaBLeoP6S9x0exKw/9+dm0Wr3myz9LnI7olGygWPs
u7s2mJoLsTCENIZrkYPHBi+9SEFWoJa2nDTlzEkHW+rKi36tlrZ4xIrBP8+fHHrh
aUUUiCHCueWBnObb2gaZ5ssEpVpBdJfmspPjiCZ2MG//RgOPa+BaLyaDkZktrglU
BRZorMkWyAKzuHgWolya36gaCYPkCq1Dn5z/FNUPEXB+KQs4JPdpgBU+XE2uEDsf
S6wrKtSljEF/A5uDTgwDqBCz/S2O+oTT2UojmqhtIhLhq237KSIayZfms1g58OsT
r62+GmXEJfrXOhgQB19De7W1IAGN0G2M0NXqKYvfelfZtvxfHeF7mBBpEmEt+IAz
+tDufHhzh9EREMXBbu1Bajo6AHK/xt6CJDlNvETa2WbktVK/Rvse7aC/cMz3j+qy
UH5CE0RN+AS52gl5FrDQ3BQmi0XRBOAMwOqK+zCBxi/tWoUL2t6NIDQWASZ96ggs
bm+v7McYN/zgGFNdspSzFnw0OOHmAsekNpbyNvdxRbhsh88aQAokSVWIRpwCAz2s
zxRSFjEpm951wHXQBva175BViOr9y9C9hkC+g3jXKAQP3gfjbE6ZT0jTT1mI0aMC
5ADRsDm56fVapKGc8FCz//QTHHbIIkgi6s4Ge2hy8tEnljhGiWA1SiCzP+F9yfQE
MM8qqd1AufYMV+EdUwh0SpB2UUoruy+C8EJyJO4zRJHQfSWpqisuCGHaYxGE9wGG
WwvMjkbkkcDtYgIUWbM+7r0jkVWeexyA1FjG3QJf5SjGw7AbTRT/F0WIBI5CgVC8
Q7BGxTbLwE1cPjhXoFBTuTrTBgrbsuCwyr5U+/Y3N4mtbyoENadtIoVnjyr/GAB3
wqpZHInW3gHAPqhQ7QqqPONvpMwMfgLYMPkeUw/JxH0SmVWNqXVijQxfQ+0vBa+M
QdA3+3UWdjLYr0NdXfz3LmMsHnFT/8fn4YJrJ1LFdANgj0g4EA+GZ0eA9iSOvx9d
5kXnv8YHp/FVsJj1Ecygm/dbsykUsgy5rrFueC90hzUQTD2SkA0vHf3RNXuVwlPl
BcGK4nURHHoMxvFujTTRbJdxbZpczKciZBNLPV/Y4WLRKgp6wZD7DtXPO3PU3rHE
B9dHIRdNXYDr+ft+9g4ShKOEtybxCylv5AEffoyGE1B+sr5BPnsVzpT0U3aqcZPc
ZSOk5FG9AXV0+3aWvqXHGkFwyNFCprpsvpiiEmYXTK/j1Xs7UuKcaYCzb3aOOYzq
tcctHZS7J646jyQ3FhgY/LMzvGmPRRsXyL4Eqe1NiwVu/O0Cx8cgN5ZWfX41Kzlz
VDcjRs82oxw26xCq5upK5GbmeQRwzDWI0qBAEO/jJqcxsfdaP+ut1/FTXme/liRi
/lyUEg5yNprNU4rdGKsLk3inhyMBFWhl9KIYiclfw/Jatq5TZBlZ+/1oQNDIGam7
M8HtoMCkrbXBC+iqy2HgFtE5KdOJfkKuZsiZADIN+0AiMYYbf6raBnv7S8ync98s
9dFrdkMxx/gGid7zaxXhQDwF+VUoxwKt5/N/5hXoHmjVtDoX8byBm634U0Hc+5s+
Lt5nR9IbjenjYTV2fiFY7nHhPInumlORMqBYa4R013WtX7NMFtW+NKZy5qoXd2L7
pxl211ozHbauH5n+S94PbX5vz70/BxfZ4DPxs7Vaa2LNtzxT/EqnvzVQtzEZW8DG
9Z52yLI5+Y+k98J07PITWq498isQeHrTXJokxRcV7wUKLJY6WqKDxNXRdAB99Xkp
W0Az/oX3Pj0cRf1V7prcc+j3MoT33B6cB9ZXZFMuq5HTcZYtuFFvzkrs67MUsQzb
/7kEjUzcInBBESKypLC+wvhZzgWbpCg5c0s5SIUw5LqHjN6NA5r+OJJFmKhq7uo5
AdJHkP0FTdoOo4hwmm+Mu7zgUMBBqsNhImykP14T1a2CfMMMheJIDmQncJwHwich
U7Dn2oouOOhJ11fV5Wz2daVqRp3OmP6iQDL6qEfBJYmhTQ/F7yCT49gvA/rxmhG9
sNC3CJtQcDViQQ3gpbSpeXSiqhAIpAgqh+SaLtmyA01+y0XIaYXWtJQxMVmHGnWs
nYu8eQqUFzbH0ZGkYqIZ+XBybz+Q5zgG0UhEJOcyOfdw3nLMS1pce6U+KN3sw/ce
jPR2SV4xmNg12WFOmRDDCUJdt9gSW2XbncLCtE0m6vwrz3ud+SRkbZgpdwLEESqz
KGNl6AXo+MtCjj3k9ghsLC41jIKQp0yELlx/TMCIKNa0HMhqkejMlN6cQ1m/f6ft
qCIk3DiHQgM1oKAzyCXKD2fBKBc+1OQ7H3nb7oSpeIhglbbSnlCQ6dIFm7RTwMfN
c4xjxcIgG7j7xM7PP1MsQ6n2fLe72RoQ7ZONNpE5MAzJBoGjOSLBP1xVzbUz122X
nHwqLNBApwRAuc+KEmpbPFZLf+k/4CYEJP+/6KDASAo7zLXT7wzMmtj5ff/sQyKG
SgqWxBf08DuWXvi/WgghMJ2NE9MQiIemm/2VPGxB6Zgd7gDxOBrLLRI+JIQsFxhb
ML8k39TgHtwTLK8kMkzZfDtIJUSPtXaKIAYnCIk6U5Mts5jiQj0z7Nxcn+yYYlHX
kAF0OuLX365IwZhPuzKICqLG608kXY0b6ByowB5lFQ8Ir+w9CrqTUjy6HtBiw8lU
M/GOc32auZ1fp/WUv7kgGVH7U7xzLL1HMjb7KaN3uJYEE4rzr7dmiTi5nYQ1tPg9
8Jlw0e/HlEH1E3fJaAkh9e4yve0+xDDjIKK+Ea2RTqeeK2O3+TuaL8YLIQg88HG9
FzX9/+8Ol58B0Gdhq/IGOiZY0jyTORVAklMovgjphkyRnjR2F3YMs1J0uOqGO/95
pBkWvZij98cGGecojDp8qLN/rc0Yi/eSPuq22Di9QIoxUJci6IsouGDXczgzp+fE
aSc01JZNueJcZmMyAB326YdZGyzaoc3oWxUGErs+oxMKje8W5Oo9oyihFkQ2LMkt
duMGYLIAyooQDDb9l0Nxm9FHvnds70orGr+sz0YpxPKu0p9X9LX/y47INJNqS0vL
/5aIN0qp0ZSoWR3jfbqkEDRVPZnCj5/UDcw5r09GY/sp05aMkLKOqeg8hXVf7uX3
OSPs9OvgWBpe0kuV0v+epwI9SDcbQ3ypaPwwRmMhCi6IXnV3cfcblR8hpWWkthR4
dvNGCWpGkXp50cseGEkeKmMirwaHkZTWsKzU4c+dX2tZsK0FKyRCs4YOEqRICQWg
gktMkTt1/azxsT5nNC+/10yWcRwdj1JsD5dV2uDx3mu/45HsJG1ag43tvj3muLLe
UC9ktKIli9J58EuvXrXGhvoADLW+hU5MBAVSOmv4jLFG0SkMCpMFe20q5ycL1iEm
ZjjJiIh3DdrsQfDBh1nHRX8gafQaRjhnEN/4oSpSiELl9ukDtROM/gDE0Y+hSUFb
xxEI/tlZ2SkQOPC6WykOGCcByKpcQOiAUAh5S4wtULF+z44+YaFKO5I8CQwUW2a1
WlNpsymrvTJm14lKxLOzj12d/ICbdfYPrTIWRk5qbwNxLgadQwzTFdXaaGM/ZK7I
yWrV+kBelun9W0A2vm4hS9xfC253d+wyPiJ//xVweA4+dPsxZy6XIxqOinVWXd6Y
ED6os0EzQ4bBvIpvKVaIPAwfM5Ohswpj/T0hzaWi73/Xqvg/3n2NqG5HDBszpv/y
P8jq/LaBEZLzR5fzokF0oEma6MMo/GYaPsGq+SD5BTJrjLIg88r/43mmI0lAU+4W
6gL7G8SrC0vhrn4qeOnHglO+ANM8HvHV12E1tNcdn50NOTp7LjQa8ltZ9FdH36K3
cIRHdotsVDyxpL2G8dsdM9+RAwHszEOppWrjPX4Z9IKxFFzFxS49XgBeaDHk0nL0
io2tCXzc8nCmb8h5OFEFj2mxNP6SnXaoE1lf6QAb0z5pZx5xgNkgrPVF5pRfdmKd
wcIK7JMsCLSO8twEAjWNXA==
`protect END_PROTECTED
