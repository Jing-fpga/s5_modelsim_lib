`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nDPOU5jfbzpMU0hzp3a4sVQnXosw0E/UrOz+pxw59LgFh0xfS34pVv4nNnR6ejad
SRk0TJk2VTpeUF1uIgo26D3pYohV/uzp5cN9d211KM2tLpX3FxlyY1LiC1fB4td7
x/cKx1TGGr+e6ae4OFMI5ByXVlh9htjrl6/of8A/NPXnK5xC8nzIV1wdoz9wG+8Z
jWFVCe1PzQZBUUfYj5Yr3pj8svhnXJJ1fDAE6cBtBjv7HE+OdJRMHymFwdgfGGHQ
+XfLw3lMixiQThXItU9+YIA5xMvXVSmNfRN6pxyzI+PgEy5dN8Ek+bUuPGdBknMc
1Yjg8zXtYKrjtvkSFiU9hGbPzumSNlc7Mepq89rmUqs1RZsGb8flUraxf6s7owAY
X1ovKwSjeQduVTYKuSOKLrCM41BTvw+Ug05h4/0XlACRsPUf3oTuqRuX0A/rohK6
gRFB+rjl3vCG7V+ILg46kUr7j2clprtkeNVtpYStKIDYuhJpyVEk+bfiIEjg5/by
pgEjuQHXyio97ujeb6Sr9RtKHfaJHiFLoFIk7Ia+cMYXfA53q95opVKKGDqozMgK
LkYSYzgvEreWWiKr0qbF/KQ8K9TY5GRF9vOkCD/X8sMAt/L0X4RsoNoe9XC0kv54
AqTsDwdWVi289McxO6gMswmmMiicTTpPvW0Peav641IezUzqVv5MkBlLN+6trm5B
NNp9XwUX/+3IqyJNzVB3j9LF2WiSOMFHfkTz401YzXBwTerzWSodoiAEm1xY1u5N
dQHhJpz8xRfHvUSflvdjsesm+iPbVo1ntmhAQwMv6hA+XmsvA6MbcPy/Xi4UAHtX
BADr9wF5jMahYjRLMjDT0BNc3hoG7oFeQq72tgzKmGwU6uLLNhJKn9czbtM74BCN
08HTbob3DHzjvNXucZwJRtKxO0LGL9LfCMkKEkCP5OQrljrAcphwTFUzKV0XvCOw
TxaSzKesfZawJ7lyFsS3Z7VjtYc68dYempnhXWHhuVTUv0n6pGvClSPodpn6cBCS
PvvfeCNu0VX1asD5uGLI3q2r0xuqy5eVe9BaesLgZec+dHdB2ANrlUFMSXAzdGLI
KCe/aRTlKkCqJVN6223/Ol832TEASrzFYrsmREixbNqc3lYmpb/T6g3Y/BdlMGTC
So67L0nNOiKzsWZ18REFUk2TNHGFGKzuh/Zlr1dqZ+vc7mn98kILLL2h7CE4xPfj
tS6Bdo/MbigP3qUPR3ANTInjif8iFmbdQkZ3qhgEIpmf9FXqPAuWfqjFSRlkwqU8
SAlpYXj632r/QW4DvLzgLn0kTyRpzZd23xaDdaqiMKHeoWV2Ie3Fyc3qzpl7/KbV
PW0MRwke0EX60gfR17goknScRfk4tvUJPMyyoHtySkZv4iXXicq3mrASepCpBD3K
lPRMaU1g+hYw0ukrPZCoIQ6BqLSVUk095ibML7toFo2QLsWZU2vhu7IcG9jX44f1
k81ib2XFZfTGKdyCIeodMnO09tcqjOt6ojKYeHSpSiBQAmpKRoUnzStAOtFgKr5y
QSmyqoV/KdAUEojqw1bwPtKxAsNk7BrtVHXlXb5QVkk=
`protect END_PROTECTED
