`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jyCKR9/X2yov+lux3TeFg2ZERCEt7mhH7kGkbwIqOypAgisxsf+n6UZOtBI8JIz6
hTR6Piy/z9b/htYYmAe+1o8f+8EbB/bE+RZhvuotNb81inGVhNUU1A2DJoURkQo4
QVZ8xoeptrTmnZsnffY3oeEtb417JPS4JRPPTI2mF5qlXfsa78MUO4abfXUrs73i
D9QHjBAF8M4ESfrIwTcZA7XoqQhAyTaPf+MUVwPmfl9r/pdppBa2dtM2QABwBUiO
ZPgO4+ktyTLnlEmq0pZ21mDTqbDBYW2qljR34BEB3fdj5rUgSF4DqWjHcio6BISf
gICuUhn5m8m78iskxFHRajwoGxfEsF4ROUBPBUlhuuuGqqkbQ203Uifiz0C8bYVx
LvQenjWseo6UTGPuBo8JgZVPFnvzfLy3/f420galcAlGB8IJRnuuBMfV8MWV6cMk
XANqxvWUvf63w2W6syw9t44ghgOw/KWlEjFbt+/utpXKrO+t7EXP8LofD5app30i
a8LL3F6IuvXdv7xh6CoQqFjuUJThgXMbKoCS+QvV+BQHfFu65VSI8hsuubiCJ3vq
+ZNuLCfp5NvebRLax1WF+d6NgJg1DySlp+Uttb/Rx4jB59kMsYubF1/W+yY/3xA+
mdX99lgWx2LjswZpjEeyLqXSwBm82emsrH8VGCleEWUbfLkG23RxRy7/er9iwrAB
MswescWU/zjWBQoltVab9ghBNSuX2wWGKyjuJM/9FLGKfVgSR2s6PBJEfB3R3IkR
Zpu04t6zMyZXQ+NhPEjVefvorc+FBPtJU8aCds43XrrJs1GLQ6FA74yUrTAsKHgx
5l/yjab44OBJugGqsnLVFoSQZKzbpz6gJ8YkU33o3dI4/qXaPVOByoZZUyAxJCdU
56upNs9MBKfyRtSvxkI3If8EuKNl/QTC0wojh6M+P3kGJKvB9n8IKl9wOMCRgr/y
dw1Kk4uj7h+eRxeL2fPOWnAfLhedAEOK1q3iYHIrEjGQleBiclmyqV0AImWjkPO2
bJhT+1N1w6PPgpQi/UJARFAOUNBFA2OtqnVqr2ZCwJAx6PNEexqp2fALpuYPfkf7
s1UA7FMCo1JVNvvz1SOcFZyBTNqyzI0+Xa8tVvKQHc1bfapnV4iKRIoSfc02G80U
itdExUUHsdc+dZIF8uAPRtIbQigvCgwmCc24RHgj9/2Xkc7odVdxgdKLWuvUlyKm
L/x/1Jl+5k3JO6aHSi48ge0ZP/DKYNn8y5Iq0QxDbxAN2TR/RBm4oiIWihmbEk3N
4PC7W+fJPICdOqyItXFWb/0u0W0xFuSQlut40O3WX4FwA8fTXy2WrVMayE4HxsbI
Ad1YsjekCcoWYfX3tCUJoM8E6AzyWgoZGjQrhvKIBxRB7oR6Wr3jQrrMtI+NXg4Q
ILLeDpTsq6ej8k9GT4FDbgQoTARno5V5EC9slomedkX3J+5ykR/o3x4NRq6FHEAn
4gaXAkp7cgP3aZ80aVLu2Rc9x3ggZgtvZVHPk4PuMjfGtrzTlYfmrCTn1dYqqctP
Ahq0CW20OwaZouxZ+C+hjGK5xcVBLoUiA5LdWmGndGn7eq7vXSPhVsGJ9RwjyIxm
eBV3/zYlrauRAZYbRJ7/9vnOhK/NXog8GdjZVjeW7raZlNm4fMIiTUkP4XIs6lAF
WtHBCjupkVSTsleylB9RjZmueO7egzlT/FM0kIoYlVd2VgM+HtPFzXk0w7w8w45i
kl/kXmxeFV8UJ/QRhki9+YeZ0/fpIa+fDeSM6QIlvM+9hRz5DT+q9c4b6jlHy0JL
J1kGJneXRXCaQji7lE6ugriTS4EGdPqy6AnCcs25RSjf43TexTOgN38hl9zrfvya
+Z9ueWsEvfCwETP7BFzKKpr+3AqBzVfsnpGmRi0zXhzFiye1vWvOI45+uF5ul2nN
PQA0U6wd0/n7DKGdbLR1eb6KAN+H8IHfC/TETYBxAoscRqXLY0YwhqNaNcur2Sui
VRRjVvN61QiBpQhfDTo/Ib60jtC4mZLnAnZXSs5ALCkw2uxo3nhoW432qKonq2y4
cwy0iSdVMJRFYX4NJVq2EGEXShKRm8jSjflg01UbWQksJvdV8LwtJIPYbfc6+C2V
IrhIFZhYJIDxDjg32s/a862cs3e8t1k8/XV5hPNVMuxcXngY/HTRLh94w8O/HdIr
X3GNiT7MwGI+mOi7HD2rq8sgCNgoafIedw5K1Z3gKRNny5sKxaZ6z3IjpZTvkTm5
P1hX5Ejzbu9cLU3oOQP+3cUnnJSkb/jbL7/NkFZ4Sb2h8h3P+WEdY2ylLIvDiQiz
EXCsOCBN3RBNvtIv/Y6CD6QfTPPXMUO+Pmn+avfO0YGdgyUp+Waua3KmVMR5CCMD
6K+WZLRh+zezkBNGlyySHarVW2AfkbuBLPZQugnCTqGPDcg/7agOaOlQ20pRRaVF
tprqpfgKx4cX8zSJcHBFdtuujVleQzfmaBtEXF6OVVq0HeDaMpPWl9Xcnwz02z2h
5SX3b3r7PM5dh2Meolys/2eAqOsdA/G2DD3XlQlnijCBoAh34OWS1wlQ+nrr6jGo
83pn6lPwrB+8WEMVcCeHZB3mdK+LRLm9RQS5Sc9fGDqVmiO8STKtLUxMd+Fzq7ox
MBZH2y/bhqBDCdOwAglHmEBB27fP3WU1vqQAFNKelZ9X8tHa+DZOaJTcjCQ+82rI
iX7qT9w/n6JE7And5Q6Oq45qNhH7m9DoUACXqThHn+HrpF99WpdFo9Qj/FNzaxF6
u9WCPxsonqhGxkb5SI739gQPc32LaCIFqi1cJdc5UTz22Zz6c3pNVz32Rc1HHKGD
FoUyXXXSPu0s99xKdR1OjX5VZxi1R0tk8VJVQRptWbWTuBpQJwV2fnDwOEXnhNLs
UoyNJliVmwTDcJ+4BJcok2OfT2uu9C4gdhBz9OsNIyxgcl2e9+Zhb3tZBIncJcN5
0Me/q6K6VJGuiFU2CdPxwpdAh5a+ufkQbwlqCih8tzXf0c16xNcHk7Ut08PJTweo
6jtERDgOnjqQKXwZD5OjBrbs5+FEBsm8qAmt1rk0jHZyz2mZVZmQNbwILnYCW4p/
h5EsZel+CjNTtpi1vZcwhdsKZSs4/OWFyT31ax9d+fopuV3SoPfjQw43LuhlgvXU
WJ0ZjWkd6pKYVT3Y6lImKqVpNLe4NfnYHx1ZLx7SiIa9jw0EJ5PuDW0ZMDLMwJJk
A7AUQGL3qLSJQ0jQZTuwYiWaFCjmAvFzK2XvJXupX39t+Qyj+zMdrGQ0pSsqeogC
o1T5GcKKXJWXA72zgFcvvLKzDCUlTlqvzK4trpaoCNHz94+7XmP2kG+R0ug0VaPy
q8Cz+ztCEmNxD4sEl5a9TQQKENdB/Y0Z32IhBeqrFM1YJtc3bd2AmYNlBQatZJHn
UHH6sQzE+PwMg8mi3vzUf2jhaUxpirEqXe+gaRnG8+YaUGGCiUAspU+0Dwluqu1E
oBtgRXqbceL2bpotJwq/yQ/Q3rYXhztVjvfXhFwadXWURThR1KlTQuLhx+cjGw/s
koPFG6lv7W/h9Zcz9ZHxsa9TaIrV1O4eAelP9JtVPckbeQDVaoj4/TBahdV0swrv
SYXiT315ihGTdgbc0R4e7X1V403sLxetaBxMVR7vY9YDFfD3kx1+Ih4e3R+NiyTj
q4XUyVvf1tRwI2h+uBIk0TODKFpa5h/iIMwVbuswOWIV1dkc3jJLMvFtRDDFymVd
TwxvG6TUzvt3utZ+UgEkuSYD9xQEY7J9e8dB8C2EEnZaD3PP9HEO2GpCqL5pdQBE
Na15Y2nZYqxAG7CZ8CBTxuoqWCPG8jf56rNxnQKEIpuAV9TE0k2uOo/AweRlBgaM
8sGUJW7JqCfX0fZamQc+OCqMzr537JxZ1UM/ugWgHWOONcQIHWCr4cZkJVBHo1BC
rbQmwnyzf65wOKm3xak3kN4mYc6OLKDkHQRRGanz8t0iLrQeYjvcgrEmUqvm0jaB
WcodXYF13EeyA8pADJWgBIH4x1tHzpgsaaXFDFVlOjDSx2iwspAvGmeFKeSSDK8O
mInwBrSC2q/UJvwNEKkB0S5qgDVvaNvNCmzRafXBM3zcQJulXCyKRG0zoikTrmjL
mPOfGctfMKYwiloVRMNHw8k16Xh6hA8Vo9bb0bHdm0jJUfvspA5A1Ag5esYdTO1x
St1hA0m3smcozGbOdJw2YQJD1+L2y7evIkOGXirJlRShGnRGjVKwihe8oibMQ76S
h9cUXt8GNhDl83rZ7L2QiKlZrH7GVxGpC2urRk/9d6Ie9VRRJUE2JvrCMXggNjAE
I2xD8zkQxYS11aoTHDCux6pJkMc3ilRxwiWhESMmXWUjiApTPwIbg2bpycfhrvdx
0MdXRUdXcOgnn5500jPJ4drsmLxicRjJIi8QfnKXlwOySNT4/F+I6N20UHDc1xrr
IpaqVN5hh6kmx1w6P3kqFXlgsFqDl0AL3qT1lFZ3z4C/A8KrC3umpUzjK99APpxI
IhavWIv4FVnJBl75LUXZJhouNyV5lApXjJU6e/NS0bW5et6slIuPMeQyvB2/cIUA
/jzp1cV1Qpf0F/7KAxPSd5ZZTIqqGJac0EXD0Tc3uDXBcSVFKmwpJ8owxEns3hYf
rNMn+Q2yCViKzxmSnDE6X38HjGCofD5agateKKxd7yo07RAe4/HzR0mw2Pbw1/ME
EftIfGUyWovAZ/XpfDVLY8EzwIXPK8Ik3VIediIqlZK9rPGTcXgWN16+1v7MC+Yi
6336U62JzXOpRZfvOoLCyQN1XHzBogKIoIJSgiXu2txP297jHH6oCBey/dt3pPiS
X5BKTPJC3tvua0YXryXHbJKR4rzO1qyq1gpyNawcFIFg19vuUWo9hSzvO2qex8I1
aPGLms9t5iagst9xtE3G3xTYAVrmIrGNI8tU1edDYBCh4QeGIlu6lVB0seMawKIn
j7ML/Aj2m8DpBpP5EWkhK2M8xYKoyzpG38ojvft3Vztkf+s0iSxGxAdpxfy0JVt0
5ymtzjhP5fQXnLc1egAnr4ZjyY2aUSxpZoDjGrjV3ujJrMriNSXKpMUWs9GlYWFT
yLdApsaLzx/NUVBdn6UTGeWiWPrfuUM3Tdw1o/GN7CudCFj+VFTPfx0XAsl+Mq4J
btTu3i09cSoZ5S2y4jHDnso0IkANk6TBBYgJruHb7se0xVxGAF+Ig+Mz7QUZEi0z
YCXrzY9NOY2UuVXp0gsuxGuGKMkLL9A88cyhlY8N8paY59rw7oY52w1rHWRL8ces
9dDA0MJzcJBHhUr3zrhgz5VfYoeAZ4kafUJ4xfp8Bup/1cyjopCrL+TAvihrDLa6
ivbaA2yPCxwvkHW9RuS8oJja3tGYrdtYSiXm1X6Vw3tR0pXp0D+so0+kClBaJsHW
oKX10XmkztIEMtUTjpo3rt45uCNiX/l0jJLA3D0MtzcMI3ZSGHTSWTOKC4QnjwhN
ENAQ2K1n2wNh2r8Ju827ghJr5AtSVPfnuc3HQ4MRwq13lCBLwx1ndKmgWlpYobde
fBQ9dwY/MmAu2hYo3DH/MEjjnsCbEDbcf1c90LuIRF5//CY3m2RjFmOTM2ySxD9/
gCYekm87v+OSSvIu774HsLAzpmfyGaTqpzR0Jv0tA0GrT6nKeLR6ehbazrAqA8tN
zA/9DCsBiV7ITy1SgSK+zcm104h9BJDCwthNrhkkt96WFrpPpHwW6IbmUbakw+m9
oJ5NC34Ofn/7dW4//k7xtetgWa0A/yv4WrbriZf6CqaSS816NZGVkhi44mjWu6A3
xojOqxwrvpCecGJLN6D0CUxl5frgRVkavV1Y7mytyMw3Lf7sK3ItqgRoUYOg4W8u
aM2K3r/ZrRtIpPl2S00o/8lEDPmcCUjaOceimT7D9FhLX6+MUZFnNvdbLUNfDga3
H21+TdbMTUXZE7IQRS7EaTPxfQjWHjM/vY45jCSV7Wd73QGz7SvV4OGBWBb32DTv
Ozd8swV/ulary08f50oefrVdwtXld7eteFqqPmGcg6Q1j6YAbWIxiO+1NT6jA/V5
Q4QmDTidFdaoOTLxgSErks4I8UAenePd0pkx2G6fL3FJ0KGAfug3rxUnQdHsvbuN
u8iCUBGOo0rvH9vc8QfPYvken1RpS7HWBPqsI//ZVKldUNpTq6wS+Vw3YidQLNYa
aS0ZL3HqfzlIqmEH0Eiok18WCKu39qZ0FR6j40BjeY0jjxpnk6pdtFWvXUnTEyDZ
Cc2eg8RuXlXtKPgIGeG9VUg256pu3vISx3+ZTYlyJeVDfFufrbb9fvKsUH9TJToB
nVqGXB2h7cJwYG8HHGZe2evd3bXJms7pcwv4VIfDUoCRGvLra7VA/Vfa9/AGmj1z
g1SEYY+PsOl8siyLCk2XnSU0DoBOsw/9psMCmfwBHsolEncCJuy8atCZIR9idxWb
k3k81xTehwKIv0qV+LNyag/OU8emOtKGXnPHtL3Wtd6YmP4LZn2/13V119urUkSG
ybg4iPYvgC3wKfU/gUlegCwNRVlAeKmzoQMYArBjFxM1GOR4Jqr5uUr04tw7uZcj
AohBQ2edt3xKexRsttZM9Jkby+dLDNo+bx+eyZOtYGd7piki9XS9vFzfyMyd++Vn
JMB5XU0scoqI4OIsEliLu7wcXaLoKRupKvJbyylf/0yhgYVtHlGmT0jkpl1fsOZw
baDlp6v5ygA3VDJOmwpxAhvnxM5d6aUcjZarYsjDJfb6I0lTn5yZ0/8A/EMy9V1C
pYdLdRa5jRm01PTzxRXJaeSpgSwDX6ejx7DFClZC5edgH8bm9cqnNUdaVTxsy3tN
tli4BK97+LXF8KqF4/LujWiJPV3x/yLIl30ZamGYYS5widPaG3ZsSbkV775Qkqti
ORCk44gY+q38Gde+6HhdNHDNi2SmEu91yEQPF7awsqQENQE86+G6cPidMtBnkZhp
Y8ZOziz5jorZtYvwlXiSE7ddZWQxHGykpw72roXJfrwT8TtLyPXCbBin0p39vjAS
MhkyxL0VEnlpUwCgduoyeyJACjtT0WhRyL+v0BE0vZUdvJmcJ1M1RM8KHtGavLDE
SnJKTGQg/0nYgkAvvFv+VLTPRMNt9NNIJEtihJVEbJYkUWHx5LKLYEn0gClxZ7TW
K8CaaCyMzLPlHwqkY5Ids5Sz443QLSPznfUttUlTi8afOvEw363KLSp+6md7CeIL
BUc/mMmi9pr1R6FS1sqSJRaawoZ6GKeigP8MuXv0yi7o+i+vhIg0ZZpgYeNwsid+
`protect END_PROTECTED
