`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hYjjyUYQhgNALi7qjPFnIMNV2WY56VD4P4wI6KT1udrKcniVQhrdq+0MNBaCL8Jp
M/XPxI/xDnWBTjKttIxGd6StukCPke/luQWleg9IQQWDGxgLNFRSKJs2sxOEVoAw
U5Zt2IaUgcW7Bg+yLEk3BFyKHEiBtb4bZp59eZW/g4fQiKRvuBTCsx5zvOVpSuCF
uDvzfdr0rz6L8I47PSCK1Dq6td7b3qMHZsMrLvx6XUFONVm3XbQ+Oj97a/YaW3tp
sLBpoLmy6PAenNByymrLVYS3Lyzwd0yXMX4f34NMqSJLMcWI1qzGTejn0bUQTWD/
HHv6EuiDwFfU0ocMCa+nPBzWDaxbimKXpHj15Qva7aZkXwxIrLMs9qGDnTDK0KME
dVgXk8hIZqV5JNwCstKleBh33ZBhf/5YIE43IggQ6CS+AMCmqzHJ+GzOQm3oC+WF
3s1TIs0qssXZPc4JHi5t4TJgy6K542wtyM9p/fRYONYkRr+K2ixIuIOrchaWffkH
cAT3m1VOd7skq7viGFJDxaJkCcLPc7GgZD3aDIrxZElcozpEKh1/U3pEAd161cMz
ZVguiYiP8ucIL41kbLfYq7ZUzBzEdn16+nZczhYtSII1TGcZBubnVVhPSt/7i/+c
oo6MfHZcnkf9aj/V9i29LSA9qrutjrgxOsO7omk5RD879B7qHMKxfPUAJhiw8oXC
8LeSP1NnD/UTSXZyHGrwKIat+FEtiDmxa5UaZWyLsmhx+NiExn9PWHUUpGCtTLu3
u2bpYF+thAfYTtRUqqcaCa0Rya5Vf6cFJN5+Rg69UmPpzvhIB3ZxadRLCtcCKm5b
G8s+U+UFxRCBH6wSyQ7GlbS52vFKJfo4JJ0sBsaENpai10TDhUxUZN/wsALjKig3
F7oq8mEUbMA86uhI6/VKgiiMTllt0KT2dWkdr60yvrwGKBDDGSlZ4mw7NahHXMmf
r5cZ5rf+EgdwbieQU8OQiigDIB6gXVSRkgfumTk5JQbhA8RHLRqfW+1wYAGrEnDf
k11VtSfYj0DYtnhtEpFg+che0mMUAfP4i2hFPKgC07VXgo0FPdg7BDIwsklat2HH
QvUfNDLyrtz6VnatJjJNmSGg/Wwzz8oNfGO0QSWmX2Ygi21iGqafJ5eAQCMM9ByU
LhmCbAMVQb30pL2Au9BgxoNfzVjTDcA6+DmjJDun+BwKHYKpDWSO58tGQYsBVgCN
40QBeDu4j/ZJVzJj8D/XxrL0WBTqwry8SUdl0KYRReWd8BrtzV2nxT8ip7VuLhLm
8HnIKbRse8OuHokXE0nU+L3BOHsftlBE9OMQQEaWlCLAXsJQM7NHG3OWnYyzUNy8
qEd2GclDc/cY/qjCJGYbea/oQbd25mHKr8hRziiPLnKnaU3hj+5GdtQAJHtZ4E1C
fq8YAmmY0Fb+HkRUEsGTYtCMK2qs9mf0sR94YcsEm2rRIBnJVPXHzKh2QrjoeTKF
ul5Ec+Wi8NwAV7le6kWylZDZYxK+0A0jQmMP4UDC6D6Y7e8XKBWrwKKzEf7fvH5c
sUh+U6Tg4U+DyvrSdZcMqw/cNF/qj0cQYUi6TWWmj2F3N1V+PEOGVs8WfPhyF34k
LLL1Qsbm50rbHNAQQTh+axKzs/mICbtpDwZ6iDzWIAZNiVvElQYkE6ODjK5tRuUB
w0Ryf1PhQXgcJbIiR1x2mKGni/CxIbFBCAO/7k1aOVskTez/85tp418UdukmdyLK
WgijDXD/FcOKMvmVTj/D/62oRRaNsBWMUgxlcIIbUNf+47ks+nyvSEoBo2MQaP+J
+dYfcOYmeYd+XhmZZFMYNoztjuTcOObw/6lWKS+xAMWsKnGeQ0fG61wG5BXXvrIV
OVDbgjlqsx9hmrhx5etaC4evfDm04rEh8cEy3q8jv4LvxKfGtUYCBOgByN62fS1r
FWfaU0iaqxI8RipD532zHRwMR8Fl0cxZtP2kFyUwNoN9VVaIfjHMKvOhBbiAYZMy
Nuc8LPuJFppGoDK3RD4f+fMIjLrP4xYuXi5PN2GYLt+iAFtnV70xYoCuVsu2j3Uh
1b0ly2NSH+uHtDUN0Y7DIHQKOgx7UoUjZ+OXPFFVn6j2jx0SYEFVU+hdRPu1BW/Z
8sG7NnFnHJ0DQLNDYKZfthZ+xSKM5nJ+itL7J/SJF5LPwH+oBpWbH18HzuICrWFZ
CZ4BLofCXe03NHiZm0x6ucO96+Yf6f9biwVcQhZ4QbN39SxI2eDbyQOhliuIVal9
RH0It9lrpFUp7j5/B++3Tc8fc0DVe3ervaAFqu+Fktqa39Q4TSxyaUTr1+aIgagM
TKSz/ZDw5aWz2J2wIw/KnMrR0H4e3rJwQfwd0d6wvD/Kad3r38WoAPwjVr84y6Q0
FE9/Cy84CT0TM/uA950E1bezgKhrvqBllHWXzUc40hHT8LLBQt/veku0Qkjjn+Es
L3exLw/UTRtNBr6pQGXBsXECMGjziZJTvP+On4y0lInTyzTIujO2FO1piykee6Xl
JLxrWPf9c/EUlTjeBTikqLfoX/++dD+EcLW/Xy02iGQjN6hljV52ar7UY7qrvYuT
JOZjLBnt8fVEnWa2yA9HOTsBz49560DgAHgkWgNRw+qRBBA37JHXRQYprOcq2jDY
bkziHZ7mHetOChWD2/e295cgxpUsxGa94kBzsVNdoQyUjStmKh/KRtj8MD26PNOf
fy0m5GNx9Zh0wBLIuSirhkRK8gKajhOs99lymQ5XVkKd8bBA9jBbeWGGMVrR4YSv
Ot8df5elFZmMyLJfDJeVgL71gjLkXeZLA2KVM1/aO4XqzESXCCMVw/QtvCorae3v
haLFSn36dPgHUl7poWex/YBnGd5klHq4RZQ5ULgud3VBNRCNQNQlTOvP5zT9S0p8
gmXxMz0lsZzAToCUSXOlJj3XRZ+rvYCPjKU280XdkCf9iSOxEoQK9BNuvjehnkCM
Z87Mm7dQhNND9PeGNuubzvITx8FwYJy3woVSBQbw69Cfp0TgEbwmide1LrAOEcsO
N2KaCpUqeoA8mdCy7gbQSjmEz18/MWyFt4G2S3BhuV7+57tZRFrhxQtvj6RDYANf
KbLh9aOQv7jaaD3JHy5N9t79Dbl89I2LyzxO2CNIGeb8C78JnwnwrxjHenXcBaUF
OQyJh19Oa1YymD4BIWuVxagO/CIv7P5U+aQa8tQ46urkIvi22G3Grp8bg/9clZER
qGfPROqhD6psshjeFj/QchJ90PJpatOmhTzVEWLc10BjUL2H1cHvnMpvEstaigs4
Kg6zQSKvyseVvF1PAcpCDodYmqkcbcArWPHV+GkYP44C8UrsGiJCc54/eMQfs2lO
lkVSiGMUYo2Ame52rLtnzVRECf6tFFkzjHQqojcaEG8k0plumdZSBxkKZP6y9QFi
HTZqXohSKhnlaiu/JkWByQFd3HkoAd084yh+haT+k9Lo+BN/YoNUrOx8BzUZnglO
cb+88X09/ytnnudC05HDzuruzRcN9ZGN4bxTDAG8DahVtE6NqBGqoetAniAmDfS4
p3S+t810wr3P2X57X0rSW23tIRIdKmMGDKIIFffQRsGD2NZ2bltI6RW48sa401NV
2uneA63tTftREjX5FFLtR538CjnAeFh/bqKPrdtrbpD0kB3CjVlVI14sSP/7NSpa
1ReiuhfxGfPW10FLqnZ9o3ZH/mN4LcUF7FGRdZsQRkL19YUx4qjcYsNM+qOjsWPt
KySdTKUPp6hgmpcX76IveOvJI2fugtv/MGpKLCNpXhYBaBxbmmSLYPO7Mi6RoEr9
6AfSNiZ0Y+kyh3K1k70DXxGTSFLx0hczLsdD8qsKb/CRFPzpVEgXLb8oWHppI8jZ
pdjL2AyuRRBdGArlIA6/OynuqvLrJnzOZjTGiVs/qrXIOv7alR/hK95BS47CUrEQ
lImgzFgaNbH6JiNmL3upl6o45V5lGxI8R4MskV0/wMJq2MeFI9ETvUzF1R7bUpYT
pjUj0d696lDIawzfjjRnJrtjJ08+x2OAH+SvXw7wP2+uhocwel1vrpYQCAiyETN6
EIiD2nkqSMbprhpJZwW3ffcSwO8LGVxQvM36MdFjwwElAm6Y2uIj5V98ocXHU3Dh
+S9WtLTi8xUh6Qwx1IF0S5ytMJIzxVfcxgJ5bjqYBhpOIcaRlB838zTPpuPO+lom
p83w2hWRcZUyAgNyD+rQ0XS45fIg1H4tyrPUG232P6eYdIFspe4Y8/psBY69lafQ
i5OCgKmEgd58PV5Ark/g2OpoCRaIT/3rw6yvMWG3x9/la4qjHag4mxDl/2VKyVCg
MxVw9chqYTfID567lwxFQW/pTurIE7iCSSpTKXGdB9IeC+iwxZa1H5T7eKS8WHYN
B37fGOYiWf0H7GR/DpXOypKLyYOqFlD5rtSoy5XXrBR3pgSVOUZDESXMW1lwNGqF
NgfmM5EIHCQRh9EhTs5txNyu6gT2ngdSw0OGHGccQ1+ZFQuv57me1x80UxYPPI5p
/9gp9qvLrYsH8sNgigHox73qZo82UB2STi0Xj/APFbLY+a2tjAxiDz3jSeVxR67P
Coyq7WJwrWO2lkU8hVjWNcu8JipEA0PjAREtRyZMGTmh15sbHjf1xLxbf6H7eyia
JfLi88DSvz3XTT0XNp9eEjlK3koiMvDsjjX/F2SB6bVmrYCjYJghj0Mtpi3ibbjK
eVJ48poTkVkfAVdHybkqsaltPWPuF6xbg70cxzS+EoqYTdcoUEb3BfXg49nvqxox
P12kb2dCcmhMEx6TlpSF2QRu92isiNKOmNTeXoNfjrd489ifhjWkCt20OX0dAHj9
YGm0Sr5a/Ktv37GqOEsC+LmegUk1zpIRE8VJ9BvZSNbPDXB4hQ/ESy2sWT1sBGP5
exfVgE8iLiC6tL+0wwzgv24Qpy6IN5bWZ5oN+nuSKwQRUBC3P36ZyjBclpkAot0Z
dmwTiT/UDYR4eLqszw+vGMGL3OtuC3vZ6mVTVf0yngqRdc4OoE2KYzR0wHu2aolW
QPCKl6kwTXmrmJn8Q8BENnqQeEmIbiK8AqAJDfgyNbXErTj/h8rog20gYK7yB4ti
6mOi1WQQJ7k09XvJVAQNOfqqZZn/RZ7xz1Ry6TwU8LCm3XvsBcmNPPK89+E+kfUO
AfIaIiRGh9tBHOaHHak5yPtE9I/lX3g1K+tkH7fdWAoI4meC6AIU9Z0L/pTwoo4F
hQ0PHwHhcNWKZmQ6D34OA1q1KSHgnhuLKl1EWdgYMEVEpAxp5Lo4L67IJ4KMbY2C
yaYUlcBDPEYVPSZ+lx90Ak6ktv3lYNgKzCmK5YEVijT6GeIQQKl82RbNGvBhlOB1
LpUrTb583EgOO2ktPcvuy4XWRGKfM8CQjaKQhLyFV6ctO0i09jWkVAI6AtO7JQTF
AAmEfOl8JoiRkKZfMLPQjDdk2mEJ6JNL442H6Dvga/esPiq5/mTkjpYzXkO7iFxk
rBKyFnRx7l6jQA1LlRC2bnp8coL/zH4UO10TFdB2xu6xij5vB+j/9sonfOi2ZW2l
Sr63XK8j5dtTqe8jMsiVJijEu6+D2ZMDev9O4EMFE9+TtzJo9Uyqpzj29sp8GBT5
7C2YnG/dd0IT/5fKlCUv901BAfjdmP9Spcw+OvMnbENg1CwIDJUMT4w7txSTs+FA
SyQFj/UuvZYqc8vH4tEeSpMi0uvXmvF6Tcp9oz0eTguSm6pK/+Ecj2EHdNxkJ+vJ
j6cX3W2MyUkPCI+9l7uelyyeZV3eoZIQQa5E1m6WHI34obcadJ6FYArEb1mClhCR
b+6UDRcaFq1HngNGyhKRBoDe/OqjQOohXePnhDd0GFePtLIyoy2OOC2+tr87ON6x
61QAMFaVV8zyiKAQJjZqe1Qx44erU+Z9e99KidmfpT3HJ6y2gCaeLSSQi5Zzl9eG
YIX2FaHd46shytiyngaEiBlm/RiCAuEzXjoVj3IqBs8jLQ1uzewiKJtue84HrKWe
VGyrzNpM/cM+ASrwfxvS9LBn7WRunHeX/oAGAxOONOiaSzcyYdiI5U3FgI0XCMxo
KiutwN9oT4IP9HzBKSrs7qklE2AjPmdsb/8cGrGjz8ZNyzj/A3otlm1TgB8CE667
VlaEzpvejgFIO9RrcYU4XNgFVnlh0akewNDB81VyWFyywcMeYrbn+0qc6kt/krO2
tngbmEVg2LT/1oiaahdO+8Qo97DUym3qTH8EWo+aNBPAaLgqmC/5elNThl51GyUD
OKYIeAejTGEMi7v3UgZnW0cAYE/LbFC2YTl/NQPRk+BJAHKCPa6AbDb7eJW8y/oH
Nwjz2233cl7gM6fnjTjuWfBz7JCxdnHxSOb6349V+0udqHViCzQfLwxza7Wi65pt
i8eKlZN0kmBaMy4uVLRjFhyvRn2hKf3slx1mUjfgPWCmd+FIbNGswXev1juv4OjX
8Pqo6H9pHJo0WL2pWyq6Js3OAMZaxg2g090CEw0c/PFvEdWEGpdhROToFmlC8dVS
ZxtXhFXLepF4IwvNXiDkpjKaiHre4oQtne2Bvp8hgkzuBedd4SjY+gkMnLpfDkHs
AU1krme16M73eeqHAbqGddHSEG7/4uKG6jMhiGuxhPbqO/4Z3jG322EFY+JLilyT
0+Sybff4SG4qRQnW4gqqog1rd352NsU78LVVORv+rvWuRgDPllg1VEaAMWQLaybn
VV+Ak4UNfcoTKyGK239FgxVs+aFeUj5JWo+RweOtClvMi1gTiWHv8HXLHWLBeeFt
HUAuDwW4Mwf44Z3CxMe7y2XRjxt4zDeUvL9s3VqZ073wgKQ6X1kz8zsAo+ybuX80
INb71AL6IZmBWIOradQhRR+zjZ01C6fLdY/h/nSguy+970/t/RUtAyCW5ztFsV88
/C1EBGC9lQMEvP48KdgfneIHNhwEvSUdKq0hpgBpMOQLcX3YaP1JuTFUMzQR28EX
zEMBMuKJZHXtSNmSJTCpvvQJlC68s3beBl6JCm9nOO0KeeIVA5LfZUfbk8cgNRoN
tlhJw9y+xww2hu5NiExxNg9MQyZ6JAx2DkXfG1BJUMOA2KcbK/IkK/kvh2ebYJIC
ZtEpQFTF+os2QoP1YXN5Oz2eUdv+C8gl6CYg8KSYl/PrEurA3ZEB/zNHMwHnX2WS
w7YS+7BB0eN6Beg7LaS0FPJgzUYHjF0RqnH7WMGnXeeHmIANtKw1aSCiMtuuruty
QWJ75Ah6zKgNZCLBuhQH7z7/riShsMUJHd92sizEuxHw/XQjDhBQuuu/tExLWUFD
BkI8dkFlUg5ep2G/1TH3wD9INZKqsUhKM6k81IqckCLOynrQe6Zx9zxLBIQnoxd4
GdCMUjQzuegTidfLl4DvKI5793l3XDSqyn5QNlLvWJCcqFeHp5omnmesJ8TEpXO0
Wn4HI31tIMy9r8qB5f7v39mhEzNveE20Kk58aZjigdKF+H1IJBQte6/oO/ojmBuC
Q5rmkvEw36LSODCUOa5d7MBpiBOplibKqtDffEdA21MWWrJDYI0N0Tqor6ZOudVF
r0+jPfvsg1BxR/eaCxxnXU9W+d0Hn4WQO+BP8nBd2szeEYxo/ecbnthJbNfY+oZ9
DLJVKCSz9yyVtOef1RHBb5d7rqGhxmUViDkCSFHwuk0IAb7eQeg3inYUHgLb0GvY
mNZCXCY7fSMAklU0Qegy4xC5HUOFYqnRxsIKdSGuE30rQqkZ2tT8JvVhfi9JeEVF
OaBD/lAXrPg1smjsVQjlrfJxpHCr8kRkABhaN05B7k/EEWm5sbojQcoRO5A7vzqk
Ck0aEtasvqctnXRGXys40JGMLFfxA6b2d1BritcLAf+80NW/20aA93ahvQV8RCF6
igv+gKRpqfFLC8Kbx1EQmHFjKWgkfU/26V42s1Fq0TmVle36iT9vLlnXJ/zBuTPZ
8nR4WqLl3mOKnxqw8PtlczzK/dLtFCpJ4jGdG7H26RpYzrNK/rQ0cKRe/fs/PQSR
QgWtxcfpxyK4x98MYDmTi2+IoNYQkOevLBOvLHoUScYOToJ6uv0dMVdnUEDOb0cM
DOqizUW7e8DGK3hUb5I/Hccx2sEFIX7czzU2xjzrTFOY2Wt1DF6hIAY237dw2lpJ
OxP/1y9pRmUfBZYt8m+BHR9mPziFyedxkwYaANW9x4hFmeIv6FFA0rt6bCdMFsO/
kslSEiDdxlAdok7Fdq1eYCb1IN3qV7h+jJGF1AeANX4RPM0gUKAkR8zoV2KaCQ9k
TsQoKZ7FPUqPO+cw5moGSTixYLTKlgAHPzkX9lmHXhL9OCYl1e8bkp7mZZ2lpLas
1STkMIgdgNdFT9yJSKZlspwR7IpQW2H69SolqJkjjZoRHDKskZyHC13ylSvv2S5Y
LTFsGmoE3EsmUQLoVLD3LyJMEw635mb+45HYGM0NpnhUU7rS+fp8owIzKGSDPhkT
qoQM5X8HW0Q38Rx/CH5ee5hPlmjo+Dm1CRa+HykCLiaZe5r3UAW9gPJedPKi2TCh
ynv4h5HMtfkDIkl327Ng0urTWGR8VRqfr9iIJPQ6oxWadMknPdfzfpnlmq2UH/iL
dkvwCrqqmpVmwNOlGw8c3es2j1B81R4Q/HOs/LKJ6EGplY8l6lMZ2+iwB13T8sw6
ryxdmOX6gx5yaiZoTtBTJ2KI+gGeKkoLsDiY2yIaO543R2xL732nCUEXoQyqXrGi
hSIUaVnrFOVjDgkAYZE+X/6pnr8F0wQ31qJ8CQMUNUxlLKOFX0W0xT8Y21ob5rZ6
gpmitqw4xraHB2HucqdccQJvxJFNkrRbh7dHfv4RRhwzG0Zk8uCIQI+yXxTYnmTl
0bFTQT4vrJLYJUQWPpsjYm3pLYW8gh1Or/9kjrrXTqzk7RDdYefqzdr/unstS3E+
5JdE4s82frUgr9077aUCaVKVWMeFivYv0xzBqCeH4YRdpVea+H9klK/+SEziTL0J
zWQDNv9ijfYRPA5MgEnkKxHb0vlzQBFZ/49xE2O36DRoZV3ypG1zvbrS/ontf0CC
s+ium/Cm+Bw5Hp5+RItYBWPy9PYjAVxQtwAM8lD5FPYgu6kfIbmtlHgNacgGtrq/
QqTCQFwP1aUU5D0HRHVwYdBJ7fVgpKf+HNksZX7rHPfglzGfeT8YfNjBBCZjPFKo
LdjnvFc4piBh9ktaP1zk1JnyPyeJ1Zec04apqKZXpd2Zn+Pd5vj3L84g+vpj9OVB
M2jzYSBxL0G6v6zsCOeYuYUtfFkGhzBATuMtA/6DZR5TQeP5sSdGa1o+ful/t/mx
J1gbC7LX2OKTtRA8WLHaOvu4waUY0Eqo0RZKPLOQObdCGonJpWTzHqKXt/ZEfdQ/
i3llVy6GgV2EGlJMfyCdWdHnjLP2JKAStsPgJWvgyCHq2rgXJ+BHmNguQSv51GvS
egh2jne/tJNpWOFWuOJsktHtqtqHcwVOqbdJuutJoCgE1vEdoHdT8dExJA2K5a9K
b43/snaNvN8NB/Rp1XncZ7BggG2NE0hT8zWIbAfFUbcD85EXyhKCzBZ1xeMIR91q
ldS5uVxqarTpfZ8oC+Mxa/gzY3F9eFvrDuPOLo7bqPM0jsx8hKQ1kZGMTaMbAP8b
tksCxFN9dpPKGgIZhURDq7/7fXEdl0+Rn2ot6JQap3zR8D2Qb4nmbzicakOIZmxa
ub6sN9Nz26jFIk15ngRUJOimp83nkNSFH+YpsUnPG4Dm40IgxKitLvAQWpg+i0rD
r6wW5MbzEd8h8g89kYH2hEPaF/8vToVxhnjh1D7fGIAr5kkq7cTyi6Yco8aSXzAi
a3oK74mWdjNx03ugQ/Xl/En5lkE/KsIeWWauMqHHKSotRlypl04DUJRUrNsycwP+
WmqAXEBgcu0WPmpYiWUd4Wk3KTIzIH0mR9vpwjdS5qkGFYeWZiV26k5r3FYJz5JJ
aW7IiYiDsGsl8P60/l3PDwcWIYqSq074n3ox/OxSWvO/BUoeK2qKnJ1dOWfoSRfY
PYCDuP4dLOTDpTLCR3jD4Jd//hmIzafQrGbWGLMthRi+sYxlWiMiEeaywmPeomuG
taFtz13HkJFyV5c3kJcwBYEa4JhCGtOazDlXgHiw9ZAMyoFHXkSQggq1KA/h/XEe
ffvRkGLbuv2SbEVmTCdWQW7qtvGLTgJvJIDeEppB4PdW5ZzEX0dyLKnXMHFA5P6e
WfJdFh6u+7VYTnELyPTvcyn5jW0exmc+htZrhzMct7hkl+qDL9ikKHdvpIe6ZgLj
t6qvjG0L4yKN4xL35sBNeA+dj8FGBbsNVlW5IsQAxGwGiZVmuuo/37dwqVMizuu4
VLOjDATLRxGc81wHkm9+JYst3jmss92xMaXebKVVIqCYn/mxPi/59g90WFQiC+c3
p1V9fhuQmXHE9hQDxdygM7yOEUeHyCde93x+ectqrfwVX+imRtm0ay7s7OEnsPn8
xQZqsww43AveZgf6JgcDRCev2EL7tOjW4rs249NtFvPZV9au7B72kIO2lFIfkKuz
dKMa1grwE4D6DfG78OClU/Es1TpTH1SgQBMXK7vvGaxeQUwIkV9zIWvfHY0oLsYM
HBL2hrh9CtQja4EeHDoxwGCUOXi1GRtRY2VAT7oni3yEFwc0jB0FUKrdYLnfgQnh
Rnv1P0n6N88pFNQtM4RAST+M9WpRRo3jOYF6kH51Zg1VTFkHsHCP8ItsW9hWggrn
lR+Ab4xcH+8qq0bri7cYYsjV8n3sCo1EvACmPDj95cotWqMPaXUCv2AWOYh2YTof
dV0xx0adFXbXOzLi8taWCiY24eqBaxA6NRagyyWNUrjfjE+4PkyTljvTvtXYvkFR
XGzYNSgMiIiKx93d3pM/ieMkUI4UrBdl/lGM/CostHImc8izgNcHPmFxqHnrsFyw
rB2X5cBp5fzI1PNeOmlcBMnxjQv6YYFEva1BXO952bUYpiHmPKvAt33FY4QQM2Zt
lq/+8tz1iIYJuMxGpNxrtR+tJX86LW2o6Mdgwx3/EKqdGcKOyfOv+eY48HgvbT20
gFoI2mHE46UUirwLvQRUWFO5x/ujJ1Cr0crz9yLU53HDytcstdTyLtnfNFGF1ZH/
eB7p4+xLNRoIoXezd+hm1bvhhjKCrTKsVtj7yxq556eOA85jzQC8X7s6mfJTJiXj
98mgmyKVaPrmHkZoggXpVJ92dpnjbTrK3/FQtZ0kKw4idhkkRNXMXqw1CczzlQq/
+dSTXJgApbk6+xw/fY6B2x0mU6/zSSL6lxvvdPT8ZLgfeXnbCehTS/Lq2dMEPupP
NU4HzMyiQ3pICP9YYTCOstYWxXXxNjfc6daK9ma5XjDObxaIl1sw3jt4llzSCqC1
u3vplnP0tJz4FQZY3Dj6vtA0OlsFzQeEZonH3TDSvHrY2M2TCV72AkS4v2o9PEZ3
8AQi0oeu9HQhkTEbTfwJ2yXIrdbaEPUiU+FuxPH7iiUHho/URxG/tUzx9ZqLmd0q
rRy+EvMIit9NyAGDs9lluvwLLXqzBwkGEugD4F2Q8Tes4Bi74w1BIMUjS23vJeht
+WOhv0Xl0gm7kyKlxgFHOt8PSJJ6dsh/kgf9PkMPoN2ida7XzB0lmpDF5vE/0cb6
9qNcYlcNqx3cVIOPXNQhaGVYOsy8RMpY/uNsajxJQedJUbsyVKbnvNjEDoHmnzdu
5wD0a3kjJkAnOZkhocXEygAt167qWXbqJPUQ9mb/EoAOx7mxYv+1Cn5O4yLRYKS3
ELTtyFDUcxaDik1iv7Q3l0ofAatkdRvGLskZeq+MDBXDLqEYqqsWjLmA/HOfaPbX
KTVgO/Bp/WkHySKrlkwgixvw5/GYKWkSl6o4v+OppWf+2Y8sbGBQ10sDRsm72CVi
zWmBKM/flTxWAW10C9uqR+dRrliv/HIkgjCMyVWtTgNsPYusFf2m6h6F5ouaXOsG
Fk+E3PiFMua59BenAb/RSNauaY9yQozgicyDfoYhy/nq/a+AYs2j7h+igbFxZO1J
5XN6P6Wk7Bbcviv5BqJqTlFXSyfDkw1NIIAWNaZMXbNZ3zc2lG32JGbjS5WvukNp
YKJ9FWOseS6DVf+P1LdEeQoeYWwqqUl/r06H2sf996MutJ+ehz/Fb+CNVksoGWMG
tol4vISWhnFrn3y5dQapX56K4n5CwxCt8nSWLTrJ8riVL2DITY+/Gr5CWq4Dovvl
R8yv3J7miFJ2RmrFCPBBqMia0vkOJ4qOrKkrhG/H085Ftlqq7IKpVH8TDsV4p6/1
i3VTADdluwPdXhEvoX7TSRnDr/munHKlDQZSMBz1+2TD4ahMn7/07NhSGXe0N6xa
0BD32Bus/P3u1N5wwQ1OnIyuj+EemmUnZTFJ91opL1ejEjFcG43C6kkEsaMfqY8g
Jjavz19YS7Bg+NNL9URfQHMNtuu2BgR/b0zStSVo/vLNc1q8HezxGrr2VMI6Hpko
zA0mvMlQS/9lhSQP2NC8nP26yl31YhXSOBgO5ZhfEl2EzFhKuyebwWE5d9pRpZF1
Vlt6zZ+NMvQperFRXlvth0U+Qsa3ueKfCUn64ywqj4++fPEPvPSbqpdQnX5moVfx
QrKtr7dxJkyjPOznkTUmhEPAGWyEoz3jYcAkeyA+7Vogm6YQMtFy0rUiLjmxDnea
3wgJx9iO3vIgWmP2J9tZd78yGNyQ48Emb74ZSf8yOWuUe8H29mkfDEbGXr+QHTVa
6DVaBVJ6Aq0Am0QTO4VlvCebpU9ohyrlqzmSm+QefhnU0O6oDrKYQMOudME2gzYR
Um6c0pwLYS8CgwPo2vlWe+1K5F/x0tz3UQwpJzbBbA4eBq0bV1mlqoytF0F9YLTO
9DoWKY6Ffgr9ucLyXMbNSLwDAGoTd3/AKqxACUl8KnTRWVUbUHFD24Xd5xDDkG/q
iLEZu0QPftrVjEZJxMw49rSwwdGyPI9qC/lpKouyBnRIuKvLEh/gLT1i1m4BRgRo
U8zc55/Xy+zZtooWwmRK+jjNcdLePXeeIwYdRRTI186oGcfR01sI+cc8BY4CMkul
NX2wzvmO/9BcL0KEnz8NuaoMuxUJ/hjGU548lu5jOLuUdKLrEfGwnSFYnW6586zk
20Z114i7i7/Vz8qDG/1ZHOpoZiJLBI1skiJHxuW54qtuRx/N/xp9fguep6t4ITJ6
4b15FHbY6trq1CZ73ARKqAP9UVaU3xSWIJzgIIQzm4Qr39wkmu0SFIlRY5Sgz02X
Uw7aytkFU65eJIxAiRpIaMVKlAr2PUHYMAFe/XhBjw15KNbnYBrAIo4I4dik7+2H
gA3/b3KuvT4M8u3bBczrjfNEloH4S7ZKx4Y7wU8kXuZoCgjR6Rzdukso74uIsRfC
o4CNqB6OJgRFGBd7ZCFbBqnCEIgWDgbgKrZMh/laKF0lXuWXRYFb+y+rM265FrRH
+2jDws4boFcS2WDLFzvTqbIjT6XHllfOqs2S7Krd6z5Vb5yCX3rdRj/BPDEIaDqz
s3bzG11jQVeXKYVVf16zsMX8UvXaW23vG+SbU0lXpH+59IN0oLhieCGZawdpnZX1
4bnYhOqaVdxn5c8AeKMQOIALqlZqSgN0BUsNurjmyKNty0WPiqftIUHYBM7CJ/sN
ar5/D7EqPaTJphXliOuAteJYCDr84/ImsqYe2KAjNspcWNh++ElBxk+ijucigpXO
VQ6dq+MEFjFFXQ+N67zw8GIVOegn7pdXS99AiJFVXYuPUyt5mqsOtmSjItXM4bRu
O5a9OWYgpGfIO1YyNQ9Hvwd2V6T/9SPTgCnF533KjQ+EJvkOyBSnAOY4Ph/o5Ga+
Z0ev1H0DuqbmfihKB+1rUdLxSm5qCGbdBhofV8JjTTYjUhkVQMrwKqLnrO4JeUg7
+Es5S0lDfDmxj9BBtpmdjriJKtaPsKP8zIOHzFucCymh/7xraOmnmWzrrWnhx83i
jyyzUGzrMb3EClXygepCDwVxAMTADrB7tObGnnEHjE2k7AAij7s8PCf7G1xBrva6
4gh8YUqS6tnriptFtV2Jh1HKKqkWtwLFmbjKI57pUAYf7mOHtwLi16EhEs1s1TOe
/6mfDdXBYK63Q5Utb6kI5VnesjfCwFN8+C2063Kx56nzmI7eAdMhTARy4LyuJ80p
/p/NqEeVum7zJ+8rrr7sKZ2cBelertPVFtAnaYXPbVHIUmsokCMGDMoQUKgq8+lD
WPVvpP6rEw9+cJa6tbs32uVFqCVaFnSfsUzfRGXXNpAEx+Y2UiL9DHzri7+MsHkz
9K9fZ5HqW6jYiF6vuQLkj7th8NbaGFUEMwfsnPH9myeOBmtqUAVA7vTx7z+f4M21
FGskna+9p3OCJgRVD3dT1xDNpkkXxa9P3zr85tJwouJYX206rKubUvnTcxjx36oO
C3XMbwaBILGqriPvqoaIsHnBiiYZxj/EfQo9IN4zeN4d/NVIsLITMZJ1t3YcjfrS
sdVLiZMkadClckh7l4Z0fCW8cLIhQQvWBlIFLkIj2tawBRx8UaIF4dBLHLxYkAs8
WbWGASViEnQosXeBZWfKLJj0GmoZMWoyr+zkGx7QGho0zT1UoaMowzxyNKAd9qs4
qRO7VHVGGOvyAr41tGspbwRJh9X/mRnS4BQmxf52VpHh9DLCKSHMffoetQO2L6Tt
1gcPZ1lku1RzRaMaOXPGoMciRkLJ7kyGj/FCTuKdqgzOgXe8nd0lFCtQIPr8uAG0
j9FcHZj/3QmzBCWDdaHNvPoZP+03RngchxHasToKBLwduClfJjqbZIdgtdBkDKUB
hXBhEIEWq3PvrOqx2rtS5DS9oztxnZFdos+dKp/V7/J/t6Tvh4aRqm9t+42B2ZmH
Vh8V8oc+VwUZ/0gJ3qa4lNUcbuUf6W3k4KlXPPCFJXl1p/ZTJFut7H3v3KpnBGDm
23L9bfbWftLbV5y/mBFOZ6kkq1x1V66G3rcTUDqsJvfEDULgnRj9r+qQjAYGd35m
lPc0kcybY92DK9icDVyNXtmIr8BqKP8N+1MovGs1FenzyeqOFVQlgaA3fV27dZ/Z
5Jsg/xNiFl1AmYuEFX3MQiuuSH5WwkiPlk3trAHrgdZKLjZxaqNVH1137aO13lq1
zVS1bajfYDVmrqVAywKhyd3xatzt5rhZRk5Gu6Tsgik0dDMV89l9QGguGseUSGfo
dOnNa+so6KmbKi9vn7sPb4+SyRdlhpmYPQGKseYkxCCB6F0GyEu9eRTEt8jkqmI4
JPaLLENS1WoHOpQZDe6Q83/OpJ5yNOGWIg0M+enHXxM1QPH0silsOwQKNPP3+zF2
/Q1nO5+lv4QA9LbwDMkGn2j85T3N/uPw6sjzOQgX0lHV1hofVukurpZeIqyMzWPY
6WcwGkfKQ73CQgm9DlLTfgVgboN8ft4O2vGQQmLwbHfAZlKQ2h8fxHZqIvjXno19
qY7fUrMekASb/I6uEdNJ35dO3h010teIyHO3YtFLLUBL0yrHN4pLWzLxlhtVn436
Jnz5Bhs1jVsTXl2UCf65osceyw5nJTZ2+dj2DKDTOqt+F1ExhWIYPLgBO6WKnwDE
43uzgEeZy6RihVr8mKzSe12cr+29FZaKYrOr0YjezskPzmmZJq9rJClw/wA9Kkvy
`protect END_PROTECTED
