`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v0I8V+tklX+Vse8WZtv0YkLk53VJqv33YyVULdL1H4927bg6ObimDPiAgXc5hraq
4px6x598rkXlkwOZlGdtwkeIFIYGwZC9O/FN6zZQnxOq5UzUdcmHwcEaIRCuiaRS
rn+4Kf+HwuNsdZX2p/cw2uz9IFB4nSrXiZvu6256Y0s6Wo29ncj9+Ak/m2mnkEWH
p/ek474d6fVBGxGoSfJR8EL0c3gOwITNuV5tUGlrDlrrwuMFjlcnLo5KbDj51IhK
wETSJ7gYDFCGF/4w8b1iKUTh3hrhbiZEcBdzI7/XO00wSheapgm0dx1i6inBYorU
puCqOShl9xEe0Xd0Qeglr76DvrrIVKXdi8+ktBwVpngt/lIYr7zDnk1klHsi7NfR
13WgSbMJPTc2YqhWc1P4zc9cuecmigpLMVFguFcwHB9TD+HQEjHpr99nOZwCtrp3
WxPy7Qwf55pqXpiGaHL5t8qF8PQQABJ7QSJixL0/OTNE2xndKDR6c7xPgiksL/jI
Jq6ZCHiJIm3PUEkeUxPiCYkA0XxSqDtxNTQbmPbC/gVITEJuUtsMoaXKobC57ayU
Fe9mr1XxcNGwOOPd/IKkzfGeLzBYUEhyu6nGALm69MdkbOilXgBmqXmdN6Iw93dI
to4tDTlRtM123xZq4dXgvbpjI+LsH9gjdy+PMECz/PLvS9KgmivwzvMvMgcgdNQh
0HXa6Bg0BDYtmDvKJAnhU1LwooIYNlafBgXNvF2QCJCpb2j6UeEttcIWDg8HqBik
uje39kK56tMyitmWYTSyLw2h//e3Qe8HKlJfI8QoEpYBdJtpXISQQ6xczeTkzvSL
bDT2f2UigTTPSeCqQtMKoJDY6ZtAAuVyeXchuH4ImK8XFn+sK6MdPDCPCFUeEOCD
UQpoebFwDzT9wShRpoYxSdmHRe21Ny2OeDSlBIDvrR5IZxeZ165fLNAmXnNVSQIQ
kZ/UR16W9iMsWJhpoVR4XQ/QHnmg6ig0caRsCJOEfdN5SlS622jfH47lpzW196rQ
Q52JqQdt1iixf7mRCPOwg1m4zkfb+MsTzP+9btXxRb08Yl9pOt9p4KuxNSc7sVwO
rVz0QXne6f1+eCrwJIcpYkbTteAQg0BMz0uo4w4Yb+OlIVfJD21NvitT5rzEBRrV
2i5iRAQaOjcj38b9DQAp2kgSv+/LHHwQOdSBpBhqa858QMVp0BbqZpTF7FIcfBji
XSByiL95Ag6sKs0dmCPzcknKRwVlZMu4YaVyRO5oE2QZ06Krz2hpojaBQwQWWZ/v
KduZWR9xJ9JeUVSP9CCcNcnX+rFKNIFPqZI8ciSpUNPQW/gq2NRR1VoPSjo8r2t5
J/DiaQaKzUM2XAkIoe4gnDsJVylVypvCKMD5XthIwYW6c0Y/UvGg6thb1YozZVY5
2E7rsb8dnQt9979tA020oqn3+xF61RlfGuQIDuy24PR2bEkq0cKROh/gXXxhgYUE
dXSexcn5DGUh+eCAG5FFuHYu94a8qwrssgiSH9/xxkZmpl5La0lsFnqjg85gp8D4
IhqGKCG73yNoL1aEwkgZLxOuyrJtKahGwIkArNwPc+d/mGolKL7GWNaAOQjJT0Gu
9EgXgOIl/164qiJbjpJo8xVPuQWYuWAJUiUTLaG76/OOVdacTgttQp6oyLGQ1/jh
e6YbokpwGq4iY43Qxf4MbA==
`protect END_PROTECTED
