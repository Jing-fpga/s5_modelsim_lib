`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2WWDgQfoOJXY0G9DZ+ehkhDVhRH3qwL0rhyM67+pLJ9zcKvzz2d9nyq7mhcXygHJ
6G/C4/a3ceJPxdRFU8UvuX9pbsjV5Knk15Yodj1bmuXLkDQEHvlY8YPilWAQ8QhE
Vnrg99dcNKCdkhn+UX5pQFkwpe3u+E8IFAtjpcY/b+SqJddLYnO1ZaaOYeFaGel8
/UsJCdOFebQ2ypTYu0lvdHHMOVuT03EbAVKILdFSBm6oWygTHER35y0gxoobbMkM
x6+YW0am+MBh4ZjtS2hkkNY/KVVh73m1BtImG2oAWvYvwd0gAFqIdAVkC9bFKXtD
Jl749yS9iZIbft5KU3WVnPH1ZEWqDH5FVeMjcNyHOVjzc2p4EhDKeQvOAn97WRNf
cdrS5KUGMZoun5WnaGPpYBD9iYKUqE2kU7kflPJb3OHgXCX70QJCtbh/q4gIYYvJ
BeegT5eSaU5l+CZxJgDJXwpPFY4cNHi7r357q1zhOMoVJlsZj6L8zmN35KRJv7kL
pWECLJeymawy7YDQxq2p9ZnJktjfT95aucdkbdZKwP1WZDHIMYgCExq8k0yaeYhK
r7bgcLfud3dqvrEWCSxnbeZVkRA3kYtI98m4hrBJ/sTjT5Ad1zZa1DDx4ssDFow7
q06+IR7iTl9LjNgSsNEL24rpmXPK2svllpuOSKMHyu+li0izSFcalM4eeqAXldP4
uGIm5P44Rd9G+vu0uq+zYF11xW1S/Sc7zB4NVFudk3PsxZTBD7n+DfAVU5FxU77h
6o9jwIUXgw7oIyehCTpk9VYz/FlCp9ZQtFFXK0qwH1B5QTtkhkFY1Nrspofb0Cl3
87FcUgZSEsvqUPdWvLxCSEUx7N7bw4fjiiLXJQBiliu15X1ugSRmFGGx9PXX/jLg
JhfFe9g0P4cSZobQLxzcRrJ249SaBHHGQ05tCFq+b2gQIVcONOxNA384QKNPchn8
udk8yxHNAyZwLRHCPCvsZPV2Ia4HBEGFrZceWu5eNAlrcIeQBFACIhaKxckMx2r3
0v+V4TF/brU2AEpVyXGxE0A9VHiXYJhwcKTKi2pqsxgS/WvhdCofT0hA+ilCQwHV
fzqv/JGRLgB2rPFw3Ys/Cz05l/xzpT6dzuU9ljLZqN8Ta0Ep/9pDP4lUv8VeOkaM
mNz6JzvtmKEYfQ1MK9H6kK7FOihkocRN6/EkYN14eEbu8QDtRcci2v9XmZL9q3Iy
1jacqdpwMpQAMUSHF7UdWn+VkjxZiSipctimVqfmF9SAEYxNQsjriiwjqLUbgSGw
ZZrndATYzucx3tHm8JIbNi0rE4iycBxNCx2Zn6YLb85IPUd8MQyrJ8NJQwGtcjNZ
HACDVzli8VZ3RSIPOYf+SQin9bFGudD/aQ0tlcobXxf3FxyWOw5d8StiIcyRI3aH
rOGrmIqKPUfrio2cvPqKQHTb9or6EQae9AEz7RoQ/soenKa/F9RwE5qtkL96FiKx
FjpI+qWJG4UxGlaQBnvyTDYgc5rI1DL3zsDbRLkxreBTk3co5YIFwNiWRRm00OCv
tny0jdOLIl4hBGWuqy6tsRzVK7OlxuF32VopSfaewuTqDRE3JAgCp+posQpyxrl3
NfFCLnWXBX11DJGYycmx2EzM3GLgl/5kbTrnCB/rQmY6sMtwGA32fJAPKrT4xwxS
dWjZRPqTv6KgnfbzICQB5pdShtm3vlIb+lIdGZdO4hRhEjY9U3ey7RhNFSYSI04d
TzXXGnbpkRwUhCulJmWwE3Z9vgG1PmJ5sanJ1c7al6z/AhOniBKgtuSOii4lq+bs
ItOrDw7tRV/NVCM+2irkcxbmKLIOaV5NlUpMDLEd7JlcPznQ7cClbqcyMSJ2xOrK
+6eYohdkXHKQYAZVGXwzGHBGb4dDIjzTKGUOoNtnCQcUerhX0EK8l52XtuEbNxUX
Iwwrh2VRDeB9yNfRmp7144HhExKVPcyV1dVlo3onaOihTHpIUoHyikfsjW0M41I2
SE7hSqL4ZJ0+Qvw63A7UDzCxn37tQY1tZ6ENbCtwoPHvSWQqjNv4SEpDxrN4p9fe
svwjFhY6l9RpMWEWaxWQEc/ylSGHDl+E06wkWOqFQfqnIN4Wp88UKgqDUQX0q4U0
nCIwf3Xe1eBpEnhSI6onjBu+yiflD5hEnJTVbJHz1u0kVPuL3aBszGruXgZAkMTa
nvXxJBg/NZTVSgHn0gOhsbL4FEnvxU4lmCV9sC5nB3d5xDURDbrP3a0rM/Ed24yi
n5klLEn6zNdessWotUcL373WHtfWP2Dn/Uy6tPNauyvMGHuAJsfHUMH6n/PQiAXr
WLcpCuwX7fDQWHNxgSXia/rHWQy0RZPAMSoPxsldsMUTa2HT8Yvl18Sg/67qOS5Y
l4jQ3G2ufcD7qPwizIOPH4FMe5dkWYvIVl3RXsAbKTMfcLN5561P9Pz7fMCNzJgp
pO0wb1K08+78DkJvFapz6HxZqQmt5xtM33GA5DupR4h5YODTqw+XV4dhw95F11wc
ww1dIIoTwEN3ndFwAYxp4A0bc9DgBiYP+fAxUt72Be9k/t0elUwLcz+who2TZwmE
0RjIZhy5lD+9iu8PhiWVghW6ER19RzRG2p0JhCdaa9AVL4l+Nz6cTC9GtMK+kPyt
QFXSVpDGj7DCfWX/SpgCLedWTsGmUbF3CcXSNvuuAyF6zjOjPE0L2TtDPPx6gVgq
Sn9Pw0KTdLIxN3SBSnxV+0cKoUbR0Lz1+he7mw/GcwGRjlAiWdEZks8qLyUezM6T
rcoNmG7L9ssU4sidoTtjs313cp0qgq6ck9yF+a5Flq5gSkb7WTPaATC7TL9IvArR
PBZdzOZFv6VzbdJPWVII7DNIz6zQQr9iauWxAkE3NnNIaz3P/9v+j+OnSggS8ojs
LOYOfT/aXYV/nlqSYanJnlwBnsQSRTBvpFerbkGdf0nbofkBZaq+3dm1Ny1EnSHI
5csf/Qto+X7omCH25UHtGEtBomN00JbFw7ujxYO0w8/tCyETBlREUReT/beCKBmM
NKT87zppvSDNpqsQGxNKrpsLRNYxM4ZJoJn5FBwxu9bJhSk6kV7hFosq+As8AYkV
zXEj8q+T03bzEeZsCJWT+6cLI0vT26S3B60xg3+dfMy8rRQv97OnyRkx3e7nSJkt
/KFyA6TuVbGhy9/ECVErM0hH65RNHddXrsjI59ptbaDtdVsgL/jJ2b5winGFD6gh
awhZFZbGBLLiZKwMX6HK15ZkEWDPYkwkTamn4L/U3ymNJLrRLqLDX7WJhN4zWzvh
ePtJzeD8RLTsnlwIRw5szC4oCSl8enuctR+X3LhV6XpW3EdV4Y5COssVyi+64Ujz
DdafKMO1R83RFNcXTjlcBh/QAuHXJ7LhYScV1mCHf6quCynDcz6284D1nS3L2kDO
nDJACsLB9klJWOrpmd/kncvuMVYlrE7Lx872J6Qom7dwEHzQVzvnHqz7TWlVigEo
e5I0KAcOI9URN1NoOGeF533oPTGaKQGJCxXFHt+WTwjXc7vL2h4OQnwSL/NYtDuA
+m299JdV7l+8c9tzNYYf1dA83q60Imyqr7OCtz1Pxssh0+ltV/x1l1wma6YbMa1b
YKYnFuhFdO2SdW5ydOOkTrr3+y/4QoUp1b79EEUxwyD1kqCgYtsZkEXHIgrFAU5v
/MXKlAZDOLioEfRxdyPVe1KSWIfrwIZP8zMQzXOqtG/b5KeWy3lp3kZHFinPAsAU
4eLy983fJi55cjEojmz3nuyjt7/I0Y/uZa93OqSwDavU9yTjVuPGjzDg0SYDgKaC
cRBO3Fzwa+wKRsEtx5TzAd5muCRnG4hsnLGgIxHEGtNCtLNTSHPEiNHxvMZQBLcB
ZEHE5dXe8NNLrFfn2a7Am151Zy2PvNcpc3GydSalOgWQbXGsyHaUC03nKm/Ujku2
oHXDJ63T7MVbGDzUKnxjJRi8FvFs9qZGrTWnOAEf2Jz8cTO0xqX8exygbkVCTbUQ
t762fiFd8nH5nE08s+guTEcQcugrafSjHaTsZSgCtPcwrRigBylaQgBvyixmbJ0o
/A/jQQBqgJLtcMIJUeGaYyJn1aXYNTMiNteal3wNh3DepxQtLzK5EkJ56KzsPL1x
Pr+HYmmYlvBIGb3d4kq4VmZs2no+ktCTPfqZuqQL3bOKPRjKjGXhZJEp4Yzf4DfO
/6YNKTSBOzFaYq2/DzQJunXEiicA2rD9xhqToDLZukx2WaJRuFN1/SRrbmUEWJWj
afs5O3z9YHU1PXnIhX4trmh6IN1WkQE5rW71rwNSXpbpbKSWnIIMesYDJ86wRRJp
8Er8DvZDLsDGPndZ7zg1Mr7SevdR24BdZBGp8cDgZPIkq8NRpj2goRKRMROaXOiO
t/jJGTfCbNNYr5DAPNJcRtkWnWGWnPsCqaFw/HiYVH06fX6/lqTIHCY9U5uQVeQI
Ullm2sSfyhVN4cP61ZSVEN4GzUPs6teeXkqcF6KfsD3cH1fYWNyvsivPezNSOJmK
nfE1X6Ybja0U8Jxmh3LUL0xl78yBxBNTpKeCbgOnnl1LjXISkjtlPaKUbYTX/1IJ
SnZZoA1eQeQp3tfK5Ik+lTyLZ17J5wujIc66tdmIEbWe2Ngg5BjNJFrf3VLSrAMG
8qcf647RQjAiBhB3niDvg3oKNBXqOee5+DB1lQQzKUOxYZgikDqMsvSxbRyWCs+H
f+daDg967YHH727bb4zBSjZ+0Xvwf1u3ATUKQiRLYKPxabMBLTjCCHkgFLbmZ3WF
ks92EN2m4y8FTjRYY9k9dBfB59WNMExPMPUrKckIqSdpc6ueZBGJGzCg13vW+hai
UKw3SSBcG95tfrrorLnyFLVDuAiGUE3tkZaSK3rAuIDT9BedrJYYkH19dM2yKjyi
n9zAszTmNvH9uHjqYHvuRBHw+tX7E18K/9fcfUs3pSCVBlaVAOlo6qLYbi7Vx3cE
de5v+SqQZlAcAmybiyn3UOA4m6Sx2SALlI8mvsXp9AoV4nM0yUq097LIez1BNy4C
5YfeVbtbXLf+rZUIv2XVKBa1bqfCtFtk1YvIjyVBeJi1FdnXZkVZzCf9WQR3JKkQ
bXx/4vIdlomznMSM8pkm8MNfy7gBqdq40iDdY/JEJUthxO0FAM4+ANVIVOMP3AiF
NxoG1bmk/g8Wp9IuQIgQj8SOjmTCHNBhxOnZcVxVhdP4FJZXWBxzG74ClqFY4bWF
LETEE7kQw5RyNW8c1Un/ZqCvkhAIqGf1UlghEX4flPkA0YZTofB03kRJnE85D/yF
HKKKT+TyeoQQlInJPzxA3MWpfV33ndLnmAhMF3usT9q9G1y5ikCsg3KbqJ8Gd4/L
W62Nf5ZW9j2nOZO2Q6+AFA4VdlNLUYdexG23DgIGmNYOQsGdp5aFYOfOGhJFJlcl
LjvOEM0Ml6zASA9Panp/L2NkQ13+MT7lnsaGJHc7pQ6Fb/kZIhllyWJc7h3XVhNi
Hgu2Qsk9/DMjjIGzQmxJf5yVyYzJhLkYfDu947uMWlX27yjAI8Yk40K//0OsRRfu
glnEvJVM6n+s4q91pk+vdfKFUxq0ead39+7o4plwFw24rXnibspmUvt3Ccl18oHu
DFTr8tjy/Do3//zh2OhrQURCCloU6+3l1xSbtDMbEaTv3qw/N7Slj4MUIul87XSw
qm4dLJToSfzvcMgnABqPynvEccm79pvynLxiNL7WMfFcM5vLKO8y06GKpk491kSj
oYQP2SSDL9PUUYRRBFwTaf1YCQfKESQaWakYAb0RNFxgY4uablpC5N5GwXf4G6FG
ivdwKJw/iFsPV9DFLh70UWuAlJVTfddRL13Sc2KGjPaoWMb0dQmqdK+lRX8YrEQT
B8caIDehkteOASff3ynKgbZdy/tplZvEQyfrJ+O7+7DPS6/F5xWP6fiYjEZOgcmJ
y1Jj+ImUrc3bMPv9G7LZwIUObUmSI2U3GImhD4sKrRpYL1fA+ldLBzQL3kKmK9fr
NYpTxho0oFC6vhgIK/Ct9ISf/DDYHSlt3XI//gTXSSgwFy4rFEWM8qQO112gtQ7Y
5RWDqm/fxzDaRdHZP+JtEmW8Y1tSz2gpB62MOQ7eKkNPI5Z31sX7GgY8lcsPb5ox
w+uq1sEcvmwASdZy5yTRkLYoMOh/SgCc29oUfMtS+28=
`protect END_PROTECTED
