`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QMe4cZGL/JcCnFuRMZ6xviJUFa1quXgMOlTCL84jhPzDE1S/W8hP5HAXm3kfbids
z0LXM7lTdIOCDgNPvbHrIzVPXFOpnhni64vepUj5DcK79ECf4Hecdbke/oKRucFb
hnjtNAR3eUDpt6eHoo/SLXYLKVxUYsZRZG1GiUyceeENk6TtdV1EN57TVVArPlt5
LsxvegHZQ11Tgm8kMZXdV+XtWwQbT1wCGk3cwqG6MAk/eJNkF4OP+wM+uyNohT+y
6vLYwF6HN6hFiy23MY0me37YIv9UEqYEIKZl7Yo9BIWh340a5BiyhvG54RH/RO9g
9jUOlYe6peXXCGkoPgyUK+286c4rns8kFQov7QUI8/vpwBag4JiYahoxVai+aF4n
YgRq4Hzd9zwCxj/zMlPPDqA0vnLFdy/ybZMqLtemaaHGKKczIfD0Q2yHh0cf5xvV
+jl/2jr4P5FBpar5SXvYmIZQoRdnOMXDrfKxtHy1tjL/FPLpaIz0vD6ylVRyxTCj
9OzGR9+DpJe5ijApTYG1cLAmO714KpuTL2T7q0xVngr5ugk4+qGLtr3nxz1Pw8Xv
qZgablMTI99LBKT9gC1MxpbMLxj+aiddSEH4pEJinsAcWt7iNF7NlOWMa7zL2qnN
IjbpWK0KnzY28jZ1SPBLDtLUQEyeYXMWtcmLPVCPOMU2CddDTOFHhs64Nwt3k9gl
MSIsbhL4biMYuqw/mi5Skh5ktw7zdvAcp5s8pjLcGsnBAdrnDq3VuaHWq/H/yGDF
w0h6RQBj3I4Vu8XDaU0vA+1+q1Djfmb9rmwH3+SOJbzSUFl2OJcQMbjgwB8uQh+F
VnvxpTqtG79BKS+q6BJKbX34xCIx+MvckFxnD9c8n5+T0+yCA6wck2SVjaDQ1Fqo
SazR3j9Y9u1pQR3Yl+n2avXnctZQrkrG9UVoOgu00bJznx4MeBDSTj4lFg2ZpmYb
IFOXCL26HBI4hC1LS/Wk0DYz9g53kEXuoIVzUoa08ivgkZ2Hj5FbcP+P0lU1mCLy
wkaCpgaMOhmUjb3966S1PnamtzTQxk4hLc+gAqXi3TcZ6+vVToGPgVJMOW/K9b4D
w8Jk+5GqCo/MKOj/0dD51hhVCeraU6FYT81VQLRC6SZOnMisGf0AUPg0poXFqIR6
YIVngocFxZIMhtd9K8wWi42OpYaIALHda5E00jkG8Rjzj1VHu6mNQCOMTQAs5FkM
PavP2lYKPYPnOEc0V/1mq5sZE2vKaO3SuZA0rJ8wuJfdnoOE0K9Nlq8s5gizBRfJ
H56KrpCQJbGBzcLtf+PMi0WRnL0iJ1kbNgUjZRpeDxoXn7Y45F0kHU01YFPCSXhJ
StdhTwBSgXpht7pC42STgR7GKWiVTxZNSWJt1IKoF/fUuElv6IWmFNFRs/LPPTKq
o/2PchZZ/Rrgh/HVOEosy5dXLCPhSa2M1SweyUReScceuNglGkI2Zl/ZfuCeVK0J
3EzS6s8lRrOJGihavq+8XExbgEe/EQiyRL86MwH2eT4xAZ6N9CNf5eKego+6sFwA
95GRDrfySFW4jsC6+NDFdJf6aWo6cDu11lScstipsDs1EDOpmpeQxK6iL98h9xCy
kturK+rQd8VrR423dmEF3zbTCBMmMV+aLhioSftFw54=
`protect END_PROTECTED
