`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kX9tsluP9ImZIcS6USpnvUjpLRkJTV3SGabsoJgGjgiW+y+ToSup/nQNJG31okfM
TGk0o/esef8BGdNuxD2OBOC8qVJnOHVwtecMfGbD7285Fm+IJcikHUydbqHE1Wac
Y+n5v+8xno/KHkXMyU4JHIKHNo0bVfCTQIslNHljhLnNXYvK/cg3WebRer/p7PJq
L6/GZvPl5p6bKeBbE+hbMhfeEktZoQHeO72ksDFO5KNKGEbkVKxCkz0n4Q9X5uPP
YmttN0YLPa+8p9zNkqHe7wAMe6REYD26JL17mGR55oOVTBfVJCkJuISbvCCASfVU
ZN9uDVECvOxZAVpprMgEJrSiX60uJnAL7u3yYPTLYXvM6okgDrYbMJD0hHeLRkxV
VyJLxuXQCtWsTiZjI6GfOoEJqrFP9VXXmJGIM3Xbcqr1fZ2cyjRlc4K4fpgjj1t1
5GI2br2tp+G6yzCfLEcMqxBKbzRfzKdhdhAV+ATvNRDIEFCpnrvs+cqQ7n8fkvrO
lLZeTJJMs1xOO7r5Zv223f/YSGeNHpeQiKcewoJdsqu2FQoJJObsm5uRsbndrxn1
RL2Tr/ejwcFRzZSM84wYRg==
`protect END_PROTECTED
