`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O+4ZGByrt5Hs4bYrn+L0qHtuo7VGIP+MxvsBAc3p+eJdWjASwsGw3MwsjFScddVX
3Xu9oe/ENeukSyjwA427uN7D/cmoUYMh23Q4L94R49MK1rIHzvcpZ+s7EfpUWQny
OHX2R4ymgHIt1SGmn7cNP90r6EwRAyu/qvtcNLnrbZZhikNXd2l16pOyQ0sYkz2b
K8mFnsqkxoeHh6ZizPvgLxYdN6ThrQjbuk7dmYbvSqrbBvXZl0i/6O0p2xhYfRIt
AsGnRpSL2b68WMpSQQWjlhjWoWS5uKUhswLVSRntW1eGx+pw9002HO+C2PegbHpj
6LwfXpo3jdmKgkb1/JuvsFxybquKTQ3vewDaw0wq8+KvDWox8hvldadg3R3LXEnN
2hgmU9fMzCuUgYDbJETjGYQIbbV2JedqlUZEONKADv/nlCfqvMaIp67VSAlReSRm
rNbQhWjYuSWdzFHjfNT6YTwtyWK6ULSmOPpFwgUtu411bTzI1PGbzZC9GhXJ6TfR
unIdz8+RNXfF4PpwdGz+QSF/EyORMYfOpwOO3kaPAiJjqQ3vQmUQUP7xuvlGKlbd
WTgrk/mStMZ8/9R37adKr6YZ2vI2BVCt2TcigxzCYfbQo2Kd4iMJiAak1wAmo8uA
`protect END_PROTECTED
