`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CuAxv/LgEg7KuwAI1vR9e/hpsAOgiiTAp5DaPZXkuEJEOxY9TGO6SjlJTYGYELj4
ziq9rxtYGoKI8i18RaoaN+dkntbbW1aZkhchD8Epu0dcyuAYQMDNDtMU9tfbnLoZ
wm++qZQOl+OWSKWXw1mu8b8vH14gfM8ub7C54DMoqIjsNUrWscE7X7CfGLw5NfkW
exirNX5App4hQjzxO5Unah7QfoEp2Cx7byLr25wZN0Kaxbb+pxeIfisAbCcH1INh
1131T5poJ3FWG6+shwqMkWYKeQK96h/L2rjb8QJsRJZrCay7cyOqVaQV6wN/Bsn+
r5xyNhq8amDxnLtIr3S8Z8oTahPTkYTmSfRFOZL7FOwt3CllW2iqpdtYe93zVUAD
YwSU9g71CG37J01PjrdJno4LHY0nE2Cx1DsqIdFEoJ3rIdJZkszJoMZ+ihexbk9K
dEerBMbqpZC6WZmhMUo4/VBpvfN9Ye0ilzGFV6ZZYudQkbbqeQhaHcaFxPdwYOzj
duJIUy7fwm5CiKz93NfWAvBO7oQm8rbP+hsXLPOEat1Q6b0PKOIdkCBvA9+WsrrL
ncOx79gosW7IfpDzpSH0lvtf8URoErRxJTkgX6hYJ7+Nsh/Lc0/6nKAgGAFf3ZpD
c3sDVrmM1touU+dyOoANPAANF6219Dwml7z+yFbWJXsqa6oO3fTbPqmpJIhioqiV
PrsvfGonk5vYT2XemgFypB+svvpScg1pn9Y2t6uqDmZoiuHYcNXDTPHnDUb4rZFy
GV9V/d7srwfLHVQVFBn20cLvCWp6Q41ZfXXqd8dEHBXUMICUUvxKwhGLwuwjIQLi
5tr1RHn7oSOq4X02CtKJ+aomCHb2m0YvcF1W90O+85vZKquOhlfxVCmigNdqP/nF
4Hkhpu1lBnbhxxJYnBXQ/15bELAFgdz0GJvGHLq4SaGCOtXRSeTGWv4GNuBN6UD3
/Vxz492Z/olfA+yBAE10TGffk8XhvYrZBZ8saa6Ed7PAfS2a1LuwOeBdqg9En7mS
8UWQHYMSLjgE+k7qDP5senrBAaTdMl5DpO+ANWXUpL/8y2XXnFwTMMEaLtc/uHME
yzVZJFsxqUvz6XV91CGDx/q4npR9qkYmWdbOwehjoehgE19waCICy/LvdAjIpTWr
g1bLbHicphE0rrtmeRKL06LSIDrejzmvNVxVAIHWjl+0FNjkyphZKPDC4OT18lA/
K/8lCDN2tk3Zd+lvABq+QKvIARMKeClFHlEOzo8KlqMZEOLWEncVSHF6oWYEFv4N
tWkFkOjlMnyRcwDCbIMInTDmP+n/P4QYk746Ox5bGEyiILRannkIRCaS7+hIITrV
8P2ZIBpl7rewfiEsYPk43Q==
`protect END_PROTECTED
