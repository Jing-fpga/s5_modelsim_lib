`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8X6HofLbqNV5HZnLDmRm5DyRhrR9s/Yr+KmssClnvVOeE6W0Iit740YuOt6yJKUp
oLRMbyaQ+QJ/N0FJ5siBQ+PTYDNQb6XQc3rSXnuvBXxnITujS/3Yg0PS6sbB6nV3
BZg6icydYF8qwW6K4nLK3UH53bC2mF04yeu37dDmNoFeMtMLXKU5Ua4tGynrl1d6
fEQ8CEqBUPvQm4PHLEoZFzYyPcAKWolamNIM9t9jSgeHSzdkqkVuOHOLchtNBkWA
Z+Hb1y56ceg/QfExLxMNSx4Po/vLcSNkp3jD+qK8Jxsl99DXQtsLa0AwC7RAU1Jx
vG9GCAI/ydSzuaeHsq9vUbh1DeiIeeObJNG4oL9vECxlpOwrYD9nRbuDNFzR1DIX
Nj5CZKUN0BX5lk/cgI/IwCNnRQTDt3uWurvorAm2nqd5vQ/HXyhrkpshX9jHpKMC
25nspaZOeHNDMITW+r1aatGsI6tduduo/6GVYWFeh92LyLmOsuHmtMRZiS83ZLSE
zZQzpr0XO34auQzAgmfY5grc6MlVqo4YlRorJGDwroGkLMpcLSpqpPyolU81AxP8
YDg78Hma2WNhUAF/wmG4ZnP1v+iDy2R83PgO0PPoYqx6S7ZRawJ8RdOuIIhV88XT
qzSexBS/1etQ4QHqKcp5rHyqVG3Tq/3hja7cz0wxMINuxhzaG9vRIpucLwj2kW+g
jMS++3eUmstOXBkF6IBDERpnz8wpnGgWRDbQZYTUhi9EC7UstGaDQNK+AddePaIQ
glbtPnAKR/YYJ5TPFK9GYkggG6lL157EbpC4uzD4/LbEM6QENNiV681OPn87GQKU
DkI4/Y86HiDoE9Fwsnh5z3EsmvV8+bu6ttAbvmN4KP0spciussGRpo9RKP1qx4gA
0LEdC8lteIspt/BWaeTBQQHMVTUYlKI7hA4drwUjKIL/zyli19cpy+SZ8E1BNFPI
OuPtw4/UFmr2bEoAuXE/z3i2mMN71kSS8StpAXUNHM6LtL5lgHi4RGhRQbKMxqYf
BHd8qE5wf0PkSlN4+CTQkYrlNLw02gRezB9o5+He7WklleFEXR9DEiWOCHcv3aJu
8SBkxl1lX38GbGUvD9Bj8p4ZQcH7qmoFyBu+iRE0bxEQjQ4XEOr0xLeoypKKf+yJ
4cC1NZwecYuayLWcQRZEIVryIoH9UVGpJsdEeb4p/dZQDqPAAw66Z5bv1gb6mpOS
hVIjMEH4eag/CVmjOO+vvrO7OG15SOhFbk/3EUok8dkioqBSosu0yDWoEDNfXwfv
o9pxYp+QSYNC78Il7YiWArLaYikOPyXCV+Wfzfu7R6wtnNxeksSWSIzQ5FNyZ1vx
NFua3PSFGG423imdwuPBYwXLTCq6gAsvj0PbJwZwGTTpbCeOyMQDpzxA8D8BuRtq
VneH/nx86PikATimJ1LsBVSnyst5LOdeYqGvoLSuins=
`protect END_PROTECTED
