`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jyOgacpgBySt2Pag4bPGHhm+CxuGsascYGSkcZao6XhzxgeEzz2rzhnd1Uh8glxA
5KUepb51gY+SBxUmS8kRp3yB8yV9hQnmWSt29iRd4g+Uf/AU60Pi2GsQyigk+OeS
ePiJHTfDs67WxkguyzY2cL4O/+qEmgfoc2q11qXUOddcGQ62eCipS4rXZjcQqm+k
94mchr6a3Ctht3ICsb59wPcVNU/MzGRi+IlQzb558PaevJqkOSc2zt91CqKNS81O
7YnUS/5m+wehC9flaocCJfYQvAyekHmOEHMPkHRFVGWnNlX4QAcOxRFEoNVIIOjh
8+rgxOKNgA3yerk7CQsQRxDnGWydWJYSn5QtLLOmosE7Hpej/ZntuTMEsC8jNalh
NFn/7NabCOb8HoFsnXI186plqJcjScZmZAz5rjOyuejSaQIyMJ9WQvTUqA+34OrR
HjQzWhq7WnRCX/1aOuD/ux1TivcTzDIkI6rclEoHv0fgCAvEmv1xSLytL9Nm4sSy
S4OgjdKFYvT8d329AMkRZizCtEbonob/BhH+A3b2PUHTlN//wB2SxtBRj374+FuG
zL0YQN/fYFyWADVm73Y+DvqfxjhHkxNdDgpIl2WaaFMbeOgwhDwVDgC3/YCEVuCV
/ugX+SF6ub3YPh4rWG8eiFZXYc5WQ0+NFQdryqje4Ah8NWoqscMaz842v8iU2BKq
/BtY8JrPsjfV/gJJpML0qIVUgbi3lgdOscdcKGb0PQKbEKOX+s6SQPLG3QJZpwxw
EW/Sh5ETgvJ7hTGgGFwEd51tARokWPCvSOtgoj23LKfAScP2HYWqjp+o9EoSiy4F
J458MH689lW8zN+dnfWjWkZse3TYajDeP4EQtdXdY7GHZakof8EgLiZVdjF0Z4gU
Q8Edi4MqNTfx1Ccv3mpATWNQEhsE3jsIZwUpoBlYSsLMw07cWThLDo9YhJv8kwzk
eZjZQfI0Tg81QvEKNOxx3jIKhptGAvy8y+00eNvETozIVFFxpUsMR0/AaE66nsVk
/DAw/JUDB05h6qpshbkSdOXKxZv3GQxGKPtmNHqq7JZf4r6Prl99QgmXj18x/tAE
M3ib5iP9hBhWCzIhDYExXqW+l9S4BdTerptCuAjb5vGuPqjRBSiVjUKt+L6IwpPg
gR6BAGfTyXojSXaftII5URd30ne2uatJ+G5AHrEGTS8i9wZHUff5NlXbC5fqczrI
x2qjMyLvArCHyCpBWucCXE1lSpUq0VWu8fliy7bJCvAPt3KcJWDOvDMW4JeyYcVW
OCx6e8IXqbOlvCcWu4ER5WFPj+5q+zD3MAQ2z7PBWbYihX/GP+KP6Oa7LxIOgp/u
ds5nRODlcFOWNKPdiQdP5cdlrsOK3doe+moNkbe13zKKi9IUHXZRcpJ2MUeWiAgr
OME4x3o69tb3jVq97pke1BVPZw0NALtSYZ3MdpWba0Vj6ZddGvZ7yTE4EPs2Wx8v
L2IpLqrBoMvTocRuXX8z5gPQ1k6JoN1q8347XzA+tYJz+RNfOyZnr5JlPpIVsqWT
XEeuuVIyizF+CYb6Kk6txJ8uxA8NKMOo6spwRDsC0f7+KsTO8yXWFNQtLxyeKj6f
0VSGBV0DSXRTzx1C1RfrhOssuMWSvvUWp3rDNFA/BJ326DZ/qVZ1TU5R0Je+lMl5
+FfWNsCPT9OPWvmyJC68pUvMYjkdnXqQu481ThJZG3ilfv1f0O3wJMZLMpznc2Cq
U3ppGe5dvaxd+ENZwJ5FuBgNfoFKxVZzlaBe3XFDQSBiIA9hkIh1TpBEMDUYw8CB
dAbKczYnsrAHwFDhYAZj7kZJWPGWYIPXkU2N7u7cZUcS0fkesXuNA8SbxEic9329
Mu3C6zgNICZMmbHeBeQpb2ugskRH1La8A4TE/OoC4fzvpIVHSgjPjYq/7QwyVS5s
yfttH6jbh0gGZqjN8EW5JKkyN1TCnnk88htqO/4wfi5fBLFzbwweskXQYlRse99H
n1vulwWredk+eFCxIRT/cASdql757UcbE6CyfT1x2E8/R44IFy5yNhuWJRYuIHlA
QbWsCPmcG6ngKZiQF6LFCbxOewlwHL1H2+/i9ZOoVEfJz1Pp0/KW0KtJXHQHfaed
6wNV+Le1OEwAoy3DnC7Lk6617S+SMc+1r3k0h1DeeHL4eZwi8WOcxXMpUYvntpdp
WVsPQCZEjA0dUAdTDm93/BHYbLhBvQR7LQ5wkMm40A+PytkeODsRNkeVoStWmiZG
IToMkGXNckhy6ad/jP6lzrDu4Jo/NN0KqeYSSnohcXjSwc5NKzJeDkNBFDfoyycQ
At5LU8SgJKGn3d0I5KZMpGplYEg2gH9NtEK2mPuQuLQIqE11mT5Ij3TTjtyTYRdH
68D8rQKtPW1kZPAmhItghxS9iAL4ggwsAHnZt7J4692mtHRfZGjD76rF8ORHhwii
GrBRSGDo17i781lbQgEAqVqmtsnQJdsuigIUXuwT6QYRbfF7kHogjHVpT/9+q+8I
bQiWm/fKRmM7oIbWgYhWp3HQ5ZMCcEmGYM9uLI379L6cnM+6+FbZ3o2W71RNfF1A
LrIx83C0KP4sqlxtQFsJ3FEBGp56Xp8zis/tipqsuygWAxyIRAZGsE98Rg98gUyw
CzGz1/P0EKEl5A3PfL4pWpLmVS+BR5T4WX2/bi+z0ANaqfxi9UZeGV+LLEd29zim
xxeZyT2Wg8HsV1Z7U+UKCV0r3uVzTFX6BowYZHs2mJ6HXrFiCXqXp+umOC73/+gz
GaYVvOhaKdY11jArXl86DO+V3VNE1Hk8fnHAUSDi8a+zGvgRIlh8Pj6TPJdWvZ4X
ArgAEcwkovqekGrKDCTAIfRwjpMT6P5+vfmiPnLO93LiOBo8moodHIOzhA9eNAz8
DHL0E9Xc5+2ZZf8TlUiKQzzC1s6C7lgdDeMX1SihuEuuuqXqboXslaqbtkhVaJEh
DNI0VvuBS2uaQilMAtQKxtvUp0pNOWQDHXkG1rGdEHU6bKc0cJMObcmPguNaxs8d
vQKrEJz5yJm1/NOXdlAy/ZbtczW+UfiKcWeAL0/EmtTM4MVujZHjG6z+/pH+7zkL
zZdZNBvGWMdA2zLWU6YWM0Ki/c9nNWqJtdFYcvgKEXYT9m2mTTyUDAYcESVU/pf6
ywee14LGrcKVNo/3439gcoHeyxtZApK6wJZJ+Z6WlZQJ6WLfmr4MV0fts75sw+zX
MIucpCwCK65DIlcEE/KZW/NSU6HaPfmH5GT2Du10DQJbMkcJE6JIc1BJZ3eaGwTx
XpkcDL8Bz/sseeltxsp9Dj7dPWATEP+9oNyecmlpmLn+Fi8A4k8C+2R99r8hZMxL
bvVFit17itxChd2c0naH5vlD6L7BIux8+qMbeLUxPpDgG3HsGUXcbH0MKKc3r5W4
HLb0m3UBWuBa/5M1HVtpaYIqXd1RnizZ365XoFEGSs5HyTep75iEIz7OVKpqnWCt
K9D39QF3uWHPLS9CvI7g9pJFI/tvuWsj1UIUQqi1GC04oqDsaODhdIi3fKd57tPL
L41IHo5tQ0eeDk/QFthaQllRzZ4KLAavTytIJRJDUY41fMNXzCK9vSi1LtWxg8tc
8vU9FBQVs4XtbHGg23z/m6riLTXzhs343B1npPggNPgvwzmbFLAdjYT54JdMRv42
4/W+8552bzAaNrtwQNc/Yi05ntOMfKueZcyku+7kS45K0z5y+f8Ov5XDZ4FFXZwQ
0mrtpZU4MjCidC2cGjoSK4Izqr6t1FEyL/Olr1nhukODlZ6WPR8MJTp/54FS4c6r
CGBFB2/wY3onul6HSUlXvCE3IVciL2Ai7jrffLD+Tl/jjifQsGzILyEZOc62n1/5
`protect END_PROTECTED
