`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W+w/e+NM8HhtIOOUYP9zD84V0uS7aAhp2BZ7ng3PAufmNRTDGIvjmJUSqbwpviV+
6vYQqMT1ctvH6WqkKRVWKFZ9siUdDIxoQ76QiPuT1n+VCSfbPVTj65gXdwi6HVHp
RF4yCKBUDz/QCsCXHYDXEXKyt4Bbxles+vkfQdN+D6qlZKzGkFxrJ9qAywTJ37P9
yrYquvYi8Kh+jEdkVzJvEpSLqpoVzpY9cPBeKnF7jMIIB+x+wpFlRb1Zn09lCJrO
mPHCrPj3K1FifTAIZ39frhaC5jzn7K9oPXA9CNBmnTLHMfk/ClxLZvZnxRMzm09y
MDsN6cbAEyyZaY6wzzFQ/YTqSg4UBPNqmAw8utH+kU0=
`protect END_PROTECTED
