`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gEj8Z8j+Y7iLW6fHEcJnqpWInl+bXucd+qG0AadKF1lNdMn3ivHq4DmwJIi8+HOK
ktVNR4TWcAQDUUlrNMGjSqU0rCjanFjyHAfJWlRM8C9UaUh2jGoEERx5gnAIqvv9
RQZQNSUyIRMXNGmxkXrAbjBB0+rRIQUYBOo6bUOvOTXMcO0j/wu8GgoQbmA9HjwD
nCIueagO5Eo3+KKj5VsYvNHK+rCG/NenqplieluZvaRoFyYmxzPpeJHwb0HaSPHl
zsLX05rYsh1VkxCxcYWzt69Cpc253dRFcu7Fen0v5wWJXdzCfrLHWSVa18Wi/Ijz
FbanPK9O1ZpXbaya4+HgkNSD1DyBcT24plnDiV1zuST1U0+X5cWw1ozGaSTy5GCY
YUfAniRFOtTkWv8DseA76jBZ6FgWsKVXAQTnk+uAXdNo7dT0wniJqmVeNrBpIZed
PzRZ81yk4ImyBSYx2JvrzX1zpQK36ie3Y4okEfziUiktOU0COALX/NkwuxaF59aA
G+kxY0JcMJ4ygpQpoky5gLtP+824drDXuBc5Ulvumu9n0i5Mdp/giCDzys3EG/7E
Rsaa8Fg8mbYceKX6dYekdMRSr7egRAKCcOztYiUyoeTNPDvRpanZGF1gqdESqCga
BQkAq9++3UHM0FZV6IAmPhxjxsjc4qBvniwumCxMynjXYH6oF9aJTm6EC7qlFzr7
92i3nYbv4s3VXvQGre19a5gppPjK0yHMZB7gmU9Ybus/JpIgHKWTUacoCUqLGZI8
2fh6bZgW/0EvhD9zWZxKSneWZ+iMnnuMPrU1ZvrofjhyLh9UUdGFewUTBbH0oIvu
FF7pkLhEV7KKBaQyuCvDCNXPMvWHlk9leQK6TzViSojqiIaXVgayclKbO+ZzDbPd
CDcIvKBitIwYXWRuXBolRXRnIUymc17AMiIxSawCAUP45wVnXgeA/GXFvBmdg7zJ
ec7iR2hXuP2UehKG1go8BaKVfyWm2m34QGxm6nbOnWKxwinroRJoCI0k8/+OeoLI
bb0kMqUNqU8sqf+ZHFtEdGLCLsEKEfGH27MOsDb2XU8=
`protect END_PROTECTED
