`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Ui0c9aB75u8mILHBRU6WGUZLXdAYXIjGV8KV8P1Nd6/Ud2kCHukI8duj28fUaz9
GVxpnyQDKSjGtzqQ5cCbsSKHsLWXKhGqtT8STEQYmT/7c3oeHc03ZGrBm8e+kJm5
EUn4ZoR+dBEPqexz6OQPXJ0y68qGJs0S7q4V5ng6LCEU/X8WVxJLt+y8pH6/9F+N
ftFIzt8KZEFz4qcsf4ROfI8UgkCb4V9WqUO9JrJJtIK2l/wSjQ7WAD53lHeJyMHE
L+NOkWBqSFhdIfdXiqtEZH84NjTESu/ZKp/2ZcbBarzRHgj4zfEAlm83ViVNx/wb
T3OopPt8Wt1ZiZFP78zNpRHJdVh27BqJO5Endql7CFWbZJSz/ay0IEoY9BIaVXuX
fW/oGgXXcUgHzRTyDstGfNGV05AIXjgSj75tFwo6knqR5JgnKXULmzwpDr7hht/X
jkfJXFzpKEV/T1HSzIAfU5qIAxZtPSqOiw282t0Ry05vdVED4nlUa7lhvIKBY6Ql
mRlAJFmWdNwDxR+HgyXva4xU6TO92QlhPq3Hcu5cgf/l11OS+7mZahxidM/b5/Ff
rSZOhEeX54zIWtAnyMtkf6KVcZ5DFS8QS7Pr+4FMPLA1jprwpfNsTm40k3HysZ8Q
9177+mQ/FTzf9P5vz1KNv40+wKFYiRZ5ERbTUx7r8Fjyx+vSmtz7Cw8afbKTzfO6
C5Y4Hf/gg3jdUTxxRtc0o5DQWeBfubYkGc056XQzifpeKYlAUlSMA1Zf2LKt26fU
W1srt2J5v1FbLwJ/Q8sXdt/U53dlrlTuozBhI57D+NA=
`protect END_PROTECTED
