`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T9229u2/WFqb01buajj/4q0Du9yN1+dUlUktMduH7G1eEQBEVL3bnR1aZfQFqQW+
VKUcYeAIEur4PEq+rcCuMkIbrqj8j3lGv64FihC2NNxvHCZ4lbT+p6eXG1KgZPh0
UaK17oX8m2AncjmfOGStnRhvYxVxYYF2Cy/cwfR0S5JRz+QzKbNdgzGj5vp0MKUH
T+H/UpRJM2HW7odZFhidyiAO9J2mnG8oGJMnb83YX1NNpCvpNYvjw3fZBtoXdNEG
B1mppSG+PasLV0az20++mReiPb49gyuL+H07PQ9VWIaKXckXO7yGTvtp52hLjrnI
6+Ep4jUdPJ3WXfN8pB74dLUHiPqdLdkmu7kmBU36Jpl2kBfL9NaLcGeV/ENOPjn9
dIUCt2XuPjjQHTx0Z11phOs1qNFmYJW/0AMoBVBuucGVhDwXha7ry4gE7N8BDZWs
HiiKFvN2A2ngv2uoCIV2ZpAVS6X51r9t8cLPrYQTNOZGh2J1BFbWws+YabMWg5LK
IAagAbxZ2K76TYWG3DpaVhYQ9Mea6oFKkZ0X0f280qbYT8+CBqgm2Yb5rx4Vae+S
QUBLljAgdUPHVX+8K8KorT7lfp4FMDQDOy7M4NdZc2ZHc/UyIpnzxCVqavUwGELb
L8LEIPfJtAMevKN+EYyKsALQ5OIct0qRjR7lJxTbk87DeYFhMhGBQtoZr0XrtUgw
EybqSzZiM+pecQzpG8eHHaWt4swmg5zZRUXoqx2WrFk=
`protect END_PROTECTED
