`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ZD5OrovADeONliUij5jYC5Byu9edz0mxWS6QQYS15Pro0DlKR1y/z0tNhrbuwuO
+sYTxHKmjcitqbqX1yZqkn9fiBF+Y+WVvygANBLAppEcj+YG0Bt9vs7/5ptQE53N
FG6NkyebzGdT6+o61t8AV7MOPvKp1u8E86EM1kjbuxYV5HvjWmozGPjOBCiWWj3w
zMYXH383yswEGaC5gpOVIKBa5ObhyL6Q35X4e9aV2EhaL1PtrRGlsXPCG+1zQiB2
aTkWWcRCW22BUDjXasDPR+yFQH48kZlJhla8/dhfgWXYs04TSbS/Q1d/06/plv23
JUJlXwXU56JcWtGEqdedyEn0N0eggSGbDaQseiS5yBTENhEuQGhtF5kZYOsSd4E6
LkiEcvPCFPswkAuwzPkmOweGmRl/W4DIqcWAC1Uw3CAPl0Q6EJM7DtoCpin++xsP
EcjP9HtvQkYGMPHdnAJ1IPDu1UbnWZ4dR1ZE4Ul2MrmYuo06dAWI0N/homO4fSLb
LzX49/nhtORqeQYX/HVxk/BgoDd9ZQ2qHbq/RCJx/S0IPM2EByb8vIJ7zJ4+PORd
/s2pESEK2MoCPJlvtdhnj0YcEgg9/e+0zweZptZ14dOGIcMGWYur+W8Jjqp7kHlY
BFc4K3DDX+wPLe5otr7t1AJKJErvo0BahLYpY6SMLEwGxsdL6BDiLHVRJD2KbeYw
UINu7+Ni60oSDJuDMxn95egk+LKlovxaeKZhjQLYPzlAmCgCJuQlNBLyDUmh0Jcv
SwwljUXBFT/pXe8aYTuAzJarCTSjZeuQn9JvunB2FxnEA9zOydeg37/XzqYzDAlW
L998JNCb17q9d77Eij2SNuMGZw3mSDC3VZ0U8GtESL5BTSIksL0+2FFmhIWEGQOk
Uniwj3ZWkxGW2E0a2zTpBjz0lKPqKXQ5fv+vIdwZMfW2eM1d+OzKgViYhc1LjWzB
/97LZ9mhVNDOmi6E34PY0++2yrSScaa5WjUf08z20hgQRoCZ4MpP0l1/BLzLgFXW
4Vj86TLNSVl/5bDB76muS8jHsbf5pjNHi0fpOM9u4kYUizaGt3UMpcShGbpj6wgf
LpQMEzkHIi/rCXXI3KIeMbRQb0YibySxRZv9i4msvYYunFGcQYbeBPjJhGx/AFu/
nK+k6w0fq9xc3O4fHvuRExjxdI99JKq1pBHaR0UPelnKiTNOGKmABphStYjpp2Ew
aXGdb+/ZjfUCL+WKBJKhBccHnnags+InnTkCFgnVCRdP+UgRVlui8j3wVZGdxi39
Yi9jUL9G7ETyz0UeD6KBAyC2wjkl4DApBBANfvFRFm1W4JI2yU5KHUGaIuLep1B6
pgcKpK9eIGWsGJ/+6mk/v9qq9S8CNZwNOWzO0+OdFCjGlHH7v3CadTSoa3z/d0Eb
C8EtFwz9LlHst5N4wdCmDXUJiXIdJi/l8pKKEPQmt8XphpYsLUFGpF2LSq3lXEa9
3jFE/WBMO6HLJbdz4q/z4aH7td5t9WYsqUcPshYWOQ/FCX+QQDokoysrXCvZLNZz
oa330Mg9DiB7GUPuarGUOQ==
`protect END_PROTECTED
