`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Zr/00w426uCInWat8Zu2Axryz2InPGx8l/NqXoHwcgGvwIRaMtxDz2PxhThwCdN
nGrhIMSrwb+V0GVTVP8O6db58Is3Jku9tvBg0hCF0l+TR2zvr708VNAE/70eyDpW
0IyZCMg3ZCncybFNgdrg7e5Zg6TykHiydk6sLgBQihh4lmbaEF4VoTD8yrLyznKl
KbQIr9jwsNvKTmnT78SPAwzT+r0AGI3vhwJTxUp9etmV0etUbC13NyDT2iZVjRp+
k7Vv9tY36993aEKNE+faMrHQr6fbA7Qo0SCWwpSoIW1L9MBhp/c7VMXZwYbRmtXj
Gg07xp1R/l104h0E9qNeQZdGxJXKHfRLhL43dcS1ws9XxitqVV1umx/CU7hwCaWB
A14qxj9iERSosl8i0ZxhxscK4zqnx7OZ+uIVpQeLNfKv9V0zsEP16k4RRluuIg5u
MwliP89mgIQscFNqb+AVZmjC9dKXLPP8QRduPdtgwhmxHXVTwf0h5JPrcxe0E58u
lX3uWOEUULmsVeui94IF0F6qvFd7pczJVEMhsZx+U+4Xw1pOax/aY69/P6uNeFVg
ZdkX3Q0FQ+q75MrIFwVSE72MHGCDkoBqkrqtspu4TzFXjFdmqwp5/Br6zdRiVO7s
qcp8hlxMIYnduUnQ2eaC29JwjRZF58cEMBcXdhsx3damP043XvTgVVCle3C0N+0h
BGzF7lV4lwh/Ud823neyfmy6ftCDcheUFEIUE0a5K5l9+rGpnkcqjWZ3S30Ue69M
rgDJ3RznWRnVJ/vpVFbOr8mr3RUQD7L6iks3voY4nI9xkElYLueomTzFqCNHHcwd
qU0eWQxlcaxyK8OMpKcW3iWRONxO4Esrg42+OGZxxYSrvyHiKZjBKK7IC3AagaLE
cxPBkwXSBB5F6yhozfmFI7X2GvlUElap+kWx1H4taalSapkpT1BVvOAIEFIzGWQO
+D/v6X0aB65ze9PkgB/Fpe9zfPDcAN9kxpDGT6rGir8Od0Yf4GxvWaw29KigzfZn
kMUYr/M47jhhPP2L/pICCnHHeFjYrmOcNB+bPZGMpW2FyS9d03WV5rUphxfPAFt4
F9sd9sV7s5ZJ47sUpGRStz7Kr3CGPqDZPFFI8eKhGB7lcPk3zJLEXiTsGFotN/kP
im5HuTUjU83AY5v0d+EBOdHJz/7rxsRxG3frRTlCUQzbPjLCy0XEV15uqSHtdOtO
zBEKNY2Oz9ClvdMbtlWlu6wVO8nbyQCvk1/txvioSAOv55CJMT3u5W3tHlVy+I+0
RmYavR4+/GzHBURir7TQnUJ5hsKHLKONGUjDJ4Onq4zL/ItxTIAMPgUiGbD7OHjE
Z6L5F9c4LzafeWJkVGp2WG3X80FXHnGnrBYLcLPclF7SiLQ4XW+8A4IYX/9l7Upe
9AshPzcdBzABXsnDkQHKEI5ZdhCtsmPXcV9fOV/hs0xKPjsafZ6bOXfV7QhPugAM
KpZDsg4xkUptMqInM5pCyYF4RR75ujNuGLMXmfqvpjONLGPG1iPfVHCxFf9dxAfN
w+53x+u0rxyTEBqAraM8e2cNbjFaw0t7oQOZE22KaDRWD8P59qLOWQ6k8VChpWd/
faKR647+HEs2aI0sAQA1foGsUiz+P9pAd1j+33sBc8/9+MPe7Y/3o7iBvZcYxubJ
FJ9FAMB3D7NMOWUXdRyY31iuuJW9MkVzJH0jpOWYY0JArVkxiHeMKnGDm8PwgrEx
1L949U7ZxQZT2r0Y7fCTzTrPqWhecghQpo5SS+hPlZgk/86PaHA+OuParE2nePCi
VcYReSpiDu3oQcMD4TG1hLREAfZIxe/ofJhmQ0gqTr1rb30bHAgC2Txio35UTZF1
v7qNObevZ6dFkodB2hAYyQ==
`protect END_PROTECTED
