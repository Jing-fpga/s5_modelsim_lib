`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ir8CaOw5lPSfH34ezxY28xLFHrWWBzAEm3ytu6KXQutHHArNMYaMwlo0bulX/Jl7
s+PsLueyD9zubz1JE/AYn0/Ua+i4jwmDv9rLBJB3IZ6z6xV8NHGAMFN1dja2UWfC
GdtRNchL6LNMI7QuceCeGBfTvuhM6fK9S9BVLM9Tt49PBe7pOQUdJiDFcDDWMUMd
VmRoUvlpHl3D/yIBinQeLd2qaRZ/3UJsuJZ2HTwa/TFJaBDFX9q8EVyThILzlTu6
tbOlUCPJheA4J9IdSopTRWKhHJBjPtiF8UafofYCjScw0l5cxOFlHxfbehS5pCWg
a7K/qRhNKA4QMfDZ3aWrNOUBKwcwF6njIxIsnSDtbb4l5kpnLrpjFLn33FryO7zH
AvOLq8My8zMBpCz3sQpL29CJgJx2XF/DSU9sGAo2itRp6VRE9THzsOi2MRbGShPR
LVQf1Q/WJZsCDtxrzgk2QB9D7ng8+lBfX7SaQWT+v74DMbHlD8Rb1kY+cd8LMELu
3Y517Pkag15VpMBzHxhxPDSF6unnFWZbaOFL0so6eOdKsg4DUgt04eZimXjBBIJT
y5VuMsgPF2h9H8q5XwXbHzj3e8idKzcZ620323FqHuQalm2Ni/EQq+7VKgY/7Cnf
2U8vR+YD4UnhJLcQeGbBi4q0vkki6EzNDgie7lyOPDjbw2xrw0w5qq9t8Eo//Xp3
QnqND9WRyKuaZWAevE9UVFEUQyvPT3P5q3BAOGDiHm0+ytdMSCD7yIkvKZi+gmZE
W0wqbbHItFFO/o41ncfLFmUcTtcIp4Sg/jzeGjLGvFEH9eOkDHqWsBxoUefmOcj0
2HHWjyzkSQPMPjlTWN8cJlo7zXmmvmrRnmuPcrq6vnF0WBTmm3WJzq/H6NiIYr1x
XV2+JRYJ3yT3ZD1IbNdeoOQ8NQ00dcWelujEmzyZoH8cGTk+HM1zpW7+OlLLywX8
OcRedoZ6PfWClNmVPYQ/R0UuIzlWtxO0EOhfBputqUKlxYoun63gvA6YK4BBem3B
vFA5PjKU50inRNTljlyPSZaAPz24iN9X0cyKPaFWvQq0gljNga4KyVRbAyYZsw8Y
aLv1AVquvmPn6fqhy1oxGYWLzCBMlps+bc9sXm5WuyzGtr11gHBY/5HQlWqsKQpa
vt5wF29yO/R/RWqNNpv3WLEfhSpx/wC4hnF40Z1VLuNq/pQkZ0h6wrOPry4k+WCo
KBneiY4NBNscREvQAs6Nl8/8lC7ZvrLb+UWHmRTx3JDewJHhEyL8fKl2fBJFRQLM
TbEOn8UcCQzhvETu548XtnvdJuvkUQYz6iTHItHX643UHStV5ntHTVquTG523lJb
dJYREqYQ94z9N3rYgNLQuMhc/E/ZGhR0z85KEELI6KruACIvNCiPmigcwu5Xpj2E
gRV6uN0kxLfFK7qPl9BKCfMqIFnryjboJGXyplQtrNUjxs8fSqxzAPhu1CRKWloK
oeIjco51cUpnv2Hg+CkqcrXYcq3zS9ZSOhTJKoIEwizAdWPKUAK64QCbWh+BoI32
ALJmcqoH9wDHc8R+qRrWz7lPhMwJ6IvWD12dyi6pDVZTx6vyGzvmvYSBdYCxqF6J
QN8SJ1JbTVDD8nWLow8k+VAOeqRn9nVB5e4DRI/wZJA1FXQR1V+AO4azkApLcrbT
jc1z5c6/MKHGtANiNoVNzMX+XdKL3Y2VMUOPbqoWVdnW8OfeXlfc8gosdXT4mTh0
UIo5g6E0KEd0EfMicnDKL4+KJt2p0MUKUu91TKrXIdtkrFh5q8J7iaT5KR3mGu5x
A+taO6Cfz7BUD7BMhLoPKH3d7OaMw67K6G8wSFPjpOYk5zNpo/EHkA4DvRrNf7Km
fekNgaWM6BzvNJv2zTHDdgIjCRa5JSteY/phBJ/+f1DMxGdDCHZM8I/awDlF8eEs
U5DmUAJv6kOVKlPoXIYJNziTwctOgpVr74IU5nZV+TOh80aAp6vmrNJrqpVu5Uvi
keRRRo8Vb3t5biz1vXeRG7wu/Q9x5BNaf4O1YYcV5QUdRyHCxqwyvnyM70iZ/weU
l5EyXzUOnZBWY+VCZU98+LUu42IoPXx0Kn1DUAdgn3To3Qdk71d59kZdljBxj/CR
er5OFPkMR2PIMlNYbwns0e+cNsuFhfQUtT+RyMSk0b1ipnzchviSYaiNFZiI8v62
8vgW7WIW8At7IHiCi/DPCO44cbx0xEaARGV0W6hXc87XWMgLzZVzPKMvEgdEuJDa
qw17mwYGppFJQ15Rkqjl9ZiQ7yIWWNrP4aLSebKhXZpMXtHEjkXIW5W/yT/kecMt
YXkRmXG+rOOaJfXmyJOynbjtEPgq6q4crOLqQCjgmMTlDtQhxwXseDklMx3AGT86
2cXYVr7jyigCC+zXMtBtdONIHAGuiuJ3bzib7iJAmDdX6qjRLzY1APl1HLH+geIW
k9gQyjZoJp1AdpC2oxhRh2j7PEiryzlmR4nSNpW4Vw8S0bMTkLTIajZKvhVFQnvV
86fEIginJsXcxOqhOu0U8fvi72jqxnA2wk4794seYgIgdfCzO3JfVfVhVh0IehzC
FUDwvjECfWHeTdiAFFTbVX92UTyg7cMH+rT0Owwg/NU=
`protect END_PROTECTED
