`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X9B5oEwBQZgd0QkYZTY1w1pbeBk7TR+lKCZw0edAFptybf1z83ja1hA3J4yu2/Pl
TePObvNtdohVR4+A7vmyFuSotZN2QfCoG+2aRwkb2Eynmixq9CDxK/bMy5DEnD7S
K1ZsooaWilkSTtEy6nOnNs8eh5xYRwdtKtNnr3IetRlmEMdIzsmIf67duY0azukx
ISFguUTaGjokV5BgG7OYSgIKhKq9/t62nHegnkEOdXvsSjDOZWNDF8jWeQeUf++p
9QszgZheEfrQJ64R1T8o1Mil0y3U/QN/X4pPfU778P6KWEtP5nSgzB14zNEx4zOR
UUb2dPelJS1zicXslPvrIhrbH5cJmaAx7ruNw4Cxdns/fhvdZX8pWG7WLZ7ooLCd
bzznDxTZeWLi9FgLppPQiyd6XD5cADHxFY9pgb41wLRZEb7eLs3SonaqslwyqqT6
9K84r3Te8QZ5iDX5ELQ0GA==
`protect END_PROTECTED
