`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E9c7NoMW4p4QIVa5DAzLXeEcTP5BGrb4YUtLqOi4gfloxKLPJE+rCcCEbFPBZegD
1//93rmvDw/dN3YKAzRwSk3OqkIhEHY4If8FYLdBIj3a45ZYTLgtb1+s5Z9OLVjq
EFsIAz9MS3rTJArjVD0r6dJDwfqpS1idm6+tcD/3RpJjOxAzIAnqAcKg4QpCtFcE
gar+nMNAkOxsWfZ7MKi01sMWBxPyQe8q/rHFj7u/UGHXG8ru+czM/CGpsK6D3T3i
Fw/FnEfsGzEXbG8cehMuzuocPCGhxFa3ZA5eWwNdVfa9aFtQ22mSMgkhEAOmR5/G
bMOjsLjUiwIk1MiFvMDIqeYzGmclI8IA7FM/pNElE6DBnEyWz9tc7P+f1hTd5gnQ
EOXvCagDn1nae61U0k57O9JD4+37DKnzvk9IJYXtyYkcRxnBWcNfOnfpySBXk4GU
Fr7QeRrU+nVOkSti7gMhPgDzcw2I3vgmN/vbXhch3S4mA1IG1X9KO6S/AzeDozjB
vAwpa7PUbbq2d2+6R4k2dI3UJwLYZewEToDtEDfYI1A4NzRSTFKgyKl6yr9mRaq6
uzSRqtmHbfNb5bdgeZ0JAwhYODY20s79WlzXLd5OusiLSgONaW4usfU8imhK/jpU
EQcjyEP7hg4z77y0pmjLkjwZOjGuWzQe0wKfzRqNN0l/nIpxezUqjRybZ8ZIp3Lk
vVgDNGpBT47/Iwe/I7WWmJZNHPds5EnhI6/O+9X2lokKblYCo0BCFt7W+9wWNHJu
GwSvDTVAkKBacF4OPCn15J+FKAWY1AkpJ1/5FAzQZxFywvPFl44GCN5HJ9u+oj3L
`protect END_PROTECTED
