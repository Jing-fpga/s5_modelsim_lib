`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
go0RbqYrkRjXPMVXcQnTgU0UikDEYxsZwQ2f4UN7V18VVc8iiDTGQSCFy1M57KFy
aKluO7XqVGY51KqEWPokb1Fzvu57oLE26QWbpqnN78eOjnnuAR98wOfkwctmAS+J
KGYnj7mNUqvUewEOSWOVaK7qWdHO7m9rXa/ileHnCGNma15Eug1PZ15YvHo9JRHG
Ou3/Sz+0zqOzR21yqGGEp+0ZlYGH0hXD20huSGcyGkfk0zSmrc3wxWXI2UWNrG5R
j2YWqrYgEuvMgXsMrY28QyZDQ9ba5YBjXMKtmVcwiQZiTYKzNQfYBw1fYynQk40I
UToUG4ygCyVaY7cVMITw8fMbmfAjjqo7p6pKxxIenhvsjnRGJImglgNfEelbRe02
cO6o6YJsgGLR4xPOxmk5mPtKPqB0Qdh+llcXYKzGncszs/bIkseQQl7OvGFYFQjH
EQ/rf/MrgeqYc0COXVE28pvn89hq2lhV/30IeSdZBgUAVdxC7X8U10SrDqI84f0w
x8omZjwT7dihODjxJMU/cKlCm+/YXdCbXCsSPcNCzHdheC6ZAQpp2yyj4KzIU/rL
qxdRDavGSkxActoX5P84LStGgvL2eWGUo0oAB4hgDlY4RaB+5nN3I0MGDoj4SMv8
rgAGjjDcmae7zAsVDmZHZbVCqKEDGrcDYKUiko4q68rohY/fDJ8u3w8H+pAZKkx6
E2+lrQY02ur9NzYAsMQN4vgtSbYpl0MjZpYXHNav8CBHu3nagRtwPfs6lM1niKKl
Z5D/xUD7Aq6gFyEccbJbKBtLJHbKimwZZap+xRaUwYMZ7RAhl+0lxkiaW1/d6wZ+
IvQToy56pcbcF4CsFh9y90xh5D2agqtWF1OXkLtt0OQU9R6OUTLXGarTUxQdY2id
kiLIPa+Q5Gv8QjuYAeJw5r/9DFckfGA6qT8JC7FoH1jO6v/Vv805lpJgdYCR0heP
`protect END_PROTECTED
