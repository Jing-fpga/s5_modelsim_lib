`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3tAd1jHuZ7rpdaDjuvQtO7IZHmNlxBQrg/zH3NNb2fhqwpHqqh6b19js7BVGJOIU
NFLwFEbcxBOXl1wHkUQ9+wYeCkiLBHXJJHtXVkAS/zi5fUaGWdsX9BPfyH7my9bF
Cb+Q2JVlNk0+gWb1walHEc8QRT7sVm4Nanjh24jvs3cx2Ba8XBY2y3jyefHKoDqu
4R8OLbnZOzNMgKfFh8jiqQi6IdIL/VI/1+jDWUo62dQrRxKh/F7JfqSpTbuvTiF5
xx4mEt7PiCFDFeT8A2uzWR4ParCVoPv87xf6tOasXHkV93Zpi14HuVjctciC+mj5
B8UylJp/PdwX0yQqDMs4kh9N+U/zXTefkFQxQwe2HV8RxdSatbo9+X2wNnDjxZMx
qQYx4XO82WCHH8c3MBd7HR2HZryce68RVmPwXKchzCDbhzPGVo3u6aEcxAmdI2Tr
YqHcNJdGRV984FQLFpN4Dz+0RxwR3LdsIXF+AJ78IT5C8w741JSk7SK/2bA9I1xZ
gAC/4W6X5S0GHkTjBGq7NSSsvNHIjFpSGR90IKs834UaGUjkVWhtvB8gej+WIyJC
fW0bOHu6SjDqMA9H+MW5Gq58LH5XAh7IrfUWptI+sVp0wkZUnqYMga84cmYO5ylA
P8Ya6E/JDJMHOJkt+bBH+aUBSjdIWiKo455Qdit2BFcl3TLj44lN5tDTVY0N8IV9
NE4iiLWPMAcCGiTfE0YpOtmqQSPAA6JhpcSAB7UK3bH+4Xa66ZNv+8ou/RpNnGYH
BKLonkMwhFEnm0D07rbVZadVJ05MomGj7GHyp/b2Q4W2nlXod0mFEluH1NPDhA0n
uP7nEzZdx6tjwke/6U5W2jDRsp/DFGYBilfnUqgMZlq3zFTX4EaUCBS7LgqoSh5t
ON0BxXlClpmYHbjxv7HsuDODxqvk5w57dwASaJ8N0cf6tug9Lp3ePAHDvQKuGKBY
VnTaZNOoy4AdNNXqVqRvjsn+ALC5Feg3V69IMAH4m2hItLogsquX+2HyoJzGgzcQ
7fI99j1jczBu58KFxNfT7GRFPCKLJokXRTgKqEFugeJAb1lmrvFhYmgp/+c1tt4q
`protect END_PROTECTED
