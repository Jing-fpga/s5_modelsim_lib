`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XvbPkkGBBIkqOk3s9s/VgFi05ePK+akUK/+TZDuSI0tdTn9JIPLyE6f8NuqHJHTn
gyq1idVneGyq6usDbd7JuBFweK8lY9nTuBPJcJ/AwE+2Q/cNJhfbk4RHgBltB85J
xpkZ5fZ47MRYz7qnLxUiLvEXQ+TJaNQ3VKnHdpAlPH4azpeSguapS4emRkIoldJ9
38dTuuOdQZxaT7y8aP425ytNoKN1kvZ14u3u+g9lLNrnjFJkMiazU3hnOEeC/ZkO
fZ9ggMZXXG808HMRLaNvcRU3M9d4lklC5jMd4TJkMqxwzA6k+uXRLtOfA9Gsc2L8
tfKC/rlnOl8qSzwcvIc/2CJZIJ5VjW/FVvOFBxq3SyQOQSO/EOJwxPIXlllFbTnC
wwWLRwGrSwUhcodCB/dSNBiX02NcSFj6Dyx+cCgZZCQnCBLglA0OIOMMpvCigPT1
X05bVRNDkNB08JRfXiczV4KH5lCDyuiBlIqcgnxBXIX7BT4a2QFHh/0ftBcOaIWw
IHY6dfM981GeM3/seW45/frYBS/zLeKOW0UosULGiY4paIUnorkFKs4FMH5XGu+L
kP/7W/bzFMOsQmLxJoLqIP8ciE/F7o8TEAEBfE81FGIBdNe4FEXletdJF8lFM291
eodjv354WCpuSlixJ1Sh4XSmPNQOZ80A3u0p0KJD/hSGU6b0UU4Gco5CV5pWQ9vy
yJHyuCZbNVCCwkNwq+c82Z6f4QutjOuYfXEKiITyemcMsSlXiHKxM5ZjfiT8SblX
4P0EcSUckbvk7YMr9YDfxwqpd9g9d6EBjoDl/3tvrsYZexEl9+Urzq1WMVCpgHGv
OMSNfzhAZ0m/Niyfv2+EjVydZI3V0aCwZ09v8h9fIWmsX7IXEW+qYH0XwD5eTRTl
Aa3heWxbNoxi8TtTne+2fGRnSeIpUvi5l05645FV8uNFfzmV6FbwAtkLVOIk0f7Z
nzMbay3dfTVVWkSCfzZJrJMJthUX/Zl0aPmE1aeDeXH3CkNeCYZy8QkNeCHSg0i7
hTaXIjZ+jzLCryxEbdn+auUko+RjBH1yu7glCLlDaLc6tcnXxmG36clRXrFVyD8h
kbxyaJb4bSjRoXoILpR0t3YwXNLY/NG+49houbZuk0RysK3wurs1KH7qIGm3Di8z
75K1RBg63vDsqxuNaU/ODRWlG1lh7nGzn7TyG0UyUUNmwK+IEdViOjpDXDbt/yNC
LsAC5uMz0Vkv7XmrbR3xgcvjnKKKXLoeeorVCxcyRUusik5qfWsoF0eY1eeyQCYK
epx9HHY56qUG1sWVjxT1wqV++5HDZDRK5Gpv4qEOh5msbWPmM3zODsokxUTBL4RA
XHTfJF3JQsahb4MOoFI2FnxPtQEPWNuXRKEAZG9K1x2tepOXkBFhzckoorWIXdRo
gkK0mg5BCP/V9GMqifw4Voh7gBeVPx4od5ZuDZgq+eQAdZwoaVvZUQSyuFri+bnr
B6fcQfBJU8Xs081EIaA5L65Pwf7YwahClgD9l6pqQbs98LjAq1clMRi38Dvk65q3
TAoFr3tBtrte9LFWrEnND5D/hnIvPbHeZIVtBZ82+8vVmnm+Wrr+nIK73VCxOk7x
puSfw+WTsJrlpMCEo8KOV/KsMv9mmhu2FU5VpJW/wprrgg+ucjpC4WOT4VEVTbcP
kQwR1Ep7HjKON5/IWdmHuV1lLedxHbiksyAA+ok7EbelAj8S/tHluGRdF40jvv1D
FaLPLHwM+Ozt2ex2SpcZcl1iqjhzsKXcDRRrEgmTgv56QZa+E+zUjizK6LudbdU4
ZAXsIvtpYcpduTqUHBR5vC9sVW+rDdWyztQqIk0+drrRqukV0mB1t7Y8VBjS8jzH
6ahrE0l8+XtFXS6sABk+W+q8QK2FBgVzdODzoTuQsUjDVhASouwLi/vqJYik29JF
1RrfkQ9f+NI7JkHcEf1o8U9lbw7CuUPubh18wrIz0VXSH7N/u/SUAIv6/SWYXOt1
nUxDIzfffDMKNX0cBIlbbljB/rWqn95qMIB43466D0EoTqrvI5pxRc9rqZ6C3put
IuIW9JPMd/YGejqp2CK5n43Ox4ORrL+zl8DSRy11/wlFaLTtzlhiMSmK8blSimJB
zZRP4bB8MS0UwQgXhCZIX9kNBScjpd6uOoXKtb2iFwBd0dbv9CgHSEQklj6pqpwk
xW6S+FHKvu+Gb28DVCWkjwAC9/n1lwLtJkWlNGJRWskqmPdp5whEWz7ODewT/laR
g3LFBvCS0ERtg98wrFX27fuB3T9TE6b6GIQKVWRZMXXt5MPtuy9NGFsmt157BIOS
lk2l14ptJlWqViK6kDAzWHz1TsGC+LRze0CJCgwX9gPDIvrdm67hsR958aXqNnFC
bmVPAmy+PkyqCaBe52E3xy40lfQrAkfMZ2XU4x8Gnuos0ImrimFUCB30USUGmfLS
Orev6rQ37CcpY4m2fgL+EfnNrnxo7HRenZxV9GKNhlBl37tzEvtCaYDVrb14rL6N
yj3GyCp+o45J+T4JYGEXWiI0Lns5iNCH6ri7AgqW7bRI6IzAMsUkJ/dBe4fOSrRP
2crtLZkpcqVU3Q4B/ic2HqsrQZCc2/De86uWqn/gzKe4CwDV2JvGWkvJz4x/c4+A
V7kDZFbnzt8NEHvQWY7WjNaWGkQamr7xImJsLwh7Ot3vZOtDy1fDiSOdsCRGAshi
sY3/CMryeq3k3a4CcoG3LuB8tsBZ1dG4CBjU4FaMyVSSD0NpfoHgBXTz9h9eA4bI
2B6qO0uMbdFynTXL+RE5b+LLS1vWbtpzZASu0BICbvIY9ICirMUPiJ72U9SON0R4
gfYN/L2BzFeNVJV/O/H3XKd8hxicoVWxJuaE+d82wb9sRno6SNa7fi82TalRUptF
M0q9etgawOonGpLSCH7vfEQxQepzpXTriJDGfq1bmnOsqdYe3V0WpnTL5vG6OeIX
lTXcYR1esCrohTpYhYXISx6TZjzejnAR51oo45v5BBsa9WEtiaUoP7PiAPb+oFfr
BR4giRx1cGulDwwOFqG8b76mtjUOvLpCktpnpWTMCS7iwvpAVZoYLv4SX9GFH+nH
w58yZn2IHc9r8wHhx72XZNortrKp+w+SHXYVRltj7n7sdpkpNYwJkY242TF4TQuh
Q2Td4jdBGmrW/Sk8ynmKUNlX4wv9H9Zh5ZoZU4tnKvXrSoB/ueaKugAQ2hjHWoBp
Z8i/PK0+LIpWYVMOQ98sZrrNBkXmFSdCaEkxwbmUTvvEg6GIR08IOR+HWvpbnZHS
mZgBEnSLGjxxqowb8LbUWHj3yZuymY8/CEBWF0WnD0mSYnlDnifdsLswOOrZX+8z
DLm2+0jYu1CNGKtJILeZg2DOhOcyz76/RMiC0MjecVmURQDW9HyxD/X7lyXQb81J
IiMUZ3i/aPIKeADbaOJjSYmYsf+Zw2ZpsFhDbkWoiLLCPcjLrJdMaaXm0I8YAYDh
P35l/nT5mzRaEBLP9eJHalAJqbfdkvngI1wLpwEJnLjaYd1slITGFEaRkg7yAOq1
vvwnCIsfKLdPWWzCWMOt2X9FMyISL7ekNROi+BZNDo8ctDr7UBsJygN4A8Nl/hpU
NobkpDJl5J5dqBELiz6OFY1UsK4i0d44syiKqqFZHrHb9WSmdDzJd34YJJ7d44zI
FRsxi8BKojNWaacx65o3Mw388urW6uMQcjcuFRL8W9oDje5Mya+FwNGj2Jxu2x9Y
2gvbcJ79J144uKI7RJJsBXHEz12PdrVwXVgljccQwHheVzJHq0+9Oh9fMRTNp2eO
92Y/n7AzETulKpNfRWc02/JDCXQWU0bhqubm5aWVHdYTPJrCCjGsRgVzrz8mffwY
MY99EEgBevMtqjfMwdGSkEF/wDBDvUFwKjJGJ8ZcrHZz62gokpDp5RIdtJMywXrk
ufVsV8DNzAxcDrdBsAVmtU5NXy7OmvDCm9VYo3AbGBw+5ZlykVHZEfveDFffQsiV
QHfboYYWSrrqz/hlSmQyDrze+nFr1IMjXGjBE49Qc0cS+dMh7dBln9W4Z9RZsupV
Yx3q0m3RTmQ9+n2V7ujtTIB0bRfscTRKN2mK7VE2sjiPatq0Gx/91IPU4gNF4vtA
URA0pz6BVWII9oKRuxyIdWE5va1CczqRMVKsDaTBLhEiYh0aP6FEy2YdPc1Cmyzr
d5KrLx5Jk9snSSdIq6GetROAZlfi+n22MZCA4UlZRKZw8VcqhrcRPzwsVuCzPc5Q
mDLVG6o69UK45eOrIAqvUqdlL2562fuvwcG/KSVkgCt6A+0be5bU4YDuTNDA72/M
P1K+F3QXu4Qq+kVx9gDcsCOMmkQd5oonIWxn0Y9czGn0ANeXUQ6Rgm3ZfE2CFgPn
2CwcCtPY3MoIzu7FZx4RsGC/8zmi5I8nKvNLvUQhdkUaEaEhCdSRZ3gaypqKuBBS
NRY7wbFM8XmKKTFmt1w7lQWHEIk3TE8wB1ZFnqzWMMLfXoWnq6Iw65fG8A30PQWb
o70NGmVQByYQax6w9mI7tafoh1w3YGTlsvWPJxL3ALkeKfPnw3h0QA4HZc0As/YF
aXXDqDplUYX83tCa9ht3zAWiwdfSXliHO/MnkZv7LTrm1H8QU0OWDHHGFtTHCgRL
FXD+qo0zhyABwqNEEdKZu0yf8VBPiCe6OSAF4SxH1V5ySKiUDwP4LaQQA4goxDOK
xSOv7orN4po8r8uNXTZXTVwrtTUq495yyIqL+ZcIZS6KjeTF8JElNK7MjFQ1QVvE
o7nILoOCHtlcsx/D/+L+GUVV13Wrq2DOK8qUbuzyXg/ESb3Y2rDP0OFYEXL5UJpP
TCTPqreyR7K8Hj+wKaPxPVvV5y3UO4NvJHY++75q2jZkTvUJ+vbckFBSPtfIgY9j
GHnaRGbKay7opeZx6VCacPpMoC0JTji2dODBHA5gxe7gZvNyD17G12vYcyN/yjmu
uwxzu330sBkaHgJA7u/46ZW+ehQLIveqjEIczWrcbfzo+LYMijbJ8e88L/cd/M1P
9QzXCbpH9cmiJq5AQ8SQLbYI14sXQ1/LdSY3xt1ajdb3+kLuFuDTkanooHhoJHn9
ZIrNEHPKy7UxhLhu85yRw810lpH5Bwa4ErGskqCqyfKBUMDBQa01keXuonux9zs5
vNUpbRqgC9MvKj6OBD1kP7Q3wUMa8Uke1Wj3RaDKvkAzj1Dpg4Cxi8Vg2kH0DZzK
UAY+ErbjuaLj3XCkTc3YUKFa9uIOu4ZeVOsr+3RfQTeQ9Et3S5+4oaNDEBSW442H
lF4VrOVRdZlTxbQc/0K9eRpA0ElaolkJl3e4OrEs9/f2MSC3lGk8yRRCrLB8nXDB
SlE3KyjhZB9iPgxz/9VAL63qX9yLSjaQ5nlnfaWPME80CP0OA3ivQ9KgIydnd5dN
9wt/sbFbVjfO23UriI3mXmNSa0p8Q4sibYEO0Inw7o0R6tHJQRXr3JNuq6YEc8nv
+XhQ/IEdfcspA+axJyfMBbkLUpq3l31MNyxcg7pJW71iAtCWkaSDlAYwI4ABdYMb
Y//DvMNaI5nWQomIomBg9AlklVE2vKdspf4+L5ixyfI6UgtBHsVPgmwGHtA27m1B
jXt1rEoP+lmf03j7Wk0KcQ==
`protect END_PROTECTED
