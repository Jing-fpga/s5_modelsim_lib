`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3iqYG6/vziT9N4DFuxiVhHTJPZviUIR8Zz2+N0Rh1XyXyUVwpRPQrisLeBAYXzNE
sKcZ4yj/touicKufwCs+BPcPCg9NjKl58y7uKMVbnfde6FsmsICP0VREaMlZK2NS
j1dR9fVJttAXJIncTUEJ8uxZhKrhyITXRNfzOAWjRJtHBdw7kAec0ItTfWaqFND8
k1U+Nv7h4xD2xi0IaJXwjEtjy7gGmdW5brmxpqHhmWP9qmJc3c99JMOpZdbLoHrj
+yZTZ5nDCkhVlm2+RW+/6lLvI0MZD+VMGgs4/KVJucpAStF6MXnOeEhBpj1B5Ghf
CRLx3psUiaH/xFpkasvKzjkMPy5rNYRRKzRbg2pl/GK1ItWyLrKqdD5B7ZgnKy5h
rhf4EratZ83wSdD8rKeVxvMBBO3+BBSRMVmGdeWrCrg1dRKnNVCK54rN0vztd6M3
50F0Af1dIyOP2cAm0shp4s98yVqnJCS1W93Hsr4D79k5YJfqlHPFqM7V0hDfSQ2Q
NrvpaO23wQc7Ug1A8fVokoXtWTJnmgzndGQS5Ig9O23PuZ+snNuaPJs/ImcTJKpn
1czCBIzJfFdIEuxPY6ctEPZcjS/6V8J13jhiK4uZpKj6YfoUtWEMviy6FOL33O02
6GhPPtPq0Xi+nLEKYt8Iys0pPc6SeAU3sMQJZ2VOiFKWI19hLKdIO43dNuHt6SwQ
hou0B3hXNpiIfBTzTBbssAprG0BJzONOI/vJNO+0tbpzDtcCwyCw4JqrH0W8k3KB
StB5dLJlQQwhQm7R1UUkrDRmgrx9E4SC4hGRSobtYpSJ2+EK0cu6Qddvs30Ofl0s
ssHOGsqERcc0jITuZCHxyLFFi4LtqNq8E5lRTQF3iKjFXA76EME20iosOmu6GFvC
nRYVdRMh+opceMKPdhQylm/+b747eoHWCYufk+4aQUSwTyR55Ew8S04V+pSa8/HS
izaxPkLC1C+oMB/RUas7p4wnEfbCV3Zx9oJRzsVMW87wgVoHZEVbSeVM6ljdJmJ8
nztauPuJ2QdbeOF/YfFqoWcp6Avmirj296XW1HwOCBRmli40l6JmeZqP08vVzg1t
zRLPCH0+eQdvYKjZjBUUmwVgBSqRcdO78SreLfbOIqinLreBikHEe1iTyJO1d8fs
BBPBbs4P3mp/qNwV7fhn4CzW8qPWaAsjIXgOQmWtDbgyOwTooAabOcElGhYn8wPn
mvAYqkbZoWDhrlg0ixshAdlt/UZL4+IrdqoJUJ3NGl+tSZSxaYYjeYJ3I8RPtSOe
+3hrtqrnWnJKWg1u3wjvVWfCutCQpBCrLxtXP+fBWrDuszowHWGvC4nWCNOjHABh
xyZ1xpAyzhK6KNfbCbVEJiAwGQD8BUQzIv6UyrWUk9JfvsIY4eu74lxkF+TbRSN9
KF1vK34GDZLbv/oahG6AFkGjObjWLy7mU15KmXDl3qbSbh7lifjlw0MCLSpuVMrq
xIYAfl4ny07MicsZ5C2+E+GRL4CtZcF0khhaccGGyFX6wHtCi+Rx+NM2qz/XUhhu
A8PdsJRiWw1N9cHf6Tq70/IXZ5HSNBpxZe0u0KejO83zCtju2tum97DFnsbO6dLV
nD9rnZyXXrDLhQsNQrV7iS2CGb0Vz4ug5rHRTPj3WZhGMjZ3EGCacNBMXnGvgZfj
J5HKvGAiNMFcAVMsubNea1WtVYQkahEOC2ZvkWbPJdBy1o2FPVTGyXupeCQwsE3U
uhh9XkERdNvc8kEXMh476+1kgBXIT7Feu0zBWt9JaL8f/OK1jmDjg9EIuMXBBL6T
LAyEH+lwF3jtJCkFJ+DA5GB8q2j3torws6PlEC+4nD31rz0EYgnTq794BBgdsBlt
O47kkdeFSg4mgdNJDq+1nYdzx7dTcEETIiOmWnCCZRs+ozfPL9ESTVvCyOP+upMu
2DgjEKtdImTa4WCZgUxCu0GvStwWBwGil4k6xivXa1ANjH17XEsuxGuWWUf0nZ/t
cSwzCuIKax1kwGPhNSkPM8DTdu6zfgTrkkGmj5mtDzYmPcA7etVaOJwaE3ANC7zy
tUCd62RH+UPsPxZznVHZdWwkEXPJ96+GwjpYVGpDBmxclouXDJhC1Bw4IA9vH0Yu
VjwKvgqtLd0OWOoMhRXmWHYt9zCQR4w2OcmAclLF+z8jdrEUh9UTDjGUDMxMHvGR
UJOkIVYxEb2MqvVfL0Yi29ViRwjCGgb/0WVVBbK27LgSFSeKDJF8Ult9U5gw9Gnx
UnyfwEZHUfzoNn3DhNvtgADgcVCZZIDB4J2injFjFhy9+6EcOaJR5CzlWNojzm/d
IB2ti7X5WNOWkU77cawM6Gsc0+NyTnemlNYCdgfRUQ/H8hQdIv3W7lpNrw+tGXhd
zz139wbQvC1Q+JioMRgXbeb9E+Bt8HuOmQbMBBgobJ53ihmIS+wkNWr5MyMBYk2n
0vZLzc7zHkzdGe6NGYX201pAV9ZpzAqRahxH+brBV1NMgXKTLQquaM2D2Nr0hIaO
ywCQ6B6jIC8OTIT3wygPmZamnIo3FXek/MRzBqhfTwIpqn+Y4aInDpW1Sd1WTJ/c
N7Y3cXrnQa7Qt6RtBzFqSVg/YWjBWZyu3rti/tLHOpiIBp0LLciffmFxpXodqGbA
jv67Ju/ngnn8rSOfCE8qs6ETlFucf7ytkCRwBDubmB3xkoSP5vG126pUBdQRj/YT
VR+BGKlc/T6iS/kY1NF3pquIyJ7WkgV7zJYNVbD/TSJq0Kj1psb/yCxq/mokv8md
8z1xrnSR0sZ+JH5vYnNbcIyiz7eEBMUmNKzAoIRikI5nQXAaFGf17p0onu27atQU
2HdfuSp9ug7RiZQQG1KGCvd7pzKJw+PdU6628MraBh6l2oP0ph5aKGZL+83+/AP+
ItNFl/28aad2yc/xaTp3KFglGwOXh6W9JIV1VUwS3IJE5wuNgZfu1iCzUCw4sWa/
Hu7/Qx9mEtSnp6mPnVJ2QJoEiHIL6FR9Hq6WYQpj9Aye3/Ov4CcRH3Crbtnu1rtl
GOCoPU/4eb2EoqNv+DxgV56jdsa9o+OyQ+o4GSU1JyzUKxnVPQD2ZlR1wRGOUG9H
TbahW1O/5ZqG9j7tjonhtrq/JV5oeLv4MrpxJHRgGGXjVupqQlwQ++i53/gILNZG
raMKenMIGzmRcNN6ekn7cmDdO4hII7r9zJ7FwTaBKD6vS11Oru0fBzF9UZRDkI9P
WlgOiDc2qj+fO88DeJcIojYyouppI2sbfGqwYXUzWyNx0AMb60ob90Pe6EZ79aqG
RypyL/KSQ6JSvvSfro7N5JTR0wSP9pyiFtWQ99vApf97uLMofRT0BMRzuSf+PyBa
TjuJcpyXwb4OrlrMTOAUOFFj++y4fsmCB6cumTcJm7I3rM08/IQ6FpOD13vVCFgB
Y4SnguDxUt/mncMOXJ4b8C9rHzD4z5LkQsNHQ9G3pWhdj0hHxiSww7f/9XUzUKCn
vo8akXICesFzvcjJSXFQJuZtqb/BYzwTodw32weVtsKRB5NBpcefikIfBl3uvRjz
E9WFo0AuZWG2eWjgeWaALHHCr/X06uqTuoGGnHxwtT/vilqywHtqUptbZC0AjHAu
bUB9OXW8CijmuH8svc9bMpAvdf/OuTJTxk8uEgYCdK6u8hDJ3ZPF+N9ANxMoB1cS
xjakkOrA7cQKsY5yR294EorCLR/4gDgdvz/AzDQMukSM3UVIjf0gLPX91raasEBv
VLpWvbwtzzkERNiOT6Gouv/+bFeVPGRzkXAduQjl3+O0wFlHREHPfJZ8l4fg2T0S
UkGvV7qOXAsByp4lQ8L3fksohtTjMGCE6tgcgxA8sWsa7EoiaxohahIcGt25x3qF
IbHT3g19dRPBnXlny3CSO1wmWGTQB6OXGH9rougn4n35Hv/fTq8C9a4z/ea7z9bi
GWHnkPIuliX5i2dx+vFW/oqTHHTs0w06h6XOZo/iipMTI5II4FTe99FyGbi7BjAk
z1hZrJfmWd9vF3cNBOrMDrkD7mCEKkXvNwlb/ruDx59ZadTqiVSwWgxpum9opd7E
2mko/OUNISXPRJiSvbMKa4r9WXNjrKldc5KjwDECOkhi8C0+tEMUXA3rR6F5StQC
aZVM404e6sVwHAdE7qkD2/wvyzZzdV8aiylNTkNH9QrSi7d+z9gkh9QlQiQK8Uqj
DHQQ9kazM98/wb1Z/HwLNieV0d0fLvTfWxSZshHVYc5YQ+Gr2K6h0JYBulf5JIN1
`protect END_PROTECTED
