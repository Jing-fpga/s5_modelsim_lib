`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g6cb7e2/fdcKlh294VdZIoLYB0zx3iI4qxuYrx8TU5hLPFP2kSuWJ32Zv3TS/sFy
u7ZpluABQogb73ik9Tvj9D8+0I6HpHbTID5owWL/7g6B2dFa6V16nB+52IyjfZy0
JkClcevfCEuSH3hcG/w5gmxb+AXuQ4/itoy7ygIBR+c3Kwuakt+mkfHv8lCNaGdo
+20DbJJEwB3f2iwHjCkrRPxtxxKZ6oxr5PFxdWk63MDhBG0KUDH8AclgPGZqCBi4
Pk5UVjsvuWxeR762vaixv+v7OzLMXGe6kFMdFXhA+KSWM1lJL1wdn7aBLQUxzcUl
/6QAoR0QhP4LCfwbcNXhiohwKJoF1HSPkGVVObKljW+y3z9qImakzvt6w9vpXpSu
ZalWXsexnxomRNO15ptyQVcNbrbia2a34UxDXBiImWC35GHjfDQgK/njlm/f8whn
qPArISJNdkUEgHLZU7fzZCSVqSVLnbZ9kEIWNKW/BGWAPih5xTGaFpcC+RDizTIZ
GUzuUWVypVwCuXsPGpaE4g9KxfUUmqWT04cIlJkcLMKe5SyBwJF/jvoesfEpsAC+
EY9fnKmr72fiElZt7XJgFRzbCTF/8apcRwt4xOSDjg2/MN+Q/x93LxkJOsQRwcv8
lIFpDoHi4z47IYl7s/6S8HBOKV6lw4bwmtpxgPt/yfdV8lAdREHGsSnQ6XiTkQx/
6Cy37Y8P8LQbzTVwY8pU7CrW7X04cwnn/BcSbRxOYYOCfglHNcdxGe9xkfnQ09HH
LO9104UI9zXCKvJ2c0TAFV9bBBEKjvSAek2Pyi4ZYcgfKPae7DqRI/XFieN4nudn
CiyM4QKYA+ZFRv3nbFHLJaewwtYYjttwFHLaoMZKFpSyPwCGS4pmQQMg0OGA4at0
nBgbTbGNq7A41pMywIfvwXM4ZVkFdA+eBSSY+PW0QuEDtCOCkjGcWUVcVA287QpD
lgz8n88uKC8CmZiFFpb0RfvHpy7TehlpLSdQt7CNDC0Wkg5APz3xoNk+FmltliSe
/q01+CP4831EFaUSp47bev+PEaNwoEw2xDcVzwYDc/qQiza25aQrS9WmhwatLPhh
+fVSqE+26mC5RutQme/ViMdOcCxSdzYVYpI0oDbdhIds2cayJLSXmfnRu5/ED1Fh
YGbspaDdrIIrENlxCOVB37+I8uUbdkiJzIwyYKJrLZPmDE0azP10xSg3PnW8OdbR
yvCWhoVo7TvvcTuOO9iTC4oUZ8I91t/IoVB/zkoWogChjhEg9zRQhWJ4XgK0YNgl
pAo/BQVnpwQ47GXmPn0X3oKM0bqxYXzmkxL8vTW9lA+2E7Day058QxoG6hY2lK2N
MrHfvEg2dPHyceYhJ3E3uK7fZTiQzZduAi6F0InVVcA+0hFhWd7J/iyMiGc8HpZc
z878YcKaNYsiGJeuuc7A0+AdGflu9K2K2RXUUdvvcwJSlwybYjpRpgoAtF/PYIqB
2DLVp2WjEfAsy/Io1qDRwuc+Y92uweVIsfcAlQ9GPfYjIL4udFLCWz69L2E+4URE
q3D3L5qhHjJrYnzaQ7l2w5flwXweOywh6fLd5AcB4W+rj0/6CGUxsTqL9j9VaHph
4Al0RYh6ZZzHXtadLNsbSqoOi6mcZtL73ARpfYVJfeAeygVkoU0Pc+4UVkaAwF11
LR3RJQbaKGU1Tm5Ky01Uh9N1rAzzlO12BEnhwq5D0DZobWZqB7f7OEXaO+a7xD96
3u5YvD5cvhNkVuUwc7MG5R65EyJ0n91ayybzcshS9vd+UjhOPhLzVVXHF7818sCe
EB2O1dRw2j1Ac4JqU1X3GJGXwAP/7SjcD+2p4JGHOljmtzn7LiIea6tTRt+PcQPG
0wT85lANAsibH0z4kwDO99sih/Ax8/F54JqEHLxpaLuq5um1A2kK3iP1xutzOCOr
oQIZNMdSzAIn+146qqWQkoXfuznjwE8XNO++ufj1cO80l8fyyAvuJl13Bw+df1a6
W+Oxc0ivo2FzvKtYIaMvkbaEA0PrYaKk1QiBsrLbbVnUZYz8su/5JOg1Q9cYomP9
cQfIxSUWjWi8GtFK+jwI9xyAVw3WIELs2msD53XhDGM0w7L1g0wvnwGHDvFUp+Pp
ROjk4BPQGRnCK0M6UzWUP1pgejesjWKX/PAyM15lCiLD+wRXGFK7Ys3V2QVJkTEr
rLKAZp9jkmqnIuaGKdbQBDhEwwgLZjUk38bXEcUMyDssvZwGGo9//gqh8YtzRYUD
JUQsiGrV3vuiPRZaPOfvudt+Bt/eh18YXNHESoGtmrA=
`protect END_PROTECTED
