`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ejzJ2MmNNm8RHjBta4RvfsQi9DiOZj4org89PTUK3etXZBVtdxMtRfVL2alOiSDJ
uSwllHMooVWJGjYRM6SM+7uAouOKj1DJ8SwhLysZSOgy4NRnRSh8+ahPX9EI8sOW
CY3qjrzW9m9qQDrs53J5kr6ZJyXZhVXGQdIZDCQUr6FfmE6YlL1vJPwBCxAQ8HtG
390zqpi5yzOVMQqHJt4A2JbwtHOPhnImSDk0mx+sDs5yNmjBeE/jMbkRH51CQngV
IwyA8oLoS9SpUuKhTCwom4FDuU/W3rPYHd7kFUhU6rvd0umB+RcatisGAeNvIq3b
adyS1kV1ptWn0i4fs8X+8x4KRI+aNElTvPN3HdIB9dro9vGBCGB8KNG1K4N5lCZZ
XyVUPkLgeRR09PO3F68CDZ7iGlF/+sMCExkP8OEiWrWQKGwtZ5H/K0oyBCdqYU8j
bipS7ag2F62B6WnJ/i8skj+8KtGHwGxAMkv0Spa7+4SMAGw/0aKP1mvlgqML5kiI
Nhnc4kxW+3wEjpEJctRk/1u8U6Mnp2u+4Y5bdn1q9TTe5IUAXtTYC4BZr7KHVfMc
wyIevyzZSJf2lD/pMykXvZD7la4BKHP5NeWrsFbSaHas/IaiI1BDbeqpxHRkZsef
mnK5riHIsRbS5rlY8GXojR2XeKg5qPsRGxLIzp7I3QytXrDoV14tARV9qkSNnO4k
xRlOVSpBNFpRd6XP9PAqxI2Epl3Ui5akBqD1E1VgTA12bShX8AhbDPl/diiPqxdB
W71qfI8gVB0uNfGorNO3aR6DuG6eQksC5W27ZXmB50APVtPpQXNud5yoCRlvSH3C
0ns2KAOf+sQPKUGOoXi1A6KfaoX8lo1L4bY/aEUc2d/X4MLl6rwV4cmSwTpnU6KG
zmTwzsEdH6LiBzQfbHgHDXhS0oEfzkFKaCma4ovAneXcDyBiIJ0pMFSga/DBAbiN
szuY0BmxNpPrr9myuGCDTo5rQujJR7T49h50I3VgdFDx6ndNhocazktl3zflSbh0
gOYaVfZaH4E9T6EILO4bZbhFOAWWpsPgGXd83w3V77bWAeY90gszyC9BBlB9B4nz
y8EHNs5Kyym8NCnkryLv/I892SxcZ5x3b06s2gGIpNknA73Szd4QYQ8beKBGFlB7
RrpS5RI4mDeBLIbQ229Qq0/LNQK8ZfgAahBcLNyJZ5GKni65pW31J4BOvsLlRzmW
vaMfnJElvo0p8Y4245/a5elZJIhSls2HMGhCUqBwlsyhcvSHsXXdxwBqN8FsceRR
UdFVyZKJ09TYP4Zkd9Cjzvt2yORZq6P+C+xlRefJe0AI0YyeRc7nt5hJPmWlNogZ
87zw4VfccX8Zr2+EU4n70vvFPwrBEVyYnJUG5m0OTIyjPw25dD1pDhgRlXk20Z2R
aMyIZX4EevHLtD052yuAelZ4ZnnO9Zb6Tw1Au27IFjn2QhydKNEESN+Ynt6ufJXP
YJtShr2XPSjOyQYwUw8hFW0Rb7Fyh1YCTNpHBViOnfHmCxkBFKKAjIRzyheXoBMq
5bZR9DyImWJqzmPZlzX4GMTO0l/QLW36RTxbFwUScFt0SIOQ5I3yqC4q722+ndCN
sTIrOfaLKwcAfhOCoRvjN+9ctWNxnErukTabNn5CV0FL6JsS1xAjrU/Ruc2mtKKH
q/gQ+xH5HYjy918gXnuydckRhrTb9fIsWIN6uRY8YMTdC19i7gUr9byACx/yicnV
FETroK+uBvaf9+ps4wtRgg==
`protect END_PROTECTED
