`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hP+1Hrnoh1QNRtWdhzx4PcYOYtF0M8ZG/+Tqvc1PBKDXe8/uqaIxkwmcRb/usP9E
Rk/vDzEkjMYP0HzqFSdaTqp13ZVPkUzETb3D6nd2aPREsKscG0NWYk1J7bsYMd7g
/kAaULmqQCpSmp7vPsnMPMHySeRlSABBvPCuDenqA0ipUKf/II/H0f2ZnjaFEGgV
zk7cWz7sK2iLiba9PJzwMHd+EMmbf92F1OQaww6LbbwqSCXtfRMRGWuPyhqRniAW
RsHEo+FOqEskVEJP/BHzdFH0K/G/m0R1StWv1ljbEAhOsC+q2ZChxoRR6vZY2j/G
4fp+6HcJH2gtUODjpcywIfWmrDWiJv7xSEBNBaUiBr5CY5WrLb6TKjQp5lF8hLmI
jLtOsr7z8+k6820NONbkhhAMw5aQiwe74RRLQqCY2Z4m2jQxxJxykGE1cRMUsbGp
D20w4XQLy7sBgFX+br92o32krrEYrFBrUnK5pKFscQ/CxJkbH6WScTjlVriJhcc8
yRQchUIJIaZ1ccPSrFzsAqEkLD1knSgusnuBqYOQJf1oPa5TX6ls+IG5OjYJuKnS
rMsb6noARj1eCOJfsSdNMFMYKceixDHOc3e7XPj7A5A=
`protect END_PROTECTED
