`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eNAcNFyFo1o5kRbvGGTkhoeJ08sJLuxQMnDxuPo9CX2PB0NiwEX1Hi4UgmPqxl4Z
hSe4kBJpisrxVW/g4ijxbZprL1RuS0EVpyG+N7Zk7cCl7YpISFJuXZdFGvpFEPeB
cbVpPN2V+Ie1OojZSNwbVjSlC+bsW2Cr+SEXQ3ZqxOZotFZcpGSzy+pvRINGuQOR
IHoYu74A3Egjj5HinDHFZsV3NXnDf5itEJWJQujWcXbKrZEJkmeahT8wa6Gj6Z3V
ilhPwT3+a0L4CAbflJ27lbbV8/If0g6F6MxVjiVNe3xmGMok3Dscz954AfvqwIPd
PM/8GcdVB4JKuSVhszcZiHX8JPMSrk4tbuktUEXsGy7ZtrwUGnlNZZxpgtFqjXvp
tLx8zR0ahI42NzhIf8c4h7oBBFQ9VCDwncj0hew+BaSPx4j8psuBvCk/SzbHfd1P
TDbSnPsWZcWATLy2Mv4bz/1FSUiM7n+pLPRBIdFltsIg+iaw/Jwlz4xOpH6TpKwz
f6M/j4de09c2oLJv0N26QvSIt494wWfmxwo98j7eIYO7xC2UHv13PoSQrArJ5UF2
sssS3GVzGrZDcVnV7uPXPZ+dL1s2yc5HyO0sI012j+a98QeCP4Qe45OA984pwOJI
Gm0mwgDSCT0GFn+QfKdoyTtmcLRMuh5RWu7A19CFSSef/MDmwE8B+7Gdr7Y3bt/s
9+vwT6FldIFArxTF6WvwrJlM9EEfx9hubixl/pbFN5+MKf2bc3Jm6LUTaqncCcMJ
XXbgScok0Gx7sXV/l/49FE0pB47kgcOuDMWDb9FvtbtNhRpi/KM/ofK4MRVQPLJn
nAY+4cw9Ut86WXVqr/swGzPYQ+z++ym+oln2sCsZvXpdG4UXzfRtpRWcu7R+2HFe
klN8zFncvkUnVQw9WhS52WTGyaECe56EZeCHAGN2OPewSMXGp1oWDbfpIV9KHd7v
uuCm6JIm1yjUY0DfVCG4oIqVlV2Pr+8vyegrbz2NwJkeOi7Qr+DwvULowjNSMBXS
BgD5xBQTY9tCzW6AC1mzRn+8r3KCevTc3G0XLcApYu3DY1MgqKXJ9MZSu0okYiB0
UE8J34QgPWHCRoZGdFe3oZz3qsmxfp7mclb1nrMuBx1BdY41tClAwVCl5PRLlJys
ixFi83wIjuthZxnHaFCahLBYiJ/O4g9O5t0ERIbl+nW8XpN2YRBG0VbKyCIC1w14
4TCGvmGU0Uj76pmDKWXLY0UxYvTlsdGA04DfwRtb4Z4r0t+iNzy25GRHZh0Rbwbk
UwFVaUGXrNA7iwiMM4+Rl45UiW43CAHWXc2h8N3aucEXuSZq0j5q2IME1+wnOrlp
nGD3CkzFLRCZfnBF7lNbzrsAPbvYl8GNhqa5brnyAsy4dGoGsmCU/FrsMkN3U2G+
senDqjU6AT9/E2mPMlKIrhBzreZQXP4CDgvSPZg8JqDlAYPZKzQsHXx+ldF1eG8O
HtuBoAEZkIuT9UhDup4ZGZ34tSjD71vILeLEXt4SSg7EJ/PzAclBlacpH5QeJu+u
gOkoJJt4xVlPjEjuWOv7IDa0teixIgL1MGV+bF2fSKeYucI9Y295i2dSK4gawHPO
UH4FIq0hBosThUPfXeoWiKC07uvKPRrNKqJVshYYuae9N+n6OiS5he91fFxEuv6o
TSuTvtOSlrdZtfAGhWiFTJf2nOJF33O7POJ/6nXj4bEOjveslYrxadvqDvbpuvhT
Y03XVMBtN5dTxYyUzO6HQLINyFYFDV1MVbhkIkTE3wscUFdOZSJ4o7NfW4f9CnJo
YeWn76gXgsly8hTtT4RPjCcZBEgn/elWnDKemIUbNiw6NomFRYKa+dZ3ySl0DevZ
j4Ome+hC0ImkbyKhWXtYFsmaBgADGWgrFpGBTkPZkwG/R8OaoCocTgKC4EGgZggu
rKF4Gw7RFhX3YTQwnKs1cmTWJl1nSMoxBxPoVsDcLbgs0VlzpV49vQIYZWQBwlpz
RBo8S8Nh1seZfPqe7+FDKlK4XeVbVzo4r75A3NhnEruF92y26ffPIvpJoI6VAEpH
uA1cS+/vJPg2JZCQ63tPxcaDFO1ff7q60eoLq1b9KVTMFaIekI/QtU10PB95N4m9
gxAM3t6jeOys5BD8WA40WdgUB33ZT7hT6bu6jrfdWYxVECn4XCKf38AwInhZ0PU6
`protect END_PROTECTED
