`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b150utMy/9a4VLXgAzDoVhqE7w0RMlxsgTjPfO3T0pYjfJ/cwYKN/eGQxnQEYerz
PopxP6EPG0N8KOK/bw6qf0SR2cgXKBW54EU1H23sDwqqU85yePsnabJIniJL//5/
VjjgbCx6YsYqAh9J7WusYf3n2jU18fzkf0LK7VRZSyieuZ7yTTY4LNjmT2G/8fg5
f6y9BnTkmXIlzChC9Ax1FcrX5u0HYge/Nf8NyHgUn1yArPMLmtNQaD+hCy8na87Q
k5bWMc8/zwq+ftWHA0ldUl/YF/1Tg3+aUVAOx2KZNudFPatrX+2fmhMp6TATF238
vSfQ1EToQgX47Fo+9+BZjOATw0mXsGdRn95Y0jGe4oCleiZwcEbSn6V8Rw2QAGm6
imoKs3RA35qlep0mCi/EJh7iJu4fPqjw25Oboqn09982IwlIhnY8IBM5h6pyDYh8
o4tU0D9c+w9pJXe0XNC5x+AELVzonxrkaBKbCaMiODo=
`protect END_PROTECTED
