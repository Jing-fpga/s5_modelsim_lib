`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JjRd4DifyMbrv29heRd9azH7TWjtWhbpIceRJ0eSBy5Lou3a9Cid5up8ZqzO5Vle
gdQJXSbEgV9jZeCXMLLwl2aSucJwjdyPQYjoKRtmzK32s/J2v8C9OBGjfP/qaP05
PRPeqlZTHVwVzw2De8C4nnDbKNwnenjVV6SNCBref+AqwVoLFe6Q2/LMNvNeGmzF
472/nbPaQ0BE2Zpm4/NSDqmQqNRpF0y6Q1QMIJNiErfuRvr1lk51esMYidK2P579
68dAI/j5Nf7ljIvvC4+dzQ4XRXjtC7yLn7JpUCVumg1JeFD4N382J62vWd7rJr/y
jACIPZBZE5erk8FOGt4XqjqEpXFcaccUKljdPGIgQRXZeXZP87kCoBH1S77nwMuC
WYMBG9puTefdPpmvhz447tifPqunz78eDFTEr+7pHCT6eK63kT6PSnWdpH84GtPp
w5CB/YjocFIhioL7LT6iI2yzTP/K5NXRl75D0HT5tvRNdLhJTdFv+ADlCfwpdPEp
OWF2sdqlQRDOT8cKdYoQ7L155t3h1/loyi+gU7wusIuvN0VXab3fYOASKFSC4hmO
M8OmtQ/KbxtXt7YnTtzGjz7yuS10kE6SfNy90TqtIkLLL1x/Y7XjO/ahsBn7WCbl
sh2+aik/YfwBM1BD2YMao6tapNZdQ9QToxbzqyHvjuowcb0eBT77iWzh3rYtvkEj
xhE/K/vDYKXiY3HNMem3bisIW6mxPuhnDNH+gefDe2EfERd2ATKSAOlIYP8/Fres
JYa9REjsKJPWpUSkV66BdqnuhUBHXQGRAXc+OiHqx18EANcLmND883F9f7/GppRP
Zo9JKPWSGXuiJwWBxvDxUi/uuPsyxizw6YuglKU6r78oNrX0O18HMqhHq+xdrJWC
6DI0o16OPHzPLaevR9qJdQ3Jzt/fO40Lla97rQ9pWBCbrOk176s+vKq+BLAeWNoB
+tuAOSKhHG/0uRw3MK4P0rb/f4UwigHdE0RH57QAkgHGfSJPWFY+l2PK3Eyi2RP5
ymMmQKS6NUOu0hwJRUdqladMZ1cQlXF6nIFMCoV9tZF65VgRAhuho9rfoC/SX14g
LX7VwoM63R2J7UjKwbPek3O2+OdkYrjKdYm+2ruGr0c19J7TpSRmdZbMQ0zkmxyw
rSMDv+/Ee9MgCA1XmZ+z+EqfEOIjUrHAo/anOquN1fUBZCHxcSeHDFvgRpESaZDx
n74qEV6v7MqRBl5ryGrCcUEM8SOsgIh3nr8YiqtxzNq3Y50PzEm3hXGw+aa06dnZ
jZ0qV4BmELyEiR9y37IF7rof2pW4j+NRRwgM7AHkhZViWK/aNu7QkI6+citZw8xm
DujfbFkDUbfiLCQ4zSqAjAd+cQ/AenbQM0t50N2W42ir/2oLxtc5T53w0SxDr9Zt
yCTgakEaehE1gtnHOU/2F78i9MZbXYjTHGUjRgqLDyGWfNFsBj5KtWEkRwfcrQ/S
qHw9GOyrt3KV+aKL0CSHgDU6mX6xj2L6fAzKTs4CVuEeMKYYhek2EXhE5B2AaYkx
QD9yz3wI80zMk+8ZSaDIyFRAAnWyBGN3vyt8a1pgdtPObs/wG6Y3No24apDQgBWs
kAuv1pxWZ9lKSbLGaSdh/2e7O64+hoVgLaq7H3iRynARLZUTJVFrXX6FjG/2LQnS
aTGe56HhbDC94UjX+/ukQ8FIm1qjt6C0D3pK+Wn37Q3cky66V6EVI7p0Dpo6deui
iV6yRRseXlfj9LCiEyl0matwHZCXOxIU//xzn7VMUpA/3STb/NRh0ejm9MIwkzFA
Q7x816pl2bV3n8BJvyuSiGOLoFJOqdy6H56frW1+ZshJd0FXNxQWhNsvytLAu9ED
icTQcfi9yLN38aCF5b7NGOGSzHYKeb5gJJjbg3AldDw=
`protect END_PROTECTED
