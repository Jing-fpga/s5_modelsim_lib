`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zmyG4a8Rmb+sKcDoCyfrHKJ0Es9/abOzXiA/rkQc6zDkqfuI7O8c6RYZXM+teHE7
8KnPhxPJQYmx6Bn6jIBl1jJaGU2uTgE4as6APeTzLcXn4EZCxwys+mRHGACmot3N
MjKKl5+NJeN/QXIiZ+zeGnFw2CNOqazp6+Jnltwq50cXW3UpNKoRws0QI+T14jJI
c8i2eVIvouPxGiKPDIiMOViVpzItJy7CaBN+KqjATe4fdScH58EhITPnXc/Zv5ZE
Yjok32msuzkztHPv9XFZ/VAnYzmuFLkU8Pm5zlHSzjhozu0D/CUduIKbU2At1/9/
7lpefLcO06j+5zVoVtXOkw4F08XeMyIW0f23ch9TN7iEWYM0u/piUeRvUn46Xwu0
fYArvau3liKusb63hrkg3T0ulBvnqR3nRgyzkPMGFBw0qvX3c++QtvS5qH3UU4SI
shkCz/Xl+8Zc64lzYr2eGfJoRFviiTUt2lLV6UTYurMYOpgsUgtyOk0z5Rmu7UFJ
7Yq+tIZCZeFAiZZ1nrNkkQ==
`protect END_PROTECTED
