`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VoODSn51JWoET9/53bX5aDr8c2D6lv4QfHaPf5WIdcJgH5RiZQE5hizmG+jkRg4R
XwCy6KtnH035YFrQbogXp946NcPXL/b3o2ATUqnEx5Kq/4IL8w906rmwswm7qnrw
6qC4awT2TUE+IvqWgT1cPi/025x0POzl6+Tw6eM6njmnq8R/3lD+LikWhZDVZeV4
TMwKDv9ujek8BPbXYzCrvIwpj4K9a1QRbDcvLC34qiN2cXU0KhM2MFjDJMas8fuR
X7voYB91yq8VcsyFL6cmbnM+RHIF0d7mUWTFaGgp7PkY37dpRHLIF5fqGc40rBl1
gAn+uei91D/STl/cMWgh0efdMyENfB2dCfCP7/eyzWMEMpOlEF3UJx3UxdUCwxMb
cyWulfgJm0J49dq5tCYphcsHUfUobNSy8UO04ZgwrPRogAHNwE+ZD4s+wwqPTMLq
tkF2Nvn10tUQ5MyWlaZ2aNVip6XlWsJuEdr2wbA1bA6IuAJT1wUs1AGz0JRHC1D3
lCdT5SUP4xI7bfEQTv9oRQzk4v7AoIj0qZv2Tu7N0U9vrp7J1xeI2N3XzXlUy2zj
GgaCH0E+OeGAtNaMp/gVv/9htY/c7DsVak44EHdFW0G1g9lzYZSvemA1qToMsCzR
MEHVoObopt5DIYCzJsYvJvwy5IiEFWdRzTCFrUFYliiZFdztz/Ycl0a4cQTm4eZQ
I7motQBYToNCf0CGH4YFwk2bfuUZHr09no6XZGpI5cRN76WM/ZAyS+bOUjUa6jMY
muNlSYJHdH7wN0Aaqggumv+en290pkcZGRy6mglNHdJd3oD2Ya20Ke+GV1mSk3HT
xpP8Jkd2qtzpRRFG+SHUdWKVKq35RfCW7utHroZJjAJk8RaNm5j8C9I6lpdLMiiP
j4pPMfV6+AbzCcMXN0sgD5LbgrzHT0VYaIbBiHgkRN2PmyoY5f3cC1h7X0sxa0ct
U2H6iU7v9lLkHYJYbBM5+WY6VWt0mlVck6TMC8xSDI41Spm5SvXEBR/kF8EQIkEx
p1NswWj4JPv+KyjhYcq1iJ+RC3+AiCAFn+Bd23NlJuH1H8mC8c3oTnRVMXCeIyBd
m7eTJvypsb98tkl77K9xp+Ak5nbZQcxOShKzxCWMyfso/kTLj95o67G5KHK/Ro91
ISZRSreqaAeYQIH9Z+CMEZSSniXl472hEBPO8EzRvApXud7NTna3IFGWghL01JqC
YYN/4+4pSUzQupCxJvLOEC2WRVQ4VGtQd4+fYAi3gfpMLGwVF39Xk0wouXHy9vPB
schQPSq4TUzFk18m39pBbNpQ320i2YpLvJARScCoHBGwncWaD25vx6+xjmAm22vv
94FbCCDw7aRjFGWo4RQFc9PGse2H8DbkpYqiUIFVMPtDrVb69Emgg9TDB0G92KWW
lwSN8BCQM9d4X5PqSn9xfQo0tjFyQCGrxzrRAdSWuodzAWBEUlgkjZAYzhWnSUnA
Von6KZgq7oKyN+JapjWm40mejkQGLUygejApwa3yZwVNn/FR48wv4eCq1FDIqJFg
cPT1Y+b0a9wgu9B491QGxPeWGdno4XhWQz6jPF0MtPYu6K4mvOAPDFUXW2iS5Ru/
IofsBDLzDrgZ8fObnxfa8Yu3dxQLCO13KkcllV2H/2PgQmdhGURt/5MQ/oZ4h0DK
DQf23AKvYsJmxYTZlYNY4K3ZR1SbiDY1JmDgvvWT2OkY3Tr9arAQVSIWaDt5edc0
GwiL5GEHX3fejvTFkjrakBc9n78wdy+wdsSkoZQb+/KDEcRxzyIvwG1PaCiMFRe3
2fulobo7sMx4O1dexfBsGu51/mEnkkCsgphxKZ5icWGecL4lnsRdf1WM8elTl6WE
BMxW+aIo4gc35YXTOrrf3HtupRR/1RNcbWqoflc1Ccx7RgXTODeGuF1OftAPTuUb
ifSw54B0ZwsiV54V/aKVHSYFODj1d6l+1VlYjvioHM+4OQFmSmHyArudP7gF6r6W
alCvX1BYG2ujHSigBUSXGJDKMlBRDfUzKKSoxQFIULbYgzfHVVUty1nEnH01hhvk
`protect END_PROTECTED
