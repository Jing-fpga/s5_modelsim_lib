`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B+qCtmDvfM/rLEOmEaGYhOCuIma06jxSUR+Zey4zizCDpp6bHnmNF9kMHLk2pYGr
8SjIAHbpUlVQrF/dyZp04mhkPNQEuuTcWIKDHMVxVtjkEkdfu+w9H9Es/oXZHQIH
LObqaVOX6AWPMhnSrvk+hevwErQugBX69JwYqGwW2cNqPajoehZucLa2aLTT+lG6
VHS+XIlnkfDlGTGwtK8fTAc6SpYnnDhdTIWmAyGYszMPkl2bS+rxL5X44nI3Z9wj
6Ou1ohkCBeXc9G3LdPUinFT2g5wcxvJRREZl16uAbdsJqVGjlT64IEXC84lXeJ1A
Ydc4AZnLFJ9Z7FhbIzF0+ouQYQe6lVHDSwtIfglJXmPy5BhIqURbWT7lHzPBYQX6
El+DVdWYYktlg8myBNbqvVIlYfynG/LBXsBbqL7Fymwf7KBoNeXwitrqIDTYXnvZ
OY2tRX/YEc1X64hgMtFSIiFS3zA9XJyEUtagIHzheGPVoykkzcUiGINpQAGOhIMA
`protect END_PROTECTED
