`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g1NKAe5A6aXstscpcekQrqn8kUu1Nir2UePBsfOfj5l0rrVLglmOBAcYmBM3jEq8
mm8OekuyCk2QVt1/Fcw4mTKRr4RBFDIO+s/bsua4j9OFDnXoGip9s88gpsN5mU7a
Xi+NvUrFPTzQ7q9ZnlnoBehKZxTmwi4+ZOROCkH8IsuDzvWXAuFHW+wsrzfvAFlM
oViVZAxQAv+tdGqp5OjhZao0giepXr1lRYcPsIW2kMxdITzhxVPISU7b/9kCkTkE
rt1Wa7xuE4gWoYGli5nNVkLbT+ILQ5EV3VE88i9Mkxpaa9RkMc8IG6O9ccI1I6aA
qq+O+He0DQLBH8JNnztH8NbhOM/pi0xrHA9sp5aD+LO9fIb8Vax964dlDs80zDTc
h1NQ7gkI8JyurPf7dmCFRcDQQu21geX23k5Ro4e1UM9KLYgP70z/GQ8gmaTaPZzd
2rqviKSJDbHRJogLim+1Owtekysq1S6jBYZM1iMOjCTSmQyD+Ro6dqnteEd2X1kR
jCy2uFbIkH0HUXlKBXgQPSzH8mGtNZzbAYCelgqg1ITbmgwNstc3pT8JLqPJKYYD
vsL5pueel1kCzEIbSSt33Jclz24hfPYWxsGiTm5zPWPtTu2ZexC//j6O0RfAVCaz
/e5Fz1cUgTRMLQFy8BDSo0mOkTh3Zi09SbBScl+MKmh/6PGFJEMTjiqcIZ2WfMI6
xAWhFqb/Hi14JFGBqVIsYrGP5jTzlGqunRUJFGwLRIP+PEdvDHKa18DDWajIux61
h6XNNqMm7q1M3pZB/HRO6xHe6UVGaljvDQeRFEcXwUnUXiGeXbxDLFOOUChlsLf9
1TCX1tBHX7k5sii4Itqa7wLSRi8/ATc6rPuNtNcgGFloFPyxMPOyfc6+7YZpvT0T
39L9ttnfjy2K54ZaB1Fi9IHyQvsWI59PVo2AuuNcx8RG6IqlbrmVysdz4fNP3/E+
XbMqTIe6A5PTT1ANkEUwA++87NTtVUpi8xSODHra/kQ4gXeD0iQpppmJerzI2vG7
Eh2AhSLGNpmAUgoSHHOY9F+k05SGnRzRZzieF24Pc/ZRsy7Qtov7fHd9+W8YCrE2
mr8in+3zmluVp70uMRyGPUJCg/DAyzywRDdUppr0qceCP+uDaxhxLSVmk5UfnZ2M
nDE1QwkOHVL0yu2APqYRM5qOaq7BCM2M6stq5FYd777PxE0SA13tSvLcsLM91qaY
5VCk35Z5LeV26A53nomYQmlIYgnFHssOFBXTjDlcTiC8dDEt3PdUbZPuLaIjNmzy
LL+TWOSYRo+cGN8TYOGKF/90Olb4UK7MC46GaN6ywo+4M5/9LWI+bH/Be5THgR5w
97Qh6LKcHrbrNsM/1cvyEa0Ewsms9vlIRi72pcB53Nw4ryYyga9hKTp1lXatGXN8
1AgwR5J9k9bobsDvsEDzRgLxJbm0PNhcKz1nYY4xOTSOYbqv380kpEUS879p0ZID
RmQ1/N+WJOyaQHxq9Y5LdOOSek++oJb0FqIzJkCCfCQb6CAvYW6Op4j1VJddzBp/
97zzwxXiXBFvSR0Y5mqYMOhUtO4r1zLOEK26DhBvMQSWLf6V5s6qDC62x+55U+53
KyqlwUYv0cxi6u23g4f8kOIvqWYhG5DE4xFu8aQRO9PJWRzdPm/kWl5oazri9Xdj
tijuA6NtlwQ4vI4T93tNY1wxKhavNzTo6nBIXkfsWK/V5dXsqHZb/D0SM2xZW54F
40uqvrSsaWhOJ6YdRKppMg==
`protect END_PROTECTED
