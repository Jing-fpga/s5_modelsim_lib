`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oulhiz1ybDx0XP+AUfFL1OqV8+4cJWGQ2TvQJtJsrxwGXI9LUjXX3VYERI/Kpoex
435wf1qpNxZ9ObWPvAnG4UJOwoPvH7NeT9wM+d0eiK9UK4T+vrcACT5KCAsDQ4NW
39HQk6LCEKG93U2VkJB7aNQIIQTEschbs0fFwdd4EeMtzk2AZc8lJQgDfsjawNXu
EBwFJTWdTerEl3bzrBaAbQMHArcLlLU79xzwaA0JRrkSTwefE3P6Cm6Bs74RRva3
Fz4RgDwelH3Qgc30I2nb+vwgEcFlBoc1Eh6/kRFTxBGeD1xa+NciokBKf5SuIALt
gLflcQnTu5nGMcVbwcl3JUjTJO8t9zpXpd+9+yy0SXL4ucVvcN/EyLDxVr4GutjA
5V9F7uyJ56aTv6B6F18BM+DijQSWmHiRRQXJohu8UoFiGib+c6VFzCHy2vu1U2Gf
68yDMB0QofnSoZGuzbv6E/HGn1JLkd+tX3y7+Jku6JL9Ydzhm5N5pXfzame82DDI
K/0fAtlHAaPfjytfy+A9mR3QoafJJpxoKv7sDASTSdWxL8vmwFNXvBfR1bJLDiyO
g2TkHSP6y8uTc7SDeR5Ca6s0S0e//avdNS3pNOEs3rW7wEMx3s7kUHy3ShS0sccT
DVL7ycY1Y8BlGxZHR9YSSLNvXo1FBqXhUZKDowrW+I9pvdD58NluvCanzcTwggL0
SkX8eK2oGDVDACZK9m2tzN7WlIwiHdOeUk87IsGImRUUCOWamGPduWQsx8qKFye2
uHU30ZLRpUq7jh3P275DEe3x2cKQjq1G08AWBPnFbWDC6Bfix5sFnYgZrlOGO0at
h1fn+a8kGr5IMvJoYDdnn+6K82mEYw06bHxfkiheJ88xUuD7lhWJ6VQl+9nek9PM
c7j0gWTmyDDWFLGn7xZqF0U1ZMiDnFWiwzWA8XTGsaQ=
`protect END_PROTECTED
