`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IRLhHkGIkNy6fErms0rFL0X4niJVbzSe9I/ywG1GlO4PmJZ2/w4Su8fLrRyaJFyt
7fC/9LxRrh9sk+ZFRbnPsZNqgCEHZh6evEWT79Df0jVhbqpwkE8eeEto2t5bUFgc
uX1g1BXubZ5ozjglruUzdemhfc3xiXldCY7iKVWq2RUj8mWXesXGCg9VBWkRxL3s
A28m6Lj/mM2mFmB+9ZHwSY8itIwU2hIHfO+In0wJ2FTyXWG4Z+UNLxYsGFL05MX+
70GO2GmrPxiYTIbM9JnGzP3ZNenMtftMZM29s/FPOdBZE7c5xK/+giOweOC/wExk
urYSibzUufMC8oMwqzhrAq24u1bZXZrAWGHNN7eGbByvU2NAnI1KPjVQn2Tv2xwW
/GqRPGbz8UpCDk/5RbIrlUSJ/9KEpwsl1FD8ZFALU5CHmdhu+fiRhM2ycF4ssUMC
1WeuQS6gPHnJ1LCTQOm64k8xmoCvIJzrMdCrTlRbII0W+2t6tP8W6LO3T/R2Vfxm
jjdsLMXbeu3C/ucMuHJfLoYg3o7el8poUuKASJeGP+6VU1BVF5qjUEObNTD28UFz
h26TywfQOpEMDd4pQiIno8oUwZcaqSAmE1/uhtPA13HcskzZk/qfMpQ38KvqYeo/
zZiGwTgpdWk084WBIQwWQ+qr6mKHcsxlFuiRTmMsGZGGLabwLvUR3GQjnKYZUvwn
+t06jAcGwPIVLO7AE/abh5qZSRQnW7HhyEHNDFrINPVMjfVqQJEUEcTtKj39K9vS
YfF12AFL3qKOAeGa2rcT+vvu0dLaYtN500wrYDQB9Y8OiSnoUE98jEgRhf5YCVok
CT83rMTvjwuv0iFwMqoISLcVXhynt1KnrTT6QcOOR2v9IU5uPhvDceyQidAOTrRN
2tjBeEKSRryPc2GE/BJr6OwMXGkO7KkU/PeRMQ0ZPpOihShCsC8hZ6OMkDbL2pbM
SonZ71aYVQ9JCgCBjpif3QrrtFbFri4QB5IeMCMwPv26G40t7vsY8KWwwWq0yE+H
yj1ILVnjGx/NpiKxARXnPcDpBzAY/O8g3TofWL2qQv2onXOB8QwkEG6d+LmUWjwP
grc05Wb3NfpFHlBppneXwGvfuwKG313zhyWREGrxQ7zpzTTmojDukNdfE10sUDie
DkfJJr8uBubtpsPKkJj+PRsmJMQp3mlD0bLycvHrsZ4QsZF4/VccCtChr5DV30nX
PrWiKj7fir51iD7f3vsomB/IGslojD3Q7lPldV3WfhtHyw9WEEig6P6oEUm/kt+e
YGnrfMYCT7/AJ8S6tFciuXjH6MNvKr2sU4tfW7T0Pw5Y1YJIlXqOywmqFc4VJibs
+stp27WyrJLh2xLN3sJCRGBLPjdKac5MMG2nT0aA8iojfukoZ6maPP3UYIxnljk1
JViqxbRGCS5VS1xukCrxNhDr0xVAZrm2YGC86ivB8OHAuO8yzrCFBPTFi+hKBMQ1
f9165o5sKIahBXxv7Eqod+mHlcRGs+/FPzOlR+ItxKA09exOoij510Pa5T3uGYs0
+q4KncXFsZcnWR8NogWoQWukvvjyoFcaMTsQ8kfvZqoDbhABxDl1QEmtdW0XnVUE
YZJbmUY1yv6AW4GLWRk4V+DcNX50z/EkCg42OcH9soztpxA7ns1HRKlRrNbcLTM7
EsAUjwme9ooz9wA4WWEvI7mOZD7Mb5hMmWvvP0l4AGyqwwWn5VnQ2HJ0nTm3xciN
ulwj8baxJ1/ou5W0epsGPbtSRjAdMH6AAtYiL4tlV25eN1+eiMJGYG9fe8CIhapf
7qiNkppZ0yY8WznZZ0Nq7FGavME+04aFcebiH2TiAaHRl66OcbeM1fWtAP6m+6gW
tzqefM/hSL9JAUWUFHapnqLUe6LihGIPERgaGj151aXdDOw/cKi4J2wCx7fLVQPd
l/rV53Payg7IBG29uuO0rzaxfXDctV/MX0Zg6icBjNAO1oYMh9VcQn7u+Q7j8/tg
L/+cK5B9ylqhNUvUanh+tVjN19a9YmAJRMY0IWPcDsv6ubOs/JbojsLaCQnsSntN
fwWkjRKJzmxw25NA0h0jHS+NUxgtdWr2PdFrWHn6xx831GOVrIfn4Ws/lNvksKRj
FdgVjZLuiFZTxQioB2OVrxH+cfpUqA26TGA7n8A3boIN4UW9PKQB1W+GkPOakheq
Afj1fJ8lIqCV+/VR53k3zsMH0tvR84YfeOtgYqpwut0=
`protect END_PROTECTED
