`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vsa+PKuTV0yhw8rlS0LFJKNbQQwJY6iYpsup22Q4s9NJ9mAY84dgkIntfH9o7CGE
naNvDdIRv91W58O1xI6COdqynpbugedV2aPYulzIrGSpGYdYEoNj15O/OFVwpVwn
E9jXO9JMe1fvW5DIxiB3Sf/7yaFJSJWRbpjM/8Fijg0BrE6NiQAdtn+AEH5JEYEN
cM2nZM0eBj3arYIEYTbgnB2SzuEVxPWihHoedvKlnCoCubM0snjYUMUhbPnQDOZ7
ArNMNS+KEvND5+YAt1PZHjVOlNpjcqHif6yGkFLJ216F1P35Lk722XATsr4PQFrH
WrZKiuxBv9LUQyy3DLdNYqEmuqEqRordApmdFsUtjfax7bGR0ciSkjUhtKW7owSV
j4+9NdSM8lZqKFd99I3C2HbnY4i6qW1Ox+Hvoa+uXrcbXVa9pW3pXrNiF95B0k0n
kXX8DRz5i6zgyMQATjgwW1JaWC3Cc5dbTaSkhYA2eW0lnN5cQHytcd9e/cqRrhlF
7tkmyA+SmjC5hmBSOgkNHdRDKNZZifFdUIhjyqh8ZCgt+4IEm1VJ70Us2GEugVAk
874GxtcTBCohWpluMaY6TT+mdgzdDStNZUKypOE5bY+knFL/g17UPf6PEvnnJc03
/kTXX0DLNwLQKOjvQvMCQk22E9fxr87twg2OQq2AGF41QgZN+FSaSc4ksvbHVHSa
OmAIxWoeHWpcueuo9UqaSuSqUMrl/ocPG1prpD6ieRYQ0lv84VI9kjuN/JSz12Bu
dQRstnATzoJuaBQAG5yiyBhaxyiC+OWQfLuM0HHrbmY+uD8mvmHSg89sd+oa7PRW
pAA44d+zX9XkdrcM1gDxKPHQzaL53X0BrABE+sfXahUXI+C/ad4ta50ywnzfgr4Z
mC8a5MUVc1//OjJV4Tjq/5Saj2iGWzHSXN/9fh3IIVTg03b3zwwENmM6cE7FKbZz
hjfeHrFb4I7D0f34YFElFIvXbtliFXbkMX8kuWipX5i1h1lviI1C1fN8FouKmZtZ
QqFJMwJ/fk/68Hr4aimvfOAtVo2GVIQDV+Qcb6udkJ8jmVyfJl+EYBRzzDOamSeI
cOmnKD88YyBJcaP2LfQueMKlCBvUEtaPMigb8a/zzOPru9fAj3+Tl/1zcb+EF5JX
GoZrtvRjdvR3ZBb77GhM7rl3SPZoz5gwvasyNOZvsoerNFDHvqPEfF2ucun3tLq5
bIjxvkRBQyr9ArAF7iGUB5yqDh6XQxofKdYYakrVtJQmnK17wYcqmqFWEuI/Vml+
tYWY7MxvwdjXaSKJXxXe7vPmXT4jPR2eJLRgIUsnFJzHPEsZEzwjxB3OIvttGOfc
OT0kZGck0am0rDWT9o4TgWJEJktdxYhvdrjBsz9mIO+sXGOn10X0ZIj/P86kbW/+
`protect END_PROTECTED
