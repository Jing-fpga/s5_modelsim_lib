`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7HC5SCfiaGtRh2b5+iAh9viIRUvlV2tw9XGglFGITS9a5HP3ieq9qk5+KhyO0miP
/LYJiFt7Nj9Q3am4rJEDAF0u84Y2T/ugIOr1lCpGzyrvB8bB45pzOb8qeblYedFk
vlpoIf86EoBN64Ty2FUhCjW6joDQIXnESPNU2CKeyRBzp/+FRK9ewByOtIsEUPVL
iSUYAUcSvwY8dw6CbC9Lz/k88lzO0Ewu0W1RRu0N57EtvYrWRdrq84/fSkUd3cWw
rXrvLy0/O6ACx+CPJg4uF7dWXWw6VvZJ7eqi6SbTpfexQ+oemmXpuKjSEjJ14bKi
1QDwkz8NKbDEkWMB5QKCEKY3y3k2qPdY4Qr32Z/zP00M9Wb6t1L1BvMCc254U5vW
ns0IYjP3GcsJn+6Nhdm34DxUr/4VJpCxxGSkrJNa/9lEljtqvrngvFqsDLj3GTbO
f8DiwCyrTYI4nGbWYGdUL3H1MKplDPm9G4IxIzuhNE9qB0bfCIZhak5TbBkFiU8J
l5yBZIqBoq549wF6FlfpTCxbg3/62/Se5MxDaD54yotrZ3dxdtCKrE/QGUvFPoP9
yRC9SWOMCradyi2Sf3MiqPZpDh08uZ4y25xkTja/Ca8BRnFKZYn11alTbM/g+MT0
HAn/wL4y7R9SwWUp8Xowiw==
`protect END_PROTECTED
