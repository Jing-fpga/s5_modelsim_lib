`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TNvBhUnSD21QMHLMWUTH4dZIEINt7XGZvEiAcD9VqtwJXfpBEln+61sAmRihBJGQ
whl5/BbutOISSyKiNC/+nKgpy9JImZ8s6GmWug5Vy66qWs/kgLdSf30wgBSc6FS5
Iu6ismw0BJmX48XuDPw+7ZwsHjkDqevx+nsibzF0wozN847NyWukHOLpVzXOQ1Kk
fYFaqVdrmm2EU0gzS4UlER78EMLNkVuCKG7IJIxlgCMWS7ajm3ikoOx20pvQ/Cr7
rDsoRTwYIt/Trzx5vn7R/RjaTLdKqum+7UEB51lNx3SSXIIZocs+JdJhJCjMaA8l
bkm4Ji/WeF288Kf+PfXySRjqv9UDmZgwax6HCMBHHGp4xR3Nrdv9GaCfVHjiKjkQ
E14MzKi9O9iYphSbOu8GJYBeTsva0scKvfxLt+f99cE6cKjdqkkicubQY3dg1PL9
5Tm6LAqkCq3qKhIM2xnTaXAGmzZMQOCOCxPbMPggcEdHR09YL8Am9ACDtv3r3DiA
h1tKCin1vOLtwfIDP+pGh6ZA3Jxp6MAiNRqVl66GK6cq5UV78dZeQOtpBkqAf7qr
1z5SAOp9AC/CPermGqfyKG+apje9yzExMAnNo3DA4rnU/fL4OdwAk86E/wDcITx/
ma3664qAylqQ/y0X6Cmp54Yxj5pwta9Ky0ufRGUx/u+rzYA1baOK0yxOUaMbVPvP
LbXOXWQQ28zkobR+FrhIsHEb9eYqLYWHsa5UmmKIVt/Y2n23/h3CszyhM1ZV/uF2
520bJyWzYSy9ipOXRB9yNz1rfbTAv8oafkYDaEsF/q7Bkm2hepLYV4QW7UgRnaXr
FX4b+d7iiKO+rbm5EkDRo3F2LlkIpEWAgjodsJwPQ/mtg8BM+91EKSRTezOxAxF+
/Bg+jIfNf3p4gGQUb4Tv7mBelgNhtRqRZfob7OF0f8DcaaxrTbeF/rnswARd2qBp
Fjb8vUhRl6/XdGzOvjQMeA==
`protect END_PROTECTED
