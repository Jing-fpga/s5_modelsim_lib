`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LZXMpdTU80dcDXkTbWVTe1jRkM0/pib0fGxG22is+vvREuZdp3usIDF9hPC8yFrJ
YI+x+zKE9w/dBxNdurvPF0CJbSpr7XCF5C0v6v+qQkj8/r83zj4VAwBWbCR9vxQE
hx+iTQlnO04OsO+U2hoAT5KOFoNafvwGnJO8FNaO+kgQNMR0MxmEOM3pwQTrGad5
dCfAYVg8LSruIOlVvWFVr0MUtzPEHuG3U91eWhdtiFRzb0VD7/bX9IuHVMNQrgaL
hrqf9+zg34Hxi9EVzx0EKH28PS82R/YRcu3h2i6AJIM7hFaqlL+JhkamgeW+RmN5
qMPkgGmRf2/Fw96jLPF0ay/O2NdwsdKrDqx/Q05kPE0KLihKT4MxmcRF6ZyifBQ7
bgOplTAmDGJikmMBrEwVeNbeoesVduGLO7LTQJ5/wJo7xuF9VXD69sKtYL/1dj5v
XJBPZ9oVhuXDjv8IkRMYqaKh/FrYA1BgucGIIM+qYc2TPxWQCXDfsrdk+PydHxT+
370TvRgsVMymjY2KzpUCU9LrCnuAIpuVoD85XxJft/ucjxqSBk7goq5/mypHWtUJ
ywfAB8teGt0kBDCWWWGbfl00nQLsNWCFBPu0ipr1dJ/k1Rwuywac0S+XIysd7CyE
kOfmT3SpCs9XSUIAKnONIh2sbw1GILD6NgHzA12q18D+dSn4IXhJo4DKqVFoau4L
Le/LgFdL6pgKizvT0TZEPjKFkB0i9qNKP3Wc0AICAlCpzpGtzrjjtZRU+yl30VfS
DybQ8+7gYvmzbMInkpwpJ9Ghb68V2Oa+fzBRMus6nop437NEPW1dQv4Nr0OPjRA0
fmd3z/R2+tg8kif4Ndd+Suw450a2jgwW5HMWox3hRI2MSIo8XmObXLvPAhQPw4sC
kWfOwZetMML7lzMIwG+F35/w/DY85YPImXRJ8bnb1oqO1tqa/1f/ztE/JoktamAG
nfollCy8FkcdxJjv+gs1xxXsqtn7JS3kJ9EUs8ACNehGf63SRbWyWHV0rcMXUzJZ
zuQ3knKrRX56HZ0XWTHkix0uWTD4FVyvtZ7yCdlF9Lo9LrdAujJ9nSMFi6W9U++l
8e8LID/PfzWVw1wklF4ZAv8a8D6fqoaQ3BlauZqCg5OsL2n/XAv4ec6dywKl3CKj
11rpf046xNiAyefp8YNWzp7fuXkn5SBFVWwv5QiCk61HhMcbRvMUV4QvqaP2NnnC
5oGpce/IJKWja8jhsW0MVDlKZcYApbOrslPCUWm8cEDhObR7v18BpmGg5JqjkSPx
7PXC9fWo72dL2PY9eSRNpRFEiJY3YedkqAYugUf6BViNtQNpkjjWxB4My5fs29xf
QlOsQMvUjp9xqGBLZX3jAQtiZ0I/kMeBK4aQLiQJnYn883Hp50yK1ym4RhdYm7U/
14GnsF9HyauutnzFq4imzLeqWqotFd6FG1xqORJrUWv5/1CH3bei2lfhxBTh9PV6
lma123nWHSGHAHzwTQEBIQ==
`protect END_PROTECTED
