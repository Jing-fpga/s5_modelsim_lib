`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
npcVgUAkwCGD1HZi8+n3fAnBH+qRmXieZaR478NKjUWTKtQYnZdOz9JsK5fo4ZjD
E7cLF8tdn0e1ENV9oAo/M2aLSl7q3HFYVVnZRZwHY8ujmnNMvDJccGfR0IPJlId0
LaWRXPfKTK4y/YIXHErqlSyf/5DcaYq7xbJhbkxH50IIGdBodob3ZvEacpvERGoW
SU43NTFtSxvJSPxTFDwzGE3YT5QhoE+7VDNNnfdSksvNkChL+QZxZc0lKRAFRvjB
/lMSae81zF7Umq1VhveqXrdXK5E9kvQCUJGjl3B66Yr3R4iTJEW9ZChlBZaQ5hrw
I2JrAxBfRsb1Blkw+dPIkMZLgh/BWe4lur5QJ9lTEVfBxTYKKmXFK78JXffxDBZQ
Tn6CztUnVS9nuex3XPK31EPwKdR+5qrOS2CWkOUYpvrUc/HBJmdS47pp/gfUaSPT
VTzB+vCasDHLInwPidAIFkqM92r9qus7mSbSwj9twiwNW+B0DgXJlrNPNsFu8Yvz
jQyEJhwBeIuGfIPmI0PqKVH8mejAfTKG0jvUz4IbmihN16Elxi5ZDsIngSkXc0Pa
SgFH7ZGj42URCM7pO/aFg22ZKli4bHle8HP+lg7I5VYPG0xqk16bciQpvQOEIB5b
JT6RcI4fi7LWzS8aEBUJx2f/ZR7LbznPluZpKxNxoPPwojZlE7w4+EuSuutZEDz7
eWAIAC56j5qh4nGE7fmstZuhpy0SBjc1P08579s1mA1hUdkMt3V3OGH0j7w/XO9o
sDS+EhBmAEHmku0/guvxAR23st5ylXyC52eu1GNr5FjcHlAVj2CP0+ajsjuuLApb
GGjUmGxoQseohJrBZKO17cSuhHazY0j6MTE6K/hmw57CHmLWdvNp8WbuPVyj2mSv
dl6NfePp2D8Q2FQ7a5aJFEeFD32+7g79WyUEtIKehcxw7Bn2OC4ZLBSXwi43wYLH
kjnwHcpJiaeVDnIwLzEmNDkK5/jSHPtwVNmBQoT+OEzW29HhYPbwgyVV/yfLqOxN
myvPCcjYkhDiwQzX/DRewBX1ZyMtJ+wy9AQ63DeXb5SqosLjFvYZAbyqbJ3Ikv3X
zLk+3Cth1vM7VUcj4mjVbOk9T/x6a9P9trH3s4BE1H12m69XJ9g4zp6EnJ3ERWq5
lPSc+78h1P3+QCp6cKWiRbHipVZWScSaodQ1XhGnWLQUFEtudPggYi7+hwlVdOIp
i0zr9bfolUQ3x+WUzaeKC1/c8I/PmPuHLR4doyJa6rnGDa0y4s0Cgl6brR0i3EM9
HBO5+rHouUtKVxLRCxEuvPUyts3qUegxI0CPJ7sQXubJsW0rgvu54h1nUIn6ENFg
8iXt2p9YpHXL81vnue/0fiq2IE4UYSioNmr0O5frNaQS7rTJu+KJGR94dyChin9Z
YpbiclAUdnkY++lP/FjnZOL1JOA7hMRgH7js+EqpJFEBdQdapErvLaFN37Ekk/A9
IWAvk8OdZmXHVDOGX8bjK28RJxXu4Ysh1jbcKHp+auexxlAFqjeKS1lzynLiaeaz
PGhLZecz/ni7Yko6AmzDA4OuMnsgXSRMpdQTSx0M9seugFwAsgpUGfblika6OLgZ
UQkilHvHTfQl1oY29QYx1e3Im2Z4o4E9aLBiSF4AnWTrOBt1AFTtDUHIla2DGGHF
/2It3tHxMY8FIkwk9ld2enEeaxDOgkP7N8NI0jBQS+aCAR1dP8SZbznku+65ihQd
vKgK0Cl4o3Ylmchcq70s/+87Gg6HDpU52J+vZKR6VvRgOTla9nq7zT7L4wpBOT69
Tr090QHNPM4c2ANdqdaUWO9ha19g39BoLYc75cVInGBMoP1LHleBTQWp6BLvAT1r
2n69IzoBxFxjEwQODYhTHqg3J4axKqCa2X2CHYJeBlkcDU4wa1OQn1yUrZdr8335
Fm24naYz3Qpj6L1vPZyc+J8IkwzQWIwxKHe+q9kgfuzCv/BCgbPf2f2zCm0hEJ4g
1HTxLC0WZkrQ5+lp/DlzOnmqqJ+lTrCAv5W8aTZFtd/8bPbg/dopmQ9d6qVUl9HX
WPQ0wNVIJPX0eERMthJq0smo8pYjJlMzvEK+6WQs6TNMwsXJjss09TkZPIoBADPr
O6i65SCbs9scb6xloXx80pkTp+d7SGALKaLAbCWQTQey4oEioOc1OuF/vZgqtNUZ
CSZfOWOF6MVMTaLN0k5w4HV4su0svlVhJjQfiHnlcp+4S3aYSwCakJGzkwPtfGaK
BvIGzkdYah+g3MYzuPBokMtFXiDvqI4xbB9UtEJlIY1KE8YQF7IRwU+qzZASo02Z
HygIF9fEHs89QKEMBgLwtX2W71Tm2F+Cbh/5AjqhZfd45A6mZ+Xoqt18vUc6gL3N
mtTRX0Py3U0G/GOyOXoXtLmZv2a//jto1nZP8pfWfgZpbxVAPoRHSK4xIZ/is0fi
V7IdrcoL0o4MlO96Np1gD59UKzqMcKg3D3IOVcZgmUq/SNwFpd5luMEqVssb+Krf
ExEUyjsE8LWqR8x0L0LDJjYrynNJ6+94pdo6MlvDrpJ7yzQM6HuoCP9pByCGhTx5
0wixONJwQ0BVZe3yU6AOxej85QZjWqDKjDyOtZn3tyq2+zI6rB3U8cfn+hdGmMkt
LRxEXVPzTsDTsPt/HFIKID+gWkuVGhPBdoZXFsnu9LKhJ4MvXirBt/fAPnR0Ehri
DzbvIEmDRMwtqlC/7h2XFi6QUw9/GYY99XKMhXK7ZHwTRGoOgpmMShe3VvaHdwAF
ARNt4A24QTf7pIirRglZtqcsGVOt88OJ2fjxitwCNjwG3tsK3y7u97pTC126kdIy
wvcEDEnlDc/KKuIL9hCylwUSOiP+W1EDLgufRJcEGG8RHCWAak5iiGrA6stnhI1P
492zpB0oAmJMSuKZSsFlLf9YeSadVjEitK6yOT1Op36xImluVDOAjSP7iO3WjSJE
PwhgJBvKj+D1HppVXvlHfgvQA2Pg8DMGW5dpHClbfOkU4EgHGS16U8Uz7v+marrf
XeLzn2UlQ/VUGfmmMw9V0ha8LabyHuJZJFBvcTuekC4Ds+f6A491SdCb/49o9m29
mLfRT3RxGV898O2sgcTyBdpJCAl3MN68wGfxjk34/FzLby7Aa74s4D/D2D1+zZMP
/wEuNvIt9jEcLUi38nt++brZ8cefuy6aEfA9EHsNK3bqHm4S+RXObJPnKO/sgccf
ltfW985SWZLyowSilUMPTK/zP4L0GyUt6e0kJQ7quJ9p5nB28at5gWCTVufU0yrK
9w+d0t/rKM8igj7PpLUxxpcgp+VPN6F3rX4IqVoe3te9Bl2yjHjHFg9g7tOwzNJ1
vGoMSVCe+yWAcc4O5F4xvHjNkJzMVCFwPuJwbQRBSuwIqFbWWXZ/KfKogLZF9gAQ
0X1cFtYOaR/nfYNcO1NaxKSUifZqrGIpfObBccIfB2uEJlzW9J4Ztk/1UY9+ldNf
7wNeZJSP9vWhGVk/ZhyemwyNxaN+WKJdYrTyNxsVAA/EdJPq9agl24VVoBA03F1W
XEx1pbLzO3VPfU09TYEcYx0dMboHS6AB/DHCfjQJQZNUoaWeog3afqyZM+z5ZT+9
vxNQW4evdxTvd1dq2lB6T2Klmox0i4dSAy/v88wUDdzO3SDH/mo1I5xMs0r12ROk
1UW3RF4vd5h57oudCXb2oJ2R+qf/uR7LUQVklSQVGHW0OsVZweVMBcqRYNpU7T5k
VtAuURky5zwtYgTAg9qA7dsGUGZbyWFcwBXuDoSr/E/r1KsqP9SzbdDkQ7pmzX45
b4H/A1Y3ykAfPrdh7q+8LT1Fro6G6eKNEQmB1T+e6EPC+xwYNHvdzM+2weERczhg
ONufUOG8U0qJLhe0PQLegZQZKfNJg1dYcrA84Nka586WW57EwtRmFuycn5/juqxV
r5oDT0xpjR54ssUu6wq95BQ9WP4ukTuMOct3G+GNGa/AqZzbwKxUSA3ujwWN9htk
/3Ah4911tFWFn+8hBIeeZOxAm1WKlqdgjwRZXYq596lnQIiT4kLN9uzc+ecNW+Hw
9U0RwBVOh28pNT5z5q4Zn4SGBJG62hHnDE+1lXmFXEEqwm8yZcD7DxUSbWxLAO0h
/eJD8SoipG4h/fwxhr1XNkRv+RhtCF2LG90EZIe4GWmx11gzKrPshAK4nxP2ofm7
lLlqnMcWD3hac7RJYnNsbAo87Jw/tv/GN/eo5gMU2/ro7ij2GaqGp1l6OqsgwGbm
BRUsBbMJFiUPzkkUR0T+L/HvktT3+9rW0DIbPODJcPK03A1rvqbh2cVBkYhJxgmN
BUmR66XP0mpwa5NN0GAg7hH8buzIacUv6uticEi4+6RUnftqU3/PW+avDDG2laWH
415se90xaZi2MShf3X+fif8dNZZ050knE7ij7IbQa6RkOLJN80IsLbupOHDSKp9Y
k7Aaw9w05cCpoweQ5HstaXeAJZI4c5GwwisuzO1un35hoTbTSEwwitJ/8ls6zbQ/
ctg4Irif5B0dPvaXh8ARFBJggngmex4ncCFt8bQ6Cogv5gO1aEmuP3c4QePr6Nra
2fcyYOQYnyO4OznG6MCt09tFPshrixdzC5tWiQNxG6lYVFiaAJ73sQkC3vgTkdTH
zwJe/h/e0eQAE9MgD88WLr0TxhzRzmwrhJSKUUX1wVbXkhsuIiG3WB3XS0LNN9iu
MGD7OeWhg4Ck0o1fK364T1qMDCpLZxgh2iOgu29JBe+aLLY1DdvLIWQZAkTnNgM7
O2Qn8kK54Ru45/6XYSsq1Z788g6ErPHwBUVpq3+07TDzNJHB3z7h0QMa2pzc7jRH
yJHonRGUrGuNjWFggWNv5E/OLYRYWZVdTTxnnURJNaPbXpev2dmASgFLHzoniSaw
qXRsHcHHtnqK/xOytcbU1ViKtqtOSz+plAe21UAZ5S2M85XTQmQ+UzBiCqdIW+it
ou5OeRNOrY2y4Qn6ntZ1Tjh2TqpMi0yEaOCBX8JVPGO528BW8+/OLIx0rkO/yphZ
Y0BqJfhtyV/mffPQt6iB3uQpjc79f0vC2G1b4worHIJupbN66ASd8EDYFAxJjdp9
iwuMhEi1tpvQdxraBHbSXjSkgZa/f7iFxu8giH60gQzJFNTg+RI/VaLeq2tCwuMZ
gZA22wsp+PYHysAtf3CFaqZo8sk2y0EUxErQPD5l9qGFILm+VAnCyxbiB8UxSSBh
ZAVOc/6Td7U/IiJJxZYph+p15rebo1MEkkubZsksIBHLLdKk1awgNB2u+RS8p9JY
0aoIsWHVbd2gApxhbr4QAnjWQlY569Rmq3GpEl57mthggT2d2KCsH5IB7RKdePWz
1y5oRFoMJ64R/LT5v4/4XVBzd6l3LQAEDdIC1eH3W0L0cPmmDyJ9gcD7n4wBFevJ
VMvpM53Tfgw2xWpZqN1r17qCfqnGDCAI9naBPmwdY2K7IjZESeicUxJtTUQ9fmkM
q0bbi/aus9q+DU8vOElre/Hvrl+SAJNAOAcze2RPj4rLSm8B01aQDsIGZHpcR3ud
XKAfRHJcSPmij9/9IKS/cAcBHUmV8E1lbZ7D2L9RfqQ7FF72k3nz2rsywUlmXXMS
OEA5vXabfqoJW1RVUEivdCNpcuBT/lZ04aHxU/u+RZ5ObjGOZhKkG4nFu4SOZIsu
1XvX9mCDIJ7IMkAsDS9UeEnr0UIUFfNbCQyQ9RcHyiLaam+3u4rP9CR1xyeXA249
jWt4kzuKMyJDCsU/CcNYZPrmqlfWMp/QHBV0NkH2S9N0ty/zgnEh7zcX8OQwxWR8
BXMVVak5hseAUdzVOeKTAMtfeqVyUUhi+tWKf8EJFsu31vqNILqc+/rFqKXTgYiQ
RpAYLpXkFCzv+Haz+H6fCO94QBi7uNln1joodT0uDasG5uat5B3tlnb1AUujaAS6
khnl3H6FA9sznoWRT6/ObPtNVe73HX+kQSkemQ31+hlbrLvJKicz+4dGDUbfLvq+
Lql0iO5bB2rCmnwiXiwV77k2tJrQDM2V+qQjdJNANRFgEAY1TPqkVufvBZaKM63z
KUzH5jn3+oyJf6RCARFHVy8ujJezfsjijQXSfuN1WkLbxuvroLlzPzwKAgtEoNuf
F+ulhPPlEpkUgmCOLVFlUiQSKvHofRzd/OFtnOsTtBm4EFrxsAENTjy0QcfIHmoB
MKd1+8E8bMijda0rjnEG3+05YtnRZs0jP+j6xdxa6jCyonhf9neDl6M7tR8EQp3c
IqXZ8iiYrS+0Fyy9MVvD2eRcyPuwwLnOAONK7WeBmfGmyZ/8pybYUWNsq+TZim3f
IYYyF/fHzzf+Fz6Hn6hGl/yV/YneuAxoCmQgB7o0iAYwU/F7NmVe9N5EOIlMboYi
5VleKRryPD5Ktdy33aPP3fNQl/eDATP7VIr2sOMzHQcCBtJ8+erO+//tlOHse/9e
6vYX6RiOtsKhAG42howxQQ+vyKRU+4s4/flaFXexRwxKN/ZTOS2YVwt9Wo0R0E9D
nEy7ZfWlT3QEnOopBQvqL2YPkB8jIhArFimooTbETgR3SFmdf8BzcV2H+eF6NXxN
Iq1T5WDbumumFCYZrzq2SjCmjYbITuSf4AIHbojCg56beN/dzqbU8RlW3cQFx5Cv
wadKfaAt6YxJ2l8zWA/MePoSA/CZushHpYPBaBri43pIszSxWKjsV5OZ+esIHgqI
elXo/6q0NqrQhfY74dVZS66LPsJlqTwsV3R0apjoF+WfwR9V4mfAn329Gwpw/Izh
LddRgRTuZOFTBfqseSpKPfuuXTHTwDLrmzenHIGiudPdHtfkO5mIw8AneykYB1TG
XXUFXlqix/XBXoCp4n/z/hbymmjBc0VukUKl4f63RJlyq1+Ole0hwms0bjEPYkdr
92/aLfJd4+E2clXrL/cSmD1fxaLn6HHCUfzHEw+8v7CSeWUYcG8q8nEh2y0Nz29C
JFgGjQHUamcuw/SxK4UzVDy8TJFjvtbEGpjqnQ+46kh5NElw3aYE++d+JUSmYcgG
W+Us0Q8UyA3IqLsZkBPQDjK5UIRm4KxAoqXMHcH93Rv4NgsSXAkmjn6KFIDQP3dz
gXIsBWu8E/FP6gX9AEU8iUIRfquxbtJ2N1APka2XuQLAusXzxbEMAZmcl3pFBdzm
iT6YSNUKEA3IXMCXCTLDV99avTk6btjJI8nVvAKwZ1VAYF91AN0Unww543zY1uR0
mUQyNR08fqI63uNDR35tn+xbfaVj+c6geVG1gXdpIGjTShq0JQhMV65EYFwcyy93
I95yMPZYnbbGAeazOBYuvi6X2syKiLJ/H4zGPlNN87+AWwOTCoLLejIpfasIhBkN
t4BlUyzd2quW1vQN6/CD2ZO+RFITftDSf077vaUtBgHBCN1cnj/8+HIywPWoOmpU
kJrW4JYT910cnWWGI2ZEEQugSfeiXuqPHOr8ESx9+D1AsGQPLxaF8ptTvANKXSyw
Xyx1nEpkwBKnLAgpRbYrk0/Weocm6OUjcwL7DkmBzMWvO1Ns4mqHnbdaDgwt+b5B
WEi011JoYQBCjWu/j81YxODZIh79ZY8vZ6JkCnPcKmWLB0auXRDgNiHTzEJtHHSg
p8N888+yATD1KJKYCaDGSgzApt6R6VpfiSSD4TU69osxloEFhsnMH5cExEMSRb8x
6PyFDNOeulSoG5SbVG/pRNUTTupO4YeHkFOTb4h82gZZKMV0a2WbuNcEUjjhSice
D09sDlnU0KhAyuXdgAHo/u/V9ricX0zDwgsfS/KTmo976btwq8vbo5FH6u0D1607
B5sbVxQ7BRdmmraF3SLu7IqlnPw2Z78JGj7BZR9lFpp7g9B3fZGpdV4pWLw6cWCf
ZRiOQWrJUcF8wUhsedOfSpAcQO46ZVM0LZczOqfSjxU6oErWVZB5l46g7fl2pMzx
7AJnOOhrTOoAWQZXRwt4shO9t+p4kjLy+5gB32ji/SMdzuv1QfP9L39YA6MXMSIf
hBXBhW/M9w//LwxMaFLW0kT7ydz8pQRCmE1thrDZMpvKh/gofnwiYwE+tZ9Rw95J
xYdyKEkpl9UpY0g/6LYI+idSWTPVvIdG5NC7v8ar8Yjg3E2aLIXqZ6ya6WzLJzql
d4YTnZwbvARyaFPL3nsoTF9StrkrgSPuh0zFBEQ9jkR+dUD3zBXL1WXhyXPiD2MW
s5NHnz8lYCGd3ImEKhE9FhzFarKE+Iy3KCPdJ/JeMojEAgeCo4vopV7ri9QWc2UA
dWbe91H5nJoxYCBweKeriMteKvWr2acrbaVnWxECdrRtn3KBARZ8TgSwrArO5BvD
zqKAsFis8yIOEt0gdx1bwPxu1XU1s6gXX5zWFp1fi8wEfcMN45kUSEaf6TxV5RMt
1GhK/X1Tt146t5av5775sw+ASsLxrP724frxD2zyQilOtTbXyT3F5sW+cEpVcT51
dOeAnlYTeoWfxHIEi9JiQ9EgSV0n0mRl9OOxWusS6msGe8eXfy0IiiYO69PH+elZ
I+XqAboNoT1tcCTjoYFX4y+G6a/BeLJEu/cA9ftEW+xkkm+cu0BvKPHYKNfwKrph
3akSeeoGt8tn4QasS+p3WR/X2ddzKViI2LBwwksMo/a4rfaIBWchs1Z49ic2iVfb
GfR62Ot5SznJABat0HEEYJ3fUXYSi3r51VH2M/3qg0qdhrV1Bj1ZPxYHbPD2egsv
nYq7Gjrh/ubmVA2MmOdFvZdzQ4xhOkdxVPEC+c7pd4KtWIROgfGd/3IqNn2dY6wO
t81keqIa9L5duLkwSujk3aJ2OeScKXuDzD6Sg8X7+INXR3U943FrRCVWXU+PCycw
d9dxF1seAhbmrBgE7ip+Jim9dzuj3wOL7zTBIL1oDQwXLVV+dbp1iUbQ+8Z/M6SN
tKWWJkNzTDq+pLi3La6R5yPzU6fht5DVh8O0zM42f08dnE3QBWOKfwyiyJNHpimN
nKhADlI7gc7bgCA90k0VE9ZqEKQVToKscYS5r/bOlfkRxMW+Gh6mVw4SdbmQnYKp
OTBflVPSAinzr+qmyp8uzIs4Q+cyCX+AQhBRQSL+uU+ptfpUGTN3fyxIpILy5ft2
8Y/QTCloDCeGtswRJMALxHNUAesexKvDqvZC0f7ncIUvBZpoxqBlP7mUa573U54y
xXcQvnwJOScvX4/WsoMIilsv6l3bSOImkrxAuAFKJZ24kARFJAr3lQYkPblnfCDT
8Tl8EIsYO5+pOAob2yp/u3ecrhF9OzpxQn58B6Cv4EAU1EWwjEp+MzOFuEGmopMd
J14Co/fDKofCQ+SEBfrI2WzW6SyOX/vf3qgzMEG9F3aTKmzRzdyfLB8Ukg67tJ5q
ffCVEH7FeaYJpa3+Xc3XUiAR0s+EiyXwlze+CikAfP1fvWUxuRXlfu8jkoRsTUnw
v3rf1Qb3qWtF8zYOMHj0yrkx8kFoqElSsG33w+jLRzs/a/U/9qx8P+GVMh/op/zk
W3VH1/bs+qzoREUiegHsUf+YLMF6lG1THYrvTs3adKaWO/vz3tKvP/XA/CHITVJD
e+BU/v2I56EnmR7TqrSJu0B2QJKkcgK+2dIs6Fzap9AhKrGc3UGYkjABhypeGXRI
wfygr68uLu1SQ9o4oOgFUCKzs+4dAQOKEFHAKwMRThI8yKC/gmIV4oDLT57zuOwm
uV0zxogL2Hb6ehLDD6/lBGiDL3jnljVIbMoTA2y6i7zBx6dwaRW4hjrxQ9RxUfO8
zfsbOothLJHMy9rzTO6md6+s/eaY9tI40bbJ2CNK9W6ywaC2voJfMOEAhdAQs+ob
F0ulqW23QbdgvqWVZimm8coKkqLYqtJzQKLuL4GuCYlOMy+Qi6WpIA1P7i3OhQ9K
hVpmEPxiZGh6/osVZBhINoLBuBQXA5ZUuZxH94O2IiqKA4aBYv8RRKB5QJygQ/q8
n+3J9tfT832V8GhnvX3jIyu9o8uDobxU3hGNQGrV/MMy4xjaK8XX87qJ1klRy/tp
IDAV4q7pfteonS3l5Ntz6Z09OH64IZAUA24tKNfcdrRyrZ1l0PiPQn0IX1k4ZtIN
4LQdkjOrW/pNuzYf1DZaeDbbuXM6oHzabqZ11BAI6lepA0Att2+mS3tU3JMaKOfh
m6hbAlPdlt4eVGU98PrEgYstHXG3cHNy34soLM07yPwTRpZ3/4Q75rdMIS6lCyar
cDUKzDt1aPQTKqeAHb/iWM4ivzerwu4dXDD8mVCl9PiW1bTzpgZmyGqe02XzBbWG
5dLHJIg5vfilmS81PjfrKbtwACDmYHazwV26a9r0xMpLl4OFHO/P5mHDwbWxHIOF
/1BtLi+hRtN94eFryh0KN3GNVb3t8FnPHwDI9XwXD337enNBMapa89kRZAhBl1pJ
fzW0sTPJILVP8Qgq7X0lYmj0ql5Hes2npcMHUqnPAlQZk8ezcksis/uBskbdqFpN
2jVSJqm88ydosgIvTEJ0OX9wMY0LTB3wGoC+7UudR+xxt+3xQ4eebjsKQNyWapkS
s2ABUR2xhTDQiDUjBJdJRL6lLINl8z83Al5C7rTAHEiChte4wBiIfwxq/PlnTlFF
qMS2TRZNcs7Vukfg+W4up+Sk04o8lb0smNJaa+3YKkVV/G5cd5lnxIxu55t8tDd3
29QgF6sGGnpfSK6aT5b6pQbYdrJ1CrfP2nejQ/txyNfwlJ/6tkHRFzW7fD0rJ10T
+87TBhoU4/gWPhCmdhmBHYNtQgIZd9fJKxGAHoOFoQm7C9jRJV5kIlKJX0WlfRLY
XmkotGCl5y+GpQePYCaKyf+7GKGl7kLs0f4jzYL7ws1YZC2OKZokOCe2JEzPvunl
Ozwd1q8osIVODKxobzLBWh23x6l/MCZEmEIE9UlmGd/1yUhafU5t9Dt24AcreIQa
8dAErIiPhywZqD2d5+7LRptj2Z/NkmTbMDlQWjCfdmyiaqo2+OO9tc7amSxGxMhH
SMPrp0xOip/w6hnjElsND1qI2y6xNu0V4TUKtvpHVHVId+nIMTnBBwpcQJeYIYOe
XIV4awqtrxGFvoqD8f2MVxXpgja5Z6gNWMXXldthng9rPDpz5mqTpsJI6W8tGBFp
n076u7X9tR5J0nW1jmLP8lukZdU/QGuzKgxhGKiqc0mA6VjAD1Y+hWQVQ/CRSoTt
NLXaLS0IonTHzVnyW0hSkX+84vJFD5o4nsV1LLfmshV/VAX9LnY9g6CkXy6ehMLQ
z10R2nOI/eivrOwuCDiCwyF/vU8s4QjgeEAApT5J6K6HXhIRUUF8xCf0nLaLB3Jz
naLzh2R+SFLF4sIQVq4hH1WxIFbKyk8VTtws4qzx8Cgk0wFYGBfWZtNjK9MhSUqn
7GCeZoyqLvOk8LA1Bv7aisOzzTmsrUcZ+b2hsuNOksAybewIRWqMbbFr0Il5zVqe
AqyADMmbdwtkH5PxKrhlmf738rCdj9RpxLcIfN98EdpVp6W0ejCKoxnC1iadjJKA
afs4l4N1GfJ+38iQOyRYBBGEVPqSgox7Q/jPoZwwDLnvclB+NmmIeKKf2GIqz+2k
rDj/ItViW8s23gt+KGnJ8WUIH0cCt3JKHr2Mggw2Xpo1yPbLqa61apVoxJnOaJJ9
DJelc1Hxf2nMJf11CIQF54oj0+QN0Rb+yNcFeFky+ylbBqISWKWOCgBdr9DCYBZ4
hWwmYrLgpJdnl6rQa4h95PKMKNM4VPBj3vARysi7DnLOkBbtWQdvMAgwUZRgnsZV
cnIC1Kn7t4eOmOb2weFHVTVwcnRHZHJIp9oUqPXRSqo3cdWDcwnuOJSd0/OpvXP3
vzE9RU3njBm0dM6UwjOGIHg9qYgBLrvOnc5iAXsGKG+tnmGfvoyp0Zz45GM+kbAw
1jjQqlqjJ4v4ry6+1uBsSMH7wTedAbqt+KfTP80jHC2ckavRhjzddg4MbySdDw74
AVMScKY0ochL2eTx+5SXLWz4FgOffTumzrD/71JtXYDZrTBG4qBwMT4uEnd4kH0/
UqusRp5vUUL/i2LH6OHblhWJdm41RgHmKsjwbwCu9OtjFCaAW1L+4q7z2p8X15Nq
ahnXbyK7uqB0ErXYFlwQrzlt4lY2lwJfIuW/3l7t+j+hpPtugvcwI8rJK9Bt3vKh
TFs/i1AWqaulv8qnydzSkqVCW5ysJGcpqVsEU0i6BStspL3BIHPvU2R/Y0QKNL1H
fx41r9rx/c2iu0LwozyCZqYWKOed5rAiMF329EBKIEtu/Niusd13F/a5KM9AnfGv
NI8U7wcf1QdCF6hLusQV9iSAhewtnXZ9/lXuuGgNFAfdmYtBThci8vITnpmHONlq
1LgnS/IBPDjfS8U9npYT/eKbUBL+RS/5nSg8Mr1haI9Q9M8gJR1TfHuWxoE0SI7K
6XPj04yyJTbcUmzA8xymMkKWGpryEqCl9toIFgfI10h3yezxoOL+nYIzqrCQ0wKs
Tg+eLE/ptabyCZ4nq+ku0Kn9k/mQvWOiEPGAvH3hGxbekhZny/E0G37EI7wPLLIW
1RR5rEL0aJBoQFg4E7op/BPOUUdAVNndCode8N33rXyapgciJyx9vhzpPz844oG7
6d9woUPYNWK0i0QcyE68DuG87oFR2ct5+m7AxipnwvnY3qHn5ge6jNwrlzxz54gf
bqxbxLM3fZFlOPMl1gGGecoJJFGxiasJLWSk1uno/sKZJeeh4wv6RWd9ENgh0I+/
MPsRoShG7QYIGKRKWFdABZs32+753lTFMWSY3oBooZAh9n8cJ3/TKEaOQEaAJdE4
X7vFzid2gQ7wzXEGs2G3v6LunPyPeLHmDPL3ljRl2f0iROooimeGzpGY8rAtVbH4
7m86KcBrN0jyrMYrPSVPfCnHP6kkf5sDL8sT9YpPfXDJ2uws09Ie5fsHlBqfW2lh
Cbn6jOMTG7AxgsIQUMCTHzUTZNnwdlbYgK+lAeVKjFbL6XAcg1iX1OLY4MMbr5qx
fSmS0vsy0GFGw+XC/jOt0JO6f9oY4Ruvn5BBxqlZ/qtyo7hyX8GJEJULQ1zaVBFv
QmDb/GC67JspRK5eLM79JEsEZtu0f79K9407W8rQWbonNrDg9y45iBbilaxgFVOc
I1GYCheTGpBW+D7pRwzMqf7XhjML/5dlxlrSk/tlB2DFMPxCrvBWjJ0FJ7hHT2qj
sHaCk2j0wXO2ggO1c80/19Ofy7vYbRF25cPJxTlrHdEIg914z/i/TSiDlDpkqg24
/P6dZj+3aQjmwVlLQPbHP5IOf8NEAlDAVwEBVMZRTRyJfg2KLc30geL1uyPo9b/g
V6RVOT7JWuTC4A2QS8B3o37adzqByGsGQzTkeSA203XpQrw225zhZbL5SSayLOfi
GDvrACq4voliyScFRx6gD5G/B7fYazuQkdskfauKMTOQ9QX7hOxkroK8Xm75VzDB
VKsPV+4Gb3wa8mMJ7U18JVd8LNPT2hlVYxxfbDqIcbMRsHdaVZ2Ni52vLVy3Yxp9
AcxUgGbHqpt2U60teLaf0oqqwQxXkednVrzAYdXaodI+AUunCK3jiPG1GIYy/XwA
c+til3rFM2bOg26swwKH2ebWcUWQM71zxuLPmlOyDiKicUXk36nHhrd53pvUOVTT
+93WfH4IyD5wPi8PA+uPR7QY5HUwKT/3aGDPCllJ/l+twvQv2vhkmUvx6gdvtRck
AcnNyMA6Qu87aLzPEo/jIjfDu+42ZopkyIr8jtu0R60UXxtjMJO4rNOMC75W6MYp
yeFaQYQq6kTo21yRYvAY3A==
`protect END_PROTECTED
