`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3VlJa6otw4guKQ4BCFWw3uZbZKpoOs5ixFHi1j9hrMa8amHiwZY3RX93XkGI4gtn
OkzcgAt1uRyS2Xz9RFUFISEBqHKm/KdRSekbwKFzqWs3yBAyAizSg6NVCWSeL/OT
S+FR50HhURBFRU/FX82s9qm1tmT+OUEhY1ZdPEh1gSWdwZUD21b51BgsYQckVT6G
7HxCPKUOSbWKOYyd6cFLpS2wp2X1IpzX/Zj8RqIDfWvyPrAD1u91N8wA+Red8wih
00LJ+Kyjp4nkNsmCX6yMI2x0tX8gMw/3Y8UMoaco1RffW9yn072YP4iN6gpbb0JZ
M7UzAuSqotjpwhH/eTJhJbGpMVL0AV4HUtgjrmBVq/aEosMweNXmxZtjcCKFWZ+w
GUnSS/7h88twCslz48FKWIDwez0Exn/ty4MhjP1RxhX8DPCWzZO560ijLoU/Kusv
Tmqr/Tv5XYGh3kVo/KujQXHqMoqKbOuEzE8cjzLPvPiYx/QhmdyUXMRGo4/7CzmR
IctEX7CMZ0PpMznqWo/2qBpt0AA0rQHPRFxxhxlY+LlJpwpJ1DFUjT3EZifw9tZ0
6R7y88Kn2KCN14ZcGhfRImL1LdLrIy3MbHxoKfMDKVyiBjkBuAHtFo8O4P/aMeW0
l7324yymSh8YVzXF7PU3x4U72KOulis2dRe+aR6qLYQxlJpf9jLsEfZ2KptKp9e8
g+xJHwVZZb8tgmWz6kSgcnpzdIiwv40RcjZC1+bfP57aYcK2LaNExMw4MPGlupnn
XRH7YbSc9LYyPiJkP00X/XcsxofBFrl1eNcfW+VMdw7PZyxmB13QsKU7ElaE23V9
7PJuxeiv6NASfwYu8WwdYNnL1is2vb+zzj93TIzjNL676KhkFkQd0nBIG1gv9aOw
nSgNtfWskV7ek9oYQp7Ju5mObVYn0U1ox7+TOBtwTb3C1hV4ZEyiuH0VbbKtZtL1
BMEFuvTdB37ImxZjyblCQhcGfSjclRBMzAHSBoWkBYZoWi6/TBUHpmaG4Pz3u8N+
OpMa+rg/Ea+OIf42hFFu/MacHhjUFoxo7j2mksflLeea2EuRNmOkk2tAq8/+gsjA
zY0419UQkBkF/poKLiZpUEoRx/EfU1x5JYKE1WD/Z9ucJYj6AaBaICoSZvunAeaa
QvilcuJKA+CFLHLwI4yjLZW1dJVtDTanfr3IpGZH0Lu6jtSqDe7cjgU/LaDAPZWu
NQmawNelDsgzuk2Bl5aPQIxBkXjlcBGCR37Oa38uA4lDVd6+s42iukcTE2F9o5Xy
YRjS3VBm3jD9wgz4P5pWHGYIMr/0vM3LmLuhLcgp+quOeUkSZTv3Am4goqZztE1G
DczRhQ9soQBBDNobqf5zMfDA0bMO5t/FR1zZP53L9D3MzWP2b9FnvmnaNJRFIbzg
5zNPI6MhRCX12dC5g6wHqxv3O+AYV1EurXCLV20EAmSKOg/iIbdX6wMb1zok99T7
ngb2rdARRLdyhxDFcjlDnNy8XAoWaCgjKcJXNhqLEjH0fYab+d/vxl9ViTukyX1p
1IJ+MwyQiZpahkknBjtitoY7iCxvqrH+o3FN3IMaOFrq1yhj44oe3rKrWff1k6DO
E7dtO3VsFGLDelzhyhwDyPKPqZdWl2gyYVXqMptGuGMmy0x5y4HfzxHhSK5CgjqH
4HWV+8LEQrOHaaVsp7p2qodgUZTEaHcuF4OrbSOuuaf3asUjKIe2bjpYhH+n87UC
yOELJMoZpJrXyx/TkhS3b9pQSx48yhOrUrh19No9y7wtjyBFTUwHsscbSkBQiNHX
tEHXUBZbp3SWm7X0r4EkdMIYQ4tfLKsppG93zKSMHdnVXdAxjRzklKOA+zX9v32T
ZQ34W4GjJuBqAzdQj5Z3IJV8z9esUemx9kOYlgpPelJjeA0Fo3VID6CTRFueb81B
TzTjPil+tB7ESym03GdcAA==
`protect END_PROTECTED
