`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bua9b1l19n7JTSHHqYRGuPGyH3XubKqIntUfx3pzsLmC9qBa6zBriIxtLgpBfEPJ
xvUfxqMZaXejdYi3bH7zYGDVUDAhThqHua1xR21rtptBSq1+tzlIs/wVspQadOgb
Z8orz9Md6v9XKkmEGa/5NKL6oRyrIB1miKkJC8FkpKI53ioJC6gu3KEouY8+dKlj
Y6XUweabirM25qCO1TTvh5QOx4iWeswLha/7UhIuns5306ZVMLLbeFdQYtQuOTRC
rQhn03qysW96SOkbJszH1C4g8VLEHqTw4QCOHVVWsWT2gebOHWud+DUk2SFDMaE0
7FFt5DBLBV6lxxe8M7iT8l31K3RId6MBUAuy4rjic/ROoB/j8G6mguUezVsvRwqw
uzZiOTzvODSmYtrulkK5AL2JBff3gSUwh3i99O69U90cvHPtWEEeWypkLRXPVFVK
Z5ye8y/30OHI6u/MoClhi5yCde79ak7hd9UkxydtdbgonowwvlUhz54q3l8EeRHt
zauLzLLOfsx1R1TVDGnTrADYC1nDa0AM60LW1+a5hjZkVzta8j1Xo3fuPbarPKLJ
VWIjBpHbE/ABFTz6l4E29grLMTe8CtdvjVO5nC9J8mjUqJBmH7KpWN/363B0JYE+
3MOeDjBMeAAhacpwuKn3lcJsPZnnYJnrkp58rfN41G0cnwHYu9PfEebc6UiUCdby
RCACer04eumQaOOSgKBoN0lxpE+BvGjuDlTQWHTocIV8wq2dqQlJr3VtOML7GH65
aPO1vcUhq27DvG8xd/iqus3MgOXaSZKoiYu/m3+mzHYETr1qF2eN+lqkWO1905Iu
lti+vUJygN3Oy3sl9gJtz8BIEzcKHCDHf2+uUy66AtDiVBFCulNgRuZgbCGI/pFC
IIGFroZW/KqYj3y5iyqUK/NWgESL6kvRuKOtXC3eB2WJ3g1h0wrYXadW9LdYT+zy
6g9RuxwcRRzwFN7ivkMOMD5Y31eZQFZouZbol9GcyImN3v65zSngT3/AbKxmVBiE
bdFsM8AbqKc9njYBAFin6SsP3J9otq2TwpjFTpVMcjYSxt2imY1UOaOpzWr2SQuu
H02lswUvkODZSQ0uVmBCCZ8Ih8NdRt0et5TiOEf1C1LV23vLV0YCIXi0Oi85/ZXR
MULVEfBnA89EWdkEosEIlbWROqlUhWuU4ZYjm8mVkhBX8nRfGIMfKJFBe6yKKE3a
QfycxK0iSTv+vdqtvG0WKXBRpP7F3TBd4slZFm+tPck=
`protect END_PROTECTED
