`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EsVs2SVi4Tvi6/vufiYqUf6Ln5uG6PQAVzwK3rCc2fF7c3FXXlCx30UcgwvkJ8YL
6pQMyfxglkT4k2dbiEF2S8yDLtYKAClm28NcY1gmYNoq9gLyYglQ0aCO9uKSTD3Z
sR1hfZ1xHWI+Rog6RI/IpeQoFYYsoyQOsCizlNb/e3S37Cw9bJCPZYwzM0P4ugic
Qmh3eHs1Uwgn9SiTSMT+yM209X0JLyNk9V7Id4uNNb32XWd9A1+U5vLHuyWbnlw8
UEkp72QhZH9lR+GSj4EiMqVGLg/QX6lY3gPC0jH7gOaRfndTTLKZYqek6Qt37Cse
Ai5AV2RR37qb7OtpukpS1QiPVRPNIP+dveXYW6kHqyGk4wzn/ns0pDYv1EIAYNdm
LWzPASgCWZDMQ+Y07U0U3Rbwm82Ymune4DCEngFhrkA9L/pIwhIGDpgm1kcb0Y2o
0OKIL1Jnj1XpuIapf3ErrBfqgUCYHIvzNMMRvGqIFXArXrXpJpUwYkSibu1onPwS
hseMP+vIBxShozsjzU/buh9PPmHo+J6kC5lKofFKVEF8V1Q2c573DSSxRPpFhG4d
9fMaLKyQuzDkXElL4PmInLfJG7Sru11XxjRXMJ+/pPpoZbL5NQWolN4TDW83jFYo
EytnFevzurPvP05ywvPVxV0PDcQJmj7iWynYaT+UIvcod1eltvEJUYxSv1vllMCC
X/kS3/h6ymAzhLga8hcOWfTp4zFh2JiW3hQSklSr26jvv0buzX66VbIGEpqkLDhS
O55qu3sQMbLFLVBq8C4RS6Z7b7ItqF//i0r1TAaD08ZXfyiRDFxcoLEkRTNoh/1o
jd3NoJiBAJmW3uXmyF8ywZ0e96FR+U8a9wzpZxakxiOWtfy1P0lXl0xWfHncmrP1
e0sGn41kLM7R3acWslvqL6adJsbhDigoGUOgdbcCsqYYT9d6D4faA7b3+C/y3Lf2
WLgQh2K478aSO+eZor+MXeHmqqYSZq2+OTu/pIbGrszyYUwU4BS8psUSC7a51Pl2
PiSXsoj91mhw3S9luDWwTJQ5DIEJze/6SAYQvExTRjNmbb9w9RvDNqlxtEWmqZUZ
OMeG625IngUIMO9kxnRLySBR5mEYRdcleSgBjpBej48+AaiYugL3lt0viJBA58Sk
WTlM02slv/L1ri8K/zBf7MxwK5wuaPJs5DvbnZ5c2b6CTYM+xzS7wSxYsP8yWXkl
pAYvMAYU/yFn3ACC/aBz0qQHRUaQyIAE/7JwVzz7JsM9r4sAue8VnrP0CZ2WJGCN
GvqEs1kFKq0yeO9ZrSCfAUrnjD7IqdX+A0QfJ8xK5/p92uW7XDLwBbHD6lzaxW3w
iB83Iak/VXCoEgQ5zaesY97LN58Zv2PoJHO1+Gda8ynzzUCV553Bw29Vz+0IgBT7
w8uyFfUvPwX9tTiaDHjheHVRhr3HVShBy89+f5YgYC741jc4k3o9YFEwVpmYLxid
Uz11xu01W1tMf5U6AzH+Y2hbLcKJV2fC6xG1aQMkhXSijdIgZgWBDniG13bCsSCv
bB5IALVJJluj9Xhcv4Ev6fFdU63MYcCXMIkwZSFG+ZM=
`protect END_PROTECTED
