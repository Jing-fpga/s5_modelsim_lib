`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vDlL7MEXlVqikye+UH3ULxeHo5+wleU1/APZsDqrYBNYRT2ljad3ortSjmgMJdjr
08qhrIb8sM0MzrRJMIjZW+q6cr5KHX17xNNwhhVohlM+K9N9nLal223z4ZTEwDgv
ayHKgq09+YZtG4jP3Opjmlsyg3XpCgIcmNL7QbOfRcEpca4fHKXaHyBb+YQYr5I3
qthyFGyeCGMDPTlgkZQMJRA9/1lw5DjwknfSzWI/tUUFFmFqO/XXuINJ59BB9ax7
dSxaj8cHsS44Zjp0sMV3aUh9feknlSJykYnvSPwl6FHZ2z04ris7zvvD5l1tTrxP
kUCnnCWHiRfgLrLiiXGezot7Pfr2HDL7BwJpFd3AyrB4P/F4vJ5F0EaBxTkBucy/
Z/7K8kN8JYroqFONS+Uf0dh0KJ7K5KGnTPlfmKCR9Vy3AaHCzq8M/zfrBpdLTE8h
sZfcsBeEy4m1Kq4YsXBUA8mq4g+T2bsHVJ5IU18UhZ5lvYPuOzz/kT/v+lBqS5S1
kk4yYy1vuRqilU6BwD/JbaDD1IYhtOX1luMpHkeFqNdhpi3BiLIBceDh0ADG6WOM
QDVlM8Bn7XJzAjek4OeVqrAOZyBz7kHih2elYv4ZenTuNDR+ko2zHLfpRjvMymji
tf2CblwqEMM/qE0mTY1Fz7dKXEIDrku0caz10hgrqwst59P4CPw19U4x1OjI8OEm
6vGgs4sDK2d3gUkBAMHkMUOZQPN4gCysZZtEDZ1VaKiVKlVZs0hBx3O1NFPmPwJo
ItxS1NHE+ezF7FxRw2ZhLhsVPrv0Ko+WNn1bPbSYrHftfyCQTnFyURZGlEnBAvQX
yKDqvaDKl6LnPC+ET7o/8nWBtnjpElhpVa2nJnjdw3ramzepc3m4b+uTybVUXlgs
mMmIf8c8i2FPdOpTbX2zP0Vanu7Kgxhb60szaOwjiXIlqyclSEWzdpo2BirjPGoP
8mK5R79LG2p7+W0saNoiQRWW/IFdcNig9F6KA1ZL0bNHHp2RfPtndRujSxzv+/wo
2SnNT/jgK6qhBmRxT6mjpnTs3nqATS+PHDt6URadAaTqi0GM3cT0IArJyLdIuP4R
h6nXvVhM5PvKdDS6RBQUeY7FU15F7IO8EF3N/98ldzpKN7/s9ew37JONPJzSwIfp
p2r0bzwYq+jyNeAMev25e8boAer9fZFyqVGCsTt9j5XveKMTgih5LTFmsuokMKQG
Tah2UOaVodYkA/4lhQfknrkAFXxBcaOeoriZO/oMUMPpnfgePbIiJ6PQ+bX2dYxg
wVGisW05n1sIJHFoZqKJXVA4EzXK+cwLtWUneFXfFRR6/8qdkYGpIoDdQ0iV44Pi
hiIauKD3NIANE29WpLJwnSk6QKOY3gDPHLtma4EdzhwBYnr1fcwp9eWWGy5n1BC2
EQ2lKyQDgmUQjJxwq4fTmdrhw6jiKqlEW6ieqg6AkcsqBLfhv8KCi4dgrXSkjyIJ
`protect END_PROTECTED
