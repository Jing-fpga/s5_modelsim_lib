`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3zjEwdT6tbwXMDFyU+vR5FTzSLgPDxD34p2782B+Q/VDxMq5B18gneLG7k3MhnKQ
ASFruw61Ksfb/eGMxhTRjbElExNiWo2zfBeY0ur2UeCGPzJXWCjYKVdnDrr4jQo1
o7qdTcmsWAlFm9lNUaaXgoA5lv+eXqv3S6StvkpuT/f2WQpmMqpOK3rtmKQ2uszD
PA1Tzn0LX41VADymaIhyf+VhhaF9gBaKV+Qz7t5fxoD1bKZ/9J/2j/aEzAN4/R7R
1iCrZo3xwSDqsoTCBDfrwEESDBwt9yXeAyzcsXUFzL5LspeKgBb7AjWEbazROEmF
mB55VG0Jkt/ZgurWS+8+lNrZ46wjxj/QviQ1u8kabuXJx3q0rsU4EHhalBl2BPF8
5bPOVPS8S+rvHULl7qNegC4EngIBBTbHuPTp1D7RJR5Qevs8ySIRd7HHdqotVyY9
6Q8VnAmXVa2mgRLlzhimzXFO0wtIoO5BIwp6XncviuhP+qgVgQvJ+PiJSoFHGHfl
P2yTXN0tvbz5MQ2jHftm9jTsUfIDFjhLM4vafnqLt5/gaPaI0wqvZopadAzIOQbO
LBMU4dQs+kuLWcoGuYbXRxJvESWSDVPW6EBPH5WH4u5nyEAJhO1+bdmmXryao53A
TOuZXeRun75tjHBLGFPb6tZwfQum8vSAE6ln9fyyQpLeUgBYEZ1ksIlzR7dd5u5Y
lTDbtbiuN8cA6zlJcEmfYY9YA4C0Pz9ulquapqMv+hUFMbk++e849511lR1DIq5V
Rrv1DS+sLXQgYyR/LVk8jfDMsLFg02zH36nrFUVkbJfWzi4dZZUKoh5gl8QxV5gB
8uUIDjDJIPXUz1JL6H55LDtC2/YwZTfsAYDkdweFgIVpdv1ogXTBw7kN4FDey1/Z
ZpeydGU8oTgNLnwZEweliCAzeYBVrgVqF8q7qUmfKKhD9c4lwJi0iJJ2OJKDpKvR
2HnfjHsfrhvyKJ730nhkGKw5uxb9IECicqH3G6q7kPDR3TYDzET9UGm5ZWlgThgS
/4x3pgXcZfFPOm0+BN5T/xu7vo48bHyp0TtdYD32ZARspLlculjEkt2wtn25byLo
xW1V2PfRrMdiVt+Z71sP8WnRQBg41EcAG5kGLsZJojHO2UosFkjiyD0AbbID3//a
Fh2SMSLpiJhq8GocWFcdkOBcJNFrq98g1LFNrDYmWOppfqmRGsdSeuSqSJTLSUUP
xlFXDz1NCJmhQEIKrUMVindkkvw8wlKPRN7W5IOk8+0Iu29NdCUfdXrC14KPMG9+
uhDB8/AQ0IV7TOia2ec1d6jVg2TJ3INQMEM2xHec0t6dDtolrqVsl1g8xrPLsT6R
ZyQ/Lh14DVEttsdxlsN4UPvlyqmccMt5XpE9LL80Zf+WppGILXilbwQ01N4Hm1QI
xDi1Z6SW9S1FSvrnclIN+fCWGLG3bnIqlJZ3LMyYamoAYeQWwGlQikYi7b9Njq5n
o4nl4EpMTO3idxnhXeyDutnyd4652fGys5t67erIGAIOIT5zO5rFyGDqZTAD5RpV
wIZDE4oNqlQB9PmXYrpAwNyQOgD6EglUuWSyLqP86Tw1Q/ke7pbdco+vxD+NQTNL
IOSY2QllxCRzef3sIZGeHKE0ZIw1PxS+eoSUJlb+jbBg0QJsMJKO3MECnL29cfoC
4S+/N36HNzROKZ9sVyCnmPWZmR2xuzGwGJWJ+n9g6968ziwVR34anxjhbhqlDqMy
+XWV6D2bU7BO/Kab2suubB2dw/yPzayaiVN5Jpkt8LGq6vFC+wfhtq3rmIQFkYyM
Fwrb6IyZg23W44mk30S0nTcK8o932/h9uIi0zlRirn36L9OyvxyGcK/chta/hiXz
cltq903ahPjmtBgmF5QDLxCi6xiPqXDjD4NApeEfqrekXor6HsueR1CFoJwUzHr9
ROcTkm6vFRc217f1RcgaV7JM0gJQf8DZ84ICRncjepVkFZIbo3jt1bWOkB+rYNtp
ttwxc4GmJIkBdM4GbkLTdZAtVPUekNhQMFEmNm515YIBJHmnSp0Cl4AKa3ZsanCy
8YMrhW0L0e2bECYf1lYv6kGruIvP0v24uLMx/8TuSLNvj49rfv9tJ1+I0AvNy+TF
QouwsdxAW7Ohba4+NdogojWebdEjyAp21mI8fwPMn0Ym0yOrqWK4TfKiRmMaYoUe
/9orrbzF+5KSKd0XMxwuyaEHgZ8030BdxTCwo8zFaXPOKowpmklfDe+WIjF45PE6
WQpLkXjWhO/dN4ahiivblr+egYp8w/fcqkuDFrAMKZ48S8M1nyrrDcVD6uhGjBnb
vIvc1r1o9/nlfsO0XUOjzaUfD2JM2zSAMeO8McmaojH/dEKxbakAuORQwBsuwk/3
HOLYfoMLSGsj3qmwmWS6n+99vvunzc+W6q2JYO1dwdXxE3RvZ3l6TLAp+ddK3eoP
DnykLPRgYw7rgCZzGpoM6Rinp9j8GOpQYC7f+zjJm7b1/WHxH0BospzCH2wTdap6
vzD/SC+jFRpRD5V+A4pdyV4SrFAxsFhp+N3mIxwWznZwnYTUut9zCUad2KpG/aCc
JkWXGByidIepU0NiyXMqtvao9+amtYZvCnSegGSGfRVGQYJuBT56ZVuDC+PVcRiP
GQSkHC0n3pcC+jQfjXZwMQ859BQs0adMiQCl+gvcnW9WL7Wg9cxEc/G4CxQV5OGe
bcAUNcgtN73ddWFcwqRxwFAOQ6/3Qi6oP+RxRhGRs8osnBa0AhH96zKS+oFsQd+Y
SmXBKPM3i0ykOhEIoou0zWubXYy+SRpBAAhSt1KVXqgpIPtQq9XQQ/wVa9NciSj1
LgOlYjbsJJkFPIpymBtOq5aSPRYXlktxwA+zY6d9utuKTZk1vH7yL5OwyUG+ibBS
1AlI/6wOyt15kKuGG97j6ohgXKt7lzS0dVSOfSN5AFXI+gBkuFRn6fRbdJQAlqbN
GEZhruD3MWC+SqfPS8hfqi0rQ7hC8fWIIMqSWH2EBbrL/qYBkB5orDdi62BjRGk4
+51wDCSATA1Z0cFQtNGF8JUlsdvT2JyTwD3eoCu+ZsrHiE2w9xpVbowwZ+HCTiuO
IjfAXDuT/CYpXYj2TbcxzU337XUoRVcMhWxAsRYS7Ks3JUDOs+s1b8/o6gO5bYCg
NMMreafj1JMmm2viBpUB8KMbDuzl2ShoZOCTOhyQ5g3Qg7atXyQr1QSY6Ux5Mszu
LYP94TdKalu+B9TnbaQn90EgQZRAD31RU25Cyzhr/ybekY+3PGKen7fMBMewRHd3
InHn2A7PbJqYiXFAfrk3ZQ==
`protect END_PROTECTED
