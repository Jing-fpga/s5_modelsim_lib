library verilog;
use verilog.vl_types.all;
entity stratixv_hssi_10g_tx_pcs is
    generic(
        enable_debug_info: string  := "false";
        stretch_en      : string  := "stretch_en";
        dispgen_pipeln  : string  := "dispgen_pipeln_dis";
        pseudo_seed_a_user: string  := "1111111111111111111111111111111111111111111111111111111111";
        tx_polarity_inv : string  := "invert_disable";
        bit_reverse     : string  := "bit_reverse_dis";
        ctrl_plane_bonding: string  := "individual";
        crcgen_bypass   : string  := "crcgen_bypass_dis";
        frmgen_scrm_word: string  := "0010100000000000000000000000000000000000000000000000000000000000";
        tx_true_b2b     : string  := "b2b";
        distdwn_bypass_pipeln: string  := "distdwn_bypass_pipeln_dis";
        wrfifo_clken    : string  := "wrfifo_clk_dis";
        frmgen_diag_word: string  := "0000000000000000000000000000000000000000000000000000000000000000";
        pmagate_en      : string  := "pmagate_dis";
        tx_scrm_width   : string  := "bit64";
        scrm_bypass     : string  := "scrm_bypass_dis";
        wr_clk_sel      : string  := "wr_tx_pma_clk";
        prbs_clken      : string  := "prbs_clk_dis";
        tx_testbus_sel  : string  := "crc32_gen_testbus1";
        scrm_seed_user  : string  := "1111111111111111111111111111111111111111111111111111111111";
        pseudo_seed_b   : string  := "pseudo_seed_b_user_setting";
        sqwgen_clken    : string  := "sqwgen_clk_dis";
        distup_bypass_pipeln: string  := "distup_bypass_pipeln_dis";
        sh_err          : string  := "sh_err_dis";
        gb_sel_mode     : string  := "internal";
        pseudo_seed_b_user: string  := "1111111111111111111111111111111111111111111111111111111111";
        frmgen_wordslip : string  := "frmgen_wordslip_dis";
        tx_sh_location  : string  := "lsb";
        fastpath        : string  := "fastpath_dis";
        test_bus_mode   : string  := "tx";
        sup_mode        : string  := "user_mode";
        dispgen_clken   : string  := "dispgen_clk_dis";
        txfifo_pempty   : integer := 7;
        scrm_seed       : string  := "scram_seed_user_setting";
        gbred_clken     : string  := "gbred_clk_dis";
        use_default_base_address: string  := "true";
        tx_scrm_err     : string  := "scrm_err_dis";
        frmgen_sync_word: string  := "0111100011110110011110001111011001111000111101100111100011110110";
        txfifo_full     : integer := 31;
        frmgen_bypass   : string  := "frmgen_bypass_dis";
        iqtxrx_clkout_sel: string  := "iq_tx_pma_clk";
        bitslip_en      : string  := "bitslip_dis";
        tx_sm_pipeln    : string  := "tx_sm_pipeln_dis";
        sq_wave         : string  := "sq_wave_4";
        comp_del_sel_agg: string  := "data_agg_del0";
        master_clk_sel  : string  := "master_tx_pma_clk";
        distup_master   : string  := "distup_master_en";
        txfifo_pfull    : integer := 23;
        skip_ctrl       : string  := "skip_ctrl_default";
        enc64b66b_txsm_clken: string  := "enc64b66b_txsm_clk_dis";
        comp_cnt        : string  := "comp_cnt_00";
        distdwn_master  : string  := "distdwn_master_en";
        txfifo_empty    : integer := 0;
        phcomp_rd_del   : string  := "phcomp_rd_del1";
        gb_tx_odwidth   : string  := "width_32";
        distdwn_bypass_pipeln_agg: string  := "distdwn_bypass_pipeln_agg_dis";
        crcgen_err      : string  := "crcgen_err_dis";
        user_base_address: integer := 0;
        scrm_mode       : string  := "async";
        frmgen_skip_word: string  := "0001111000011110000111100001111000011110000111100001111000011110";
        txfifo_mode     : string  := "phase_comp";
        crcgen_init     : string  := "crcgen_init_user_setting";
        crcgen_init_user: string  := "11111111111111111111111111111111";
        frmgen_pipeln   : string  := "frmgen_pipeln_dis";
        frmgen_mfrm_length: string  := "frmgen_mfrm_length_min";
        rdfifo_clken    : string  := "rdfifo_clk_dis";
        crcgen_inv      : string  := "crcgen_inv_dis";
        scrm_clken      : string  := "scrm_clk_dis";
        enc_64b66b_txsm_bypass: string  := "enc_64b66b_txsm_bypass_dis";
        frmgen_pyld_ins : string  := "frmgen_pyld_ins_dis";
        frmgen_burst    : string  := "frmgen_burst_dis";
        indv            : string  := "indv_en";
        pseudo_seed_a   : string  := "pseudo_seed_a_user_setting";
        avmm_group_channel_index: integer := 0;
        compin_sel      : string  := "compin_master";
        gb_tx_idwidth   : string  := "width_50";
        stretch_num_stages: string  := "zero_stage";
        pseudo_random   : string  := "all_0";
        channel_number  : integer := 0;
        dispgen_err     : string  := "dispgen_err_dis";
        dispgen_bypass  : string  := "dispgen_bypass_dis";
        tx_sm_bypass    : string  := "tx_sm_bypass_dis";
        test_mode       : string  := "test_off";
        crcgen_clken    : string  := "crcgen_clk_dis";
        frmgen_mfrm_length_user: integer := 5;
        distup_bypass_pipeln_agg: string  := "distup_bypass_pipeln_agg_dis";
        prot_mode       : string  := "disable_mode";
        frmgen_clken    : string  := "frmgen_clk_dis";
        silicon_rev     : string  := "reve";
        stretch_type    : string  := "stretch_auto";
        full_flag_type  : string  := "full_wr_side";
        distup_master_agg: string  := "distup_master_agg_en";
        ctrl_bit_reverse: string  := "ctrl_bit_reverse_dis";
        empty_flag_type : string  := "empty_rd_side";
        data_agg_comp   : string  := "data_agg_del0";
        fifo_stop_wr    : string  := "n_wr_full";
        pfull_flag_type : string  := "pfull_wr_side";
        distdwn_master_agg: string  := "distdwn_master_agg_en";
        compin_sel_agg  : string  := "compin_agg_master";
        pempty_flag_type: string  := "pempty_rd_side";
        data_bit_reverse: string  := "data_bit_reverse_dis";
        fifo_stop_rd    : string  := "n_rd_empty";
        data_agg_bonding: string  := "agg_individual";
        del_sel_frame_gen: string  := "del_sel_frame_gen_del0"
    );
    port(
        avmmaddress     : in     vl_logic_vector(10 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        blockselect     : out    vl_logic_vector(0 downto 0);
        dfxlpbkcontrolout: out    vl_logic_vector(8 downto 0);
        dfxlpbkdataout  : out    vl_logic_vector(63 downto 0);
        dfxlpbkdatavalidout: out    vl_logic_vector(0 downto 0);
        distdwnindv     : in     vl_logic_vector(0 downto 0);
        distdwninintlknrden: in     vl_logic_vector(0 downto 0);
        distdwninrden   : in     vl_logic_vector(0 downto 0);
        distdwninrdpfull: in     vl_logic_vector(0 downto 0);
        distdwninwren   : in     vl_logic_vector(0 downto 0);
        distdwnoutdv    : out    vl_logic_vector(0 downto 0);
        distdwnoutintlknrden: out    vl_logic_vector(0 downto 0);
        distdwnoutrden  : out    vl_logic_vector(0 downto 0);
        distdwnoutrdpfull: out    vl_logic_vector(0 downto 0);
        distdwnoutwren  : out    vl_logic_vector(0 downto 0);
        distupindv      : in     vl_logic_vector(0 downto 0);
        distupinintlknrden: in     vl_logic_vector(0 downto 0);
        distupinrden    : in     vl_logic_vector(0 downto 0);
        distupinrdpfull : in     vl_logic_vector(0 downto 0);
        distupinwren    : in     vl_logic_vector(0 downto 0);
        distupoutdv     : out    vl_logic_vector(0 downto 0);
        distupoutintlknrden: out    vl_logic_vector(0 downto 0);
        distupoutrden   : out    vl_logic_vector(0 downto 0);
        distupoutrdpfull: out    vl_logic_vector(0 downto 0);
        distupoutwren   : out    vl_logic_vector(0 downto 0);
        hardresetn      : in     vl_logic_vector(0 downto 0);
        lpbkdataout     : out    vl_logic_vector(79 downto 0);
        pmaclkdiv33lc   : in     vl_logic_vector(0 downto 0);
        refclkdig       : in     vl_logic_vector(0 downto 0);
        syncdatain      : out    vl_logic_vector(0 downto 0);
        txbitslip       : in     vl_logic_vector(6 downto 0);
        txbursten       : in     vl_logic_vector(0 downto 0);
        txburstenexe    : out    vl_logic_vector(0 downto 0);
        txclkiqout      : out    vl_logic_vector(0 downto 0);
        txclkout        : out    vl_logic_vector(0 downto 0);
        txcontrol       : in     vl_logic_vector(8 downto 0);
        txdata          : in     vl_logic_vector(63 downto 0);
        txdatavalid     : in     vl_logic_vector(0 downto 0);
        txdiagnosticstatus: in     vl_logic_vector(1 downto 0);
        txdisparityclr  : in     vl_logic_vector(0 downto 0);
        txfifodel       : out    vl_logic_vector(0 downto 0);
        txfifoempty     : out    vl_logic_vector(0 downto 0);
        txfifofull      : out    vl_logic_vector(0 downto 0);
        txfifoinsert    : out    vl_logic_vector(0 downto 0);
        txfifopartialempty: out    vl_logic_vector(0 downto 0);
        txfifopartialfull: out    vl_logic_vector(0 downto 0);
        txframe         : out    vl_logic_vector(0 downto 0);
        txpldclk        : in     vl_logic_vector(0 downto 0);
        txpldrstn       : in     vl_logic_vector(0 downto 0);
        txpmaclk        : in     vl_logic_vector(0 downto 0);
        txpmadata       : out    vl_logic_vector(79 downto 0);
        txwordslip      : in     vl_logic_vector(0 downto 0);
        txwordslipexe   : out    vl_logic_vector(0 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of stretch_en : constant is 1;
    attribute mti_svvh_generic_type of dispgen_pipeln : constant is 1;
    attribute mti_svvh_generic_type of pseudo_seed_a_user : constant is 1;
    attribute mti_svvh_generic_type of tx_polarity_inv : constant is 1;
    attribute mti_svvh_generic_type of bit_reverse : constant is 1;
    attribute mti_svvh_generic_type of ctrl_plane_bonding : constant is 1;
    attribute mti_svvh_generic_type of crcgen_bypass : constant is 1;
    attribute mti_svvh_generic_type of frmgen_scrm_word : constant is 1;
    attribute mti_svvh_generic_type of tx_true_b2b : constant is 1;
    attribute mti_svvh_generic_type of distdwn_bypass_pipeln : constant is 1;
    attribute mti_svvh_generic_type of wrfifo_clken : constant is 1;
    attribute mti_svvh_generic_type of frmgen_diag_word : constant is 1;
    attribute mti_svvh_generic_type of pmagate_en : constant is 1;
    attribute mti_svvh_generic_type of tx_scrm_width : constant is 1;
    attribute mti_svvh_generic_type of scrm_bypass : constant is 1;
    attribute mti_svvh_generic_type of wr_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of prbs_clken : constant is 1;
    attribute mti_svvh_generic_type of tx_testbus_sel : constant is 1;
    attribute mti_svvh_generic_type of scrm_seed_user : constant is 1;
    attribute mti_svvh_generic_type of pseudo_seed_b : constant is 1;
    attribute mti_svvh_generic_type of sqwgen_clken : constant is 1;
    attribute mti_svvh_generic_type of distup_bypass_pipeln : constant is 1;
    attribute mti_svvh_generic_type of sh_err : constant is 1;
    attribute mti_svvh_generic_type of gb_sel_mode : constant is 1;
    attribute mti_svvh_generic_type of pseudo_seed_b_user : constant is 1;
    attribute mti_svvh_generic_type of frmgen_wordslip : constant is 1;
    attribute mti_svvh_generic_type of tx_sh_location : constant is 1;
    attribute mti_svvh_generic_type of fastpath : constant is 1;
    attribute mti_svvh_generic_type of test_bus_mode : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of dispgen_clken : constant is 1;
    attribute mti_svvh_generic_type of txfifo_pempty : constant is 1;
    attribute mti_svvh_generic_type of scrm_seed : constant is 1;
    attribute mti_svvh_generic_type of gbred_clken : constant is 1;
    attribute mti_svvh_generic_type of use_default_base_address : constant is 1;
    attribute mti_svvh_generic_type of tx_scrm_err : constant is 1;
    attribute mti_svvh_generic_type of frmgen_sync_word : constant is 1;
    attribute mti_svvh_generic_type of txfifo_full : constant is 1;
    attribute mti_svvh_generic_type of frmgen_bypass : constant is 1;
    attribute mti_svvh_generic_type of iqtxrx_clkout_sel : constant is 1;
    attribute mti_svvh_generic_type of bitslip_en : constant is 1;
    attribute mti_svvh_generic_type of tx_sm_pipeln : constant is 1;
    attribute mti_svvh_generic_type of sq_wave : constant is 1;
    attribute mti_svvh_generic_type of comp_del_sel_agg : constant is 1;
    attribute mti_svvh_generic_type of master_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of distup_master : constant is 1;
    attribute mti_svvh_generic_type of txfifo_pfull : constant is 1;
    attribute mti_svvh_generic_type of skip_ctrl : constant is 1;
    attribute mti_svvh_generic_type of enc64b66b_txsm_clken : constant is 1;
    attribute mti_svvh_generic_type of comp_cnt : constant is 1;
    attribute mti_svvh_generic_type of distdwn_master : constant is 1;
    attribute mti_svvh_generic_type of txfifo_empty : constant is 1;
    attribute mti_svvh_generic_type of phcomp_rd_del : constant is 1;
    attribute mti_svvh_generic_type of gb_tx_odwidth : constant is 1;
    attribute mti_svvh_generic_type of distdwn_bypass_pipeln_agg : constant is 1;
    attribute mti_svvh_generic_type of crcgen_err : constant is 1;
    attribute mti_svvh_generic_type of user_base_address : constant is 1;
    attribute mti_svvh_generic_type of scrm_mode : constant is 1;
    attribute mti_svvh_generic_type of frmgen_skip_word : constant is 1;
    attribute mti_svvh_generic_type of txfifo_mode : constant is 1;
    attribute mti_svvh_generic_type of crcgen_init : constant is 1;
    attribute mti_svvh_generic_type of crcgen_init_user : constant is 1;
    attribute mti_svvh_generic_type of frmgen_pipeln : constant is 1;
    attribute mti_svvh_generic_type of frmgen_mfrm_length : constant is 1;
    attribute mti_svvh_generic_type of rdfifo_clken : constant is 1;
    attribute mti_svvh_generic_type of crcgen_inv : constant is 1;
    attribute mti_svvh_generic_type of scrm_clken : constant is 1;
    attribute mti_svvh_generic_type of enc_64b66b_txsm_bypass : constant is 1;
    attribute mti_svvh_generic_type of frmgen_pyld_ins : constant is 1;
    attribute mti_svvh_generic_type of frmgen_burst : constant is 1;
    attribute mti_svvh_generic_type of indv : constant is 1;
    attribute mti_svvh_generic_type of pseudo_seed_a : constant is 1;
    attribute mti_svvh_generic_type of avmm_group_channel_index : constant is 1;
    attribute mti_svvh_generic_type of compin_sel : constant is 1;
    attribute mti_svvh_generic_type of gb_tx_idwidth : constant is 1;
    attribute mti_svvh_generic_type of stretch_num_stages : constant is 1;
    attribute mti_svvh_generic_type of pseudo_random : constant is 1;
    attribute mti_svvh_generic_type of channel_number : constant is 1;
    attribute mti_svvh_generic_type of dispgen_err : constant is 1;
    attribute mti_svvh_generic_type of dispgen_bypass : constant is 1;
    attribute mti_svvh_generic_type of tx_sm_bypass : constant is 1;
    attribute mti_svvh_generic_type of test_mode : constant is 1;
    attribute mti_svvh_generic_type of crcgen_clken : constant is 1;
    attribute mti_svvh_generic_type of frmgen_mfrm_length_user : constant is 1;
    attribute mti_svvh_generic_type of distup_bypass_pipeln_agg : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of frmgen_clken : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of stretch_type : constant is 1;
    attribute mti_svvh_generic_type of full_flag_type : constant is 1;
    attribute mti_svvh_generic_type of distup_master_agg : constant is 1;
    attribute mti_svvh_generic_type of ctrl_bit_reverse : constant is 1;
    attribute mti_svvh_generic_type of empty_flag_type : constant is 1;
    attribute mti_svvh_generic_type of data_agg_comp : constant is 1;
    attribute mti_svvh_generic_type of fifo_stop_wr : constant is 1;
    attribute mti_svvh_generic_type of pfull_flag_type : constant is 1;
    attribute mti_svvh_generic_type of distdwn_master_agg : constant is 1;
    attribute mti_svvh_generic_type of compin_sel_agg : constant is 1;
    attribute mti_svvh_generic_type of pempty_flag_type : constant is 1;
    attribute mti_svvh_generic_type of data_bit_reverse : constant is 1;
    attribute mti_svvh_generic_type of fifo_stop_rd : constant is 1;
    attribute mti_svvh_generic_type of data_agg_bonding : constant is 1;
    attribute mti_svvh_generic_type of del_sel_frame_gen : constant is 1;
end stratixv_hssi_10g_tx_pcs;
