`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rhmXIeK/8QuIdxrEC2AH+CQJ2dg9GudsPlj0Y7oOKHNWdMo5wcviQtU5puJHoqns
b0Gdr8ufcq8+WY+XIBLqcCb4gz06dYYkZB6NTvOwB7XWVa5t/TrvEj01eFIYW3Tc
lQsJc67jIQPHct/ALuZw7zwUpGHyAnhWyU/pxw7ZXNQ0JvtmUzxl8ZBGQPsbwcVI
BWsrgWQp9a/AcosC0Tim/z2lrsXnkpzgkrrjLVbh+X95+Rqn3xpX7kKFPX05BDDW
ZlL71Yo+JMJBDqZewH1tGIit/9NT6plCIDhDV9+BHHn5JcQA4/vfJC6cQBkT7HCq
VrDGl1HCEsuPhdmTuB4hd9bT6ksnJXkQvlh2iePAvTPFm3miwpXpE8KX2XGzqW/P
enaKPuTs/ScC47A6euqwPeIQOPsrvR5SbrZ6cyJKnO/eA/CazpcxWoAveQHyn/Nz
xtbSaCroEoKwxovaUXjHj+u2gJFpf+bLFvmocL8tq6SmKKQ6tYXtmZSPGUIQ02Wd
8HWlb0yqbEjr/dKP4UODXUOYbzwRetHpK2NMltYFa4EVsAVNcHjLfx6jVj5h3TLo
GP+4L6VOr851HELfHhR2GsHQ7UrPU9g2ys0STaRmdOHKcOTEAGdjN5YoPS2SpDRM
Fa5C1dcHzB/fVLw6wooySLkCuNA5oJNnI1xBER0pP9xWErvqabGUA5CFzjQTRBzX
km20wLPq17KpGjPDm0cWHv0FoZGfwwvScBfCIQQDyEaTVGE4ADeoJNT18HZcA4uj
S2C/nctVxzTh82d4G+VTXVN+fU56As50u2SZ1vPEYHgLOIoQwxDDuGvEAdcKHNDz
ydc8nFANEdc9K/4IVsTnsrbvSigxZWcb9znuO5z/jUf1taFA7u0E5yIEiEkP1aYj
/IhbxXB1SzRvNPze8UzoMUNKDrK9zGN6fv/fHhVNSVDp7DemrypG2PuWyVfiMQgL
Vmm9XJ0rL7q+wsGyTowEza5U/GavmRYPm5dw9G5k/5ClVqtK95Nw+f+p8QIadZlo
ewEj7VCpWrxPzACDHtWE+bPrewMS8KTb6WXu3NJBJBuNg8VaKBWnO64UpRouG+1a
xg3EqtbX17W1FdlyWRITxAOqS82pXHux/jxVTUcFOA44kRCvlfjqT8hmo62dWSRz
9+QBmI7/GiOGwT2YQ6QWDsaqP1nwUjnfmleK9yjZlpxQeRCakzKuNNujBQPxXArM
TeP5xJXKAgK9h5zanPcAyjG5cN1dJ4KoVM1Spu7EP/YnOfce4gNNC65wS3AA+Mdg
SfaT+Kz5w7JaGzCHZhq4tuVlKNIYUvbzEr9GZ1EEQ6vfEr+dtMzGjvSN5N9j6HlK
aZ4/NJdue20a2Ze71si+6ZrozPxzzXzbWQOsLXqEieMYnzSi/1wysLu18d1ogdsg
y0/pRWV1WPZMU37haOjGc1a4AFhSQzaW6EftNbKHWKkq6NQMTTmhxh7IPTcPIAod
8O2vAdT29cqGMh/hv+tYJklwWzz/hO/KSwbNO1yJ/jTjM1GC6C4Wo/TXIIFSyovi
5BvUjbGIY+VHFYTTh5w/0UnOobx++GP9wtgih7Tu40cTZ/qtukNer5USKot1BzSV
bHjVlXU7X48SeauaHFeQDm7kqfbJzFiANXpZZkuQUtjtFrbvM5iWCCvhItJyiF8f
gUg8bYP68YaWNVpubqueCQ4wgUYpi/R551bLPqqdQvxm6ZIdsaGZpyclHna8D1Wp
NFYwT1C0BKi0C1V0JjQUzUWUsFdnUStqBF7cW4w8IAqSKEHnN93MGZIYMktdLMoX
T5wlhbeNZ9H8Q3/pkJzXK4Gwrpl1yHaIdbxnTTQDibDjnZyI6QpnTX9kWljAMIc+
ZxdKuFcP/fIAXgcUZ/CkiQ0aCgxrXxum2BmRJyS9zEvvMZwek+TVLD0uHvQwGxuH
o09OiO38YiF19eTWLroed70r+EX2avLnvPnXbtf1hB8TTk9mepwENZeP23+Hgsyq
mWXcBBFksjoeoX9MPpKOrnMsh1w3G7/tSGojDqq76iqH3AbgM0fHQtXmvEMWkTrc
i3d7JTVkas7smptqOzYvVuIcX/yd5J0ZNmwq7LBuxgc9tO63xsHLY04n7FdmBPHA
TJgVQqKNGvzOR62mrjrJJfBopdgnBY2/TUpsfkpHyFZUOjGqhop9MvP5EarShPe6
KueVDkf28+fQT6XBS4H2cKW7DqtSg5zYM+Rj7lc2E9k5zYv8ix1UlrD+IUB8p2iR
C+bvHINPbHPQLP+uhSNA3i7UD39c+Iqt9onWxhlSEJx/lFvnf7W3Fz9q2l5CxKb+
sp6ctPFJNomZIIxScYpq1LmYIT9zaj8PGk3qden47Qozj5yEphaXqHiYnbCVPMkS
aIntAxIPAwCMDLNCuYRns2fTA8gVN98XQl20v3kUxB7wzGksl84NikxsL3awtMv4
0MoeWJV85bRvGnhexxEE6i/9Fznn8kgRNMUpXwWgn90c1G/u/PfRBHXCgGRZnF9s
LxYpkRKTLpOzHlBHEh3e0Xek/VNhfSUEdZSpzlB+xD0UiK6WpEJAMTSzlFFBLJKD
bY8pIu/UVezy1svlnt2hwaiA1voWH1nBmvizcCRZSVuDYFQc7Q2pHsn6ZJen8CNu
s4XqTu2vrI1vghGQueh3y1XIkw+2RDbgmR+R8SV4QbvsJZDuyDUDgituQqw2XIzs
VTpdqdZT/+eZYyEu8wdfqXzRhJMquW1lw26kok/5LldwEU4US9GvSlNK/70mbVvP
7idgm3CUC+c8tvPeWkF3wKMwmnbKr3kmmmWPh/9bn5tEHbc8LAhqFdp4DBKyBpL6
AjH5hffVSvT7oLOWlo0t8VGQ4k7W2lOoFHyTR6EbC5imrL4n+Sj5mCrbmV164Bha
QCipINH1DPzhdYQr8x+JRK0whFfav3nftNf6Oo385G6Q5oDX47CGC15Sz7fWWzZW
lVKh3nATnIoQzDNf49JuJx0+XOOVep5mwxyM8fpmodD7n//cgCzajLbQ5qYbC+yN
C7cTSD//Vs6ouzUrGupPOafpUYQkRuCdSJjrWYJLHP49u9LMaOdEHaqc8NblTY7P
EHMeplooZvEpS0TEjl9Wtq3EkYgib57l8TSMXJ5P7XrV0NsaRKPeOMaVicV2X/+a
OQf1BqWqQFjEciurYfNkDlB933RIuJEHA2CNEUi2p3i7Xixc6pUqGTS6mnjNllJ5
3wNJipp3R7zhFEGL1N+w6M14faVJr0dokECwAKTE16XA0XqNfDXYZHyjuo7sro4+
fj/2X/xtdPEbR1SPp6YFueyxdBPM7UWV9VMonuEomUMMHiVG4uyspIeTWdSF8JkP
9L6AbQ8TEXr9Gizcs6kXtypugD7B8gpZGr6WDnb1JiGF0W9j9+nvEwyeLT8cdvZY
zKsW+MR0Ti5ADrWnO2jAUXimolBkkvzmr4iOWEIuKJk37nAxMpjcgXU/NImdKH4j
C2GeEmtEYmMbvAuaQUyug1KP9hMRfkOFjqwW+f0dU04+DjiSxEgAi082jIPhL97O
FW7FLEOhj9A96ReKQf1Qn5NrFRwS0+PaLkUIPmim23CaBGnO9633TT40/VwkJyO3
HaWMhGqKAocs8l2eVKrtOR3zb4mURO9gnRgY9XEplmQ7/EhJMOs66zGXMCJg42Ly
CGujnn8MILUc63sFUe8KPnLQoBi3IjN/oL8Sx+a+vxOFBD+tX5NACNJdNHTEFrq/
jff0fjZhCXGb9JZFYJOx0ac49yxzzbmn75hZZnszj0bJrvypWbvg/f7vL7ZYSPkg
2q6PhdZN56K3/0skPAj41ap6dWsPhiyf0E0zxQM/Z4sZp+0kFqOMbkpOXzVfDIOX
gUyUmJSyDyQWonjZxs/9oNUM7Bf4A6MxJ/yrhtRN0syChb/RqowIzjLEI24aI615
tJ4aWGzgIEoA0ROu5AWSJUhCzJkGtfNainh4aNmSvDO7OHRrHVS6Z/Z4oiXJ4rnF
m5m/3iZQdaZYz3eGBr8S4gsFho6Kt/KggQCp2oDGjOUKrqal2ho++ky8iliiCj/k
dl3Z9k04Ph68UrQL7StQiDaCg+I0WDrn0KkVSSUBjYTPTbTL8qvackoMl8We7D/u
D/IdBj6fgyEs/FTae0F8Dwb+q+JfRwDBXAkYt0R/Oza96u37rv9UGh3l+lJ7jMBF
wJ/uZzJ+qaYbDokhNdE4ZN3lgf2K+r5nSjlfTHlRsFcfuxrpZesdTdXKmz1cRrSn
yrqp5DKBA8hYnbN+u/SL0aInktd4VQwatAa24gZKyhIJ9Dh9FIrUvOpo7EEIAwww
PDM5F4deamEu6SihdaazPdGAepBe75Y7uSXcY5kIVOVcwelziciS+xbyt3vb3q3V
zeF3h8VQ76idQypvB56R6Z25nsiPV6Bd3jn4qfr4BueuOS6115rCBngCoH5MuTf4
XNOWKxYkKSE8i+JwsiyNUfIME59Qnih3xG+N9dmW3xg9TyzUibkZNFraniwdA2Y3
hOnzgayB4hzB04MQBOlJikTdlUxr8OpgEkhA7gostFofKC5TpbfqBxyL74DkWOJZ
GXVZ2kvxwH/7ggzER0Whz+zmxKm6ChmQuyAcKVlh65jPUgoUeKEVTMitaGKKH6qA
F5m8kXcWtihOl2XgY7Z//fNBSvognFNndbWU0JeuwXThV3kv86CvZFqfTVAVeOGC
W0zkX3Kxx/qamVng0Ah6eSTkZDXJLOjot6Ad1fA6aALhk5fGQoQSTE9qI7SbQFA2
kVFeYDq5oTjEVoIqmg7OUKvOBif17X4WwAw6YH1Hya2e2bbMu32SqWq6o7pZUhP4
6GYAldOw1fqrMGcmND7hyFynEr09+NIR2IALl/LPrjjUdyAPoaHTNLVQCSf9JSNo
1C72TzUq3SiCBDLLH+mhkJcsz+HcVKps/Dd6/kHU6vw6dxGzxZcyIolb9S4x02H3
/tuFw8yYvpM6yGGF95Cfj0aVyWS5mZXzP9Oo8ZsI8rzmf8NLXz/Qmw4S9jKK9LQz
0j0qomHLcS1W9Wal9Vv+dBExpsEUoeHwkfcdcLWIXzhaYP5bzbtlC6M3ABp9ZMn/
pg1BLj7WMNk9JAegxC1/grTu7qpZViPh8mR1LocfX8UBV+6ZEu29IgwOCdpRDwgC
rZbVZogBC1u2vdFJ0ajhWrsv15KoZWh4j88q52wQjia5vwet6QiDfbOdOTz4t0Ww
w5xqX8eZ5NnfEUqbLbDEy80dCwxwfnS4gjKf8+skDj1pwqJ8yMMKFhZYMYcXBtLg
HzlQXWyY93nOTfyGUcE0jimF/0OqTGE3LmdgPe4PHTtfv4OCvjV/Yepwd2roKcRT
OOubinXJMaFnKEvZtL6EUtcmAKHEHsBm0jpos+2mjhGk3eYrvKY4hdONXAGvI+HZ
0fcHl8RFdNSq7q0VD8MgofsyKCjIGKgw4WQfHqX2to3DvFhXiTbyuOPCF/VLtM8D
MdJHM+HZopb+rdWL3etYxNJfspNALmBWw5bMkpWLNCH2O8Zmvp6bJZFVlbjUqGAj
qP86kkIrc4sGQXsvazuJMwSTIraVMZl1v5XRSmnETtyUr55H+rlY4WEumAHC+G1G
fl9ez2m+oZYUNLf5ukoJ4ELU7O42nueIOB3MrOaMARiqnauQjmmxGY95zfbp9bQQ
uKwPdPjQAW8ZFo64V0Tt1k0Crf/JY8rrZoG9iYMPbCvqWycXjKvq6bMN78ABhqia
ro2B/tbCRG+0VchiM2xrKVy3vOPhZ9jeHGYWX5Og9ZTe6n5b4dZ7kSeUJD2Wx5u9
1TdrflwEfY5rVjOxzbOdN35/UHjNVSim1P0NHgAvhnIKwSE5RMjzDj6L82LbMEVh
uH44gld5umSVysiSmrnLA3ziJQxDGW6z54xZh9ZTh/oOxt2j3bqPNjP+kzY37jQF
hwoeotZ4cMHznPap0LzUl5Yv5eRL8l6ZzIQZyOVKRxFwiKydMdgxQb4s4FkOW0Se
HhLxoHTiQWbIiyClzNAaYq/ETwqSp7zXQuktvF7ECY/tGMrWsnY0YZ2C0eGmVNxN
2ltq/zNquplyCm41ytqaPuf3brB0tn5CA0h8uUhhS331vBAqkyaO3XWmAcpNc22B
TTz+uLaxgOz8V3BBA4Jo4/Ve9QNN9yhrI2aN6e2WJCDA9yJCP374hpfxw8xToHDi
ZzVBI8wIpYj556ohOwUAjz+3oKcqy2fDmEsWeL22GNj9rYhsAhHC1mguXemjcCu3
z+2/p4o9JUzpvsfSWpcbFjlI3J95uHvUDYO5qjFdEjeYp6pFtxa0X76IYlVqNmlH
HdddnhcOd1hfhHahqgQI0wjv5LmSdcIOMatS4Mg5CVhtVLoiYRmc7drAyrg7blnw
gF3hGsKaYDcgiiSOr/Y0+rub04vF02v2z1PHJXxZ1jfdaJFtmetWo7o1zgIX0XFv
Ixf8AD0PgI41CMne5LlxbxcM8u07p7MyUtiQ41Lj+8etgBHQaJUPkfciXFIQtCWb
eRQa9j7PV1/VpTDvXbq+LWlexRO515ae3myx7OTUkbH+vwQEcymiSDGydWs+3Vg/
dGBmQCJ/nSL/SGhi0/lgO1mWGDArxJKmKLq5ncA5/HdQqLYa5AlzeK5+cF0qtg2x
dfts6yeZVirOBHMwjsoAxGcEAnp2L2hcysG+vztTVavzb4dXiZv9l1f06bTIkLD5
H0vT5pZ23UNbUILtPv6O8FBl/3+BYnxRdzX4oAYdDgCpi6RbEiN9P/WC0ikNuL7w
MeXAE8CulJcrhZrLB4CbhfzPCNgkTG2qE73Ypqo6j4mw86CXG7v7D08nYTSfyoLM
XLLabWZ31o+mGkdRyJGYJkSYio4rLj/PgnHEBzDHQ74BBQU3/003GnL3EiwTKwdu
4F5LC7SCPIx5MI4Ir1xPViJcyyyYCJqBNPq8WZpwTnWgbc3B9qdqPVt5tfgt4wWu
HleHZzZVMO+6IQXGfnaeIC17Aa7ydMlqPfuTauJXp0xHQZ7vp/WDMjQO58KA1zAt
p2G6hXAc7EW0Ndpxw3qUs9VWIuFGjof4ZWPnkfpmKHiJLkDYnaTcL3yxju6cKj6e
mrvSoj5uuzxK+N9ee7ltZ7fqBjUqI+X7vg8G7Ge2RoGtQwkvv6m5pZWFqoI99vpL
Z8jBaKsseoMqqO8pjjY5V+hRirOgROVVZ2If/vsnXF1F4s8Nu6xQN7KLfSR6ZVQU
Uaqg4MsN6cwRs6QY6Na2x9pepY1R869M0H//y9s7xXLmkao85XHfM+pEwrXwyyEg
RH0Geho28DdXUpXMaGEZV7gcWSHzIm7vUKN/XnPBpyxDDx+JZrGZxMmMmBl2/iCW
MPQ6Otupzqm4G3TQJX16Ag+4GtRW6XBRaULliPTMsyvplYufd+hqz11n8MjFZ0SK
815XMlMgtWyoIXR5jndRTtVfjhmKSgVAxY87THVOj37zXhJAa5AZKcQ7nNMhCOXQ
FzYHHAIQzcoBsnFRm0KRkVDJkr5fQjHivhLPvATQSDG5Um6KdCiBY9BZUFf93WO5
dNc4HQ7zVwkZwFE5+AiXuPSg1Ncg5gbszOCQzC3k14fWzD73bYDMw4dzzBPJg1i6
PBDY1SBH0Cdswf/VszIZ5prILLwdXM4F+e4hIqxiK4Q/O8tWKa9qruGebjO/6DPY
sYVMSMdMfUlOHoqcOwV+UxfRHl+ME5NNBfWdgHlC24nMO5ZL4/bPnOszFm5BBsjm
itwTyPKn6NBDqD6SjgRnlRmfFBcrZMfpsLywvIqXO8S5LGJW/aXp49zAzRpoOrIF
UZb5uGlJwE6Ov4yT5nPmlNx7tiEt6jYzTkB+TLFvjVYK+ZQhXFS371fZ/UF/oQ6/
RQtJot0SDN2sXQtslDBY7BPV+xJ2TTRGm8wI6VOrH3td9nuup+kSoJKDJZnI9PZU
wKr8NPJ/J8rQ5AR59Q8r1Ibu0IL/GLn1qCeBtjciAHOkiDzny7fCNtDidzW3OR4C
vCA64R6ZFFrLfDZCghAHwd3Lb7s3tDZgcq4InTNlzHFkSjRsHyMoKXbE2jMuZNT8
VtXD5p2T0bjhgSivujTRBUvhB8CcMUtiD0W+tl5b/c6tW1ya2MjjpSyuMLiH9q9k
jOn/Br2BOaB+cNWf+vc+uOLBWCLzdFgIwAs/v77qgRtNyah/qAL3SHk6xR6VSES7
baqY++1Ntol2+aJ6UAghXI3KHBzfRr/FHMTQDeKSxMpUM003KHUfDnMgwItUudzE
sYopUcORp7CnfESYm2dC3m3zCxUHVvWdYfkxEj94EFwKWWJqGWShfgKOMIa1Ndrw
78+nsUGsA2XJYJQPXgQJO5CqNwnhPaxLie9NCD4t+T8AjtZykYbQZeqm2pMZj0XA
YJPNEwkt5RwqFWiu9tcYxmjBGFAtJwV44oNtzREC6u+zAEWuFm/g7OyyY3G6srl6
Nzz0LSPChSZd12IKD1Rs/PnHJqETJVFKFhIhZ9m7B7qGogzzh/qG5D5RMRPY19w3
4ov7fIb7NCV2hTd0QVoIa8tR5uzdhOM4agnzXom8ve5NJJ7kqH5+KcHTstlK0oeG
/ZnFEFcU32MSaZAftySinwtbDnB9ADXh5cEx1gqDtwcIVdWU5Q4VLidxNULSjW0n
me3cpfsCxw+z+ymDfTr0iOCGVLCmYOtISfDAfve0riCboSk4EA/YNyx5d282/cf6
oUEc9Z+ahBr++RQ+zrD5FrpbQYdjL5wPdf5AybH6gsJYEpmxC36dONQ90nGarLay
1qnPsfvpZyp2QpCrshEE3byam9PQTbNVIwmED2FcloEX3DcpsJKfImh6Pho+GPDd
WW/mWDeOLJZw2NIo9+4Z2NVpBGOadDz4xgA//5de/by4a0BEP1We+Y7lh/mZ7zvZ
PsUfMLTec5ivImx6xw89RJSnfuiyZFhO11nwrMJHgDGsEcnOpjSlJaLZsPQpuShx
vw9zItQQKfhgc4wogR7lB1Bg2azDAuQIvWHW9RKt4juJE4mJgDUcTQERU8jdyfk5
r/KoCpoCt9wtmrYjx6kmsdJnIUax1Tseawd6qFBRReYXsLoD1xfV/CJ6bH8azf1+
3FMPuJfzvaofWexys3kPV+HlBEOfj0EEicUI7YfQxQCCqyCvzG8gr6aUb50djUlQ
g7h+W3rjwBuTx956zveDMmiMBhLPf71m2GUUT79krsN48ZydMN8aCUmZnRKAxCSL
5FAvtZqVjCWpBPYkqJuz69HTBrob2+GwqeCgV1H7BtrZpCC0xH9cGJwfHgdvPLIF
V/Ija9dtt9pupMmQ/M0YjJasMY98HsYQiPmd6I1vbeq6Tb5yKYns7e0/r4ytWbzn
p4u8rKft2DeBp5YUc6rJykTyt4ZZsGI/oUltGmkeD/vGwBYPGm7Qf8ktJAEi/X1h
4Aeoge3+GzsL7lOCgIeWlwt4mnfxYIdqm2yBZkiJSP0oKqQj4cVEP4MhRQWm9mEV
O6vIHQdQqECRf1CWBe7hXTZ96K6NAuRdKZMp98gwkzs2liqG8o9/yTX/wy38IUem
SCO55PgY3L0Jcha6Agk3eR+3wA5SRQ0Fm0zE3yjMWMjSLXQ47RbtAbERlMyBq9ux
Pqt0Gf4gs+KB9E1XvzBy9AUtf34sWf5fiXT6nRcCNhWvoaZadRQ9uoJn/+2h/mF6
63rUaoshcScgiN2WNJU4rUOe7MgmaadSbSvLudDtlviedT8dpdMxfYL6ohaUAypa
18SoL09CuYfS7DxLXLk5eVJwVbtQWbTjj9R/tEVoGDipLLKQS70dxMo3IUqIXz19
GROo3xNkxa9vI6UgzfFfLybtBRzwyNgnzhmFXCj8d1vT0sM6pifAja22vGmHdNrF
hbCHfmTxkjVtRpwifXsLFabLY8PwdyDHO8SDkOhKmp27mF+gjWeeO4XUIosNiutx
tUu1tqknd9jBVxVYYRXd5JvvEKx2Vp0DAgXalkY8Hve7v6Q6js1qghBe9RmdByr6
ZJzhl/44Z7Jh6/Em9jp7J4/nXUHB3qyHjsnSjy41BzGxC2nfN0HGkIRysqne7dBQ
ID/YMVd5tDNYG4LSZcYFXKTet1ojJeaKU327O0hrBW3tcWKUUNDoz89EsaQjNLEr
dvfXrN27sTUFfYgTLrH7P1BjYbXooyBqDxbvHVXUJtuXNacpXmeuT1klfstdyMJm
D4xswp9Q7ehBM2hmfDtsRFsJYUEZgjEDJrUF8oR+TxiblKfK55zoB9Xbccec3ZHh
z1CPitT3pcMBj7zsoCU4e4S4F8p8I4Alt1pG1WKCxYTEcxuIME6Y1ilZso+iXvh5
qCK+S9yw1/jpds/3If+UZxoHLqswquAx+Fyna8sAw9VKHgA8tjgkwrsK8qXRuCmh
Z6PR0rukqs//Z6O9tGSQ7oicV2agRuftepD/1wUuCV772DOp7K7xfANRL6gCYcXP
B4WUmyGqviBF2/pYzpgGaLwWolweG+wGpf/3DuWmJlAjZxPcaPjnfASD4Wbdd03r
G5aAd3hNDS6B7PCy9jZyh6EhR0SRSawOoPCwt0ox63/HMJZOBZ9YkTgklFLtqezV
ebv7Ic+Z4F3vNvLWEXdE1taQBeFr32OsKvXB0KGoDvnW8iRxEcUTzXDbBh+PVSOX
WpIuSV+ijQqf6t9wPtYkE+Vn5WOVPdbFJRKIkhiK4DSxjV1I++0QfEEvsSKRKaCP
RCwEBBywUv9C0IOdEI7vIX3A+nen102isGxDsq4b53i1uHaN6S41whdF5G58L79p
fi5sS2mjC01rcQOS5rAH33WaUw3raRDkFXyHx2RE3QFR50MIVHNyQiLVRyxKFOvZ
HCMtVDrReaFFPY82DhjjFG3axLgnzCi8gkoUZ4iHNO5nCd5ynwTbFITCO/vQln99
t9B2Ib7iOTMtdN7I7DLaKECsCZmzsc7y1o63lCai0fo8zZeoyw/JXYJ0ylHZbjy7
P7SEoSjHddJ6uNd1XXz7OO0vxOaCgwa58xh+97fxUVeawyw/RaOeGN+4EaHGdx2a
aCGuD6o0jJGnMLN7ORG/TvWGrQJGYUxHiwaMwtJUzjHXeEoTrZMHt2Srppb4bC9A
A/Mv0exbe3xj/YEpI97NEVbbk2BkPmjmI+GtqSqZM4dYKX5naGqsj4D42Gtl9WVb
MwQQ3PvGpWjYmsACO0NzAesGXqmJtX6A++G3VaFDvY2YKJB+xynok2bpvjcsEpwu
7co8+0+IA57Ug/YmfxawiHyOxL7Nxdmp6Jrc8H3lM3EfJNDHHfi3GwWSnDb1z1WJ
2Ej/L2RMIBglBc11G6JBpUEVNtGDjp0SK5jC+RerF7roR3w1ZaUNiyLcu3yioQVd
FMetDkv4QvVWHFxH/yw8w1KEs3f0MESVSEc+JB6PqGKunFLWOhF343DglUekSHm/
fS7Qfld4Uk+jgTZLiFd4Oi66dbrn/xELn209LkqEIq4Kf9L+TgB6umLtsJRPnJZ1
vOu5PfgemkPuG5xnCcKlDEf1WYpgkvP7f7olewYRjRUdkxjhOdJs0HINOqm4riGr
iHMvGTxqZJrFQ6JfO/aPtrzmiQRPzXwkG4t5t1yAEfCNr4wrEOapTNoRrGJT3LNo
ntRyPCf/5CrKZPobicM6H5AGFYs0oM9n887IEKGO7LuAp0NHpwvAcXB13orkL3TJ
iFkoR7xct+pKDnCNVs8MJeMI+YVxPCPD7cbVEJWKcsstqT0NX009daSrKuSBRAP7
ZsMeZBjF54FPZM6TVxvKA1joiRQFXLIoLz1z1KvjcljQe/0o9Og8nxkS5waUzdqv
HQsxYRgY/Z3Fpr1D+mQOBmPgCw28rcqBGd8suG1mvemnEOYwYpWas7NzG3X3SfOO
bfDHUzb/XZCY5pLAS8b07U6A/18DpxYPqPHsJtTDAF7oqHDhCbabo0zxM8RjZlRG
GUji5GDEdsfFx9VHt6ktMz7kiFkXgSnbOzCDBm4jawhrTKTh7eB6oJBsMgzBTAHl
suJ6jEsljiIdmCcavXhdUjWizMx1ewCKn5RpHYmYuW4AbDzqiESpknZaGdL4Xpxu
9NBq6LRy2aHs99fM+acQPaSqRIA1ILLMRBGxUeOEN6L+b8RaQ3qdpM7jLviZm3hD
17WlWMNvlfhB/6tbBHZjuvhboAl5K5TqxalOk+NU4wAQ9+eOY+1CL2wiK8D9IoVm
1I6Pr2RN9hi4Wk30MhF0qt7sL5IEUlRcfi8r/mN/LjUnNam0kFdZJv9jJLiL3t6r
/SogNROkZ4c5ouUvxaTkevtrwiNKVb5f6GW1H6EjMPxwnOK7CMJ28D01NuzkucPY
KO47L0x3unoOd1ohCYdEXb6tkIPi9VdLvkGWLy+zXaIHmPIqB4V/C355cldVbRt1
ZoivIJpBWHHaLXUwBzGjzbxK31g07LZITIHizLnQCETDLjvQbJ9Swooj85I1f1SW
io1G5TSFCyt1pKskAeyfP4Qj6e2YPqpkUVdXzqm/44w8vqJnw2nudlFBtT2yO4iW
c5hlOeMuvqhUYgaIwg/McLW+1LuksjaHxLvjcexDTYy3XYadHCeXmWyeC12+slha
3Nh8Wa7K+6fkF5xtQX7qJR/L8YGA5pj4L0r8Lhr3Z+ScILBE1ogml9qmbBDseoUz
nhJToHC0ETNcx3uskWW2SO00amcsE2jj0X6MiDsLtJGsWrcdrLVT8C+DJIESAiUi
mgYLjXSFqHd5z6I7TRcKo5cL5QbUQ0Dcx1s7RgHw0LcLcQ7bDCcDcDIzd30ocyQJ
pb+w2nnLoPGhwyBODgg2NQoSg9/PmJqvCwct4vox0+Wur2fWL78u0AAHjVb/Iw1P
GwxooOjuXdZQt7k6ftTJF0yo/F+G01z3nAdL2boSLuOrWALQXwB2ZmNi7cnecqFy
9lknHXLbf6y1hzYK7Eun41LX3IrN5itjilQpJYIPnfCXAb4bVIYgMQbnCXKLeGmN
ijaEGAPnNZ7rZfD+wM5ClnoNswwTytDOJdKkDNQdKGy+D+DzU4M7iCXiyr2MAC+R
hUPe/xKu2368kNpQUWN7Vu+b0F4k2WS1NGs6ChVvGqmHpAg5LGwWqLDn9PlDJQ5V
xLcjebuQjmO/wyALf40sA0tsjwYSzdUsfo3vW+fpWcEivy81JdkgLtF7ZBKjy3jV
ZCsxnCwM4lsezzeOwaucN+RDDWK0qDq5+6G8fBKxS1chu5Gu+1iydWdh0saXjYj9
FY5xQj7WEgUFTcQsuEGYn7nWUnli/kbK5ycuZ3elPU8J8L12JdmSxNqXT4YCbz05
Z1//bNkGOTQJHeBDyP0MbH4R1/U/FrmX1JXiuj1d4Y4fxZ9Wn1qP0w4Vm2SUYytj
5vAZRVdiuiABzwwq4hnGSU3S1mZmLCasB9Y9DKLbgopO2UkqYx8QAeg23/hgcqxS
nPGG51Wb4xJaM6ysZqJ1yWYp72lMm3+RAuf7utuaT8Gf0gP1L3sTLgIwBcGUZR2A
RcNrxzF6tMTyYv2ToIswZHPZwp6UsyM7b4VS9JC6fghvQHPf0sDyzj/8CIzy9xbn
vBImfWglYyjDyJa4+P9XTF2IEbIyKu36jxuumYX7/fTfn4zCJMoSQqsNu7uP02R9
uWH/BDdQ7hbEyQBtITLaGa8XpBuRXjEYChRfkGoij/V93u/S4xTB9Kn7JYAXpWi4
ax5sfnHTJITmNF+v+TPDHq5NqpR56hdQhph0lrq1fsZVwHek2SRbtubLcqXkUD++
JhNrskxMxuN5pQtos7MMyRWLkh2PuM9OA5XuOMPnUQu3urL6HH7uY4oiHE5YbPMb
EguUpQMsiZTlbWCz3Yr7TlAIccu0OQWT1hWrZ7h3mICx/QU0vUfNxiidPGhiCdZN
ToFFx2Kp/T7cwekdXbxkWlb0xekwhCIMYMUXXvAQZ5gBRE1EMD8+1YbUWwX4naOG
vENI8SNlimwDrzRepHbKsGIXX7ZQREh7mldA0pcMGE9Kpt/6iOhXcykN66ac4enj
tURAqCmfim9RPcBA7q3M1/3MczmkHO6TwqDIj1H/SQNMCDYl33Gz9kp0ANNiNWXc
gxJhSLV0YU7T5mBtrGutvY2cRIRyn686DP+AQjs4YUphGT8ZlrLxutj4G6X6rUta
7YfIzgJi0PQfOZLcD0fx9Q6V0ZE+nS46V62Y/QumknOnGTN5COaZ2TgzeobAmg2i
nsIKSYozaCmQScQ6nh1WglsnW53ipsGbQwQBV6xmxuDFaM+ViSFwLt9bTJCTr3b/
VmMTaVcBGNk3eaVJ7Dpl9NCFtCzk+QROl5w/H6/TOptTwHAxqhMSd0bDqn4v3Xxs
ITmSs7IHrbtWJHyOZ5dikda0jA7VGeLSvJnEDPu5hfFTFayzL2pVvFxbVf0ocON4
g13ylyra0z7WMAtHZTGi7VZXDNYumqWPWy6jGhzV90ttbTeMivqvMlaASY0DT9qZ
UzIp4TTI0cugTej43VsvaK9fS1+HerJUC3kZCFpAn6ch9PKgwResPqU20WsubW9s
mWuhrF2AUQIbHkGaZocbIX2xJXQB+KleiHHxUL3l7lcX5VR4mEXOJcyZwl1D+FB3
4W2D8DAvRUAYzem1hyJ6MpBcPLf1BrDAYe38/QHDoIP+pOMsMP0Z099tuuDmfBos
TKBkeJbhgMNvxVWuaaVBOLQkAuvraP6PDVyrBqIeommYvBGmNNMM60dq8a5qryZ7
gGDLH3J28VKDfblZZbAueYDnGUUkvWIbub+f4fwdCcRpPyD0qfEeNt11O+QM5xuY
tNSatSGZskn1O0qBmZRPAm8b2Mbexe1RMJsmUrN9RJDmUWfeNpNWXtzLYbjc6ndT
kJZz87+PkeTy/rRRYwDwuqCU8gQdsVcVniUHaJbf2nDiHmUuWKYcxBrwMh+rKJ4R
Mk981kKHvnmrwsDuhFgXt9ZNFIMR4e+UKe/HJybNPiL54LKvQZtGpnY0M+MMCQYP
6s8SS2FC7L2BeGoxoOmYDu0qukzajshNMzK74gTcdwzYYFTVwHss9VoeIii+a10c
z0JIfWIrMuCyrA3Z0oGyXObi99an9xaphx9FwbVeQhTUjgnAZalIQ3UBKrhA9HkL
bBf7mALaTxdite5KjWrxsXAb1JFfyB7PIjCJysxS/U9NTqWFKYABv9cgOeeFcIaW
dVfxRwpWi75NRUmg88FeLN5DH7wMHku1dVIRZ7rwd4JUTpE+ez6NDFPr2qcpT+Li
9gM1EXeXbqz2CHMo6ItSPVmK+5eVVNuRACaj3435tPUu3ZiMnMm74IHViB5FvGjK
0O75tpdXQVw+kQlhYopbZL41BAR3c4evhsUJ7cRF7A1gm7PXlg5+NQ2cK9NbpIdJ
eVG34nLiTtic6Zz5Knd/QQUn/WiZnpq9rcCZc/vkdCL4Ek0uoC/nGG3bZcCIBR81
PROCdy1bB7hrKhd63cJMU8e3V0rXtuKRGEnfVtYdMpK1Yo4xLRE7PzdhN2CnFx7k
MqB62rmFNrbhWTRoGCjk+fOW9Q2qxb2FySonOyh36aOKETgdRIoJIe8xs98t0/RO
/s5ZXTd7YoEr5LDnkmVDM4Gbaekvd/lghYkEaQigMWRb4RKpHfFajdD6OGpe9Co0
iHk2ksYtJLYJ78ZZEQ1Q5hCft8+HB1PO5dTcv2CPWmZ3diJW8vDteGW+MbtJQsed
kfapQcff56gOJF224BC+hKb0JHVYVtwZ3mCDc3tIbSTQmiqQT3N2rDdNOvWHHyc8
HYMJBOV3XeAP280RzDv4qNtY1ivf3g3KsrPlRzBvCF8AkB0hfl6VZSvZKRyxB7dd
WhS1c+xEZKN2d1rvszBfrZ/X36n6gvdhjZiUcWoZt0zd5AviTxFcNppJ1mVk1+Us
XwgyBLQmtozOkc1c06T8LS/30jEBQJl2DcTW8ecGwv7CDSUln3nFItJGcnvqDOhm
nKGqN35LoUVaRp/8H58QgJcrvH//27Zbp+KXPCyMZMHtUfB4j74dkTzmVil4Ef5+
a8et/GyTqLb+Zz+uKX1xfV4AN2Hh04nwV/6rwvBz4pNkFFOIxdEtSE1y0TmfkWr1
W2a9iRZozE0R/+uX9gsJSjinIwfx8R2Aw/IIYcpRzjg+/ZJ9t3yAZqxFbhBv9366
Ahlh9mbISJ872tBno2zOyn6VkWpfTl/NeReOJUPLyIlbOqdcLF/Ulsit5bOYnhPn
cgVObhnMzq2wcIIoNng9MRQnSKCtHKAT5T/DRsL5FRqUvDIv7lMUNSw+78egA3Jg
heqNh31muQ5ejDfg+AfTHFnEeF4ccJnDxXRl0ls7sFiD91k01oUXa1E/IwM1bqh5
pYnB2QitPe3fQHJ/YhtOW7gm2YUGs4fe7U3sz/TuNEBkzJ/vvOzsTaxpnB0tnrvX
2zyC4o4mNfDzlahdBTrI8zM8LL4E0aBEi1XIiSgpy8jf2XznX8X/t0zFiWfsijQ1
YNbzVCW2te4sKc4ZZZhgN4zTYLh+qICqlLvyf27mkoNYRvr0o/Gb+2cBlDV+APhB
bwMOfDX5lVwJa+cn5tB6+xMZ2U3fM0jFQjWmx3FMcIDNjCnU5wDLowPrgx9RxA84
LarxWXt24RacINViMlCGMfWICYSobg5M5O8kYPpLHpHAOz629UYOrOLOnQwbrBWy
TggY/zRSXisnLQSf7Fl9wkLQVWlmbWeGSmj0v332sR9BYf4ymgrZp2ykeBHoUjMf
GzpF8mScyhl+xBNUfYPrUxaKQlK3TtWfGqifbDF+tFYAMk9kHevDR9bCKddo+w7g
ZKvMVVtGPrEw1ipcEOyLii5QWLZ6iSUcdW3maxnPOb956iHaflg61gFWwEMJg9aw
O1LYi0kIE2rOKX/ktX81760Sv/lrAIE4y1ZZa2levOmQIpMWdclCsJveEwQ5mmZA
HESIfPesAFLFzqvO7w5QVUStiJQpaP8X3F3QpYKxLMURir4VrRFqNZoRBSw9wySa
ekxFFibXGshDI7vne6cK9cy0VpaZTlTiYHfT97Q0dM9TKWWzdkfo9UIxnHuM+aSm
8kBFfoadD+nrmQP7GXma9MjHnPIf/A0OWZFSs4fM3rBM+4v9nl57WIDjlkFCtdY7
zPUSCHZdJ+fwrkX2PtYRsMY8WtTzO3B7sukpKV7UzGKj8og0xia7WWhlhUC/lcFJ
Pp1oDbuDJzjoXIK6fkzcdmIWj0G6LIbSwUbAUuqybvltJG8JgYusrQsQlRlOs+iK
T163auX/vPQZf9HTgLO10gwe70+6F3znF3Ky576VWqUn6K61c6/UR8SneTOyEb17
29jP2TOMb44PvBManfzEhKU+4MW6PWvpvVhQsyKM57hj0BJO7adst1hzNUaAb39H
ZZB1VdoE/hby0kGxUK0edTWHvGaiLS9s8LfSEP+W/bLtzHN2M1PWoD/rwU+PRx4A
P3jWTNI9qhvHYCQua3DhIaqkJWb7npmphNq/bUWl+KDjoRl8Mq3CmtH+VRawJQBG
4pIsrVIxut5JursxKqh3C85cSZ8Wu6TgKXudorlWKoM/ZjiiiRkBZQwKvbsUABF9
II6foC4JS+77SHjEOQpzA/67ENZHtPNVCVp/OL/FbHrtQqNnUYc5LFoHRRKvSYnz
whh1EBNYM0hnzI0Q+c1vJtC19nBdvIUCCw40+5vGRutGFp+Rh4lgWN+lS0jewat5
ntoikibyNONgCtvK6nmj1m56uJNx9Q+3a9TaM5MLS3FpMNfXTWjPSEuOyyy8u9Go
4xt39OvqdmoxXvRDfx0XGXJ/PTjiQjCMJcdLZQV1umiBA6EzYBBwbSRaUrdbYRQ7
/S92nno0FCcTYOmyv+VYORZ6RO9bA5/c4PTA4uSypss4fyyMxtzd90TT5vRgZhsk
V2w4dptJ+k8dANf6CDzVOLUpXx5maWpynuAR6Eooah+Is12yLxrZTA1qweOrzKpP
tc9i4Ni7bW2+X2hEp1RwhcEH0+6f3ROu13CC9UVnp9p9I1dJKPKEDqpMNSVmHUEN
K1Qq+tfinDhZwOaT4hcfRZojJ/+3PAgVqKyArAUL+gcGdK/P7aRHKsLIC/qqVh87
JKwH27yqbg9VGDu1OMqPJFhh58SYaqw1xAY+xP/u6aIxTFr8uKTx2e2QPzSpOxMH
KD+75EViWm9u3gS7C7ZtZSRkmZQVScGvSfUk8duGKVZgchiTGkL+8XvgWV/blG/7
UHvodmDWDRkuiO93TJvYvG1FgBDanRfX/nsmtt8oX+ZN329ld8gx4g2Wc7rWwGQG
FEmXhDOq6g3an+NHhEiAWlyMpn6qsc3mzdpcrgh32z6zou44M8NL8rIqyOT3Z9wg
w3XYUpkN4O29sN62lopjlrh6aSBc0KULFt2rEyPbnTAFUuJlZiyjNVmLbxt52vEr
mW4BUX9kJty8txBh5yIWw41EjJMa8SOLxkq3LlsQtGv0Go1J2VTNF2KaF/Csez7g
6w0lEEmqY6HapRE6msQOZnPpiqcPko1nuo6tXCZ8k+LVOWja4AaOqeuzkEzZvNLB
8hkJOH7/zrnXCpSVRBUIvUupvcay+VSURsMHxOzEDMgW+DPkMr2ELcUOgUCsCNOb
e4YTE0PTg7hiQ9HNvL2cUKp209TDD7CqvTXsjbtiRrOqI4ZCKtX42U1slwqwYYSD
kSijw/pOxnA4DbJZ+2Bcwcda3LUZiR0fiSWPLdRS7s7I+UzaFE8UeqXNkrtlo3ap
h/ogRYtv3r7cjl5vOswD5rfFyWBqYAa0xWS2pWAiEFCPUdw51pH74bxq0BJnEKtW
aiiTgp0mnwCFPpZ2DyasprCbPjL8RC3Ld2hi4dNkEWW8MfJO7UkASF5etj0z7ZuP
D4ECnGTDMBgFayRSd7hqGPbRcczCWLn0DylOzcnYwTpsJirZrM/H2CsyQnZdl8rM
Kf2uw2JkboT0EP+77tjwzODyx1Hz/Q7phzMMk84GiSy4BYoH73aU3wHYEQEvxXsE
i1lDaocSgZnSK/PAq/8XjXo+O/aSVQoFKJBpKBjHYSpmC0s+SSaVTHXZQy1zN/Xu
FA06iYCqvGtqgfozQxRCpHnaTrcP8wLqElC7synVQh4EYeIiuiDWrKTVKmJvfSPM
uFpn9tSsHv+kWyV22+PZhOpoOLuKW3CjCAJnu1IF4UNI5gvH+nn2H2Pg1GrV0Zro
6ug76ceRoUovzqHDad+nByTV0XD9rg8wI9kP7YbjA3LdPZB7jwNr7GXwvl2olKMp
urYDbaqlU/BeC7T3u2oPtbs44Vvve6RK1Ljdm70ZJJFAfxXiPGQ44FBHlHwDsK6i
DB/kygOc8PRhcMizKcyZwXO2MmSkonBn+y0kzYSrsGwOpYWw/FnW2Z+BOVgFCRrr
q233vZiZfPlTmdsnXtYcVjMj8GKkS4UXZknjAWt3bwHjFUnZSwd4pcYYoGkvaFjg
6OgdcYPrQAjN8FlYLWvdaxVx2hxx1/lMk2bH7uQd27PlDV44Tgrp/yR7ufNlBOLw
Ur/ZC5bwSvteOurU71Cax93Xnls6IGTs4v0j2E1JJBKMReeMLTr/aJC/t1nVhyDB
ivcMaphYFSf1qTCCRJu+4y/IxfXQlUqea7AHWuxJq9jKdBCHJH2kkZ2sdSq0Dz5X
pl9FDWklBeyEt+qLAwl+Z7cIP+OcmPCWmFy+bIs7rEJKO9vpIvg+ROQl04/HvewF
w97X2+Lr+e9WpwJde2xRVvRZaU5vXeg+CCR+A/H9fDKCCNUjinfsIwrqTL+KNW/1
DpQI9g4FLIOH8iZHllQtg1Q6io1V3sYijMyGP7jp7cs1E+Z4PAqGyH9Fi4e2J6S/
gj+k4/D+Ow3Mc8nAy9CJKIi/W683uQvrU3u2EJAgqsBTPTYXVilpdSM2qfSiHvVk
wTJoUlQMAU9Z4rXDXI3Nzk1y11naXPddcfIzVikM83rAbYspLswCd9jjljN28LPk
kP1Yl2FYsq5TlecgHZ807mP6fAjJbO1faYLBnYlCZZrl04/o7e/2bZ9h9yIenI6i
J/+rA1v/olsXauUgcmtFxA0jZXEPw814t/LaWIi1ruv+PW42hjg9V7H27TeODcbQ
VyIXcflm1NbRKkm6QEIT1FwpU/mk/ptP5xY9gwdfs9qdP33vWofuLWmlX1Ud6ShJ
0pITREbGNnbCQiLrPlwzQgieyPIO6DgMJY7qpWFSKe53WJehVLNHTfQhPjUWlazP
Kkog4KeZxz/ttspgS329eAXWpxWdmju2OnlJCzjmMaxSDNjUfxJnuiUtrLePgUrf
Nzz3RXKUV8+tNFGwubCM21fbpO5BRIdkSbWdqj2Mly7GT0Tc9tYli0JtDsZTz1F5
NzYetZkSkU6gIPwxbY2UPP2pr4O+sGtYHmHy5JCwSfURx/iepKQ2vkvI6fu8Gj9o
oMenCqmE35ciXk/+lUq4EvxZZ9KSB1GqzUb/6TTcXCuGvXGR3XHEKnNwmgLoIyLM
hA+JYbXDpPN/p9TQSIR3CCNjHj0fVBHVgvNJ9xdjq6u05Cg+6V0DaLyKfRmCpaGS
ZUdnDod7A/XGT/NbIY2q0fP2GqnDpij2XrAyaSbHAfsBdryEzQlif9guRxdf2+xF
vjj8Udulj3sOTdBoXncEUPGGL7ITxCBnhp2P5ABwy9ovirPRoqYk/YyKiK96o3kI
ntvAkLKwOZz+HOT84BTo/lXSuTnmk9jbym57pftjegB7NMJ1QuuH3CBc82oTa0IF
L+ltklTJMqkNcwDbxCwdUhmoVKrvmykqL55u/z4IMygBICUkZhd1P9+YBJ0hYAs0
4CuNxnf5aPDot84lD8Hw+0KwekzTcvJeixnf1I9my7zcnBisLvWmrgUC6zX3S7UP
8SxN7cTFJxkEQYvPV0zwc+REnOdwsA3x/5DJCVfpl+epv06vMmUl+FkEB18mCHkT
IDy7JVYTtrUcyllHrceerAIdZC0CqX4J4mDHQzSWkVeYoyrqu2mMBp3A/SgBQ6wg
LWyu05a1rH22uNsuMbTYnBdYJ76j7XwARMOljuUl8E2XgPkMDv91Hf5v7bqI0z+t
5xAyu+OEQNkcUb2IsctLrZWJFSpbxqtIsimGfn5dJDJ5jxsRW66F98FF0R7t2e1g
Z4DyaL7Drb9yP/EBV0RclwavEOcneO8k6SD22YGwODBSJups6yjE26ayu1amKCM+
z0sWr/lfhAale1IeeSnYZwXxThSL1941odA7Ra5fSwWS+ZmNsbFS/4/MphEG6bSs
6L1XltOqJhHtvC6lfQq9IKj2PfRXjakBpzvopTOAtR1VwsIMR98TqZyyXzh6/n9M
Ys4fRk48Xc9Fq9vC9MbTtPt/Z365iFzYp0g0/cGlDE4=
`protect END_PROTECTED
