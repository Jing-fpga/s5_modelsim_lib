`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1GUPb5xGlniJ4//SLymf/eKTHEsUZe+4fZcyIXhsPBbQFnMINovEHGemEkhMdpoD
ctKwhg9Sy3VgpJZWbZZFjbYPDvNTP2mQc8fdwK//hVk0BKgulf5mIkBJFxXGXJfg
W4E6wT7Dg27q5cL1tOAneuGofZ97qmJhpSZlaTB5HT+do7hWaSwMP5InupnzxizN
Nur2/LE5SB3tZHKHYhQ8wFgh6oMM40YnGThjraOSnDzm9GJaZFhteIBEksM347To
SXUvs3j37Do7DwuILNXk8btWJE8wGrilUgdkTYU28Hu03QH94+LcZfZnvFgs4T3K
nz8V3WuE9rmg7clOWQZ+QvZuiG4EB6sAJgcNw1HuLnHbtsnQfrEMva2OQjd/XYKm
TskPLkTlZlgxzL3kx9J7jlMMx56OrNdQvons2/B1Qjl8gWKw9sE+UW3AGJCcLZpJ
rhoTveKiDgn8D5QOZkEej2QpjDssMbBSzeMi80+h9K2IKxefD0JsgWVGaB445M34
Ic5TA0DUNODEJSFbTb0LJhe0soMFmm18rnXWh35TSoc5aXQy9+tBIsQwgVk11vdT
Jn7/DDFTq6qG/N3BCxkekfqockmJs8TcCZvgrfDMTq8/l0V+LUIsJxEYgFE9bgWt
l8yTh9aC/kvOg3TqmFs7K6Uo95rw8Du2uXJnh1lIye7PZvOohTe/SiG9EM53YgXo
DcAwzOQcUf6nYL/3WCnvm1suMRdCKwycORJ1rcxUysnEat4k/5m6YY9sK6ELp5tn
hrm+8t8sXwfRXa0wTnh7g8y9uD2ufNI4FoR/DPyaQO1USKjd1JBFAVRbRiFf45hY
3X5KN5bD2wvws63kax4lktWQBEPAgXXyOepwaIekqGQL196aZoftJMT20HlIS1yQ
Pa3wtih+b8YxhWpnX1aFGEEbiYmAUfXa+xBpSAd7JXoZT2/0OhgoaU300NtNZEPG
Mb5lV2dta+wruJ7VCadvh0mZ/Y85tprW/HCU/I3JMHNp+m9h1Wzbkw2Yes8Fo7YZ
/TEstZNjjXDstRlUZ8H1V+HOV/3dkiOPdjdC4CT7Vf+Z/cRHYsMmnbc3fk1Ff5aa
x4wroqgoynOWYNlWkLYJbBNBY1tgisgjZA6QhS6tRbKOTW14se3pJopG/haHzsfl
JNMqm5xOTVLBtzBocnMswE1zs5D7n6iCKHQrVuD2K04Fk5JqWKXmD8uE3gwOIZv5
iH8xHfKWE+j5b1JtVDa4nsY4KRqXHnJodBNlL+xYGpD+hworVrp4wMtIi//IR367
Sr9tDI+/dQVAWL4IHftVQGNFe/fiICaQiqYHU+v2USFgK11aYuj1JZyrLPrYeYHr
vmUiHjASngl1Xpu1fQsqqw==
`protect END_PROTECTED
