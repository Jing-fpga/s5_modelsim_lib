`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wVzs1qMY5Ur4CBQZHYX7JnN8/661mfJbyG2VDOQhV0bPAie3YMJRgkJWTOPihfBp
Izky+GxdronG3U/2WrzUjLwvE94g+yZpqZgH2dMv52uToFW6P7gsz/kesjlgRN+8
y/03644riyCTiDBfVmjUOtm4NUnufJcjeSYEz2oB2g/Qy4eWJgH9aVUHkZopkQCf
lyiaizV8aODa7QRAXZm3WQ8ITq++WqXltmnPKaEg0W5Xludv2EdmC9LctpcNJ4dz
xzLwzT7FlmHGnaLHvfPZQgBHAjO9mwHCFY3OpIheZJgVv69lLwVMoh94S4zhNZ+C
H6L79RzWGVaO1ptmrWhSGaki5zWsN7Zv3xpOXuNVxVu5kse3+167ehKUGoNLtpxA
WPuHjPxAkDsYnAccAiqRF+lT+OxJ2jWiL2F2Cya3l/PzMUSM6UgS46PHZa/mk+Qf
jX/llRHsTlzuBdCp08aeyCkQsH4KQLVcOCFa3Q4HYhNdy4LDyva5Dv+eB/afRc/l
ZLQkYE3fNGDia9yUApY7bD3RC2ltvXP2jt6yh8pCqmUfccFmsw/6CO+qE8bm3UaR
LwYWwmhGvn78gwnjeILpmRni5ywbL06TEU0HxiDvIac7RvOlBQ32Tx758+rt0NuO
Eb3dvWK6POA1OFMvZ6rkdi/vLuVZl0X1i3RxNafx9NL+r1eSSJUdEeXUL6X6WyfB
aFIDDNWHlAuTSjmzUb/5KrnnBFCJ6Idc56VeKDTFOWNmnFWeVLkPbeu0h3Bo+/Eb
s5v2+vTOE+oYt7us+vXImwPjQ5hYzt3y1qGB9JoxZFbJWIPX+QKXtoNgINFC8TbF
4b2wbkFYrZ4tOSDkaalfgxJP6+jKytUGo5JBxjRTUfDMNeHDKmXf1/q8xtSZbXlq
h3IOSftVB1wDkFEoZEq6lW0JHkFScu4ndcLLCmmojVlqN68r+SdmmTb28whXL8B6
UBDAh1yu+nTyOUogSC/PQHoLhN9ygcD5EO8FYgkh/aRYTYhvM1AUxuGXNA1y7B5i
/HiHlaMjqmghGsbrhbRV7t05BPuUX6TtBMj9UUyF6xh5WEJYH52hSK+G1ZfrrtQ0
rwJyptH0IJijX5VG7Q7fRD874oDySWtU0KFm8gyOiLc1MTvfvewkGQ6whqfiYx/T
TvXyXvYLlIwTwJcq0msppUYkERv3ziGnXGzr24dQWaqWamZeLc1LC88vPtW0UeVP
5VKoxB36e6u8Qn+UC1GH6BFqYs0wQlSoTm7nZqz9cB59S/CjolPqOcp3gm9UnUcj
dp5zL5TEvITavxM367TpUzmZqZi4+EVW9vpa58uVTaAU1AM6h0+k6njLf+pmF3eR
NM+NDUIb2JfvRR1+OIaTHMl2LgTFQ0N/HP+WPlNVqTz+8TkiKxmO0ZjE0un/KfYS
1fwOt8NfPRKbO20RdRckKacpVi4h+7mwDZt968GtwhcEH4NsdpwAQwBoSXkMFYf/
ksop4jQQytYfLUobl6boTs3uYtfkZJ8YwTxis5RANqMDZ3CUAxKis179KTK7lUi4
sghEVnh6ESclqs1/D1P7SjZmRIy39+sdz2NUnY9J5IrKaxZvcTL2OH4NAdHc/yWw
YyRde3+QZIf6mBy0LLQ+Idbs6EddezE0Ozzroz9qnN/fenKfjDsK4SkzDoHRhT7x
2nvqNRzRHweIDsYEJyISku3/kk2XogqlChyQZDE2IIIfpIaQ3EA3drbfnkXeSywq
Cmb5cWPJSdGTa3eeSPtqbctyq8oKtRlFhNwy7QjLF4j55eHWgIlpWPy+TS70Ga1z
7AVTWe1MHuJX0/vb2Sd9vGHi8aVI+EwN+Un+QJ55qN2KDBFMF2kdbr8hn5Tbzuej
H5ZhjNOcrtEN2pM93smzGDCR/PFq6sU+11XCiEJF974Zk3kmLqgQS1Ve/p3VHyWK
w6jYNCJ5s5AZ23xmhM9tD+3rKf+7eq8njUM6FIcaxI7qcipDvLrN1JJpUvdgs3eD
/iXzfbkFVbgbSgUCrbwiCV+TEXqXRFuoHyZSL94RmYCAwAhjkOkiFE8N9FX0/YqW
RV11KQa4uVo8ilI13DHXzrt7X85Fpnk/JP8Gko8VpRURneTl+yAcxdPyq8hLQP3a
6a7GISH+x9fBNfz47BSjZnL0eOP3NNfItrXvE4BdSYfIEYGsgodSGM9LYkdrrvY0
Nah2nmA6TitATKl5J8WEchSqNK8lO9WhtXOg30Fq/JdQwQ/uDt2fPsnhlD+qetpi
k2PzhrDoi2W4LAtVHEkAGWfu5zDaFQt6nqcjtasJLvPtt8vjxeY4TJPvqMHJSECB
IgeUst/yMDbmy7h7gTSQzeuKGL5Fa3v9EsLM06DZjARL44GjfiDnwtHRLBnVa855
Jmj1IJ42uBA6dRptJ+PHfL+coSRHO9R3jIuBegDdqQ7ZjSVorDIA5X8Sp5wlOSIP
gwHuh9qdu0vt6CU7xJObs/TSKOMKNebbxt58PMlk9WfUtAaYL1Glaoep5NTSVhet
QSEDCibSDgU2fILMi9PPXDvBVtmOXJWS++0LxutNuB9mNaF3SUOpAH8HqdSyERF+
ClKbM3y0jCXcStkkSmHiRT3fVMPETaWQXMVWm/kYkRM4wGwst9HV1AmTxvJw96vD
HIMUWK2SiJT/ZG2FLG9WrXEPkhNRa5sQrh1abcbRuEa3AemvqA1yvm4XSxXCD2eB
rU+YcyYP2/31ZOhIiOKz6wtpi2SIp5wrKz1l9KdmL2NKs13XBhlJBB8pLKeRYYZR
TUnjgxGdw2r51/bjCSsfzSuqaJhL3QACVJXSZ7w2qwiOGRqNXWvOQhokTrYZjcol
Xc4U7QP6F8KTHvTEYo8UMPZq81YLoy3RwU/NiF+E41o9/8BDfuzokD3sBfetOftv
lMtpJs/2+crdLCuhxsgvpK320699EcjHJor3akKo7fXz8iBY4fRAnGtOqAl5rEnk
bngC4bjzyvXFnZ7uQmMdI91IstlROFoh8e+veExX51L7NFDbo1tUUWV7SSJtWAVb
rJ8fhcie2mrwcugaJXT8lDgUrZdPQ/ARb5i9AiirmPppLmwAlSXVp9/xHJ9I4fXJ
1voVyRZhspm1nS8QbUnEGUlHQXqf6j/TMUY1BI2x6r1UukBaZY79/8c/hWdXvyz+
4NpFZosw1jtC/i9iPY6ms9qEl2zeITD8cXyFU1WeETTgcIn59/toTASsq4Mb+/J8
teAk+K1I7Y3FZoAxjPCXtSiwPYhpbqYpE2xtNtoXdCsJPnrcZQWA2CUaCGGR8P9w
BdGGYsRs2/Vn7iF1u334s2b3H76pRQHjJEvZWo53sjt4NCKmtr0CHYxn4C37FNc1
9dp0DY7XWNwGvvmGKGGwDLxZdzBq4hVY0rRK6lldYq+J0tHMZqsjnZUM9VwqI4n8
elw7pCbKpRyb74pMKHf+ZT5eyKodpx94va89i3YSxUhtnVgBtEzDbKBHhDHyDw3S
CEwpqhA0HIixS16y9OF7yQ28YCNZ7uXtovM/5FekRvJW6yWri/8FGY9n819+Qaz1
DLHpGS4FOmQPf5Jr/ezdRU5x0VUoWGL5Ij9wGn+3g44kofnYJcf/gy14lXxn9tcV
fqztAitamqGhC75UHLAicfAZVQT6jSoBVu+9dUFN5tqIn0GdsETGPIFFUqXvOIHi
aHy4+Ibw5b9M13RzTSqVeYsb2CYbPEw+6w65Ya1Q2Dqc0RAmDYvxTNOA6XbAR0aW
`protect END_PROTECTED
