`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9FRtacCrR1VYK7frarVgvrzdml7+k/R4yg0Krt6by0TjSHtaxwH7CcifQfwWDhME
MApYM7sDmuahqo+FukWmzB+odAUVRopt0BlS2WvmYIXFBfifIK8USAOwjvBlYIDN
QXuT+Qe/8NCTBoTjxblr+N5cXj4ssIhTTAva9BtnmlCISAkSZauWVXezlkWvCwdI
HKQeh+W03CzAWJlTOieJLR+NGYqWSx+byX85Mhlx3EoHVefk/I7vrn2weRVEwcZC
2bs+bn4r6JTkIY6bbIDOY6HQ/BztcZxmj0fXqOVmtM/gq+w0s0QUqcwvH2OXZR3Q
fNaOyQ8u6c6XJuOJxPeHUxQzZh1ZNNJ/uHs6mV9hKsw=
`protect END_PROTECTED
