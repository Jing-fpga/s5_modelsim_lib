`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RYbfuXaP/UQSqHt0qtHvdTqjDQ+QGn/AL3xlLvyviSfChEGH8mP4OgyUvcT1P+54
x0VCwsbt6U85fg/BGUk3zETrQlDfmNad4X914k7ye9iNGM2DSoNqItM6jEO8cgaY
A3/BAh2pz/PQEb1D528FpFIrUIIXukcAUedUxg/s3SYZlpPlk2uKLAv4DOVwxUA9
B4Qisob1BQo8YlnR8UkRHWKjPV3WrI29k00eKKi7XGBH5R6zk0thxyEznsM7qncb
yRzdqFzmjDmLO4ltN0wbTWmkHspknEsgn/421jdHAsr16zSa2jHfpD4Dp7wzShYX
DJzTNBihsVzk1FhYNDGhqMVde7kyfC5q30GsYNWQRrkCSC9l1lpYT7znYRm1x0dQ
ZO0DmhXq7tq2aZDsvgRk5Qnp3wsllYblUM6WIwxu3uho0hbVsfRpXnzgSjusrT+8
B+1HBUvLDmXikoPJWodu/pluF5sFa5BUviYE5bdnFjkD9HE5s4zyduBQAB8ziI5Q
mdxNn6iQeRRqeGjZD4S891NG7vZ4EeQkAneDTL56/b7oPw32Dtr89DFGPywlzsWb
V8unLAhW0ZTvnnR4nVXNyrpYaef6/1uo9S9lFdfjaX7GCJIj/B1OEB4UST6VY3uu
O83BLmEC9s265VYFH8tm9cg5TZ+fBkpJFw6dk6XqUHNwxUJ+nOlHjTrhQGJzge8i
8q6chQRs1f2qelwRoyysdcKngtMLAc9L27pTaIyUrubfHVEawp/1DdYuSqu7JbwN
ioA0MAM/TRQKy0MVx0oLr85co/iONFJ1L+zJu0UwM4B3+0nCpiKSR1p1Zjhe4WAg
87nQ3PsP2J2PqAypAykmJe+qpT33xYlwYnKkikbItaFm58cOjGqmX/XCMtQiMuC7
ppTAtNv7G5GrJ0v67RWGzK2VjxpxgcCCSHEXyV1em06+Ulq6cs1wXrFTZrXoBSO1
ILgWVor20MGZ+eUmziT+D7YyCU6A+9kqSdepMSwamAo3jW1jMyU2/7Uvqvu2wDV/
rqfrZOD4TfL5n5ZlpsgdA7LeZ7tFCkrw9cFD2K3/rtZ7LGwyYXePuxugxfBNFroW
ZA6fpR6/7IzJbmJtTTzU1RhjaUM0/eBA7DgR9qiel6RgJsGDDkJntkecKxpU3e9H
YwvxhknCAdp6RCt1viYljNOqUpFC/mTCq7k2SsFZL+FjAQz9kZsuwyd0rriUV0w3
SHtqpxLbYnZJlP4y9tQwohTjLKIDDwPaHEW31aQmiNqL/zG96YAt6JkLnHRigpFT
KYKbtjBuHeqYUbrv8lPDEkAEN1kTamcHWc5VjH0M6ytH2Z/ILXCwMqiRLTO3En89
z2QL6iPfzPzIhkhCzmkLdExKfb1SqxiHOTN8S14eZGrmXAZzvJIUs94Ed+pB3gfS
Kp0yPYs4a1abzIDTwiVgsftkVXGXN+3j2G19rscskBvHpT8RCqECBsEELFbN66co
W1HGKXQQ0MYFOb7tJXhOhg==
`protect END_PROTECTED
