`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BFHX+eK1B+9WUrsTjg1C3YNybjmbl3/PzloNbsmU9bYXiq2y8S5sCgLJGhGKX2eV
/XESz9t46uMPAvDHhcV5jk+35+PKA4r25QCHZymFDqg8tuxB5MGVnSRPCyITresb
LTvMrfQZAXdgNt7WWp0WFz0WaZXKoS8tDTAzXBeMl2CAWhE1ES09iJtA52hDnFfv
2JnV53NKp9FehwA+SE/QHFlD1IRR8GwwKKrwCDAfiQTIVlwe4tJebtyNL1huEzuL
0naVAAA0p4WBgyYva2epeuZxqoORzCx1z9HAfv4uhEbQSOLyDoGoAVwBDQe6m6CW
wWvYoiLtAIgwRDfQFuLsw2nUWW+t2/VVw/tLBhuFVD49nI8+9DIVN7Fb6DzUDnzx
1R6ddc/bhU4bKrQzHxUSde/JrsVZPIYzN62lvQUlmSOahLmOISBBIvewwRrWgyU7
gRSMwAMSls0ZNM1h2FODCx+EBTX242+qg+k6AgxqAOt+d1riHBCp7w4/zdkYgIhn
hA3c6hu5WqgNXO10OXJoKkRdt6/OED2u+SiC/foDI4C936G/KkauuP8xhBAxWeMW
6i8/yJpAnDwn+/SZGQGhgHSOwNk0kcHkPJIa1wmt60wrPIFszHG1h8oKfWp3jSDq
stqepojili3TtPgLOzTA97Hu04nOUJAYtbgQNSg/7MBWlPQZ9tKOJgutKunixQdX
u+MuOet3pDNkv/0UH+L3qfOvDO7gNBjD5xFxQdW+iDLGR85cjQzgmkrUVfo4D6UP
ige+vkZhfnORBtvyrrvndgUV+/U5xb7Kyp7AxPucx1aig0jQxeGAm+ss5rwD5kM2
lcqO5+7BErz4M3Mt420Jw7TqaXeF3s1d/uZnhj/wLVmusY+3pDEUSeT0/BXxjXKJ
gUvKeRG/HT3Bpab+jamlJSME5nFaH3oOgg3PIg1pBD99AVoDPsssUK2u4yDaSGz9
0eJ6T4ok0452AKG61nbDOhCruwu78WXySg86EfJh2Uc3SEkMej1sLqGhVhy3Y+ZF
3Ak/gxDy134gcvjco9ZwN9LB+BRMrF+4r9PdAxJhCCDo1SqAGC03CvCWzX2CBTFO
TEA3aBzWYtSEIxwZMpoo6UxaMgtJvc2fn0dSASDo06ulYXRh2mvz2dv9js7JCPE8
3jKvD8f7/jJx00LWGm/vFAzIwOEYHDGRP1POvDMGacpZNzK2MDGF7gy3YL2E5hpr
DsRRIor6oRpxAUGTylqmAjNzY1NE3/pFMdZIXTdfRdu1LSwq7uJtfn0bS1oxHc05
jHe1hFNnz1V9Khjv8ljFTXDAn/5j7OLh1pcsak/8p9U/jCr5HbgoYsZv/V5o6n5G
FVSyrcqhOKsrwnD7yXQNn74rHZmgZoFpbi/BgNicD0rV8b8NaV7afda+3eWamo0b
dYLEV6BjPC14PXbW8krGOPa9dyHUzKfg74BXZ8XvoNPYZXK68YpwjxGRef7hYh7q
58hJDDr5JDDHfsBq0WNvl5m8z8DEA80NKWbDRj1rIVq5L/xogy+n+2+DyZ1kx1Cl
+TSNZXcpu/e5z1Si0p3Z+ePToWDSknLrHh3toYx1PmDvjTXUyA9QZCuEE+LancVQ
ukyFZn/zoMnHSp2kv7r1ptHgHXLCPcMnlL0wy4Mza+rtrDN1L3lGjp2Fjci9e6TA
V1og5wIMCoUunpbvn8FQjjXTwthmyFuRm7md83KjPcw+PxcdP0TiNSMI9P6ondt2
QzVIvt+DV/1dAMXR3WpwVc4xdYZOmuw41OkdOSkVLLy1UbF24/AAEPQbArFcVDj5
VY+960KvnIqVl3gFLj1l7pmQVLh/Eyt3xeX6ushkfbcL6aPi7HXegPxL+2tEZqZ/
BwYY1IL/EYbfpi0x1PuxTkX5O7t9LkGHcUNl0sGK2qrWl90gNhGZjvG1KoSnXCUD
WWGCe+D39N83meF8FepRrfmQcluVzMqSyRvGA9G2c6Qe9VXdFQ8dvK06EIP5ErrT
w7F7zbtPlYSbPO7VwpFzOA==
`protect END_PROTECTED
