`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kE7Bw98NSg7xSZK0yzba/EGnaWGrL2374YXcrlosOv4Iyu8/H+ZTbZqofyCUSilv
QS7S378MmLOGr6UoNNmmx+MKxC81oUysmf77BplHcoAVMDass06OUcnQ/0fVK303
vgh2oDA8m40iwWno+RzC+sXoW9U5V1Dzc5+9WkNh8gUP+cc5kKBiDro2NQJCDg9N
Ap2/bZ2dQY0AG5tEfbCn0CC1jIOIfEBEg+EsQOYc0wNI0Fh3DpAHZ6UFuWRW6fD7
xijhobSwgnCYw7CgTWLVWQhOX295J05iS/bp8hbhenyv+C/JOUIWQrjNPhdtDYNU
CvqPJ0vr9KNJ2Spsv2mkaTDOINHAtS0U9uh9sinj2JBR7vv4ekFBQsqTvpnwUOfK
REMPBCFe2jttz98H8NTlBUJmHZcId1vWQEH6ax8JI2ARmYPqj74vv1Cp9jm5n1CN
hOV298m+wddQBRHavKaqqLs9UbS9jLiKiYtf7M6pGA5qiOm3XsD02wU1Dsq0j8dV
0yEafBqmS9hrcgFrLSmgTxBTKWznWx3E344kfYydz4NvB3i4MDKAp+vQLUlG0VjW
WJaMUhlaixNJISyzy8/PDPk0+f6bjJyXyUw3tImS+gk5OTK2BXyplhS++V0WgMri
uz1+7tpAzZff+TBwLAuSbtaf5BUJU1fLlTHiCOKMtTQUHjt6VyyWXcuPGgpbTl5h
iEp/ZCeFzSprRGbf0qpMZ3+rUOvNT9MOm+6PvDTX/adKPuh1xchtj+NXsOu6C+t4
l19E1J8S7XNzc2eMAvc/DX3DOqVXmUeJbUxpRSR0gckkDRGTuCKigsRezD9gNE0U
Gv+N9lF6f+sOF1iCvUoenXA28Om8ULLxeP5HoSusgdtln9fYux0kXw6OwdUITMUT
M42Ho/NjI5JJxCyQiryZHpSZa3kZidJxqn58196CZ84MBPBX2v92gXc9NHI9i8BN
p9M+dm9MZHKjv8nC7XkRCbUuNRG00bp3XMxTsrIqFHA=
`protect END_PROTECTED
