`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+WQwXyLvkBGe/+1vKXfp9rFlXiIMQFq9z3jofJvc6BPhkE8RpkpehTZZ/Uc8BYB/
COf7lnCNEAJg3vePifgCNW4sQC/Pfpz3RnI0dya4JOz6/S8L6Oqvjy1IboqUkv/l
LKXp6QBkp8805JAiwQg185mqltJKqFSnutRb2l5NREvdyhpQgkejpQZ5QT3rEowS
V205Weaq2SJ1h8JKuDMSqDZyS5o1y06xtuQSUHDavy6IsJ9DM56V9Q9BeVz4vSBG
k2dAa8n/7mjjy78wu2S/aydHYrAWcLYOcoLDzdRY3k7xjBwmLVCXpSEAzSkj2SbD
Gl87FwpJG0F9xPFMaO3zAbpCpzfcG7XQR7vglU1Prnk3opWjFJpVE2vXETbFr0+V
c2kffCnPfzVpDAYqRguNVjkyXIxGJPPubWpFpF/Ta9YIxh1JwNNArVUIjDi1J8Nk
pxxS2HlvcjKUanKm4XJJL+RQgQHm/TFuJ8jA0bygsDx6XAS7N6wdO+OLOMjnN+AJ
kB8RAXcV3nc3yn3eBccUWEIJbr3vX0Sg/OKLLnLAS2YorERSlQtCLFbe8lu/mRkI
iwCpjXbJx9l1qkSI63CmmT+cH733/0sPVIn2YfsyoIhaAZNXCC2AEsMTIFpR0DTf
uWQCBVYj7l/E6FVIE0apRZ0LnIyJs8RXXlnIsqckBdQ3BItJZzyVWNDJQ+tz6AfZ
xip+v7PjTat495LehMxEE44FLDPJYreWaYwH/i36FT9F19x4+VHUAQJ+81+/u/Kw
EUKkuZaxtnzR9eHt3wd6QiGra4j1nafBqsBW43+UH9oKMHzTVKRVx5F8RgeIeksH
VIsnXJkhT60yG0tm7Hw0v4iQd6z5M6zazoRmQoibMI9HtfJ3NkK8UtHvUOgvkrYt
z1Ra0n4TGZIH7VKcp7FCtMN2I112EdI+9Lrsr74AYxT6xga/lkhzEHH2cwiIl8c2
c58CPw1FTvyYQRXUk7Fm2FFeQYtQ9Z8ulC6VIOA8b8Kp20d5GnKW5Ci/lqaDDzUf
PbMzftc7iQ581Fw/a8pZw+NOPWkzHPGmahX8HVqNHNoSb69U6p0AQrimQ3SmVcE5
bvS2baTZHBlpitYSrdVRcEUOB6UzYrWktWU03vr86m4aW8KI71KFkXM4uMIvXTTR
uiTMc40MqQEkKULltZ7nq1u/VsaP9PaLorqrjF/jz+w4iCqHk/O86zEFEwXLRWZz
TZqcFTcGPLLY4yP2OaQ3YjBiXcG8InSPl2TaL3MWLj0+h97UvtapmkOjyufwXxOw
A3JAmLPJbOWyewtgtXiq3TSQxksDhGDunVvY68moZmAPik6/8vRsYQB1WBEVAjOu
BsdXjlA9h/b9gOe4cCqbgNK4ZEGzbftPPA/6YvoM/lflup2C3Xfol9NJCQ8RquYQ
Uu2dz1zuPeWwqEIkQsIC2+Ep94ab1bSr7v3hyy6alsWhVRi95yFhmFwyxLN+k5O7
6me9gLEaIJAD8ZV7Ue0dI3F5PZW4P2PkAY2oHpbMgEvJYVfcp5y0SCIoiSCiM2bq
ilacGA3ZPvPMYb7wIyUw3WOy44DtOiuagyuCgTthvbxQjnnkI8NuxJJgvuw+Q1UE
dFt5RJ2TyviEYo2rJd3bsBAQgdq4MENdEn1RCq/kcDyEfHbyLcXJ0kC7rYSNnZPb
B2VojSeSedt69Lgu7j+jDV/pLPOWszuGDf5iQnkMvlsHZ+o95UEs7rnY2fzj/olc
0H37XsY/BpzOT1Xe5KTN5GBUH2SliXDcdLEiVp5yIbrK+pPUrmtTCx7Teo2/zMn8
xJf5d0BYQxQb6pbLo7an6E+qxS36e0GL9eZroZxpcBaGj6+EWpkQFw56EYs6U5jC
B+OFpu7JKK+PDyOsChYNWra7mGv4qqUN/r8DM9tkdd8=
`protect END_PROTECTED
