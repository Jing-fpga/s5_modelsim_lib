`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ilAZYhbQMLsbqRYyINHBgEQXjKAJ8EP0VSAtFNb+BPd/Gj4ziRZDVsVjfoQH3UWz
4ybpebeWCklkoANBrhXauFjSTDK/04UgCXlZHT6/z9vOh2vuKZlmZVYtgpwogD99
QsuYpj2ERDXDNTI3ZJbm3jRkF5w4BUZLFOK4ka1V+MsMVZ09IydL+tAsvWtIdFFT
6aA8cpyNWKVtLmAdyoUjXO+xA08AOJboCYITj6ulf/KYg9Vid7zm86LHof9b6zJQ
l/7ZjHJdJm7Wfi9tyu7WYwnqNqBicLJcZhooYmhuh7yAsRLfKedI2bF29y6zNMPK
mf3fZTIoTvm/FWwAPb9FZ2jnZPxa97BkGsgMxtJmEnUWz2r8Nj0nB9e6v5NzY30c
imRHOCPLk/Op6Xa7U/TU13Zd/NwM0r1G5TOGJxD3fp98bDir854AKNxC30xC5ywq
lKsJyRENcz5Cl3+F4ORPcxIMMmBdnFENtgPDT0V5O4LHBoaKks8K8u408jNIbnkA
QEN+ks5Q5keH+a+ik1KRbbbJb3jF1OB7GS/tLFhxklHptt/ayAyBaKHNUYj+AKIs
WP6h7Skzji4K+SHdJ4K0bg96hfTkJ7hIacwO/8yLMOPPVvUuHmPB/7OjhgyuCcGz
Lo/cM2SXuYzvUfhOEQezL0h3yO69EMocQaJh6139LsJEmWHfDvW2l4A3sfCYdCY1
S/Fz5D1KgYX34q8Zy18h8EFt1ukCxg2IM5n1ozzvK6QxcFsMu/aazhC583E0HA4n
UN7k1+RhscCLD7B6+joeYgjqFVDIsCkunVxPqhhxlFzjXBhIL5mZVKvb/dWhlaba
5S/+7HRO9WI/ezg/S6uXc0J8oLE6ANmMRmKrSG4A8NZSJC7li8KYrbLgQxerIVeQ
C9fT1QufDkz8k/u0uPsp+3Zr0DWOGkKUFDEnniSFqBjiKiAmpWCcfUCHppjmyNw5
pS0dYNCxZzBPRBj3ktF1hInap/YRFVQ66LEoevstArH9pp8H6rst3NG77lwX1yKm
hk2ol9BH+7AL3LL/9GEUeAZaXid1/5dm6gB8xCiFUbxvzb8wX7ldmrXfof4+GelW
ZVo3IEYqEXslPi6N9kfG1kPank9VX3oErmFeW8aZQJzbptzKNi/3PAC5QtauiqvR
CF+zjeVrrha1mb7xA4cuWMea1S3HE+49jszWtehfOWsybt8l7mFicjUE/92wBAOd
9/KLjT7XWZZ0iTOZPwjd1fxOVb5zQreH6LfMXeiGKeNq0QpFLTtMoUogu0b3/7V1
oL+dDwbjhMw2J9QwJ6DuLi9J4hzc9dAc9ib8kQ7cCUmleDrV//RBWqo5HOKmnX/s
7bnHmITmLGSGwKvXTr/hcFUdNpl0CzUVqrEeG817dQvD2rASs9VrHQrMJ/PONag8
XYg95e84CoK0SDLdeJjPCRq+ZwTcJpJxuconJ/J3m8giLSuzgl4M03enHUN2op7o
Q8I+K2z2vtnpu4G8OrwyQ1kgfl5Q6RPFRa1R4OkxLV4nHdrK2wkkGbOWfM1I8Qpd
H4Nghi8rlyp7Ga6i3pb5oZiYEmZCmE3SuK/1MrI6NMJnQvHzDowmQVIT+NKn5AOU
o2qbCYBLTENgLa48TIgxWvHsHJpAMqQCvPuzHx8YmWkQbs0V6nEaOHWF0awLey7K
mewWKvN34mE3MIK2qdiLZIK9/gXU3ITSj+QrA2sR4ia8PrxHWpdlYqgcj8FuwRc3
CFqLZcKeL0JTHBJ/Pq0mHVpWYSh1mAJETqBkioQiBa77sbmlk+y7p9BjiHpyjbE7
9J/PKnLmdvfOiPYAvtd3KgHR4xDB0jNQF3I80PTA2qoiEc4mPDoZg0r3H5oC2h+2
bHZJoorm4vmMOvow7EqgQmydywWe6gSpaepePpY2vbOP6MmUV/eXmS76AfbLVntG
ptAAaDPbLm4ttXpl5gE0mdXoQQWMkCH4rtX7404d2qTXhLR7kzKZCWl+Ymh92PNL
FgAYURAZJjR+jqVt7yiSV6Ufk1+Q5JF8bOBRsrBS7fLl2N4zdYU8hAeKuEDNwsYf
pxoDnwC0Y8Zpay1OMMgwktyxofgxZSAQciFFTfje6PMnjFKkHym7xJgpJHpi7bRs
Z4VJVRst2hf7Yvudbb6kH9+Xurt2SS2bNUiH2xdHQAXIyOtTMbCqhBeGY3J+fptJ
2vReDrNHKgFEXEPexY0pK057n2Dt7y5GfaDsfHb4zYaO8T3PXRdOhghnjA/p/nYG
eeXZPowrV9eQyOqzJNcGO/jhvmcNIkdYksSBixdG3MA=
`protect END_PROTECTED
