`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9mgB31+Id8rtrVnNDtpMkYRX1gzq8DO2ScGA4Kbmcj+Tl3sj2iGHwuOOQ5cpiH0v
VJg7yeI3L1ypHobksGfCg5TV9fuI1dduo2AKO5/5ulq+GtUaBHkP4Psv20gEtI8o
541T8YAJSJhD7AsNYBtbjpDzWn5sZhE1jcoetqw7uZbnp8xMZxyEuzLEbP2gpukd
eN+QoEEnKefJz2ytecHhdlMfPp1DwDh8HkWjA+ojwo52No15my3B9gWsl3B+dLGG
tRsBIXlJjTVFK9lhrYlPPSxs0tldfQvsK3erT3KD9PQkjeYEaRr5O2mumWuEd+fd
Qp8A3SD3NkzGSmicwHjZQUTTv5ylY9hU23VtwRIAD4h/u9vbyyAiI51VD3LGNK/t
5xQnMwF8LuPmoooudDmbRvxzhPuHRHUClM7tLBtIO56btFADE0+8G99AKB1OJnWE
fM7Wuk3xdkgwHMgVXFVUc5pc/GgPf58QruK2lSpqWLWwxbDDofg3FzP/YmpWceOu
1V+upAV6YU04deYFBBgnrPiPT+DEFZPIV7XPZLFrJfdjL3QS+0q+WdnCl7Hn2X14
6ThFZVWUqz4652EJEFyMZi07mes+z419OhMgdKbQ6ZJh6O5gNm1oah4mvwXO2xiz
9Go3qhiE2gWU91Ch2UAtcaA3WbAFP2wm0H6NiQFx8HY=
`protect END_PROTECTED
