`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I6QJGPpqjwpdrSttmIzm76GbF/3eaTpYRPr1jPnPyyk8iI8q/aPSSJyV+N13U2sS
lY+B+8rwnqZLSdI9z5iZbs7evWscUg/EwBCw0L+XBJVAjhAkmBfWpw72uObL5SZ4
GJ8MF7sledpuAK9ig/f+0ZUtK6aQzOKSO6ccuV6C4z0qUEzAUlPblyf7ixmXUeox
Acp+RoHb7RIPE7+LkDMuwmVYI1BTDV0k2inPDMDpPmvJWy9YgrBzT9NbVTWycOue
fNIM6ND7KJ+gOIX0xIjFRCnqa+tHjXuPLU/i0jUUoa0PJnGv3OLhn4BNDNmAcgDd
22WyCHu16FPFYboKHgY7Nd0Zz7q15Ln4qizmkiok3yuYNnJx9vBLAdR6EDWTjnt5
1a0jog/uxBJGeNz8RbQ2Rn+1U4NjsX5dzxrpeAtLsdRmUp/ZO1ZvN1iKKodmGiLZ
4/0quZgldUTje14C3xiBya8UWxvzosBUq5LIpTF+d7RgEcS5QHmiGqyN9mj2i/IN
huwKuOM7Ag/xtwC86ipMid3QnGFSov+1CL4AV+SomJ77jloSimVQGvh7sLWujvGm
ADts7uiXHDupeIyRcRVeGOBC/LxUOt+FLjd+bENsl9OncvtLyuVd8JGbGKXkCeD0
BdKHFOj+PMFGMusZwi2Tv4BOsZaAASVMf/eajQVVuvg8w4l0Osg82dJJG4O332Tf
WpwG05hX62ar7NJ7vlkopzyi+4KXTUARqMeCM7oUBwwwt5LsFokDkctZ8D2CXub5
BYsCDBPhVYSHkMYlxZPqqHxXH7iH73k8/8+70CWIrJcUFYs1CCZJSjt2yTBfLol0
6hnOvtT+H3QOXU37rdaLpA==
`protect END_PROTECTED
