`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OkGaeWkQE6IWIfa3tLYXL1yrN0q4bBC/+IHPYrXw15r98QFyYFVtokAf74g4PZ2W
Ce/DxFUoSCw9EOIYodxrFoHe6jOQwCscXbIdC+RiSUGwnQ4i34draoC/UAt64e6d
1lcfeg1a0y6hsPxWZRX/uwet6eerjQKLx7e1UdbDMAL/0T3BsIgGPVm1Ff0B/SnL
n8/2PycYkbFGjv8ZcCtqIB5Ms9XZKgSj+Z0wv+av0pdpm9GOWRE5qn5AWxRetgiS
exs8T4J0fVxbalTYC+NvAjO3M5uCDjRldRigyIa5jt4Sy79Vy64WgXacsI0psV8f
8GTIq5jwFAnU0+NNyDqrDt926qJPHojvrU9JuKGCrvY6YCg867JL+MperaTdxTM9
BVGgzz+ay4ZRS4c3lGTQLXIa/6npFyrvGEAjuWa6IqJunaJHXtWj5FiIBLfcZO/1
sdUqbV8S1OJQU6jgktg67JjrLip8i/t7gDen7nw389MpgKYky2xTU5VxxLVGozDS
ZfVGBu/UfX+81qdesTsy/sBwYrByWFbDCBkg514QsQBo2OOmaGv7thaCOosXvVHO
lusWgbVLsam6ONf644GEKE6ZqN3UJzbJd8kYJxAeaFSJP7riLwPcSzpTXPFzabCR
Sszymcmwxtek2wqryglV0pavHFbYqg5Jwqm7lrXzu6hF/O0jGZeq9S9xq2WCLlc1
WoLJNqoqRab+xMX7LDCORUPGvoD1wRC60om0/vRltcENdaGpThRkYbb2IccPnWKB
2A0FEmoohl4z9Zq2TVLSzlVvHYSm/p5RDaqT5KubKpJHejcJEDlZFj13BVTMplpO
jeFqLvvkW+Dxx15gquYI1oriRMe/RCwUJxNv9cGvqWWQ2wh/ZQJmijdxXq9o61Pm
qZXAOjOtvwU4W5ef93HYpfF6rCTDhVj1uaL9THGTJ+NhmFQVk0DNW7WRY9aaYGos
vfGI+YdNtwdtrge28IkHve2Kje/D2O7m8RVPvx3r0P6xt1DypVgvM+a65VRFkGYu
1e/4hV9lyX5skZgRH38VTBu/tjKqzfVKei3r0QPuYBtxBlHxXQYj0kDx0SwFXy2h
fhy8Qgg68VE85v8CF8v0SRl4F1i3hB+wvyG4lnZQ274HXlH8VXTjJwgBIHfxzKkm
u4FAXinxa98rYOiSYmc4LGcbjW3XQ1Ha1Rxn2+Ai1PrljttaxnvUOELQkqzlhtLf
x/3kuoVzVeL9X95pNNGJju1xjLR1cR6cul4ABJTnf8uW9DQWNfQTQn1rHSssf+dJ
Xj1c8MQjXGVpOzvzWfhDf2vbmJRXpt07ImGbluqIQX2/zzIJQFfnimb13AY9ShIZ
7vlZiQBNsKJxeMKaWBCDXuEpsHZn5/r4XiUMgCGmPwJPojZr7pa+0ezcvyzPMRMH
CP7SiGI1YHT7+dPJayQR6qGflSwzPfpuNisbeNDgKwmSetuSJPR/qp0hiP2eFvdl
/wP/1rpIeQof4RQafYL69rt6Tjy+jxpuMnYg7pIq1EWHmiXYNlbM+lqz+KrsKAeg
XHglF7G3oTeigK1zhI4boiCj47ayC59MI7j7g7Hzj8figyqRv8SuxtruBr21lVxS
y5zhhsKi86p3vqaUW5X33X0X7DzjiZxk/Jnz1pKsLSpmzAv0WEo5DsOluzZhjzyn
`protect END_PROTECTED
