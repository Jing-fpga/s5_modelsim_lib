`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/TA5wGZJ8G7HUTBwOd9StqA4tSX2qAy0ntk4JKnM8kkf495BFitVgHiI502D/RiQ
oHfq2ZFE1KoDa459h3HU+OJkzKk5Km9gwiQUNPI9C/PRdBLr9mRo2Wr8ayiobmbQ
nv44GBaXxSYMiaOsqM9WYfakonR/J38zBtDiX0DioS/ukw9i5lyvVLPYq/sGJPq8
+zv/e5Mi1Z17tgCcU0xwqDYz+THxh18ysX7Ihw4QvMTeUFkKivEl7galdIAnPKgN
s38SgZkoEAp8XGmevVUTiXbHrgYnhBZQvL1RzIO5lB3WFAne4Z1a5bi8+3f6Xa3M
gkPHJelUjFCppx9PzZTAKPBqUQz0eyFb+cfhZGiXwYm3IcfayCc5z+DnrN4sohj9
/nW2KnuugYz4B0y3tLKmwA6GGCrjLQn9/DEh3CDjaem9dxNBJdEdYUWzZLG40u0c
/adHZVWTto6Eg25H7zY/JfmMN9SWMMSIa6zxcmnIPzwt1SVJClk8mUI8kgFZ7fGJ
TwZybAHXhufa0Rjlq+Rp0KRBGmumz+AAb1WE1sWPzifqjgkBQzWSk1v/un0E86mP
AI+dXyTFhV9v40kwQmR3fcFzb8He9BO89OHv0tsNygwNl5GWRrynN6Ka9LmRXo73
3iuIwX8OdoSHPeGXcHKrlBFV7qRb94PnjccvRslnH8BKIqBCRqwR0lQIYMyhO616
mAB+kzFbDlcTkGyVKEP7wyQ/WXh7kwwBKz91AQM0mITE/u4ufG4PxW1Sp9ldYiFX
C1qsIyAdgjC3frr+QhCTBzg6H2VvTmLbGOxJyZL/sTF5spwcWmm6p8YxkL7zMqdE
XiiKu1xmnlFA7TYddmH7mxO5OwsLEelZAvrg/aiOGBjqIzeQZcW9ErvG9cd7NUeU
yf7tEf3TkUo8/GaSOJU5XRdXFgRfX83efSLMgq+8ds63/d1uOnZZYA+Xpq+Qu0Y8
bafjGEB3V48gvIW8koNLYm14DH4a40kITsIJu0ejCrLGgRlJoKP7dRz1WEb6SX/h
vWU+ygfIecriAXWKyntdhsdPiS/HiFd0+JTyCVSrLnz90tSVwV7fAHBc2GLbQWz9
lcP2K6mNfcQPIzZjtjL6IdLlcJYjOvrh+TsUTlDN1lPa4GEOYar//FhdP4jWyX5T
d3Ea+JMrcerCUOo0+ihLGq2bc2z8+uQQ9zGi/FDb+pHPw5Dt/J1MJaFxE+Epe1Pb
BdkMtnz7VOaVE3dgoDIMrrFUpnL1tK+El6ktgpblvhv90BAzkNK1TGNfSdr3BarN
dtNM8yliDw0PvfN7SZHu4EVTegbjhwHc2F0y+aqXWoWTEBI4WakGSYywVGkN5IfY
tORJN7xTmQDMt1m3AkAvsmqOgHcOBPF0Juh6WtE/Q5A=
`protect END_PROTECTED
