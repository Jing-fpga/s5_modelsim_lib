`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pFuCUT5vNxpG6CjQhMYSqVBFuz03emQcnw97lKOrHsMYPUdgOaTY9liGHTtQn6dp
oCdsJDfPi73P9t66grYWy7P71IU/wfh5eYrm8Sw0UQ/TcMy8T97rLactovR8iUdw
ea6guCqb1THFXDOpk6m5JaBIrACXgQuRE9olnQI0pe6H5OG4oCMcbhQvvwSpYTl5
TVqc1cIXPt3H23PmJfHkkzbS31hwbjDHTyhlWzfDwnYPPM9w4nDeBpZWyHV++JEu
f5kJGYcqEenVd0yZ23ybX8cja0JOLtq3Cm7t+LyXYyANz/JNKoW/lJLlKNqX2tKC
CDU7kt/AXnlHk1WAinZKUWeXf+kQ1sJqmyd2RXUMLEEVkOUGBPo4XhQy5yk0ajMB
V7QPif2vdWXfhG9GYF6j3f+FCFPlIJ4hcQrlUhrU3LfPjnWSjRPh+VMUh8LD5Rps
WE3LlbADp/i4CVvHxDkPgFiz4ADkJ0MvVG8SLP27KvXXTDoSVn6jVnxqLQg1Olkj
j81uP3AGcAN57IhQmhOB6m5jBJLP3735rOzMsV0hrU6IZQAawo10zt8UvKC49JDX
lqIIX9z7juKr/6Edcp2mEcE05bJpOSGbQRSEI9H8SmR7LlCZ9HkqCs9ZE1/x8aZV
aELZgkVg6hU3B3feuf5iXexUlpDq1eJSWwkK54M5BGYFYPJDa6zqcadKhvu6e5iL
DomKChuv72FjE4wy6m4iwURXZwPTIK5991f2bAJSWY1/UlTRnmuFlDzWbafhj2Ki
QUacyhvCpNs6I01NiHp88vy1IZqM5j7lwB9QWvKSjE9FyAJ/EcP+uDZVqyhfixI5
o/6+VkDv3bqjsXL4LqvPHU4pXUDD80cWUs33l3bUvFCtUCS7DmVulA4u28n6WAaY
pky1KxU0n+pkmkNov5QfHAyMxatA5jGwjjGli7isJa7z5IBuOupfaSDun08iFPRi
ih+2Zk2MxJME7Cs5Xm4RGKQELxutCXs1lyFAL142Dki8dtTDkOXKzzrra4DLrcDH
uH/w+IRnC/qIBUcWFQ3ZqJZ3ZRwuu/x0wsTDAAFPbeSen1r9Fq+d2bEVsdNsAyNb
rpactBis7nyF0eG2NO40HxoKjYjhoUbNR0JCrw5EwNluHHrylFVEJWwBI8ApbCFA
MpmiL49a5fNPjPTPpeUAGuoKI1+Xox/sNmvFFUbQjIJ1d19xx0o16VJswB6VBkub
OqAl260yiONbJth51JwTvvG2LYqF+tLW0zUPx9w6tURxBuSYu9bPXCOV7XyhOBrL
YExsbTG3wVmtXqyNQ1BfJZBvGxO3sdES/16BgoqTrzzw40T3ljzK4HNfNVvbab41
jxIF0kiVwvJdvDlix58KKyiS3QZwvSBVQUMz3BC/RXiNp7725uKpMMW1VDTJg/4f
rkiShXMBvdAYRoks2//q9IR1BepWK0LKE+Au1a40hwfTjsPcqoq2puW7Y4AQOONc
mfwtD5E8AzdAIgW+DCImJoEz81qW4YpXkFJrmtOIk9cPNH9x3aCmCHBSTj6kuvtL
5e30nooSMkY/+y2tBflzm1iutpEef/ZC1kUwBUmwX7r7SHjobWBOrv+ht1RE2WiK
`protect END_PROTECTED
