`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xd0V4dy2Mcp75LYi594aVXoqbwV4VOYlVHtKkP6XkpHBeUOei1xd8gQW+UkzyMkm
2T/+dsh5vmAccHDKKY1i9Gp5wB4A1SN9DNxtPeB4QmqNyAFSryt1albXzOKzHfLb
kaypbGDC1yaunQO+WSW1rErpHq+zr/hQ+ufszfP1FprIa+f1LpKGLYMqMNmCI731
VkLfcVj8Qfvr+Ja7/koqDb36+/VuRwqRAj0jNTdp4HTQf3CtdvV+Af44Rw9zn1Vs
ftMl4SJN3XiWBWdCdajy9oD7V1JnOBjGkM2pcVwaJ5TG9RpTEyN22D50WUOIlqGU
p+FF1F33ZbKAcS3JWnk9UBq+Um2C0vm88RMQGuLeFBvC0BVgyF5IH+/mAC0CUB/+
rwUMtUYVzjV8bVpNJMhX9yRRCUQvQ/1WZP3iAGsvZFSNRwwpkb1A3kMiPpw5/0Ao
4gjEsH6fzzLICQqsjxNK9ujviFpNQ/Cn4ApT/LVCymBF7hD/D6rxNZhPts2OGJ4J
KWRdGSlluvvySb/P3JBBkL5pUere+RS1CG1f2PC+Fump2AMU8ANJa4q/CaOpQU26
CFPvtsOi5u5keRxqmfZKg9OCc5mWRb2uS3G7ukm9QBo1g0gX3lMnSgx71/Agwk05
GtKNIvqgOIWYKOLEhaaZTxQzwtoVx+h2zf91yBkhcrube0TqArXo00qmzP1IIzxy
26LLUBm+3Z8SeX6IpzHe1u4oTRvUtMP6bg/rOqTCyBaeOJVkTfrkoykeK5q+JyxM
ccKu8pAn4VSuayeCVUXtGkHcOIXi+bbF3UZUPmS2OzF3viej1xqIN6cBZc1VzQvZ
U4131rVXXOni0Ev+jLBNLhyOBJaGk4LO2OvBrag+evZerRFQMpLudIxe1NWiq090
WKErZb0qp6Ly5C0nJWErvM+0f/IVDWaxZQGkEGKJqM6v6J09g/aTQTV0PBLsCnkz
YrLd2SyUB2cNd68zpvBNBLRSv2StudBJ7SJTf7fVrrDCvO3p9mTVzkeMJBT2xKJT
ymBgndNxhwl+YRp23OcYuyns5XbDiPRQHFybfFGk48n1k6D43inQyVAYzewX38Ti
gZ3dgzuAbmYxZuAPW4D3uX9Dt3ZSSeoBfcCWDFaLbep7vyegTQma4cl/8L7dNbY6
dTSchoIJO/GYPcM+1hJYdFNgrY20X1k8sRx0JeLAEY4aBc8lGSCFg09raU0e4K/b
F6+CtnThAaBcHObJC0zjmVz7NiDH74OdfjP/uIjUHZSvmXO1tl020pG40Qs0m02U
1Fkf22xnWXmCtTrlC2iNUtwoiNRbP0dgzRyczsLrRyqtXZ4CPDUM0zcfBYHVFp+y
mGm8CIoJwMYvlteRqlKaoJCGSIQEfUO3qi+o4h1DkGAc9c0Lhmy2xYQFf98tWB65
hIvljGZSbhrfN5TlCMVzJEnEKFcbUFGIaPXfp0Cm+ELvZua0OYdEGZO1LM0OZNC+
SbY41Ro7cPnvnaCEsuHzux1rgmj8cwgBHcVzTzTUgKE9Zg6RswrIzt5DiyuVHl/T
VepJ8Oiw/XOqY+K7GbCHUZoPCbs5BcQ6FizQriRTcvkV71RdE3l3D68p4f0oRw5h
aqmFoLp37m1OpPToilF2zVFzy0Nqs5769kit0KQHitFidY9Hd9aPK2CU02/JdZZY
`protect END_PROTECTED
