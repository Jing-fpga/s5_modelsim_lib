`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WDy6PqoUIJnET5HQFX9hm5Z/SJpN1q1OG+8m/qWPF7cTpulIIh+EcmIH55Ne5Fm9
5rxSp9tCDoRZnU8lJFLTswvAgVTzXvEv1f/+AyNirSNEo68bY+GW8+O+WMh8ojGg
RDyEGvzYwxbivYEoPYSpHR1PQBUwzPIRBUOHN0WO4D0JJeqRp96smrLn4QyPT5Vj
lm4dSNRVpkuw6YUgY6XLxQ1Cwe3MYRqAnePekgH7YbbJHYeXXs2j7qlfLClCB6X+
bz3NsKscF+pQTxBO3+ckdhZ6Z0WQ7f150fc6gilbiqdzyyk3D+ctScUr8vdh2xLK
4IAvrdjTbOcBYsCZc0N6zI8rl+Vh6LzDb0UUHmCcLCmMqKSBHuaQ5Mt+GpCHEFQX
818dxsYyccaNNtw4JuYqRtyH9I/umxfrFTfqng+FD+HY8mLllf3Ejn8/dnNW4J3d
SBhQXe1jJDAT6ACq3heeF8Gfx8vDrCYtuokj+HPH4OkaqmLgLIF/5UJ9nJjp1vR8
Kb4fRMblpfA3m9f91hjqABZVCMnlvzx4gYguZ4zTmBHhdCsraJwaMfLeIO3361o2
JP4Xs6cCtT1ImNGtVUrEEj8pSubWnV+mqZGKtxJ+BzyYadhYrtf6oGuG/YAEBA2c
DlqGNEgF9HO2mSiuiXtPESyRHI857vZD2dVkDqBsNCvTifi/XcN7zKeyMczgHljd
G2ZQG14oUuB5tuhq5zMZ9c3dX3luyjIZHgw+V4L+P8u4clSXAsR0JdRRTZJr8pSl
cqPOI+nor+zqFxFl41DqNmwgHWuAai7NLhmqGm6M/vZAG6f4e3Fdi3ccXj8CWxp+
Z+vgUQfAVO7nfmH5ZBaCxvqNOxesydZ1opzO0VENbEHLfLuXX3ZVCAiiBjNgNAZG
EjQqAZsuKU1kmaZtZ82xWg==
`protect END_PROTECTED
