`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JMJPcVNqhqH/HkIb6kSE4Ax6dqyDp4T9ZS9qxx2henRZnb8MKjwqIs3Oh8wsSdj5
K52zwEwGY7yuftd98Y5mgI/W0KMKBGCcMN0uSDzLcNymrr7yaumyOXFQmB7nkkhg
8z5R6/g0dkn8Nq2CKD1o2YLy+C4DRh/Y/p2YB9I2ii/E/8+yTySrUekI1LhhAg02
`protect END_PROTECTED
