`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O97r8Djv5tpwqtzxtEkMR9smtoXdkt402B+NufB3YeAIczSrBTyuTZrpMquK3jRG
hB8gyS2ZdWANcC9r9phNokBOrw2z7DzmQP/0egblbemZuOxM4zVjFb77eFvDkm91
MvzurE/PEXuRdbfrgVaL1Xsxkwis1KZoRkLNLcopBk0D1Q/Pqaq49M0P3Iin1tjU
+qq+6RuOJfCw/wR3XjlD9Ld14MCjngV6nJupWr1iLWubD6dncPe3rqQJ3f9eJNBh
mZWqxtV6CbyzJ1bHhALWUZVzkVn4W/Ihj4SKe/M+VCFRA/UOQvCsIyp7W02ebuHH
hgk6kc9IAPuv53Xu66OzR1ApQYU5lPMsocHFAOm6EVHLbDYScqZZyGQ16SrdFUNN
nmbyaUmVtlWs0F/x3yLbhESwjSWlDfSup/TC42ZXaKZJiX3XOMTdkDzhvS5+plXg
RmeUe8hn/L0G2fwI0jCckWjM9r7qZmkJsABmHJUhPb0OsXeTCrPVuGESDHZeceJ3
dZGj+sVkHfq3mv1d6aA2iDNqXC7iXv/lKPjAi/c2aJ5hVR2K5Ld6SBf9iYvMuNcX
1x3+02ZbFPD/FTrly5F4ho3z6EjzGkmQHe2a92dqUMgNu5avqMgShRBBRduUQ4qw
4gbknx3Szldp18PbzJX+b6KGWADwz8Mf7iBiUzSRyCXSuM8S/hQESZN8M4v2ePxK
7ZlaAYHMVGPmxrG8TFfI4lPbLYo1BSsxadzK83Tyn/iiH32XPtrbL0bGqRxeiigD
hx0yaFFbH54enb37cKA/MxZaKWmBNzlNGz+3Fd+6uMa75kPAFDU++YDefc01Vn4g
C6NsNUrLg99ECkJOVgXjLd3AUWAofeb1PP5wfTIzrXS+X23jg5SJriHhfMXmTXsZ
UdUpsdeF4yL80ZAAvlJCjo229nyKBdgSzUtZjNIp6EV1NGVAvLEmdy+nmzlfGTTz
mm27tvm5oGHj+QljCVqlhUftZHYnkjP0levrgimdic9NNO2fUJptg6yXuVKp3/8b
w8q43P53rvbZEUU1eKrURAjr2ZUUOgyzCWP3xK8Nr4QHJGETFs00CLErRvqXBLHs
5JaYLzf1f8k+Tzyol0HRS2Hdg6HrgaXhvpy6Q3CdKwSCoymQGhbBNvEvNWCD/Npd
QLUjh3SL58UeXN1AvUGza00CG4904PoD3GOXU702U9TTYufvZV6c424gfkSqxoty
fstQSv7Jr4vA/ObwftpnrrdSqQHKJVqLYKqcwWheYlpX1PU/Im0dYeYO4elhmsGN
YdpQve9JQZu1iW3qcwSM9dKM2AVaiBcrbmzIaFdqI5A6zKnOGTFz0sfyVa7Dvrn3
YrDSh7YTw7f4Hzwz6pkaWefszvUGih3E67xHBaWZ5LTf3b9yohfvxEfW+iDMXkHf
hSf3K8Lyv7zy0Ju6qt+n8BShV0daVUVmEz4FqhwSSRy0MfD51pU6MqXfNuDaUZrp
jh2Lg49Lg2QsTxKU/8XW/AJFyvylcvEyR7rfL7WOxkM0mg8H+v3E2MC0BsYEN26A
oEjaGfUQb5Filx3BMRdtcWiVXbC+rHsrBcIHToLXntzCvHg7vD4GxZ/ubW5HefIr
UpO/zy29behWPMS1BKV8uBwkr8ze566fQ47bKZCbfoFv4P4uVZUSr89m0FVkylDa
Bk8kr+1oFHl2yZ6E3tMXgGuF8538kYiTcVwO6ZD0GucOOprLkcT8L7BbVaiTdb/V
m5meIMbK5uo9idpjHcRSHyx748wAmkHtDh5yJceb0hwKqKbTxWqnEApj5M8IeqMJ
xLw3HB7DpS/OQ5Go7jOz8PaTiHIEBYqUPnp9DxIi6BlBuHETA+Wlzm4YMQPjNmMk
l44Jer7TFKmCZ0aaRXJjkIIf3zPhyWfzRhrzPcmhAgaio5BLvbyCQAyP7sY2pDZS
+1HadVYQVJKlE+rJtFY6dVd1rOKBnM4DCes0v3FA22WAcQ2N0W5XSmaEmz/FdvPL
kNdc264/kfQoFxBeiK2qT9YIXjzsQRgDJ2RPvB9BLToxoPQJmQhIpkzk2tipG8yc
qeHG19eqW3IbELXDh7iy4vgKL6psAjUZYTop/m32QNMFZIRGXJb92i2Cm5DlFj0Q
Mf1mxi+NslBjxtmeQAJMNH0ZzOhSXUrMKKb6RRSi694wcu9Fb5/bT71+K1b6kKiP
82xWGH/LzqoI6dX2dPUDJ/YC1LcyuDAlez7AJIz86THVfQAPBppv+Suht1NKsThI
B9rs+pET73ERMvLTqrZylpXYOuMKathVlgkqYWMf2LELE08Iroz/rYipUcp3UjAq
qXli9Ur56/1SQFEGFx8AchyDboPgr6MYK8oRengBMuyZcIx2glGY2BE9eXALeyvD
WOnnvFx980Z/UrX8ilF7Nur6Mn++Y8ZN6icn0Y8YE6S/byvUguG+SOKQBH+Tv4pQ
QEol62w+NHqXvSa8NOAK73T4Y0usWy0qw0EPvmZwquQoJlH2eCySczK5DQw7N53P
WEs1vieCrinBZM6LQAgv88OpMLWZnB2ipY6daBWR3J+VjHQZJNwqmy6VWay1QaUX
6+XN65AzJvSTAK15JzKtYSeFBItCF49338oUwAmbGMijDOPlBSF27pLigTmwXMKO
jPR/kF/LWPjsXCrqPHIKWc5UTuxf59BTEoKT6a/f86o1i1ZF4wO9/BFolTsloKV3
p0GW4qHIqC9+dtDVB/NZKDLZbHURPCKhJgpcyDiA71bMOrFpO1j4KDp2RUn+5ji4
kR0bmpi5h1FVQAY+PQBdd2zXxkJPcyCoQb74GwxzbPdrbW2ounbE6Zu7RvvBr0Xp
3qzsoVGn7Q0cqtholXFXOv3KvKD0Rto5Cf3wQ0GJhHveWab+XkIe2bGHOW2dcj+u
HBjv0X3MGLpBAOL2NiVxK+ZMGCEM5qRBzyvooHOsqx5+PsrS8aX9UxfDGzdxKbxn
8dBrX75feN28xFxvb5MHQj3MFd2M6WA+U/HtbWTBaEDbPxwRhBoZCFtyD/fb8X1h
RFIZpkpeKgUUe4smBy69JeVW+b+9kiVuoy6tXDshUrHMu/PwPBtpraAN7/evpLeT
Km2Qc8aMQJq6o+OEL0GJuA9tYStveRxBbhfPvl4ylRfDjU3oGsdQz5YL4BNMAist
faH5yS07INURv3MBsaT5/6QyJRkPkZhTFvASK4hnouG5uw2+nuW3ppJ1ocFCX4Cv
5ZMLxK7XWAGHlL0KIaN5OITlu1oiikPKOPa6x00TQJOF0t+4i33QHDXcPjDQbenf
qvi3SgkGy278A3fCi2i0cb2UPl2cPl1b0Ut4zrnh9S8G13Onk6cHIMzBptH9hKGs
k8oxmPt4BH+qv1yHhPBzFZVzLXIlQmEKkF/dydJCg2+hxCKIDjvp23qVj625VLAc
hvd4pj7q1GjSl1Q3u2y0cxMh/u1XSPmCSk0wOODJJMLEr5syZCikpXtlERa4yeIV
irZnp16A5REkKbR/oy6H7S1CxQAZXD955kQWB42+Fo+hXOhNYdks6FHmST2tPb7Z
bZdIzyq9nSODWy0psn82Zi8Gq7sjhcJd+CT+cqzo+3R1rg6Qogu7h9BkZHC9uFYK
6C7xTA7wFAMgL8loSlyD6NUrjb6gv7Kzg3TZRDbqlKusGZWQxEGa++jGIlcbcE0W
gdjf8ZZhEDAYr1sXBHmeq4qjQ7KVOaVT+QdpRvLfcboYYhk4K5HzsyQt9/AAhL3b
mZsgN4rGONCI6JX/n5vbSABGivrUgtyf0J7vq9GYmEw31M6YyBRTzDP9KC886OlS
A6zcUGgDTwPCgqse/2ccCT479bpXSjSyt/E1GlCNfwa7Sh+oJmLrhgIB1SAQEQ2+
jvVhMZM2HfPYC7Lw64JpfZjRNwGNbqZRqkmMH6xJcKunhOjxckawWxA62g66XWVy
gd5QDNDwtHwvcymv6xklabRiho9AejvUaFAXOzthb4/TTkUErG8H/Tz+m88bmr+y
peJM+wRrnZaELFfI5h69OvFAVtAKTqYeJRjx+qfpDHU=
`protect END_PROTECTED
