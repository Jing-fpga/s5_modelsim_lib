`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L+1o2GhNYj0d6KCdgQ7kSHmtwDhNl6q/XoR6g/jvBpGlmiuvgCgTRSgYkJ2dyxsO
zjGec+O3m1fNoTLbmwCvR5+jxCK0wO2sfFyt22c1QruNN0pBzboU3EOq5F/FKEQa
wHVOiAVsUqUa071g/+Ul55eEjG75F3Dz9QQpaW41mungS73s1BVo75iN9OaI/8wP
Lp1Y/fcIO0e7q/LepyZOfFay8+51BfrWJtXEuXSHEP1Awpymj+ZLJB/OmudKxvsd
DPLbyhlQx4L8Q/swoSr8ii8P6axPCWEEyyIVB66rCy9w83UyilBfxRfU2Zodj+VC
wEdj2feEF9Set0tD1UW3apjGiD3OwC/2QTgaefKRQR2vJUr5ynAtCsNO5D4vq3sO
NlzTjbQwhfGaf852vS66A2iJEkdzJFNxu+2Vr9tcj7+/Kdj74tnuMeZEw4i4m6n7
bqon5DzQ74247MTwzg9cgxglIH9vHxBDaEVqkqfW3LOxNo4btlf9enDoITPSzCe8
kUMaM46HaevyZffoCVEBSeYphR2mqgKDUqSShxr6Btzosnfuf/jBV2DVMR5U11oU
8a2RN1r3uafOGH+e98o8Bm/cFSTzqEe6iHbswjlQnWstlDUmWgCYfNTtkgBbDo5x
LsgtEBqp1bKA8ZVnrlTafuoyXI9jfPe/j/C/ZUQIlzIPdaFouXOUh47fUAXY2OHc
TIcPC7p6PJ3bbDATs3ESzmRCTw9vClLqKmBlL+Tr+97FZFqTEMYJN+dnxmeHJX9N
R60O9TudMNEmWmoFVjXweT8LiQq5uZi9FBAVWt8dolegV/je6Qa84Oa5uBGepC/5
C4GoWgh126v4IfU43CDWEv0VZK26yyo9VXPYONkUXXqHAvfildMRGaI0Cm/2wd4h
SvPk5eCYkHcgQN036NtH/+eCV+uxYxsl80nVGbNvMp4hPzo1tJrYY/DV3kPq9b1V
U8RLNLtsF3SH0gsNzKj4YIWeMW4s3EDpCj8zRuLt7mawHSHopHbPoPvoTSlLbsoH
tLFQoTcW0QyaJrkkSsZbtrk1Jc5iW8tOF69OGWrRQ7nR4pTvrmvmpWm5i6/esFqZ
m2WHKn279jRzCBE2qAutedOUh2xsx4+1I4r2AXJOPCWSGzb+WxdfQwNGcVdpQu9k
AphSL2bolsYh+UQt44y4i7zz4dUm/DyrMy11AWS310XY4SG6s9u2CJ+cKa13jGQ+
nqxvzMWhfnki0K8lkyEKxBV4mmyJHVTb3r9wrGHGrrA6lMknzL2DL5ozvrIeex1w
2lpXmFDwV6RnjvbW0S/3zyu8x+cHcCvUMX6Qed3Lf9DVvuPWdextdhcf2ZuwFomZ
4D5KI6UlpElwFsXvvXMxgGE++K+oGyJwPWdTOqnnRoXxaazudyNMITxmhQV52jKD
DOkecvAW80KcXY+XO7KCYRNyunzl79la4wi8gpblYz8FaU5IvyqAfngy+0BKNfzr
eY2CP/+c84P6TEmVmV3JFknxLuTOMT+66ZUpdNrEOHtfkOVaFsFU18/7dwQJPnN/
7C/goyEx6xWotSYQNn0HZ9G6HeweYz3Y3XmCyqODfMhuJgaBYULcgzIZvLHDkDPC
XHVElne+u9rVADdnNZKtEo8F1iuCnPtlaFxHEnkxolr5x28ZVDfnprzWHqTltjXq
1KjCEyfDCa0uahrxBbGR+h9iKz3VGj0uJbyj8lH575YU3weXrznDfhjgyJs604vQ
vwRwlpAQTnUgs2XwVrDbRMsYPzLumJXHHJkTzHZkb48Z8dQvLkDjnumuUCoV1bEy
mEX1f9BoHDbJ0qJ2fCUNbGNx1dzRwNlTEw06ZX/JLqNMslzV/Z3wluAPf8dy+Auz
7qQ8r659XiqZSz2ZH6mbLs7oV719m3rmlw78N1mqFqpjLxetvhOfM/H+hQapzxvu
81VagXMbyN1exiUkCKa7F12Qhn4B78DojSL5Nu+2hf/3fdHlhXYyuSH1pnblqN4d
zaC9IbSKTa1hTZESJy+aCOjMRPva48OpU3kqBTCyfcT8EWZ6qGJ6KiJlnHANIEZE
VWjug6TeDCTQz0BWVGrL9m0o0RX3dEP8gKgfS8xCT2732GkqodLXarOCHm9JZmUi
eyixWGqjVojbVY+S8Pl9mW9ImLcLzU7Lh547oEgjICq55go19OhgrQcM5TRhBcKP
PNXCKi3/0WYd6sqGBDQ9H7Q559zit5C1lGz+wsHr7RbGlCxwSXMAPlpLN8KYveoP
F0w+eBxSIfdZDXl0UULcQIk5nQjHl1MYGoiL0sf8XQuQVconBg8XpsCCr6HVYUc1
v3jkpHzqH9dk/gOrCBcViNwnIhcESl7AxkHUNqXGw358gtJGptCxn9S/bHGtABq4
AZ1ZQj6dxbkch+fqjY7onD+/ir0ZOjCbQqhEpuemo8eZxrNmcUlF9LUw13zZ3+ud
SMFkM/ouBi5VeMzkUzfR6udOh4GDrVrY2NWsKRYHGwLOP/ytafvdTVA0pUoMdJoF
9jxp+ZkeV9+ip8CP5tl1DGMQBfH4kWUQX6zGMgAmcT43STphmnsPcTQkjEdI34eq
+rzuYDL1BP/rm9r8PqcgqS04rIL3PkPnkrhJUx3go1cMCiwDrQeRfJBsVlgUIap+
jMhzIXZhFcn4QVPaXOV55NGlCc7Ppe6GGpOdmu43NtWshUxvGwfep5tQi/oY969Z
2SKs210akBQIIrAEO/WNMBFsVf1CKOZEoPnACS2/zULUiG2jBI+OaUDimmSOL4EG
xyqiFMbQbox8Ai8IGuyUj3TygyRv1ZoL7euvN3CouKQpYpWRAlUDE1mn3JzsnB0y
YKh9nkivPIZCoTKh+9kQo1UUWysB84vIvfPxsyDA1RFDFR9qt/Xb0h2RGfVw9TMm
dHYTk7aOD4lC9JjgtmZBy0l/BYatFA4214V3tQH5NBpZ+LMxfykU18DVIgUDcvhP
vCDCaoQHn0aeC9a4S0Rf/UB5jvSEBbIMEs9Qf05dKLFssXC634wocYYfjj0YJ57G
kb1VzZGPocGD3FhtHfJgWLpASQrSSwyIx2QrpLk4HIlxLJEIONoDk5Q1XMwsSMmn
U80YAZrjP4kw9NZ9waMpm7/XY3w1gxg2hhoMAJsv1q5UhDaFeUvxEgKBcN3YONHO
+Cy4sbNbQZOqyb3axzLlDOhS7BAp6C+z04v7q3rAM5xsCJDAUDIIqrg6hMlliv1q
TcYO1rHSu7WPHd0scOJx8A==
`protect END_PROTECTED
