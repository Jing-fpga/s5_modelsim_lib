`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JF++/QgiQYBz3o73d8uARxhNX4mp4QfR7MWLhYCw5vs+k4pLHGwssH0bsjcZBFHg
MeR1r4Zt5VUyBlaqi+tCF3sb1mO5zNMm+PTFrcQvNNblzygaQj46xf27YS3JlzaL
Q/6QfAMXBXf/pLgFABvk/iLXRtq6wPfl3trOQLyPzbu/OSpSywt17CxOJcm4ozWC
hjfItCrIVuQCjexTQGb9PtENkZLEBMSuPS/HwtqNj7l0cz8IQAu0GVl9r0Iweni4
H1Nm8BYMmkkGuZdevXDnwj9o0yXB3bYV0ZIPIkOjh9d7RwmL/3zVMn7JmVuQcgGQ
372w/50s6lURMKWOnTuHIGTGMbrOsNw85w7MKxlq7on76yNN8UMh/4JjBs2wW0oz
/e/9dCZc9K/4SUvbqSIocYG+ZSFV0HlPf//YZo35Fcix/BNoS7K9CpGUMTSs1eVb
lFOFq9raZqlg9V7M60JxLAhPmZkusCNVp8lN9NkTX487K5pvt9Vz1v7PMmP6Uvc2
cibGpBIgdFCM+F7IMAY3h5NJGobtr65UZi035E6YT5P83F8uQCvLhSzfO3/J1PAH
zqoGHMRJTjdl8aagyZ0PxYnw1oq1DUoSNaB6EamB79XvRYhqi3s9Q4H0foWJ0U4C
vJxTNtPYv2dbgB0B9F7R06oz54kUr1rDOho9chpJ711z+hnTHDUbPmZwFIMAqzGw
Vvnx8kMqdE2SfZfbyno/hNdmeBQXkPMAGRFXbKJrfy/7V84vAt7hq0V1xIiu3+rJ
JYMERY/lXaT3iM8+sHZrdraEzm+dKIZ2E+mD6DMdmHdkbr8HoUXJc5Vxf5HAppiR
+/DKzfz3SKj0y3wPJE3xiA==
`protect END_PROTECTED
