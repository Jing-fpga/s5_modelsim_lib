`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u3sA2Vzig4+TTbn3f804Xi/aKeHCXqYSaagf1nKQOw/j+10f7ZwWHh7gVpjdf/b8
JAkPr8GJ/qzgXxgw03+d5u1nY2fWHFLaVb8yWvYn6/g2u26zSmr0FG4auil/esjL
ZpXPXTJFV4b+O2yJGcoBpYSZ9vFg4GytH9UbJFRRIibruwseCBnadgrS2jkqQR1E
2HxJ9oUJ+RNXFrwZL/9Z6lyjZ8jVzOQb0RF8TWhWvYOuYyjVEW8k+h8t5xvPWY6Q
twfKpBbMWWocyrOcD6cWxQqlU+pO7zYZ6h99Kgw5Ic0rBWK/LgOr+z4WJX5ME2aZ
SxQKiMGOTHD0pmbYhfGdRk7ClB4yiIOJLpUg83yp+D8QuBtkFv2TIix8ZMYM4A+j
Ae5NibrP9kCDFP5zXzARWAKA/epQza3eqwtRbOhSrnsjgWpux5jh+tcNToLTwrvp
FzRa42R1OaBsi2wxN307CRNHfPMmDzyIACZOuV8M3oneqil9kxc/LIcYCfaBhbGL
ubhW49SwvTmvZCwIa9NAY4MBER43xFzpMsL2fhuyheLxoHvP7nENtek4egqIUo97
xc2cyplwRbuhLfcVsb1xPCfdrS54WheBXsG3zRinbQxEJua0iFLemLhzujjFvI/b
GpGil8ZkjtZui77U8uo5CWbRyZd1lIm0IjepXoqCCfYuiNmG+oOeJ0PkcMnA+97y
8D1uU9/kQm+VHQJ95Ilw+ytV52TFG18NfeWVIrQf9/mRK/2Xh+EMXb/TdtG6uIDZ
ZyrkqzHVgGMsuffnYzNm4k3M1NbIAnHXmEGCcVVCNJ81L+/2++2qZe3U7hHppFcj
Xn7qxRYu3aEn6Oi9oR+rd9tO5D0jtnc7Vs0B54R3V/1lDiRY8v/KILpZ6X3vmPGR
afYzBftFVvr4n9n666WPw+zjvxpx6u9PnZks73sBXv1/FBEEc4/3zPtTsP0lPWEf
XdzBffjKwDNVF/mxtAnRZWVxmU+C4zmMVltDKiVoKY+B7c66C4g0xJhQt3ehzI/T
jspKVkDv3tWW5YYN9sMHB+7emxpW2+V2v/RSHn3BBFALoC3oU7y/2Uod+HBEmXo2
lbIcnw++q4x8PdO7wZAzm2JU7kybFgnmgeUElFkGkyYh4Fj9OiTYecRmN2ARhDeT
4QdCXrLngm39fEpUIyLFabV7LqGPakV6QryWnA290KcX5qBDDGqTwfOmXDbzK39K
o3FRYWfclN0RXc2lULGBud7TsaoEX2FkBREM1XaELSREAVvBIrjROVhresPbjJrO
/VEHbrJ5SLmol0yoU49zqGzzQ0zOJKVz/devNT1eHS4/HeGrNWGbgeQ01Wr3JFgG
gpH7DTQ+yCb2yrq/MyGzk7ffKqtVjz0rhvm/jjYJ9LUSLVs8l+0VwPPSe+rHgsOT
ewb4HNV2FutgqTJKna7P5uC0VLaP4KgzMD2621hylrUtnpoPvrVSXIPiKBlzDiu4
j1onPWmHmH9EGtomFflnxmHktg7g4IAK0QXb+0HvP3RVX0zRupVaNkrAZzDh4zu6
O7JtorTuMpArrV+Ug1E/yctqExjOh7VcC88X7NdZG7mdCVb6q6DYGegG4dF/Vrku
Y1hYe8xAu3S20YKblBHpM+PM2YnZ3mfQcJErhGP+n7nNyCMoZH04GPo3DLiObfZH
CbGtL6IWpNtkln1DoqoWxj9vuuvNS1SVntjo32FGan3mILBczJVu1jtj5LBWmc8g
zC35/K1abH2oyO1FIOkEoFJMDpftU+lwGyouL4PsG9YNehd2hbfAG8auoZ5jfsbF
qY8ZbD3DKkjJPR9ynAS6zQ==
`protect END_PROTECTED
