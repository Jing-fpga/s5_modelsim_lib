`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EGW8l9DuZ8ZAEip+A7Dn9Y2qyCZYOcYbULicev2ClAxgLFbL9JNKD12h0pP+5PNd
THCYJ69G4LdquXVCE4KJ5Lv0OSPw8llUd5eOCXwQyiY4L3tQP1BVY2fH5UuCqEqI
dI1uCortZC0fk2g+FbpfvKk0zETwZptEtUZ7N+QruptSGsaa1yt2ijPXDGdRfs3y
ZhisfSpgADi2MjTSVAzVFIQfqOalL6AYynz3cCEWsS4lNd5cQ0uQOMqZp2A7Ohfc
vlNQL2NekdlAdT4v9zP49yvmZ2OW0bRsVUPK9AGS0lmaeds4emFtyZajcvGwjAHB
0s4h/6q/VKbzx9EKbW4PR8v60rNb1vhmLmyClBhDFS+4YTHdl/sT5Ia3hFNfjUp1
kfjNceq87dMpYi70uYsWL/vsTGjbnSnLPFNanXWGP7I1ufjK7J0MdeixfFa6HP2j
WvhA2lVoKSuqgoyfvasHPTATdKFr7pXvxm5HL25igf8S/Rj2SHQUziK8o1F7DEqI
qs6opTVSG34wKg+HRwoQkWzrB5BqaVGBbRzYNx2+kdM8djyjZhIpWuqCCqAaQwyS
v/ocgm693Ioo6wfGevacjEKcP20W0aiGB8FWoGMbzwguvIytPrxhyB8+6yzVD2VU
nnFXd8cDdPMaRwhOkDoSQGVeBJClAm1bB8RqPV9q7N8Dk92ywDfaOL+d9VfTFVHW
fpSEwbfLLrOpAPWQ/W4SJZyvAsrphm/FU/xV5bHaD9ssEhxSIRxQSzUYpAfR/wFG
fclKj0PsohhllCyjpUs1UUOvng8sXsF9I1vJPi0Eb8wNvqHMkJ2E1Oqf0aKP6gsj
KLbvKkdbqmOyKr+iBnzRXQfDxwzFKEVWaaCfAId9VxmYnYqY6Dtg6KsbgITrky0L
0hEn619MsGw3IovEzwB4qTWb5mRFmKZsCDAGLBf+aRsvEfsI8wRB43PPk/4q2vlL
iThuX0XEjYJ+iz3x/8dTlg+S5g1WpLsdBRFeSe2jGI1/aWSj6oHyK+T0I8M9xlS/
9llJelnp8xD0RpOQp3lnA9c9m6l4YBSupitQmMuIc2ZUVouf75H1RN3iSeF1G37z
HDTqrg4DKSfE6Pv/P+3TfxjRtMPnrMGLT1P8yOtGkGmDeLBI8bEichFJe3NtLPQU
BhGw+ajjXeZ94jCpxCxE5f2skxSxXEExBmthnMuZvClkmpDgcToFHQ7/8ArZyJLk
cLBCO+VlHp0wu46UgWbWian7RcPS6YtO9SUl74CkmQn5A7IRX4dqQ/Y9BDDaoXWx
m/y/kUxmuduAvl2L6tFx8MsI9+vfeAbG/lRIrJQl0f72Ttj2KskKGyl8IT8FmTaX
VVHKaaFAxyeH/mxGlRrAR2RFTSdHlF8WvuW8BKK6Bqu4SgfjsR2FjhUs5sv5dlnp
XiJSxrSHRG24b6xmseiagII+E6XZfCB1jOh9OsTXqu0uPcKkhdgbah3sIFoDvlSL
gTT25nD+Qjz3jn1z5twYg0Y0BdJMHjPRxk2vHbE2ACMgAvW3SqLH89xa3gAJgvWK
HYftSzb3SVIHMrXpH3m7PZ9Zr579lsz+xoa6iIQ9yj3ya/dW2vjgwJf36ji+2fp4
ETi8dMcDFqfN8/z6lQ8RqujJmul4vG1Gf9nGq5+Fq1i2w68gZTn/cVyDfOEB0sIc
a3UrniILvKwHeuYQAbUhgYh6NSNrRzuKambiugzhXeCZC3I0HEIt6eNyfmuCOy5t
xG/cdPlK4ZzjuFVguyJDyWjK+aU8qn2TfosB3ioDqax0YXwb3tBtbJkzCKJlC8nS
j8UcWAmARKkHPGui8RRZDtL39YN/K6mtgEUdRsb/s+A/pqDLBSsIJosfr6L9neBY
XXPXFOTle66lqII7YND55Ksu/1ZVqsye6pYwiVOPXe0Zqa1AeOSjJdylKkyoSZAh
WHuO4hOOMDlO666kLXB/eSfQvkZJTDBW9Tk6fH+Zj2fAto4cE20JVwCjt/x8BFPw
KTbtyzuUOoOMQxs4nnthtfQlOC07xZWopj30zzAsaFezjCXbJqW7oqr/KnrM0FPW
ljV+LMl2qO+gAZ24bSQz4d2U5+TrRn2wiKu2EumpdMEfzVuk3dWCWHd/PgyaoAZg
cDOwyhCse8ENXjNJ8FEXmY2HOg4bU32z2e2VhEv3Y25x64LbJjpxsteZffDRQk2V
zomzyeClWyRDvMpcliVn9bd9SGQLMSfbxY+Ku1xjrYyniZffC3NYCsk8uIWJUh0j
DPCVwzKmZNvnH19BWaztFTiZ40MB0sOZtvxn8pZCVx+YRlNVWCjexYN25dTTHvVE
117RAXLb4ukI6DKNolfASSUiKlNvjBuSsmLoRfFSWYKv7QG+EhaKwidMaDCRTAuJ
ghaJ7tSF0aEu0pdxSRIw8Pr/mwSr4MnT8dn7Fvgz4FJ5MAUl8sBunu+s9IDnan2d
WQ4Md5rGF0wdD7AOqChm//qZKawRDqOEC0mKar4B8eOyvKY2mq4zEWXEf2lPtzE5
`protect END_PROTECTED
