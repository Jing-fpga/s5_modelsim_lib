`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c6/0ul4TB2nYMEt22rx8tsqxzvHeqIysXPGrDeFc1ZegAZoxUhJtH2WVOPIWfPQj
m05UgQXvU4t6AYBO2v8ou8+NF3smVFoBeIKvGiS0LH623k6wJ5DVVAGSd1priv0Q
aE1PLOXBo8xXbE6eUeRpuAh/8yzPtV+8mzYJ5yLO+/w0ruZ2DNvVE6CK68WbR/f/
RzXh7/pfXMEMjrBjFkrO+EOxinuTKt44Tnx7C1THjQwo+nYt7pq6qjyFk7CQFldU
SS2Qo8nOVI4nuicrcPn/uf2tgXGJq/PVuLfUvMjmDspqg8kni6NKOs37AekWh+9Y
aCKGD3PlM8jrT/7erAjAZOcVuo61hiu1yxoj+mXnvbt8qYQkq0omD+GiErvGFCSd
hc1yqPI/+WKDfVUrDBN9pGOHJ+gqEelAJ5UCIiU7rWtAjreTeg1Uaj1nXEcrH33R
e5kgQnuC/SQpaZvdDxHO5K1CwrHyxI0xQlgZYob29chyRT+6JuRllieGTxjx5EAb
ihpDzCIsLg6XLRgYf3bNi2HOrXuS6QgN4zgTj+bGeucXX/R2sSGQqSzYzSlQNDoV
6selnN0yhtNctq6DpUUdzKJzX1xHrjNL04ePweylRRLXH2OFGV1u+qDUQ4tyNYp4
9A6dv4vpfSVV0nBHJcVTRAnLEbEhYevjL9Wxg8YIug4PHAX3eGqydXIqqj5tfbDk
u1H7Ed0FuQ5y1Qb//Yz5nBvhv4y1vylt2tAB+dCVAJqObWzXtz/CpQo8X5OuwJpV
Jkyx5pdCCT/IT9welM5QGkuy6h0ZvFg5LTb7PDm/dqBYmF1IUGUMQfv+I61Btb4D
BpRYPx8fTiDlXTT2AHFVVJXNBLGEofOnjWVwf1utRYbvclpoQMy842Ka8QQNHsmu
c4pZ/E9V7gY+x8oNw9dV96LgOD7d4PB2E03HhUhKlL8gMKRiSek7syljCfLywygL
JPvWTrG5qfOz5UAXExrNb+Ut67LauGJB5BOxqC5xR+a1tg1WqhW08UOeyKlsqzsL
FiLmBeCGT28jg0sfy3JpMVjCBm7MznqKM3diEaIUq1gvxI7m6RuSFIjZdvcAOJpf
7XR91MYE+2rTGIqQ0hHQooNVe+7m3h51KiZQXOWZTwWLdfKm7J7DBFgxiX5/mZru
FmvgjHPqIeOBlq00MkvBJDK9gFJY5SmDC3L/OXzXLVGcz53ccy8itY7Cc9dQZAmb
W/Oz6Po4thjxjdb8BixSKf7lVMomoJeLfyshwmW8dUamixuR1SfQ7kCS7nOJ4YP3
5ISR+OiOcM1ZSTKs1FSY0s0V64GxIhq47+5FZKc4mPDxGSGB1mW4QBzFCfUADzTc
/XR6ISrscY7sECC2+D6iKXlI128qtgSGpcHoBnDIc9JSX+i9/GjA/KEs9l+/a+FH
anf2eyXbq5r2F2xhj1jYXc4vlM300XzoKz2PhnWIz/aevVS7+jHQLVXNIQeqLsZW
zM3uajkGRpZS7749uYud2NeVhwrsH9jDhqDGlGgUZdrSe4lvuuuPv1tsjELWnoJB
0VdB+Xg9wf0sYyrNR6fE8ZDo+bUAcryoAZL+g0usih0rkkrOt/p9XGPmVzpTlcj1
n4LJJdtijdjV4Fq0NMyxDjx7hMJgBnQNPGVJWs3vjVyzXuYb5gyj0LxphcH/V3w/
XUem+N4IjJb7FFF4OpM9Ebc7s/gSf8kqsSKB3mQZqjx4SL5jVW/Q1K0UMc7H1ntO
2tSWjmXKJe+plakDCgTVYuPYQVgibQmxvft04Ev6TQxJUmL8d7c0mK0jmaCEAhbI
TrjbP/S/yiwpkwv61aPF/cknt+VisdQiSZ7S3x5mjGz9RiR/bD2O2pUeyGigzuiO
K0e6U+LbatJqLoAsxTdqY+DV+V0avejN47oTcfoNo9M=
`protect END_PROTECTED
