`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x/SHHULdMyakdB7j3/XR5ti8L1Xqc3dfayNij5/LQwqU7nbzS1+nhDKxPy5fTwP5
yHiat4gOjERu5ADOAOtDvNwJT3xqhEZBOaHcIXWwW3h+9xGTh6GJVfwRbMmf1RYQ
ZBIjNChbwTY/atTHUd5AIHqURzP6zuAUxOQBSMlTz1qQCCNi7N3VO4pdH47+3MGt
xgWMuNULc77wIBEae+gu5Ye95wuBegNc8B69h+k2jKf3Gp3NYxVtwk9Pzut9KpzD
2VCKvi8MMNIGK8ckd9sHaPWMMlwDZeXJXppK33Nu1Ffy12ZYlVqSC9YRrfA5GQbJ
dNiH1Az74AXP5+HI5+BRxvvJe0gV9igaGT5RIA1bVVtq1ncOgAgfR3Sa/mw4mxsI
EgymJtds76teoC7wmCCGM0z0l0Ad9DNThy4FUYH+ZPjMPjHKYqG7cIChJI1M6JCz
R11hUbofjxkoOGbe/PvBqlpAPgXiaI4/eybpztdqUHEoVfpn6d8b3OeFg4AQWtrI
4g6DziMduVbZ07byJEe765WiwWRUgQKsSkTSpRBjZb4KtXyTOZnH6u62IeLgKtNI
dzQgmPeLrv9R6X6o1YHzgfptGOYQf9GpWVfWjrin+xC/LOW33Mop+d/Z8110YHZj
/60NhmqdcRfLviI6YrTBAIndeM7boYthNSMAP/DycmNfiDkp2Gzj8qB6iQ00i/Xo
3+Y4B27Ruc3ePijKJeU/1sYxIuBHXaN7OovFJsU+TZPkZ/XZfYyus4wxGsCA8wMF
xHS13qRq29O2TMpfSS+f0pb4yXfnh2Rs1OvvVew64OYI7AfLXIBmaznayrKswTX9
G0SVMr/PleO5SxqhS8kBh6byFvDhRho2ao2xwBDxMUzxZtXEW27zAGGJCaX+/zue
qPGl8N6p7kPqcJ56Y96Kf/GH/CSi/jGXAlkFXaIzejm/IjjFIJanuGAhPsW+QazX
KqQIISWH8MZLo9r3MVraWlLcjcRkbYSKMKBhq9ohs2+pmDI5cYsFVw332N7PDd6Q
S200V8IlqRTcodAoYmkBuFUnyXSYMaFJnOyPBqIWgK8=
`protect END_PROTECTED
