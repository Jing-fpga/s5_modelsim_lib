`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wh19lA2GgSy/bobGRRQvEYrkptTbg/oA9fmT/4ZUU/aUw+Wh+/iFn8/UC1yEV0PQ
ngLkbT6c9P+RupQImKsBPqb8q/1FwL4caWGRYe63UiO9iqx2eP2zW+G7EqUJUeAZ
E+F6FGuw7VNbpPcMqTnBkN8ov2dLxGfFUkNHeEcXnRT4W6zMkgSYdw3EFmPchz36
+tk+52cp5c7WIfgjQtzIxyoq8amFogr4ELGcjTP2ZUhCesjx+7Rk/XixXaSoEnb9
zN/td6U4yrcZVbQySTRzRZ5gR1Cwr40eM9nyBWBu6qImK2+J9aUdmDBMS6fCw7a7
sVw60/jFZXrtGg/rsXEBeQLX0lgmaFLLb/buimoJKmblHj5jq0zy/7MWpPHE3oXN
7FRyZQEcfprD3WgfXqws+SnRsWCOav9lx0vyE5TND4KARIzunSxUa4BCxYDJz/ak
oa+iLZ+z8aPN9YyGcacgCg8o4jlcmZHHBuXobBbAgUZ2xfcEC/ciSBjdsdWZRLBq
iP4l++C7B540Sas2XZIcEgpEFteXsaejEzau2cAMcfu7mVaJcZRb6AgXa+uMbcLg
xWqO/aBZHQbQO7uDTmGs2cDYCzu26O2V7mEYp/yjMRfSi/E/SOUCddUkOlsXAwcg
8LW7DhnRR2Br7pyL0snNl/b7q8hMteTSsjJasdKI4o8r+RBSW+DanpT7Va36VNnK
tEZEP2S9jE39fkb8CGmkpGClkWZUSz9/oa0dxXDw0xGJBK2gB1NPkHOiM63QaSP5
Xlm4ngP0WfJ6Wz6D8yQTHqQYd3o07j2BJFiICcCYdWCRzmzOYaz9qfecddVWFhug
/xGIZkSOb+nx5gpwWQulixYvfB1bpxIf2u3mdE7bkkJaBQDdJYA7VPCLgJWc76uJ
r6lwAp4db8ZGWESvDa38fUSfcvF2RjZ7N6NJp0mlZ/Lk8xLavsaywGNKdHpQKAeV
9jdQ3ixIVdeADM6MGBGfdt0CYVU7G5L0m2324LoyM0fsFT7FYgdAvut4PYxIF/tH
KA6gdTUlLNZ1vXLyRnZsMk8/+PsXZ15fNkdBNc3TF6nmSx7Zs3OFKW+S28xrG+wg
BtJ0Wf29gIxuwa+porJtFZOVEkuhgMNajTrexrkshu8=
`protect END_PROTECTED
