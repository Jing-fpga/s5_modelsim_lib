`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
62+CkHNjHLOnPV3163nTnpkgJXSOThb7Ywir5QKMkG/d9kjXJ9O42pPTYeG6RxSs
Zr+Dx66FHMFIGAbgsl+L1LiSHJ2VVMhdmI9IhmraJd+iRk22UKEgxGVoeVR7gKYY
cb1GY0DNb1xzXA1TXkVToxYp4SmHtCTmEMR5CeGjctijDFbwW14shLLDLqvNX5Gu
D13D30XNsnMrCLOXfnbxNqCotF8JqET9jcCisa3s5Jw9tnItTG38UiQ666Sw9Dtr
9smOjMC+krK+0KmpJOXheMlTcaBO/mmnN7BJFpFM3eOR9l2QYIqUz8OBGPghUjDe
Sh3elnCNlhD6cgztw66hTJ3gL+E+zsX7iso7WAKszWobP9FQldPDY3ec9jWBrJbz
9TQoS/ihz8U2n1S+WXZD2KT21MZQqpswrcfLeIL9ANMtBVN+GtKLjTNm+H00gbGm
le1eJ8afmQ6L6HTc0rrsvv/j/swHdmzbChfjsU/wmXFKe4dniOYmUKjn2rA0vQ1t
EO/9fIzWz6OC1xxTtEQPYcuX8aoAchTQjToiVPoegAd0totGh8tQXpRt9j1M6UM3
U4dLgLsER8mB16wKf2BAphDHFyRxNVomFtHCPAcTSezxb0ZtoGB967zondOIjPcz
BcTrGObEtafIHWdp5L5UgaeYfK8GcxOxIW+B83koLqv8uJk6NgrI/2TsXUbs3YRI
EdQXjVilyy2Pm3arSWn7PMtYF2yhOpfJxJyUmTG/s38uPFXvZbEGYoewLYdNs6Xo
LZJGqOs4S7NF2X4E8kHy/0GcdUFHGAna3vheOHI4SlcNIL0IIIRR4R4hVWw3rTK5
pOBRo0XNBbnDPLR9ptcfjkWrbkQCUpLoUEtZDZwWOe+11F8A9blvdjIhEcb94U2T
v0WjnOH9RQ7839NrqFKwXPA4nmjllxWpuf9kXsN0bwBO6qRw62SPZTb1UFwQlLOL
XNSnfVT8uydPfOeMyc2wZiz93pwJpGpJlqtPynt1REorDZ+gxxU8/r0TcM2ULdIy
rJPNpGKulBHa6d/o+h81caTjIHE2i4kybK2lt4bDKMJfvOtQT1F+90nf7VByZgZJ
pNx6MEcy88cJka8Ifn04Il4+p9c4+NZfg69C2iJZIlTLhr2Ra6pZvhAFmkZTI5ij
eZ5kDG4bMg5lWFEGjfSixSSpz+iUZtnTRQ/B7D/B0xZNU7CPfdOEaJAQF26gFF5B
fYOPBc3cVbnClgZGId2ySdRhgNMHZWXADr1NFU1Ph+Yu3H8Xw8m//yWyo5w1dnaE
Z6wRlw+WKeKow2rXAHI9uByE5KaViIgX10t5qUGdYuzftCqTtVQwD34FFZzwjX9g
facWlkco5jbQhi4byaxteO9a6CN/W7R092YGylBF1N1mKe9W0JnjFE9JPtCpunQ2
eT1+jC3Am0sgsQNO4GwBxoDMhj9+GWvaDA4M3EKNOnzgZN5jEgyjNrIsU2FgTQ1I
rYdzv7moaOLoeqyp6X8xlp243kDJaixl/ufvtsSZwEnFG+tuxrV5+17NEumbpWqj
f78gJGLA/9Yq1ykvaNxvqQnwZ4eKX1RtGpsoRRyJaLpOqVUh2e1Cv+WVb33pVfTb
z2yr6lvauvgqdK03FL6VCfjHL2xZt6XdB35pinGRs7KTpgzA/bZKKEJjIA4h53pF
9mJlxAcwFyUwtIOWaw9lb0M+Zf9RkdIr2/an+abaJXZ6PSzhNS0YWrMzkuPFGdZu
u9/IOnab+fZFmLeslh5ikiRRSblvRVHXNRcNX5n2yCLgreokUJ9xEbNla/KGhfGn
LnEEHcTzYMFg3LOCZk/3Q2DnXnYqNLqezK5Q5DnyCubhwFElOBI/ogsOA6LUierc
+Yze5SPh+nLnCq0ZrKrrlgWW7DFPGWBZ8kCqlVr+PCaxp0cBuXxDl2FcG8WVzDYT
5AplZZhXS2UKxoyO15CsXE8Z+OFEXMiFQy4TYHx8EqDqzjmUxbn6t1itBqLt7aS2
BauKTyL+iPZgfEV9jeCK8I3BK1eJ81iGfC9woP/x+jZ1bZUwlJIwa1HBk/uf3LEA
kQLAozOTihYhkFaAcC/SrB3oQfdIl7yRUVjUQopUYq6Mpyo5CqfCWutsKU840JRj
tA3i78GrFyXL2d7fN+giLR150cgrPt90pqqTu8xW8lHIkFrx+cHwlNdbfuWKvqje
dtBiYRdfDRmRexIkme8w2leqCKgkUILyAWCud+sXcnJmNfBmEssc8W14olleQwuW
m1H0ElHlejvmKnnxp6m/JOTSA9NXrL9XtAzFtGij8tl6GRRoHTf7ZtHfKD20tssz
mSX/o/SHpACk/p3haH0R7dIYVNFqzH6gGKkXWLhVqzQ9TEQchWlM10tBqkrwCbwC
jOOsbrmzDbPD9o3sVWvQEL+TRWGYaHhwz3BZoh1iDm0Lz4GykFh4QqDO8RQaEyTO
HTw5tdc3iDoi1DK6N/a41p1Q1F6TWMH9TWKg/GQrx/ifD0CxKmPfKHU5ez0Mvtop
vYGAE6GBEMmJnbcs8VIw/uyPjDeqmti6pN22yjtbPxlfWuoBY9HgS7OrMVMdNjm/
65rEHhHfP9VPe9R7EJe82JCsMDDUj4N88n1tRTwlDSV1Kml6spFf610iT55Ve+xo
XL4HRWXdjrc0uVDug2XDKLJn7yfOMviOXwZq0nb77SEDc1HNY24zkD7/Go/yeQvW
KQonM7d5+a6bRcRvAFk+RxCf5Sc6Tt/3sVFqapPgckAL3Ow+5X1EhT3HBktAcWj+
Rc6DLXUkTHAawTjCjXkZl3nCnBkhbhXw7ZsZPeDrCpfMchUlzbE7u5OzF/HS2pAw
bpNYNNu9R1e61z0x2o61wbPcch6CGZl3oAh1DXmytAyWgLcNMozzk0wBoyM2TVi6
Dxe2p6ACOJE5QbKk/wQtnhGPXhMZ06yojJqrrUsLYk3h6iiy7on7YcGuwGWky7hF
P6MY7eWDlBns0IH5UCWaJAIrkyGafduqbfbcHpRBZg9BpdFWEjBGwqQLRX+m/Odo
/9ifHw1R1oQkrO3W19KX+rURUL4ovD0A326V8lNdBa78PT9Fu/R3m0UNBO7dKWiK
X+GQ3ZImj4LO45dGw6rQYCAHthedkWtE2Qz1K8gIDfE8da7CgyFAsh93XdaeawFr
VkXo8UZ13HhLNYwC2jF2psxBHY/bEmDNEQAq1OGfW5HMNRzNgnjZo805p6+ZbChh
ccqFirjkGz30ThJ7kFrlOjeFAZsyBLnPMJ1OPayg4gN3P9eO/MMxCtpHE++sHDC+
l455iD55mLrLrgxhPuazcF8dJHxwkEeILXKe/X/AuLQOcf3YwWptJU6m3NVZuSJH
gg0nu6P/VQ0gThbA2vXgOQbgGW4pPn2V57e6JJ4FCdb2yznsez58S0R7Sw+uWnmR
Oth2gqW5OwaTfsCoNYv2mMR5hkHZovPusfwjCaE6oE2l0aBmoPFpBqy8yBC6i9t5
RvT9eufarcgqYnc0KUZf33rPwmP9kFrgIqTcaAMQh8o3CAQ5rAcI/QnObRJyEdhI
IjS3ej/CbvuoKUzYxr0wccIBuuPCzD5Ji1riBy0tk0o0eWj9TGHpfdlqo10Kw8+p
fm6mNFPnw0xVVYuaGediE8BeuVKoGWBDsnubcdfapfnBDQRZzD42NJjAh7xiSgJL
wrvfsAPO4r5vadYxypRwrPKavJkC2xJ1zf818+LuJx4pJRvKX3PqfPSByBWqktv0
r+v6FTaxe/yX5aie+9w3J6sgjd3OPJ582BL0gtbrnxGpVRFKwIreP23SRuzINpF+
dFIJ8E33z4HhaSKmLiLxhqMQypqP49pOlUiUUnUbmjkvm4V5bM99SYgpqd4/o/6r
JkTDnYc1MrGfdWRB8PwxZUTJ9orAJ4dKYdkCRUdxKBFEu8bvWCYWlq2G7Ij41Gd1
RacExZyX60h5NFNA5B11Lv4ABJzIhUDul5/bUvpYf04o1DhfgikuGVJWAFLrI72J
xXz2/lylCTrHGStOa8u4ckkMnKamhG2TjwxVs9hAGc5DClNGuEBSWbOLvLDINDB1
HjlmMW6zqd0OPcyBq+nH5MprJNAz1N2hCweYkojmK4jN+kXsuPHjhq4W40YsYP7X
r9Wp1PhbD8PYMhSyjZ4+1Z5AJHjwHDkZPZ8WgJ+7vsfME01P6OnGTGhwHLqdNuvC
eMs2Jx96RX9xVhUmIBh5F9BioygBFcN5Zs/OBy5oMMeqwxRKU/WG9+Gtxd/8ZwgQ
EpAIX2o6VOlqYzWUl+mIMqcyGAl7mLZS0PstxRtrQh+OVYcysry3l0a1g6yuM5oT
OcbfRsgEeSvcYyTt2qmIs61CIWVRgCJwdQTdUwQJayxo4dd4OqG8xxbULPpaDW5m
btOktUab2kTW2E2OPBZKLgWO32sI1TUQjnU1k315eYA/y+GoGxgE8fS04eHUYl8j
IzKN+GCeavRInhU1nvC9dppmlo6+A+pFTWVQqkW95cUCuiuDSB2LPcTLbGyhqTmN
lakR7wNmdE94hf/amGAcNzNRfZWp0xVdyckI/Y1MXxdR8XOYeOndmYL7OnjmWiFM
jlewFIkPy4Yl0AcbuHNOeZPnJd/Q4gXStoXdZ42fmI39guD/2JAEjkvvNH/90HRy
8bgwpNUUZNoUrcje+RKL0w/aClCmMzSjudqSUZ3p7BV6l0eUxrkWNWfs1waNUfs+
W5ffC2L1Kt/6f80IYokmedhNU4NjbGnr9dAdIyjoiKrZVRj8EQu24gHHBR/uuk6Q
8PN9a48yYbC5PArg4TssacmH25UXcJZZD5aUbk+vU/ej4b6SOogK8Vie5+SkYvre
jEqWzK0vtPIWOYUobkEnfqR5+JeAXssK7BRjYicOIMjHl9UlATJpwKJgX0+bwY9w
ETj/1UOgu7AbBz8Z0hmdWnniwbkzgK+eVQ3G+LE1DQhqcMROCQPmUgrj+Ags2tNH
K+V7m0cS+hV34wfHaWtEUN0/pQ9cgPw+imb/jv7WOfm9ltkpnKuM3Nk5iT5HF+ia
bBWzCK/nkvtgQLEC5TaXuTPgm5W0cyy7tJRnGhpYeMaF7+pblcLnq9d9SUwOVkfX
YqpASAmi8f9sXK+DTtxD56GF3eAaotMV222dRnlhAkjW3vFfZGsSYD7OVtS0c/qu
xKQFzMSJVXZUm08Jh+m6X54adiXOKIBF7O/WvWJEZll9ikqlidhmnmYJ9pvDbtHW
itQoMU6u1FFJghX6dvSnqJ7wqVji+4x0Ax0oEqCT8Vw1p0dBIQjZ4GpFrDrCMj0+
ywMvmxVbjAPRwEjPuQ/yl0lfXFWPaDSGHx8n14+dbfcUr5fFTLrpW6/Q76OIDJcB
DVRujznyuYZUNcHDnSaTsX9YdjSqZ2bocysawFALG/lhNiIJrBmEdgwBBnkb5ZfB
NGkfseiQ4mtov5awa5mRja+j5BnmSUfPPWTwiijibmTOqzUTg4AKsIePAJX5e3LC
4LdFBa0jF2a4ZSvWWq2IdH6bDO03k6HFWHCGBbd8yuOVN6KH8WVSslCn/0BlZU/r
spPxKHEcHt3d1fl4dQZJE9d1E7eKLZzEx/3AHhN3bAZffQNok6o0cU8rPRiawzYn
KcF+5aLIO9EGM5lSLNkbTCVZjrhB5u8u4c48TChnM/OSi7m1YNg8jR+3T7E4giaS
MRj6jvfCO/QEsP+zA5mbqxMfw7UgcJjEzeTCa8m2O74sE2kA1B67SN8VUXw9Mblq
+a5SRnniz3vWpQE3woeqSBSn80IXhSGHruIHUWEA2dZCvp9KvPbYnOgcvehTLeFl
jcwBAqJe0CMu388wGuqInNpUQJKK/DhoKtcFzWSpKlBSNaFUBJ7VooWzDMV7CPFL
OB717NYBeLNxyoryGvFFU92ZnzS91eGBvO+wf+zMFb01g1Ebipl1Vjiy5jF/FFh/
/8/XJmquDjXMSm87BrhR1tB3F9OSkjRnxD6EVaM3Wj/TSlh7TD0zZOtkqe/9IAkY
yuMH2MeCGRAHtQWL4KqWFj5MkDZMGdCDk2z1oQz3j34O2aXl3roGh7U/dcAD5+MI
djB3yLtXOhoVYzv4ObVBgTTbiAwJAyn3NOJMoJ5Fk0ya9VtThFkkpWcl1BXShsef
u5DJnY1+nJjcuvwoLULf7CWK75KNLYBiqmmrS8VC3QE5fc2BYr6n9GaNJmDrum8C
kNgBXpSV9PkIZsttfoI1sQYW30Kpo9j4eSoPtFMVkpHDWO0u0pvMNaLPGo+sLzaL
xwoRakJQNZlGSnaTpAkI5uCI92NgkcgpsHDXN98o1KNFW7LQDWjRh8lgQ2rTn7Xt
uU+4j+weprq7iSkL8ZSN5CU8scN6PJ1r53wNd0bHJ/SmI7Jlal9huHeLfhUpn62t
ySn6wt+u38viUmQdPOnnTbd4NObYHaPPKqd+TtJcuyWsjoGv660RMk3J4uKxcbzf
hJfE51dsTZJCgswXcL1KdOFOXKWhsmGiSanbz8IO4TtBOKB08UI+HRLaGpvHS6dd
IReMeY9w/6gbAQ9spOzG58kjx2cF5PyYsuHKUr0P1hAjz5GXa5ufsyx2nRwQC49o
Ov+hxwVeo5QRSyfeSqJ9cKnpi14ymbPWT5TcJ/cgx8Oe1FXKXj1RfuCbvKmvODJY
lbhbfDW76ercOy3IH/v59pyyJyNSBxGvPRtnsEKKm7FBZQUVxgaFnxGljDc6WPcC
MIjrWa7r4qCerAGtOwsu6e05eQlqRWB+GOgOP3oGN8Q9k3jKCodWaou3FQsa2qpN
0qBB460tAltVT3V8b+LMJ4VhLglvRvFfyFLxJ7kY7Bx6vhQG6mqxA82c2PWpAH6V
xJixVfgxzGchsdB+PT8+RdUENPCRetLvHBBTueYvw4L7YKQVdE0qiIzI1mqTuf9x
muMieOE5fh7GtrikNEm3XJPIYpTwaNWp4bvh6kvs1GykUKrz54xgB0HEw7TE7JDl
Ey4MgvwzxCpshgArsByfSw0vJYqQs/I+4uKsAsyyygsCG7oijkN6CLBi1UNui82F
19eAZ71OwWBOjjcHOgadN6yG9jYfOtbCQda5+tWjf/7ixH65n13n+m3Uess7ybBT
hG8nEJi8Nmqq4pyI7GXChc0MDGeSuTivqsFwblVxPLemhv9oSZD0+01VkrUUuc4m
P5o/+OwSKO2wu2tVbDPdHD9BSgmU0QgHn+pw0RhH9ju6rDok8wXA0ODPbyaJtV0+
wAIShHU3DZVQmn7497/ngUzHZch2+718DF4qzG3C+DU3h2Qa6r0fSgiyctXmKOOb
rLkRvRFF5rjGv06E/hsY8OCCOrVNv5UM24Aid3CKuI4Go+BqPkSL4uh1f+VPFXuH
CR7WkuqZUw3XVEyrOKMuwebletj/m7/uDcxFZWZPtfMe7R8lSNjFN778du2wTMeq
tE5Jx+MbiDAw+kn3yjzry67taCXQ1gQGIheVAmaA+vV364IPg3frg6lB2gZwk5cF
0SifKxmCvxR6coMtRpBarSPKlSMNX7JMay59yuYmfhNYPvm3rEPquT1V5W1wfhp0
4l5/sHR8rfonU/k3wiAULTRU53PmprhvKQMGpvqhqlMC/T2hE/Sl6r541yuh+hbQ
UIF+iTzik8T4iyqAX05KH6W0KhPlM+9m0ekFOYaQHyHCSqLG4hy+Oh4oo4X+hey+
dGEUclo/nOC/FmGecNYeKyEVuv8eCCqJ5BBNrPWf4g3OfvbHRQiQsc3mdbXgU5gZ
tKcYXypxjYII+8r6BvrGD57z7IiWJXcXEK6ByLyBiLw0QhL6spUUqTnUx1kwlz51
1PtxHy9TxLd0oeLCo9KJ1a/8+z9IKmtnX7reOAZJIRLXcQYzvtrSi3xqVaMzkZRA
TQlISPoGTz89aoXTO8+sCgGAP6/uNngMUicuZKH4ejxj2AbwmOk4U62oIEpy9t7z
Cb4wrbhL1gKwFTdjVHB+mZ69/zT1RzMPLggKG4ron/GB0wsayxyUvbIJibcOVL3B
zNsjuvYPrSI0t7Xa9g2ub6rqud1kXEvnWXOU987mO8fzmU+C4UhZRBAfkuorTR15
glS6YJUVkqxJklizcqWUIZhZcXfuD6QRCvnPjBNRlEDSHKZxmubQg85LHnf+4H5v
vRX4MBR4T3GW280rx3FT0GVQk2wgESxV4Nh7UA3TaKM5bhKvMauATotRcF84d/mZ
rR5Yk4eBKNYw9SLIexswR5WK3AzzV/fsxyZetOsz8hfP10BlacITvunzLAeKzIQA
88Rqk+jwHu5bBPkdLGNb4I+AjYX82sUSz47jF18JoPXmfRkcQJqrUEVD6pfr67+v
86muxwg3qIXtNmmdWHY20awoHaXgexg+sthfkuCUglMcBaUuuU+r4Gm7Tybgg1tN
1y5igkqjuk4tSoH56SzRDzsOGs1fG5HPJyWirtXUl4kad6G8WODTbuwrdbQSuqam
WUsqGOXNqJmCnEJ/xte7iGte/txYU40SeDRjimS1M5EUJTOW+V7+x1OnJSpJ+TSm
xVyDevkmZKqViySS9s2+YM3XX5GbgKPMRYa/dorWBa29Vxr7I/gWj6Cap9nHB/HI
5LmyhoYCgHYuyfk5oh529szXfnesfGbHGGnVWqZRij7wweIU16WCbuPVFRbLS0SF
emYN7MK/nH4/XSqPvI9xUh+zvy5icXBDwMoJjOrzAJeVjAQbYkw7jPHbyK5GKOGC
daHLpC8IzBQd8XD+nh3P8c5M448ujSdVlE0CGuJCg3HyeX+R6szsm13cFuiCfcOr
YGsLA3hYvTvqF2rlS0HTIXqbISp2X1HhBCPm38MwTr2x6DbKCVQFReBr4aDjz7j1
6I9V4p88gLTHyzjiUtNTT4P0E8RwbevLNObwKpKWAnpQK8rJ5fXOC83QPtQC5966
l+v+Lfm1KnG02x8V9Yvt+PJDv5QURSUimldBjtK4M95xZ1aMBCYmD5OptOUSaMrc
7a1YKFmKHcY7DL4cfn7Ug57Y3Si70TZahmX2Rq+wqfL/oXwO3Aiar4fdbOhjmcBw
NkF/i+jpHGCY2TIFRp4XfbrsAQPLGcW7bCRF0TR7D8lpy0VbAKfSbOLwoX25shPs
aYVwu00XSdWa7Q2xb4Fxd/x9+P48l7jxeG3/+WniaeMhLf4c7/JaLtB93tdWdzi9
dIkl11uOmQ5is1hiNvj11IWLgbdpp1bF1X1FCrxFkpHo44th37cMVd+7t6BUlyEw
nioNwd/rX2tir4vVG1793KrpM5UvRfsoSRfo9bR1aeLGqXHgDk0c4hJ4bTccPiNz
bHRWeONz0GaNEpngtR6BY1wqNrYRXCk+gRVrp2UCs9ZjgRcTIsJXrj1yOr5M5AV0
UlspuTik86u9MCguWlb1QlmqCuST7ZYJY322+DOUPOSTHxf5adHswya1rMQeOsJ0
ksI1D92sedNEa7uObJdeJ6jF5j67fgYjIG8yRnJIyYcXIJp2kwZnEkOetkSWHKIm
mTR5AtFhCtdTzZBJ3AuuMQ6VaRQI0FU3C02Sm1/dzby5eWUAX0VauAGeOwXampML
xkX+BYlW12C/0UrMQynZT5z6pECkYnWvjXszwFYF3vwXj5gh0GA2zn8h2XcvPkjE
aH0AUHYPA67zeyCK1CQ+GLlYOH8tx6HDrdbxtf1hH640AEjsqxsmfYb9/6FCa//A
Q1Pi3Jzq/oLXqY+VwNDBnIDsPYL3J5DQ9WQkoN+mHNaj47b+I3FbOYbfIxonvqx4
4uPuYx1eM8Cg09Qq/Z5vcuoisVJfztW+KqoboU+vtR6x7pVsfJJ27gZS9LdidPVs
QYyeqQ590Tz4MzpHj/OraMMLcQwDt36pD7btmHUv7D4IHzsOidSQe7TtddfF0bA2
65Lp3o906Sl0nhsZ9eEzSEYsscnbNdsxnScfNn8PKMvLkEL9FQfUlrb3Y7OuEeDr
L+Xgp5rOHdWFydwwnwQ0MkDi72kk0IHLf5cOZ7ZvsP6iAGj42j/WL3ah5JNFd2Y9
o7BdUuzHCdKo5i2hc9BF4uSAWJkyMuQOBqRkE863vmkXWHdEqcW9E4Pijv1PS5hI
PN+Oz7TH/rfyV4TxToq9HtHMmORXudKQ8VDwr3x6OqzTRft7avhCcv+DDsXFAQVT
9Bb5xIk8Ymlp58ZLvqk/Ebzw1UiimUApqPR/OzTm0sCTnBuUVxGU2ZDARo7Ttf70
R9M8S0vtpbBb2uAgc1f9TismFtio7jA4eMt4SKWH+rIrUdF7D7wssb7tsig5qZ0G
fyYtj9EkBSRijevRdZoRFJdaZIxbqs6VH8t4ejC57DTKA4Qwxsrdp0KyKbGFnovT
Bd+4majvm6O0uZ+cx0RWSh78tdRVWjvTVBPtv+VdefFSdWyDhPhi5lm7Tj2d7LIQ
lKsPFoWiRtyeUWvdpUR89RUPaPIOOqSMxa9HIJBDu6GssL9uF83VU/GQ80WTZpLS
7wFJUE7lITxKB+vWDcW4bt2dPhbZFDCUDxfsZcNb4QJmWaBI2syCokoBB8C03S5Y
mZtc0NRGfpKxhe9VqH0Xtg==
`protect END_PROTECTED
