`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ISZMtToszO6/RzsdrE3s+3xVv3XbrAH93O5swqWepzR7Jq66+sQvSCz7LLPElSrQ
hJj/c+uIqrwa5ObvdCwgyW97QdR+jedIB+Q7chQkcRNzCHF4fyPlJfgEr1d8ecjD
nY/1fKldiFXsYzS8wNatUcZcOtNUttODY6VOMlSZyiuwYKJmDThLTbK/kfiSVsUq
AhVAQJTZqVQdMkLk46Nh7fgP9X/gEQxjv8KTkwmvU2VWEO192JvRiVrtIVoZJsNo
dsqN5LP2MzvyOFFTRg6Z1F8KABeEmOXAmG+Ad6YW+Tztf4KzqU5aAk4H/OaPiGfL
CJvfAh3K5WMDyIfhSy+VgKJOlwOnzYIFwwiH+Q9iUe6GaGuoLKI0GBFKiliBJ3Ek
szarJt66vGyt2FzTeTLMvnOn2wauFor6Xsroxi2pErdMWxG/LIy1RBll4SgE6DGL
29eQ0RupVIPA63//D21yRw4f7Kx6w3xeuN5l2c60gzneNz0ZmmXUcPGb9Ekz2HCt
tsGi1AY/kU6kcxzvf05OkFozGW7BXTPES/zkQud0cmuFRF5DQ0ldF2JFMa9E3I1B
Q0ejabBOaBbw5XzoRDAYPGR9gca8cvqIryVp6ZwEGCDl6z7x2XHumczqUSZjTQuK
tTJx4+jbDeBjgQBw8vOTC27mpwcv++Tsxec4PZX7NbA=
`protect END_PROTECTED
