`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6RUk3fOSQHLDtwJh3qImKzjuEnCm7QsGFEzCiO9iBIf4Nj24qo7dWDdomjvPoGh3
vbfPps7aOW85HAlWimf7fUpL/5Nog1vt2f1JgKgWtXZQTVl6syewg78/UBMsYmQc
Jh/JWpyETqQ8lMIZelWqXEdNj2fjz+0LNZOJ4RXajlUwj3UAB74pJoTY6RVMRaC/
EiJfZL6GAf8Gtil787alQhfjcI3voLqI4sOlAHGG46ELjZXhu3eRLUJGp17GRBIQ
JHVEs/7GH6FTECiHYJ62L5DHVIatV6LdjAB9dFFcQ2JO3OVWuxejC1SKczuRKiiM
b9KY5DDBXHQV51Nu7gOTUTk1MsVIHTQwRZfJpmAHpwUNq+kExtE6aBREVg4qfhQ0
0o9w2RHIhOGb+j8upJrf1wl7znhcyTvYFQaQEm89SsyNUwcqKx5DDgiQO897SZc3
ZGz0ZdL5cqbQmiMn+t+3o8Pf082jQuLFK0dzyR1+4I0f3PLpW/q1VVcNDEiDAT3Z
n2SRIptYpDTavRB14aLQV+ah0B1lY9TxGwkPPo3xr/RlD/kxl7xrvYpCjeCBDJWr
xXVzovxnLp48fbctfP1KkN1IlgLZU4paIcFg6CwQGa/yRArZxVWOgRfECXwih/23
2GrwuclcqB92E3l0L5rwwOLBbo+ZL0WpiPD75Oq3VvfGm7b7Qx4iF3l5A7D+oWyH
jLiKYePtPujN61P+7Wyz8sZHutHHHhtznOkdTLSajOfPAZpcKHQAhUcx0lo/+LBr
uKkNubp2ceNnAn9rgea3rzU1LPOhM+xqbvdNPsL67KOqNK6Wwl8lZ0bi8XXXc38l
6k9TzIpy+/ds/fzDRh48lbPJFvNQGhr4Mel5PVddN9XUMhTMlh4CsXvWS5KlGC9L
iFU8pEYnTjVA0ehz1sYJb9I2BHeov+qfyTqmlQCofeVig64Z7ikJG4wSlAPPOyLq
Ymu3NJZ+nrvInxp2IrvxI5LTtQwZ3QiMTwtcA3VLxWVOiEsdGRE+XFW8YVBe8Hol
DjYCOJNFQWV6dOA+MpDFTFA0HK6xOzvdXNO37FSl3Q40VwwXMDUzsApgHSU3Rd7k
Bt70Cska6Bbr00mAH9DAc787qIyoqyhFzjnIup7y1tID5VrZxHXoH/309JJ8WhvJ
YJqdyZ34j4MhxkRHm+A+W7lw5YN0w4K7MNxYwFrr5NDn8czFqUoItWt7ZEZmmUdk
4+yGSl77KGk2DG9eXxNGSnwvasUgzYfUGjq8N/QEeuzMStgEnpvwlm8TIxZ2O1jS
Xbi5hNMVb7kQhyHKDN5Lkso8ynLpuCB1p4/C8g0SJfZbhSaGKVsCMPaEIrf8se1Z
`protect END_PROTECTED
