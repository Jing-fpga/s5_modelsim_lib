`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nA1MtXUqYEB85L6WgekG06Ky+vZE99WSiVHWh7zv4pkTkoQ8v7BcewVf3pmpf1bU
zSCAiGcsidkVzpEppi8J3MQsHSMCWvv8LPWoEMUsi4IbvPYhkvU+iDc4LrAa1FVG
s75c+5TGmss8XLB4q5Kc+oYb6QEi8Vl75DvS4AWms/F37Dbnztg6pP6sJsN5iJVH
o/1Aaz9Ni96aorHP0+XuPuA6M1RSDDI7Tn/K//SHLiCgEWKWP9I+sdVzVPZ7TAzw
7zqjwh04fTJUb4UpENzbAB5u4Zw/DXE6kZXEPnCVq0aoHboyLPh2DtSSQt7T5oHJ
aY8zb45nqkugwixiXjdxzbP3onwiL/ifI8F34X/IhYvBqLyILgrgXLxQSAfxzCJT
0eSUmt/CyivJMOkD0X4X3XQU28uevxhThklLKP8vZ1GHYPcjr1upYAZm9ZzKbx4W
m9xu+/bHY5xGl6ol1Mmdl1cBAl6UwbxSftUQwO0j8+WuMYMo3VOnLiBfp9pbE8ps
nMMKS2Oej0Jx20v3rB5hspwPKz9HA8hrcnZljvQEx13SKw/sO++K5PFXnO69fHBy
RE++mNfVYJhc/+yoaSH9mD/9H6KxbpIWnaCFOlbctYEYa5XAbsNMkCSFPZNe3RUC
wEkXn0pZNzpwUyPCNUQ81JHqfDGbcbFegwtULylshHjaKrd6TsKq7uF3KXDq/ebr
pr1qf/W/s/yf8DdQZh+mZWIldh52MwvFWjrq+GxoBxgpiY2uNUUWOnVSQOtbyGVD
YefP3B8GvD1b/eYygxGpWrdj58WnzQ03mTNkwBCZ/IleLxvkeDgaC5QRIPP9CTaQ
1MntW26na4cfxmP4wB1a66ivjmm1zpl85d9wnjJfnIi0isjaaVI9ZVReKa2ayVDz
mQgVYNAog+5dDmyzzUQZuDCRlzdM4b2VweKSJl+rJ2tBCJHeQB9sCLoGHVwcBSq2
u3tOQOEq6V83zJ8qSdNnDLwlYdBhZ9/ZTv7JND7E0vJGPMy3VfjbMwK+y2ZujiP/
AV+427Z+PxjSYdKySDU1LrW/YGB2s0nFd9px1JV/v/jOkNn9W1YjyMAFLAT3Ad+V
J6SknQSDiA+PudByoXIxeSW9H2tAsGIk8zWymBZVcIDxD1l9F82mGeWOlURVBXpP
BGFaVHmikZRUOe3I5UwYp2jh/RzyuUyHRuB3OCwoWf/6vdtFReNXn9XWcrXOxcjy
hI6NAJqXQHDlp8rCquWOdFmiePD0dhJiJ2XaEyA8dzOpg8SC6PTmkxGWsEj3yDHc
GnVEGnKOn64SeTx+cp2mSAS/oPfpgOLgzhTe95B5Ho3SrjB4NOLUZOMz1hoM6mqd
vDPtnWoPcM4hfWfb+NRTtRVXVdd0l9PAjJH6VAECLmwk1KEbfbEI4Kq/CTpw1IzE
PkomUpC8rPdPjaRpqqNs0EA7eedCqGN6w5q8vtC45ybR5YY/Zk2QympguBr/Rp4c
ADd2GtHz8p0GC5rGfWMYSQ==
`protect END_PROTECTED
