`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aeR0CDAK5UzNVa847gK9Z5jBjUSbczCFvuUTDxkPP84o6sdLFtx1ZHs2yt1u2zsO
xLsvX77rSTPRT2GEaVv6Kg6rqNy7arqAigtoQQiyPuC1wVeotVXOvhXUnjrSc35O
5r2eslJTV/uhi5wKQZj+kl7Yhwg2dnXj0bPHFfcv8+eomazd0eHw2ZaWUpk0E40i
j5hCJGTdcsgkaeF3ycZC+3743iy0QEL8Z6dxHGyZEtakZozNjz6orrqlfgZF8KD+
tBibHEnUiVUgGP6ixGsDBweNfnmNYOBf190g2go8C3H0Dwiii3jW/35CL3C/CYaH
P3xWo6kgyagAENHIieDQM9EpUqrvPZtk6XziYrw3zz4YM0AlMm0dmKm1H8Tyr3iK
3iS9pxkCxRvFjDrcb24smyLhwHW80xLk7sP6wmp8CSRGl305tIrTylYxgf7sjwZ/
2mkRji6Ee+qmOuIguz7H4dGTR543bxjocyjl1x5s9MNw7HsHWQck6xKFnU1eAcKy
6OICLcYjb53qucnOZIoZfWNZrKcA0OBlTDI+2hdQ+NgiWgswOhm5liCS4yjP4Ntg
XjWcRuEb4aifg+OgT/jrmIEtUUpqiwUY+Fq+oOK3g8UX+hBt0H63lJEFUnl7fI8X
QQg0ml9G5C2YdBAZ5p7BlOoxxEDp+cAColE2kGXPGKRkVGpvuohyMBQKrnt9IT5q
yqfi52d3Tm0M0v6RB6aDWKLwWxnoZMBpB+TEFBKyjtJq02UYqWPavWI6glB+Bb+4
`protect END_PROTECTED
