`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Coif+fydMINLm67ABNKduH99kDz6hXY6izUIrJWotoRNWo5aWpjRHxIkYVmyLsHC
g27TkWkhLiKk39j8BCS2baWM6jLohLZ3CIjjxlof0F7D+wr0irNomjeSC/2sVFvT
8hLJgusVurNFCLbYSo1JF8vCnT58GWZLnLZK/mBJsA3yXQgMCzztGeLxVwN2fGIg
8W6EfkmBry22Ge8BnuvjlUDnY8EO1Fea5+JPYsVp9mbr6JhL4c4J8EANUWxHL0yv
JjEzDPrXdHeNRfkNXldHL4lX/sh9pcmT/So74Et/IQ+Bm4fUWWjRucttHEpE5a07
C7PWT1vayEI+mt/E/B9BWZMV/SHLFVZFpmLkal83JnN3k0nUGC+W1YR8V59jK+ik
5hbvDRlGmJsbDeaiTALN+1IoHaI/0vt0PfnI36zKCepecuaozj9PgCQj5LRQoRb+
oCv8uY1RPXdvXPE00ldOrjmzm4+KzmU1Hwt5ant+2J7Z2LpENbNHM0SrAzSTY73S
DO6uDQbqWflRwR9RqikNSrihn2Tak2UMh1leKLgSzi25mYVh+XG+KEXfHHWMDzaj
oUmY4FFVbWjk9l0JgQhAsJw3WPgInNHxcr0lsqFwBWj+CR9kAoB4laHrM0TwWz8Q
hKlEtnpqrElPcn1gOFJj+A==
`protect END_PROTECTED
