`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jM9e/lgy0Md6tUitzc8xHyFfvVayc9J9feDhiY8S1TGJ9Rc3P0ebB5zVr9N3PSWI
hpONWCidKZrEcBQhjpgWOhIklMYTred1a+O01QpasOpdGEnvRna21fOsiMXv69oK
KPTbQbIc/BoW3qNCnEYM8ndYrSP8ToiYnalb49COHy02qsRm2sIvVr28BEJo7+mM
Zx6TWrTRJ/xuSwHPj6Pvo1oCeRFngp/xEp8Ao8v8hZgfs5mDWgtbOtrUPvMwfJRg
PkHKW3Wt1ONeJNsa3ZZoFxuyLsfg3+4Nk0zu7/rvRPL4wYYHrn60NOgB4Tq3OyBz
m2wAVE4G87m1z/UW2uWO5kB/yavX3AUkc6oYxHOdfo3zAAxuUhObiSwt+w4IrR+c
3Y+27cxMzKHu1G0+Hxt57RlQynI4RtdnNUB/3/9ZSs/jgz58hINGewq2gZh501WF
vaSIbf+ECm4OXW/+Dk0QJ2nS/P9BZrqSgT7s/Icdjf+bmQEiwseH83L6r2RW+OUh
Yne6aOVdyGUDQU+kJ6WFSU5aKuX8njwsduFoXFjkXGRyQvV9mGR8OTmPTxjmoMaL
coZmISFX1LbjnzJkwPQvPBWjzfOZPPKmQy3OUXI5Onn1fNkmhQI5ooaRAuklV1MS
lvYNq1gJ+3MyNz5+s6Ro02gJMOgoWRNdkDQgsSwZW4WVkgOJy+h5cQKYGsQg5z99
JjxxviH7q6tWU1PZe8kCQHnWW7sHAQOgZgfntxF0BKE1oDgfjQqHPx0JueOEzjFY
+7sSTccEyNDllTeXvGvt5jwHlFQRcCMWoIp3OA679867BvyvVow/gAtkym7RcVrV
rmQvWv9NpVn1qB6OnnR9HfHl9HtUXG3LPbqUun9XwlHBQp5PccFQXcwIY1Kj9EZV
7W3ns/TOc5atqMuSlqClf6MAay/t2ttaJyaa/GvhYCB5Z6HY3inibx7NRlyqTFWb
7YFBcBCTM3a1SoNjLCUF2IWbHsl24s+xuBXWfp4T24XXS87O0GxO0PEufdTn/+pp
j6jibpZSZ3QBUwrdLjDtCZA+FQYxMjo28xN3m8KZOvM0fnR4CK9Ox6KmashkigwA
Re/cxYpBsk2m9XppcRi370sZpLLDme0Dv4viHxcXZtUXGpiLcXeZXzWw9iur4UPF
hoV8Afnk+i3VT1uuZ/J9KaZ7Nx5kV+BhmgbR2KvCqPn34fY9H1UyzHe+K/OflaT/
E80CXHswHe08ME7QI/xyEgwmfASgVbpzqcUXI6PJv7/QgzVuz9fPGA6vwIxDfRMk
yo6RF2rVFHbqojWYNiXJ1OFH05qKcww4dWl0f2CDxjZt3J5K/xsA4ynqTLUlX2+y
7f+mnNAofjbsQzrIop7XekzUAQ6RcMKewxIyqC5/SJOkIaP7lK1Uwt22DbQC8lO1
OuJGVbOLHTQqfbfTeyj+ckhzz4bPthHKYs78zz2W4uJwoLlOOnRyAtFoSD5ujb60
gzVw30yJPQvyxtRfmZw7vYDW2Xmip8ZfwgTTdmnBSnbXv+WxVM62cheINfecUvnr
fJ0RTiIQlo6T5wh6V27gXZJvu+DDbZ5AIZPihpt+3sNzGFUhKtfm/nr2UXbY/sD3
xAeVWKvcAQfDNsCTr3AukCK+Mle4FOUIrza7k3Ya77Q+w9r1T8z97qtQVsldvZog
kZg9ydqhR7WYREc0bosw5ow8tKDT4XDu1N6tNJoxZZin5mRpldFXNMd7q0jlkz8m
wl9s/QWzuvb/cgxpes10fA==
`protect END_PROTECTED
