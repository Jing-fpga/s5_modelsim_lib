`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f9vcalaChvjgger9a5TkIZmoIDCFmWbDmBN9mLczwrCs4f3Q0TwqhR6B5cLbIqul
2iFKD03AQrb9eqzFFU597Jy95kYPwprcf1Db7xN3T5YugbxdaCegx0OJJu45/kca
mf/VEF3S8viUEmJ3TO71IZe51/6QWIHMZG6gynEnfv9fkGragHEKmOXiN0guxQFU
B+A3OQE9iFEk/oeLSrdmmFUTjf3muG9GE4gR8wQiK4NgKCFnb8hwnVGiTr7yvz3T
5XvkZRhEsFu/lHBy7TUPNjRHNssBTGDSbHQyNVaCxIsrPZI5LuE62QTptFS1ZIXx
x0q+hVM3SNQrnMA/2aJC1a4GdY/tyuEujgyOSfW7uKCSMhjF+cIHuH0tlJcgP0N+
S6GDBk3m1fssdHBLCuTgxXNytnSddpz1kk25qoL7RhQ8EQLbJCyaJS1t0CsTbz5w
`protect END_PROTECTED
