library verilog;
use verilog.vl_types.all;
entity stratixv_hssi_pipe_gen3 is
    generic(
        ph_fifo_reg_mode: string  := "phfifo_reg_mode_dis";
        phfifo_flush_wait_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bypass_rx_preset_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        mode            : string  := "pipe_g1";
        test_out_sel    : string  := "disable";
        asn_enable      : string  := "dis_asn";
        ctrl_plane_bonding: string  := "individual";
        cp_dwn_mstr     : string  := "false";
        rxvalid_mask    : string  := "rxvalid_mask_en";
        elecidle_delay_g3_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        phy_status_delay_g3_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        bypass_rx_detection_enable: string  := "false";
        wait_send_syncp_fbkp_data: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0);
        user_base_address: integer := 0;
        wait_pipe_synchronizing: string  := "wait_pipe_sync";
        asn_clk_enable  : string  := "false";
        pma_done_counter: string  := "pma_done_count";
        inf_ei_enable   : string  := "dis_inf_ei";
        cid_enable      : string  := "en_cid_mode";
        phy_status_delay_g12: string  := "phy_status_delay_g12";
        pc_en_counter_data: vl_logic_vector(0 to 6) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1);
        data_mask_count : string  := "data_mask_count";
        data_mask_count_val: vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bypass_tx_coefficent_enable: string  := "false";
        wait_clk_on_off_timer_data: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        pc_rst_counter  : string  := "pc_rst_count";
        phystatus_rst_toggle_g12: string  := "dis_phystatus_rst_toggle";
        wait_send_syncp_fbkp: string  := "wait_send_syncp_fbkp";
        elecidle_delay_g3: string  := "elecidle_delay_g3";
        sigdet_wait_counter_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        cp_up_mstr      : string  := "false";
        pma_done_counter_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        test_mode_timers: string  := "dis_test_mode_timers";
        pc_rst_counter_data: vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi1, Hi1);
        cdr_control     : string  := "en_cdr_ctrl";
        phy_status_delay_g3: string  := "phy_status_delay_g3";
        bypass_rx_preset: string  := "rx_preset_bypass";
        bypass_tx_coefficent_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bypass_pma_sw_done: string  := "false";
        bypass_send_syncp_fbkp: string  := "false";
        avmm_group_channel_index: integer := 0;
        sup_mode        : string  := "user_mode";
        wait_pipe_synchronizing_data: vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi1, Hi1);
        phy_status_delay_g12_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        free_run_clk_enable: string  := "true";
        phystatus_rst_toggle_g3: string  := "dis_phystatus_rst_toggle_g3";
        ind_error_reporting: string  := "dis_ind_error_reporting";
        cp_cons_sel     : string  := "cp_cons_default";
        bypass_tx_coefficent: string  := "tx_coeff_bypass";
        phfifo_flush_wait: string  := "phfifo_flush_wait";
        sigdet_wait_counter: string  := "sigdet_wait_counter";
        use_default_base_address: string  := "true";
        pc_en_counter   : string  := "pc_en_count";
        rate_match_pad_insertion: string  := "dis_rm_fifo_pad_ins";
        pipe_clk_sel    : string  := "func_clk";
        wait_clk_on_off_timer: string  := "wait_clk_on_off_timer";
        bypass_rx_preset_enable: string  := "false";
        spd_chnge_g2_sel: string  := "false";
        parity_chk_ts1  : string  := "en_ts1_parity_chk";
        silicon_rev     : string  := "reve"
    );
    port(
        avmmaddress     : in     vl_logic_vector(10 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        blkalgndint     : in     vl_logic_vector(0 downto 0);
        blockselect     : out    vl_logic_vector(0 downto 0);
        bundlingindown  : in     vl_logic_vector(10 downto 0);
        bundlinginup    : in     vl_logic_vector(10 downto 0);
        bundlingoutdown : out    vl_logic_vector(10 downto 0);
        bundlingoutup   : out    vl_logic_vector(10 downto 0);
        clkcompdeleteint: in     vl_logic_vector(0 downto 0);
        clkcompinsertint: in     vl_logic_vector(0 downto 0);
        clkcompoverflint: in     vl_logic_vector(0 downto 0);
        clkcompundflint : in     vl_logic_vector(0 downto 0);
        currentcoeff    : in     vl_logic_vector(17 downto 0);
        currentrxpreset : in     vl_logic_vector(2 downto 0);
        dispcbyte       : out    vl_logic_vector(0 downto 0);
        eidetint        : in     vl_logic_vector(0 downto 0);
        eidleinfersel   : in     vl_logic_vector(2 downto 0);
        eipartialdetint : in     vl_logic_vector(0 downto 0);
        errdecodeint    : in     vl_logic_vector(0 downto 0);
        errencodeint    : in     vl_logic_vector(0 downto 0);
        gen3clksel      : out    vl_logic_vector(0 downto 0);
        gen3datasel     : out    vl_logic_vector(0 downto 0);
        hardresetn      : in     vl_logic_vector(0 downto 0);
        idetint         : in     vl_logic_vector(0 downto 0);
        inferredrxvalidint: out    vl_logic_vector(0 downto 0);
        masktxpll       : out    vl_logic_vector(0 downto 0);
        pcsrst          : out    vl_logic_vector(0 downto 0);
        phystatus       : out    vl_logic_vector(0 downto 0);
        pldltr          : in     vl_logic_vector(0 downto 0);
        pllfixedclk     : in     vl_logic_vector(0 downto 0);
        pmacurrentcoeff : out    vl_logic_vector(17 downto 0);
        pmacurrentrxpreset: out    vl_logic_vector(2 downto 0);
        pmaearlyeios    : out    vl_logic_vector(0 downto 0);
        pmaltr          : out    vl_logic_vector(0 downto 0);
        pmapcieswdone   : in     vl_logic_vector(1 downto 0);
        pmapcieswitch   : out    vl_logic_vector(1 downto 0);
        pmarxdetectvalid: in     vl_logic_vector(0 downto 0);
        pmarxdetpd      : out    vl_logic_vector(0 downto 0);
        pmarxfound      : in     vl_logic_vector(0 downto 0);
        pmasignaldet    : in     vl_logic_vector(0 downto 0);
        pmatxdeemph     : out    vl_logic_vector(0 downto 0);
        pmatxdetectrx   : out    vl_logic_vector(0 downto 0);
        pmatxelecidle   : out    vl_logic_vector(0 downto 0);
        pmatxmargin     : out    vl_logic_vector(2 downto 0);
        pmatxswing      : out    vl_logic_vector(0 downto 0);
        powerdown       : in     vl_logic_vector(1 downto 0);
        ppmcntrst8gpcsout: out    vl_logic_vector(0 downto 0);
        ppmeidleexit    : out    vl_logic_vector(0 downto 0);
        rate            : in     vl_logic_vector(1 downto 0);
        rcvdclk         : in     vl_logic_vector(0 downto 0);
        rcvlfsrchkint   : in     vl_logic_vector(0 downto 0);
        resetpcprts     : out    vl_logic_vector(0 downto 0);
        revlpbk8gpcsout : out    vl_logic_vector(0 downto 0);
        revlpbkint      : out    vl_logic_vector(0 downto 0);
        rrxdigclksel    : in     vl_logic_vector(0 downto 0);
        rrxgen3capen    : in     vl_logic_vector(0 downto 0);
        rtxdigclksel    : in     vl_logic_vector(0 downto 0);
        rtxgen3capen    : in     vl_logic_vector(0 downto 0);
        rxblkstart      : out    vl_logic_vector(3 downto 0);
        rxblkstartint   : in     vl_logic_vector(0 downto 0);
        rxd8gpcsin      : in     vl_logic_vector(63 downto 0);
        rxd8gpcsout     : out    vl_logic_vector(63 downto 0);
        rxdataint       : in     vl_logic_vector(31 downto 0);
        rxdatakint      : in     vl_logic_vector(3 downto 0);
        rxdataskip      : out    vl_logic_vector(3 downto 0);
        rxdataskipint   : in     vl_logic_vector(0 downto 0);
        rxelecidle      : out    vl_logic_vector(0 downto 0);
        rxelecidle8gpcsin: in     vl_logic_vector(0 downto 0);
        rxpolarity      : in     vl_logic_vector(0 downto 0);
        rxpolarity8gpcsout: out    vl_logic_vector(0 downto 0);
        rxpolarityint   : out    vl_logic_vector(0 downto 0);
        rxrstn          : in     vl_logic_vector(0 downto 0);
        rxstatus        : out    vl_logic_vector(2 downto 0);
        rxsynchdr       : out    vl_logic_vector(1 downto 0);
        rxsynchdrint    : in     vl_logic_vector(1 downto 0);
        rxtestout       : in     vl_logic_vector(19 downto 0);
        rxupdatefc      : in     vl_logic_vector(0 downto 0);
        rxvalid         : out    vl_logic_vector(0 downto 0);
        scanmoden       : in     vl_logic_vector(0 downto 0);
        shutdownclk     : out    vl_logic_vector(0 downto 0);
        speedchangeg2   : in     vl_logic_vector(0 downto 0);
        testinfei       : out    vl_logic_vector(18 downto 0);
        testout         : out    vl_logic_vector(19 downto 0);
        txblkstart      : in     vl_logic_vector(0 downto 0);
        txblkstartint   : out    vl_logic_vector(0 downto 0);
        txcompliance    : in     vl_logic_vector(0 downto 0);
        txdata          : in     vl_logic_vector(31 downto 0);
        txdataint       : out    vl_logic_vector(31 downto 0);
        txdatak         : in     vl_logic_vector(3 downto 0);
        txdatakint      : out    vl_logic_vector(3 downto 0);
        txdataskip      : in     vl_logic_vector(0 downto 0);
        txdataskipint   : out    vl_logic_vector(0 downto 0);
        txdeemph        : in     vl_logic_vector(0 downto 0);
        txdetectrxloopback: in     vl_logic_vector(0 downto 0);
        txelecidle      : in     vl_logic_vector(0 downto 0);
        txmargin        : in     vl_logic_vector(2 downto 0);
        txpmaclk        : in     vl_logic_vector(0 downto 0);
        txpmasyncp      : out    vl_logic_vector(0 downto 0);
        txpmasyncphip   : in     vl_logic_vector(0 downto 0);
        txrstn          : in     vl_logic_vector(0 downto 0);
        txswing         : in     vl_logic_vector(0 downto 0);
        txsynchdr       : in     vl_logic_vector(1 downto 0);
        txsynchdrint    : out    vl_logic_vector(1 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of ph_fifo_reg_mode : constant is 1;
    attribute mti_svvh_generic_type of phfifo_flush_wait_data : constant is 1;
    attribute mti_svvh_generic_type of bypass_rx_preset_data : constant is 1;
    attribute mti_svvh_generic_type of mode : constant is 1;
    attribute mti_svvh_generic_type of test_out_sel : constant is 1;
    attribute mti_svvh_generic_type of asn_enable : constant is 1;
    attribute mti_svvh_generic_type of ctrl_plane_bonding : constant is 1;
    attribute mti_svvh_generic_type of cp_dwn_mstr : constant is 1;
    attribute mti_svvh_generic_type of rxvalid_mask : constant is 1;
    attribute mti_svvh_generic_type of elecidle_delay_g3_data : constant is 1;
    attribute mti_svvh_generic_type of phy_status_delay_g3_data : constant is 1;
    attribute mti_svvh_generic_type of bypass_rx_detection_enable : constant is 1;
    attribute mti_svvh_generic_type of wait_send_syncp_fbkp_data : constant is 1;
    attribute mti_svvh_generic_type of user_base_address : constant is 1;
    attribute mti_svvh_generic_type of wait_pipe_synchronizing : constant is 1;
    attribute mti_svvh_generic_type of asn_clk_enable : constant is 1;
    attribute mti_svvh_generic_type of pma_done_counter : constant is 1;
    attribute mti_svvh_generic_type of inf_ei_enable : constant is 1;
    attribute mti_svvh_generic_type of cid_enable : constant is 1;
    attribute mti_svvh_generic_type of phy_status_delay_g12 : constant is 1;
    attribute mti_svvh_generic_type of pc_en_counter_data : constant is 1;
    attribute mti_svvh_generic_type of data_mask_count : constant is 1;
    attribute mti_svvh_generic_type of data_mask_count_val : constant is 1;
    attribute mti_svvh_generic_type of bypass_tx_coefficent_enable : constant is 1;
    attribute mti_svvh_generic_type of wait_clk_on_off_timer_data : constant is 1;
    attribute mti_svvh_generic_type of pc_rst_counter : constant is 1;
    attribute mti_svvh_generic_type of phystatus_rst_toggle_g12 : constant is 1;
    attribute mti_svvh_generic_type of wait_send_syncp_fbkp : constant is 1;
    attribute mti_svvh_generic_type of elecidle_delay_g3 : constant is 1;
    attribute mti_svvh_generic_type of sigdet_wait_counter_data : constant is 1;
    attribute mti_svvh_generic_type of cp_up_mstr : constant is 1;
    attribute mti_svvh_generic_type of pma_done_counter_data : constant is 1;
    attribute mti_svvh_generic_type of test_mode_timers : constant is 1;
    attribute mti_svvh_generic_type of pc_rst_counter_data : constant is 1;
    attribute mti_svvh_generic_type of cdr_control : constant is 1;
    attribute mti_svvh_generic_type of phy_status_delay_g3 : constant is 1;
    attribute mti_svvh_generic_type of bypass_rx_preset : constant is 1;
    attribute mti_svvh_generic_type of bypass_tx_coefficent_data : constant is 1;
    attribute mti_svvh_generic_type of bypass_pma_sw_done : constant is 1;
    attribute mti_svvh_generic_type of bypass_send_syncp_fbkp : constant is 1;
    attribute mti_svvh_generic_type of avmm_group_channel_index : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of wait_pipe_synchronizing_data : constant is 1;
    attribute mti_svvh_generic_type of phy_status_delay_g12_data : constant is 1;
    attribute mti_svvh_generic_type of free_run_clk_enable : constant is 1;
    attribute mti_svvh_generic_type of phystatus_rst_toggle_g3 : constant is 1;
    attribute mti_svvh_generic_type of ind_error_reporting : constant is 1;
    attribute mti_svvh_generic_type of cp_cons_sel : constant is 1;
    attribute mti_svvh_generic_type of bypass_tx_coefficent : constant is 1;
    attribute mti_svvh_generic_type of phfifo_flush_wait : constant is 1;
    attribute mti_svvh_generic_type of sigdet_wait_counter : constant is 1;
    attribute mti_svvh_generic_type of use_default_base_address : constant is 1;
    attribute mti_svvh_generic_type of pc_en_counter : constant is 1;
    attribute mti_svvh_generic_type of rate_match_pad_insertion : constant is 1;
    attribute mti_svvh_generic_type of pipe_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of wait_clk_on_off_timer : constant is 1;
    attribute mti_svvh_generic_type of bypass_rx_preset_enable : constant is 1;
    attribute mti_svvh_generic_type of spd_chnge_g2_sel : constant is 1;
    attribute mti_svvh_generic_type of parity_chk_ts1 : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
end stratixv_hssi_pipe_gen3;
