`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r9N5ZbXKzYhffNV8mvwNa9O+wi3k8UL0eZUaxEnhgIm+Hd+WbozSwr6mF7c/ikYv
y/lcAoadJzO+Unaur0pcdeO76R/3Tm3P9x4BL8AthE2zj2dT1JhxMg9+75iwn3AP
WvHRMdQ5KrnoM8yMu1ioKn37yfajn6GRI5eSys1srWZPhZcR54hQ9jrCElrgMw4+
IJyO8PPZJZSiyuQNU0f8OsEhEF+bFrXWecYRDUE6GZfhCPNpSgnhcKgzG/eVbl52
o/ZFHHS1FN6zPQMTY3+Xd0rEzGQvp83QhoqnW1Rdnf7oAff+1AXzBWExo036qll4
CW5VJ1h6oCPOnsaw9/W3OhXp4WpCTUyKOPuRhtMksMVOpkWzP3x21QWz9wDADR1v
sLWJiKNStx94qQ13RA4HvlS0VfYqlGBcf5OmKOkkIYBM4Skyz7BHetHVSKhv7Th2
RnYEJTsdmAe3KA88ULA71Rm7b/qob0tDWHTKTK2EBQTpMkpRwgMA0bRc1+vuHAMh
LUWgHpsZT5Xttr8DZJun06oiKmVKL/ER0Qx3JX0SubtPv/hAm4POfD1ACTF5j4FY
66nDAoAusV7+S1bkktiD2/cMo9PbWJJ3NxxEdyXm57GkZlLO0B6xOBy696VhMDw0
fPVifrHXEgmtbIDLYtZo9CLxzpeOqmwySYbbuKHViPJkzqaP+CB7txA0VKTjZCxh
M9NVxlAPtpjPDg0KlLgnuBdmnc+LvP1cEsk5IOYFW82rIhvCV1ih1qKB5s5SvfJ2
07Mu165JMjUw4kcHX9XYISVHXS/my9G4z4AJMnKafZ3ryvxuaMRSqV44Q7TfOqpb
Emie0acFWm57a7aZopNNjNPyS4ftZHqfTxw+n1PySinKGcfk6gJ/yBJHJMz2Q/RH
7KjJEG4evdmDMprhp+qEmTzNE+MueqjmL7gndDrs2iQVXWpAeaaPOLH0XzDQlPdj
mpzQG/vD5TMy6QPmSbIZ5JABTmzuS3nPglwPgoD8sLGvGng7QDd9B66tEAjmLqPm
PDZzae4/bglDTX7Waws1eYssbTJEGGcf726T9Yx/LX0M0QtK43vCwBc6W1vdJ+Fn
8VrWysSalcUp09J1/qwEXc1avtAI6iYTxnus4NG4KHuffaPmNDameOlH3YN/G18r
q7yVgUFUhogMS5Zwgcnzx6SXMFe/4YfU73AMLx9h2t/zs0NHVjGF7EHasLb4Y+cm
DpjdTfHJsCsMBoVLj6VG4d3yMJRjLKgpZ1U1VvledmP3Y2nh8OwQJHZ5zytzI0AK
vtd/g2+4W24OCtFc7v4IFyNHdAJ7qvbSfcFpi3Im7w/3lHsQ70sHhbxxBM8wFjZc
c/awkLxjpjr71AXdiTtho/EsG4LWCRX89mVZt9UCfKx8yHeXmpXPvqI9LkzAJihS
5PLRuXDQVLyX+swRlkd0ocWKTCFfp6ROiTFcemf2T6h0YW3TP42EA9/rZn9KWyyb
XmqQdpIl2D5Hvc6aurLLrmnS71SKdIMak92haRP9fqaKizobcMpi2+51o9kNP4VM
5Jt5RSbzkEd/9u2sMpkUzjbTAOQviz7KyDFYbutvYdpGxMPnkADIY6szubJCwis2
6CODS/9JDzrQoxns8d4/t0wAk+67PTE+bdvxtbRMNKqTfIU7fl13Ko24H/EEbcRY
AZqwR4yY47fj6KbW0z4mWVAvVyE0prMzieg6cFgTFTwVlhHKOpArgxrQ0Y0Yej+J
vb7ke8h6fcN17qlc4+UpaU6019iEGpRYtX0rMMBow4/GAV6JTC1k/3XTtxlyvAWX
OdWBcTpvsWJfH0wAiDWUhuvHcYJR72nS3VU9KiagEl+PQoLQ6sQF9DZZTtOJwG1s
DVTjCtUOORJt8EqqqmmrAQ0VyKyVLjbMPcIGF/BgovdqHlIMTEqgFFBfiY1MUvuW
eeztDJdBDOgQEEOHArduN3EuU2EJ4T+xF4ur3+Pymzov0SXg5M6kgpctNHQoWP62
jALhQpFXFsk9tZQwnjH+Meo5H0L9/li/S+S38VPDczNLwY9yb3WU5ZSeLUg5id9c
r7/dpj6ZL+8YKjYaWUwxiy4iiVMV5SMRo+QIv0Z1JUq4gpnSXlnqzZh1qeFHOPqI
g65rkCwGXI/4mDDsy7qDPOkFdYHzNdmlOw55pGAWJgksR6YLRvBcBdCw0gfvu/Kw
HpKxqvPlwjGMjOUbV5bDuOCo1+WLJ38S0n13wnxmtv2gZc4Pzhka6ZB0r3wdXDpC
iELHugYf93bpu8qp44x9S7OLNrfj/ZpuOYOTPpA1K0nDzAsPpSUgFHg7s/8P2kU0
E+DBoER91JldCcrUciPcplmh5fO0QuV4aNILSnzNwARh2SXmsCLhjwk1uecyxmpy
12GLRJj1+mIwY5Dkl6P+3w9v2w06W1lzmvWynorccFJrdc6Ue+/HZbMu5dkazdub
hJn+eSOjEtaWg8S0kHFQs0W8x6W6HJz1tmpclQYVDZd/Sk+p67dIuxYnlpMK1KyU
vLrMC7XBnr5k2BeECZKfmXOpiQesW4mXnfzuOeUlMuz03DQNTzLUZ1qyPSos+/ac
26Up66vb82jOCfXRbP4Py14tfKW+YQLlhRFEFrmBCheKGjRXLePPTPfzYsDgget3
3yYqiwCCQZlpSU5fMA+ejNcaMAewP51EfhmSrvQDmu4pW1y696NV7X0gcImI+zM7
3zXNZ4pGw2h5fujtpa8lMBR/sHdR7+ZOFnCLQuRFkFf5sPSd8tiJXXRQnSZe6ygi
mivY6OgbbBpohw91Gx5FdBLZA8+9wyp2U0yqZE09z86+oxHZLcubkV6VBVVsBdaw
OMJky2OuXhhP7l3Z7wqOsqDVQ2LMGntQX95KI+a5iG4arCYU2zBjqiKljIEI79Tg
duY+lSjHZjcwBew98relwp620NsbOganBJnQ6SFcq1S9B980+p29JagFamNffFLR
8kXE++efxANc083xl4M0NoiOCYC2EHu0J3TFwC3PAupez/NcU57oCcx32StVBGB8
a0b52FYvtzoAhWqmmynfKp+noNDeaRTni4Q2OZzPi4izsmniYY4vmiAiDAgXTvsb
ZEn6qqFG3PCtO3QAbl/NPaslDN4bXfeVTcXr9lfZpJ2zEqktMAswCSyWQ7Xdt/pQ
VxHGPO5zO/dXfZM2YUT6ZiTsxuTLqePuYXQPC3JF8SYHywEIdzvVmeujm542ZRHa
/sZprS0h6jpbNvLOuK7VdON7+bmD0FHUKV5zxso429rjufUZi9cMmA0KLEc/baj+
2oS+ChvCEorxJh2n1scvbWTFZspYb6ZCdXxZ+ed66Vlup4p4ChIp82JCadRk+4Pg
8IYg2cP8Gx1NQ5TX2RAm9xX0L9arxmwscpV1Ank5qlyfzzxK61zcVus7VpAB0Yd0
t49LjGLuvaOTLn12WU94onLumtz8YLV1kLPeuSwxpHVykIovpXVx4Cg9cFbEl5Nd
OKEjjT1TmdCWb2H2hBhRg/JtB5t3MPVjMpOVGrhX9kRl4PN4HzA7ckxtbhLyGqXk
fmSNGXNAP+/FkuCmcqE7NWF+n8lTLSjdN8zv+iNaGop2xzUYfdbq+hnmHv9hggcQ
snwj5m9ZvYLnIqupIncC8ZGtMQsIOMwez6prQq8a6kVgKYKZ7ZYIybAUZcJSLeYL
G2orSsUghdwzxy+UyQLOunhu3GKJJk0X0MBJSSzIk0cgt5x3rkprSgZessxopYHj
QpEClMdwqqjU1mHEpIMw6dtcmxv3wZoDKHoU+hlTCMrYSmDaq6y8Tnpw8ak6zmj1
iECWikVvX8hhwqP+AEgkOj5tUCAyLDV/PxJGssYigJZUckOSmm71zx/BVRBTgV9K
U47Nyy+jXaNzbrUgmL1vVzXil3/qISbyjKIdrS5t3U9iccgv3Ftk0JEr7Sik4Q9U
2OGMwQS+Os8fhc3MxucjUAbaPpTPpJhwR7BbASUbtyhyJ+hOCwnILJYgtXsk6Qhh
abrfQLjrlqfMJ0IKcfTCWvSjRXlIDa6G8DFxIIPj4rOiDowPns/YU77/BDRaKNX9
vlo2LvS59jxvvt4yzEPz6NdlObQQ4xZ8MBAueG/fB7towUQLwerP/95qK5ua+5Yb
13Gp7zHKSiS+qrNUrhUR71K73mztdSmh94P/jr13VBg+8/M+uUQoVnnxNn8oaHdh
+3SsiG2Gb1YiJY9VSI3WDljxjHBIexMQ19bSOQ3Zy9C1NlJfX6HP2pZQ7HVacUc1
xaryHyjjQoQAZZzP5d5htGfyUTPh8p5fBxa0y+5jLGsSSe+2FjYUmyqGSqwm8jCM
j0xLHrR3XaEZ7nwYam3qcBRdW4vaypIwvifuXdFUUyBoTrvhkJMxH5CsQWwXOkbz
kkAvkTJk+i/Ylhi99CmGyRSofgbXay/MMZfnL2duRt9YZZt9HRnFUpPhZuAeWd8i
69IuxdXrY6Kd8ibULat3jQO21ly2SGepOU065ISgBjE+Kzjb7yo6m37Pjuv+7E8q
9brQzhLXL3LWR3ro/UkEB+cNSVoLBznUTwNYpNENjxSjhNjgoTbbwJgiNpSCUyL9
7yiKiyoE2LzC6Ukkf2MgSGVAngPXEU9HguZFKmPlwq3VYQj/Uc24cps8CNqhruEF
mvemt0nUc3bIasFd93JRYZE5K6hRxwBwaWjomyP/6j9MTYj34+woo+VnC+/U4h49
vf44KQadgCHzBIWwRhHA24B8ihJnzjorsu3lDW2BklC9rrwjZdJbqy0AN5A+zGK3
01daOtetRVTMghNtC4IBRAfnQ7dXbIgRoaZzITV3SOAJGTSBtuhd0Tkm+WJEZqlH
BNg86K3n81VZ+2Bfiw97ZvPJNumgBRHI7CNGSNrN+phrbBlIITuEWvpviZwIrz36
7MY8JpnIEjMyujws88xtcWRpazAbL5TCYReFl6921LRIaAHZUhYiG3rwvbFsIL4J
6Tlw8ALhT84MfH319R7Ic6hIqagKJJu8YxLU2o5IiW8r7l4wjn6WeF1hSpj7wne6
DkRiDMzE7GBq3VkWnzn+NztJuzG4moh+zbhFAozT3k3/ZaT5cFs7kSLBB1i4bSDi
+QY4mV9DKTAop51ZMNr7B9koeu+qcmm/eVGj9/RrhKTUCHVkHe7pi/XylAyes9DE
wZtGbIlmujDe2MUdPRjZkRTdKbE3zSWA9RgdLNG2d5ixBb7wmiZXkX2bvKLGHEy9
cRevOEOaz1RXfrTFPwTboG5SgdDnnSZOkfs05fUY4nFKRzOVFO/UQPagNb2tOrqN
EcEhHYSp3PDP1qwTqQkIMQNzB1YseRjzIFtZ6tEI/nSy4YKUB5q4Ea7TdO1gK9FP
v7IyXcLmjfgLPnZFSFDpDmmne9w+IyLcqAukcljhETg2VFVj1vtJLg+JFet4mfvv
y5emDHTOvzmxV2Ij0fRDoXjs6EtbJM4pedLdIQPFQge8zt35iF+GlUrfpbj1SRm5
UDZdy65LwWUAXF8AN4nsIdCuf3IJsQXVTJ5D3znjNW71DGy9VHKwCHYQGJ6qN/Qu
ky6A/PKykWXrMCp8ifUDplWyNUnwK8qyoaICEDTTrUT6cJA/FyeuKcbjHOCMAsTl
net+xtxXYStNcXhjezKiz5E7NVnX2oIj2gDtAszzutj38fNQMlTytCMQFTmyTYId
2oMKCbk7wqNfIPAG/H7QdWPmd+fnqslTowQey0llrEVoBYsslx5kko0JfCAPIooc
BI50LxJ8+ERoVv/0UvDdHrYgdEZHFzZYVih0SXICjoBzknmB9jV7g8itNrtvnnhh
/TM5FYhu9/20sltTZOW+s+WH0FWOnzRKZl7KStVJRSdduydCs2bqhdwEkSM20fxt
VxA0hHKDoOPH45z4D5BPi5E/dsJnVHpD9OjVPMSgY7k7iuwv2AmMSalp4+Ffc5V/
Yhenp3L1b05gy04ORUHL9SBWjtHqMMTPrNdcz5rChd0/wDfOB7+Cml9jDQIGlGm5
EO+ZV1BZxEkn4aloouvGqyqdpFpCWDl7eBS0U0D6Cm9znoizTZVtwZFEat6pptHc
jZ9vlZ1NwA7TpmjOdV6cKiqsUhTZ2CMAiBtEgcZUsdVYtZLsml8thgk0QrE0KjK0
ziCqDoMOf45GJsrxgOkbdy7gGMZ8tCoLJcubuYzbMXSWSRLLnRaDliwbwUyzIJJG
LBEJjS+K6Em1xt+J5CnHG/V5Fmg6i7ZpLVIQfS0fSD3pXA2qwMHrmbrwuHI3Udp7
dW7ZbzcoZ10o/VNVO2yLQANH9lyBNusyaqTy1BQ+fK77TN4SQ0SMtDmhOGh2xXD5
D/r6dZ5xVrmEIF8lXp70VD5av2Atxj8yPB0sHF7wpkV48F6tVhLbSNkrEfZ+mlz0
pHVkhQWG4boKQapSN5lERahcAY6OYEu5qMxXuKCI1jZi6uhTDOaohCGsng41fAj+
6r6zi2o7ag+tdbem1WDZX3JxvX+hBwhTvEl0JCAXEPDrxMHViVwvOU0N2415VZ4O
B/aC/X1y7YrPEOC9REDF8caQX5EBDr3ZNyQ8oLMpgVLAuDPyQJzC1A7SIZ7B98dW
/pdfDTbpbvvNAMwszJ1fxqbwjwo9T8yqYxbS4SMgME2g8PnoHK/nqd32zCMwg0d8
KT2efO03njjL6SOUMCm5Dkue/ihCPum79mrLiUrKpJYpNVHm7rKgp3HV5UCZEL7c
Glp7kAkw/beUmmcfIy8l53V7NJFx+l9h+KtwQbzd4lVASfdz9kBhnEelFTerZpTH
L3ulm4FfnqiDcBmVp/zb2ETehBDMSxOgIYWXEXffwUU4nl3hL8FyzDgawvFCNJZl
eldxcshwoNFht+S/o3DzI7Xng+aIlafsgaNXF3H8fuJD2JjAEDOZKawaJk4zceFF
/7QPdhJjjt0L06dnwtuUML7W6zESpik05mKLylk62X58xFjubLfDtdqA+fQUQWzE
rcEruTTFeYefSxzr+6cWpXIhRWiWsFUX3AFKL/vc65IlK5S5jb/cjtRoDJIz4NjZ
pkIlGV+rb1CivC7EWyFiaVQF+nS2/o7bR4kWHopapi7rxxX9r+yqdL+rsT9tS3Tw
oSemjMH8Q8RXFfwDFxrhkx9ot5qMHnlzlTj34vJ+V8tIy+QYgwDfAf/RsfetdUjy
Jdo2r8LVGz/KfPcF89GcI8Y+HE4reoJuzFTFn0jCZMmmO0BcSaY31BY3oyiW4C7p
A5fi9Ad7curCD707/F0c/PC6L9eLwn8Q/RMTIQr4CaK6v0dmE+AsVt/CXB7rWWtb
mnqsJsuWdxPOIa8YX6Ucp3ssJXhldEVlCO9+AtGm7/6/LAaFi1k0zk/ko4W+cXFc
30d5BT+FYWHsTuen6ZwntpZBNEQLs52iBxdGFoedsjwD7lwSEJ+0qwN/5Zt8bSC3
KO5iqLStNteKfBHUjkPkKUMPr2MFLUtpvYn9OJivKQQs5D5thWPLbI+h56wwZPYE
6zWG+IcmZAiDKdZBQmqiG01Jw1G7AexfMEe2Czc3jDbHAQ3+yFiq+ieMWoIwAa+u
y+eZEOfUhQav5W69kya4utp50dW6cYnIfZna2j3qhOnKwgq/VA23MTKCBQXtAUuV
tKeDsxJ4sYeYuM7wRemkbXRRXEJiS9Yzt39rsDhKZQNGx+SAgezX6cF7YMecG2Zd
f3B8ZRefRx5kMazfEc0Jkh+i93nM5I4RCway/ZmYNxmSq1FlB8z7JDYRX6g/HUV/
aJZbHrPUILqeSQKViS0dN5/0WCF9gQbAZq+J6gwrjclhCy1dApwoetuLYpYm73gu
mihGNL8o9nFCXRgwRBdCRSc9VALPb00tRs8AYx1/h1QTtcrj2hW17vFnjzYWzXxU
rj0hNIGyuW2o2gLKEx6u1YK2wwcyU4uYsfsWRlhJ0kf15J8ouFFv+efGhBiwhIuE
wu5XMLfAeYoS08bzZsD8TU8gCQX0ggeDzsEn7lPJtUI8wjkYXAv8ri4yN+qiHJk4
iZSz536Ns+Jd/BNrfVDnRHrzlclCQsSCqRKWYymvA4MzdMBUuxEgpBjaDJKPcHr/
RQOH3Vug1n6G1MB/xrMTteUdsFGaNGrl5mfpgd8GgjW8aCXB0iEqwUHq/Ds1PUv6
CO7bWMosvixlJKgF7WsMhM0nyzXlOgU2TR7ZBxyCsIElzcJvv/6Q7gPV+mY1U3nR
K877ebfTHQGxC7x73V/ygCKVcRcy1a4XEEo5IE5IfxTbSCsJiXBpl3wlSb6jV/pn
yWwnC2HI95ZrrBePGJzBavwyTKqLNbx7dx+gBLRpt6MO35Z5elIA55DhjlgiRgMq
/n0WP1l36N+fkYrgp5goWHOavDjkSKAHb3i/hFznR3+d2DKM34+EPQwLmIUwcEyX
+Tt4J+egvuzgG+7DpAt9JEycuEDJJImAxfosjEBgoP0wCJojI0ezbTr/Mx5D6nRA
fThFOMMLIKIZno3E5NRBOQEx8Eh7IKjzN+KSalTuHOO1sL9M0bedbNrPbfS6hpNs
oCozR0nyHE2Tvomi73T6R//wIiFYiEM+d5VaqAbIlmEYq0qa0dpoQU6je0C0mzIV
dGoo1N1pTOyYLpSfAqSKliWrwFk5w38+6fUwH7BDTNSeUyANLAsHQZzeY/Tyh1Gz
TchW8B+/VktPeR5Z0D83zxnoielYQQ1I1zsR8cbOszbEppgvSHPd5Rl2WzANWFO1
7PhjGXmcJQWgMx7QmI547rM4IwwKR7QGQFvJ3mXs10U9ntE920GvKlGaMpxamW1y
cx/S3xVSbN3+IAhmUVk8r+cCuw9aFSX59g/YJJ4qa9Cp5uQDaOAxHMGx//Ued6+H
K8XjavM0RB8kfrphh2JnA3BIoBMy1RPHyLQVqFL18xM1YbiFTvcnrwS3RZIEWK8n
NYN/zIX80IYSIOfvyN4kWkAFilk+VB6nogSoLXFvDg2mor6xYn9ZeZF8z/oVs0Ci
Rv2u6Yh/UcALEuREtG8ssNARu4xOWS0oyreQazCdIN9TNPu5yQXo0FVcki2yYszp
uVHjfbcPqWhUThDHgJPTul53+huZz4C9pdbNwDG1CpWWBzsXtrPPhggSsDQWptts
NrClo1PK114HQSzXfrGrF632Pt7Y8zLnvLnPI3GhSjzHC9bvYRQnYUl5/Juj/mZa
8n3bnb2D4QmiyqmoCUjv4lcNbFT+kTZHvK5/TBSsW7wq2BLueV79UnOcGYXuOkjz
ogk0+JXSXJXUZ5fbjPnC9wg517b1kyvfcagB7E77ub+ux2gNYznYxwrtY+sliDhq
Lr8Z2kvPS7IgpQ53ioeRDlKOsKl0Gn1ZNd5CzbMZiPFuc0t3V13JYuKQ1ken0obH
U1VGxiAIjBwlATgCTPoszBDjUgW3bbEN+V5bmeaE1w0T93ziaHd+qrVofAy8JBw8
9uYH/LJTRFoiWXd1EnixR2zi5pLwjMIvypdX39aGEcpFsy+uJV1igzqiNgxDrrle
R2Z0nQGNY9J20lLQhihHYEU6cBQ7V751wjF2J0gfzBKG5LIeqSUgT63OCRE/h2Vq
aXACJm8qiYdaFbNthSNiJ2HrtICIU3CM90KTd9iC62Pkw+qPN0N/fAVXppHXXrqn
ZzqA5Y84Rqya2kaNjK3dyEMhNtDgQr2Z2Y+aq4N4AHikIxHVQ+YXXn5+1BP65FlJ
7iOP5YEReNSov9cTDA7h3CrnCV+jQQz936UY73K5JaOnjlEmT7z6KjXkuvJYjQ0n
opBGvK6EcUpNw1SMkIDVVwGtsvJGTFXJRD4xcTGsnxAWDelKkVjwMAXmA4RrQr2G
lS7TPAhDu7JbjzNXR3MPUY5zvlv7qoPXHOfLVI4idlXihZbDgyyV6tCke30QL1px
dy07VPMd33XcJbnw+TRcnE2tBPe6VtG6f9BVBiLxmFVwWNdO627jOykcUkaVfA/g
fgrI91QvvjgZn8g8vMI8sai5VeXV1WkgaxBamPoosXD2YuiQAxsgRCSNNbEL/Eef
X762Vjm9dDWZ+VngPHd7N2NPvwhhUwCza9KC3QwSqV16ATIH2Toh7uCH3BrhSU+U
6s3h9U5h7kZdjomEPeilDcD3hHiGU4SSqWwbdrSQtmgmUEDBrVOH+LPPi0Tf0yJD
ZxqCZAtX8kF7jNtte4rTz1anhn2fqZPWoV8COZjEHHREdYaZs647BgqnT3LiUycw
c959G1xrpYuSJ7Vm8GbYTJ4EO2+WL2bSHK0P/j8NxPESbPpJMv1IHeuKgO8NAdUl
bz+CO/myRh7ql6H/9Wg1S5XUU4JxaYhy4Zdygav7BlvPg8gRtoeSruSwTdW7UHhQ
MpUYKANIp3/SvBIGxIf4J72lIT+qTXca2VSbY4CQrHTDjjC7VvrHyo5j8qjsRnmo
h2plJC4Eg9bJskDQFuYJRVt9bAqGFjGv4V6LbJ3HfRE1yhZjyR1CFnBKskQ/ts39
cdw22k4rRrOn89uHJp7CsdaALCk+UjtUcmEj4Vr2eEa3lvsDix0JEYNGPSLP2zUf
5Wzw1uRB/1fp2SuIrYIbaA3ST07Jw1oqSr0bT+kmj6miK9heXxNh60fHS530BjeT
Az4a3uGRVim6AQdeIJchRqhvLaw6BJUhdKMDjH6MZIgn69KlgRBIa2Oye1cA3F8k
WAxTAwccYFwU0pdjTgd840V1A+NbvFB4zJMe75m/luEGPoptUMDec2OVmqUSqPJY
TvfdHcHo07t10dLj1zDYl/NalXU2gf//pT6hXZ4QIelg31GpfArcJWSxHXx1OB1j
phXYVAmLZLXJLz7DdLU/U6VuEHxcmiNdvRWerSv1R+fmT74GkzDzNDvvSGGhDpEV
b5UqPbj8N6v48+iHl+1XC1rfrLTREceFqI6adXtE7I2oHrLvJJiQouxZHhvw6n80
ZqNhUjJxxRgPDLyC1u3h7zKPUAOkEMI27XBaeVaLJEDvFl2eBTIisT5O11HGgby6
N9BamLffFIF9EK8LebZD00ZcrQBhHiK4n39sJmUjKW6TjYGB2t2p0n4P2jaqYIyw
XlKVtjrys4BtnA7J10UL2rjbh3Fq8K4K1PC8wUl+UXmjvj+L6lYPRS8f4cp73EFi
ruqDYYtbZTGTlbupdwxZlglQmyqCC1wg3HyAKTWArtBbCkvLFAO7ruPkkY32SELG
nOXCuqktRdb0yczPS55d/58V16cps/YuWyqD9Buz3cYKG+ALPCAL1TtdS/VEbl2W
Io/9aJE8r8r/suuDFQLQ4w6/5IptkDZpB11BdNn+O+kXdUx051mgABuQrLRryLuk
s4YkPGcl9mYdUlquab7iRAoEoW/MjWi7IWNbOIP9y7Ia/ver+Qzspsj+U/Od58Dl
flvDr9Oo+VuxUo4g6hn64g6xJJMnp0Mfpmt5ZpNsyYXw3sGCnKlve0Dvi1hpUKts
/s2RWpgzks25jNazyNak8KQENVoNDeS6RK9mmjmIZDbAtBThn/GhFJ7DhH8GL1wJ
QsMtBiLtSRjGoOKliqmTSclIqIL2VEWWw7TSL50XE7DDtKt7rgJPIErjqOpKJ2ZZ
YLjb6lxhI8nKrLTpXKEeSCpbNiPiBsuKGeOpBCpfCuecJpm5y9trtpdggXxrUqFh
UQCHSMILB9zfon4CnRdivfERWrJv1h6etmSqtgi40dN3v7O9AfMdQ03kCkAIrBwo
pLlMAt50fCsYaId6+7ShF5bCvWv0SxDyrdTdv0i67PFKHqZTb8jbEtw9FGNklTV+
+BeDiLq6DzGJhjo9n7RZS4MB3EPOmaSdOcCIbXJs1GJPVpszdOphixCfaZ+xqnCB
oPr6Jid+Woh5cxTOFziExYA4GrjzchM4QrhOIxUzwtfYSG9kpLki9kDtGTXDlLVM
uibPazN2zTET5FOej8us1UyAdYsuqcjmWzUaFYW5Lk8UCb8rt+00VJM+WszXh9U9
PY9evi8H+vRMQUxLLBediZSp3QWeQzCyZOzsd+svuVjRQHQBYjPOlJP25LB9+os5
oai4PgoXOgf0AzqvFIe4HXPo09+fzFrvhK1R3w2NtpR0ifK6nYC16+PD4t+xOfK+
CwmnBbXNxaoKHRtXG/5nkajn4a2AWF/yXtzv3YSttYWaBdt2mAcTn5ncS5a8WPgv
j72r+TzPKciwERbdl+Z6ROsz8SejYsf/IDrnAF162k1YGfD2WxEsaSE9RCKJt43h
h+n9k3GIhWvAW+MKro8o6p9nIWLil/7F4DMkLdIOm8ybBENzkXgtLfUyfjPieLwY
BwUR8zF1W0NFQ09XPeqQAzpKuAQoVFcGpk2m6vKxv1BL22Sj1oxV0tw9a3DZGhhy
Y6Jee5CVUf9EUIlBphK3poaqg0AJjmiKwnDSnmk+tdhEA749VuvoXhQqoKK1lkq5
xEMSh7P9/NNWQZqoADB0kt7pDfNsjUl407alBydHiHgg+xisGwofj1UVT2tcezc9
4xH3/HyEg+nLjMChvgwrei3Qqn7f4lw3kMmu7TAdTlBm8fVX+W9tb8muGayUlr/j
BvWJxoXu7xV0Yd8SUG8zVagyk6CfeP2gET4ELocC6ppqK0VJm+WyXZES7cs5b+/k
Bo6apJ5f852GEV2/zU/0OQkH4/0Xl9ApaZuoNLZVyENwXZx3ggrlCSliXNsmkFpn
iJlyTLKXNdmxBeToWY+hW7NiIk3lQAevJTOVCRd9QoBNMQjBu5BUP21mjaZjQbUm
IzVSZfiHW2tYkbYrF4BIs/I0ff6KvRFnypH4SoEBt5uMqI6kmNXUHqlZ+pv65WUe
7g5r26JagcQUTOOoc/fk94BTzFqviLzHgx61QC6QowqPT4s17Ick/etpksvEOa58
vug6Z5+mwqXRIOcZYRGk/xBpoPdIKUG/5CsNyK/C/CISvs2lpwheQ13F9B4FgcAz
233iVe2uBc4QfZ5pFMPLR/ojrqre9l7mYpUAXBCVHSyeSOgsGN7qJzK9OMbqiTwC
DrraB/gb+5DGBDxXIz/nOA4TPfunZIEDRNlN90oC2oeuufUrOiiHV+kQOL0xINGa
9f6n6UgTSLGEQWfqOwUXV+1/jrBJ1Dddmqiw0dnGNo6ufmAC/hkxPmusHA8FaL6c
HiryXj0KlNoCQo18u9mh8uO48RbkIhiOJEjrOW80HbxgyAyXabKzYZomRqJTLvCO
XuPT8q0JijkEA4OZh4f2S1Uz1yAlMWBj5VNJq6g3/zcq+Ge9o4d29DJnvoEUw/91
MRMIfqMWV9Ni+XBHNVoqeCUwvIS/G216CXc7zQkfxD/Xl3sadVuwaKj6HEWc1s7b
V6HzLn6dviDun7CPo1gEy0+Ma/QzBtlO6CSnBbdDNKuu/vbDFf1y6Ygw0OKEqRK/
lys0EyHSRIWpjLuRmhaWzz90Is2FvWxc5xgyBKx35ul5g7U1JPCkWnhOmZMltuRR
d01NHoECc8Ed1paUBesrCqd0T5TC9kNGfSt8xegS2IZwwDpSfHWfWS4/xp3xvGTV
70sE7onBovtI0OaFsX+2dZEv4cEyJtmaVfiHKoiMtDB8OFScaqGSDcLAnavU8hRE
zPVKWW7kIGxdfSmFcGnYtgdnroZpUdhsvcrZ2XG4+poQfaQ3w1vlbkouJ/q+TqZN
FH5jg22eLKj/S/o4qQggVAEl1AXme3wKh6yk5cMgbPZRgO3QWLSUPAA+Zq7Lh+km
tUCkq2rzZVKwJL25ttMriEyTikZ4jgGfbKjj9nd/dCplsMiumHxCljSQP7sD+/oe
ub7UKCfwHeUUKz8Wu04SifA3Worhh+AFvTYDmGQ9SZOc99WZOY5py10fPLNivTN1
5NtlLJPcXSzlrD1R0h4fx3HK/U/lxrddQSm4zyKgkQ/MqUuiGhhKfWpqIV/3jKns
1vad7GKZPS+fRSTGeT4AQq0KbAqVcFJuHbyBiQ+KMEYmdtj6ajQk4YpwvKBzyIXn
vL1cBO/yKr9y9eDGIG+U/KbXbscM/kHZ5t23luiqYym1TG751EfNZFmXyJRsheon
/aHC+dDn5YpDRFUyIjqtUiUxF+G+PNMnUZL7Q+mSQxfNTQ68t1z1mvIyJlsLtGgl
sZRN0fYrPQFZ8VWmEGFuHdWog9LSdA86EXwje9jnG03KY8+Qin1SXmXx0qwVBSTn
KLgp3tc6qUWxWbFSZiF3CIhi1SC3xd39tNiRHHg0yueoMS9G3qrv26dID3pw851G
NkvNqP1+aBxADBYfR7TtlxtaYe5gvitk1+e0tb8/1S10Qx1zR41qzR9+UK7JWGsr
r2TIBMpOxhiCI310pZ9dQ/J6nzNdhm/V7dD4QlbScESkXre9t1EFKG3sZL3WVVmj
UjsNGbPLoJURuKxyj1BkAIZGXoKN6RIogjqY0MhxltQPls475f4M+hcv/XPTk5Db
3gonh+qqY26Fggemjrt7clnK/RPGVqGItY/dJ3AkWPmaUSVciJn1p0es0lrANawc
mRl9v0qC4+tS9Aly9deE6R044b/dHBBPdvt/3TTTK5tJdkLaaDKlCHxgGT+3Nwu7
PsuBodtVDeLMKsgtpg240ZG4hEKeSpFF55tSqZWYcO0u0ka6Q9VsA+yfSsegFSyf
/GuqOrzHykvZGM+F0sem1kfPiqZW8nDwWKagYq8fRTuSyOPrdLeJ2bEk1u5+CCUz
BGVNtegBAbnr1CkatJoN9A0dR1nloxCJ4SJiraWBWme3pa8MK9QofdhLh5bTcFN7
6jPdpNlis/XBIFiSlRLPgMrGdCzif8bSO/PLb6trtU6By/jMzCgecrllyG7UvUB0
+MsHDEeiihx5ZTEHIxtUdlz3V//55KLMwU/oCWhrUmF14thzofGsKXEAZEh9ovhM
ho0TF2eutNaq9AIeE4+UPVE6vAhwrwKEMFkEM7oLDexRqSVmwUhdnuXy0SGgWq/f
KVtlC4PTwafeNLx1lv7Mrn0P/0+JoLryydHKHhkZmwfE6FrCyZhIeTlkA4kjoLzc
fr8YXCYWXtup9XHIRI6peApZAGjVy6Pxf4b9SWbwMFI2a1x5U97Cu8SHizHRXJNd
MKpCdVPIMBDoUWUv8bKBs4Ir1dr1i+UpDXNEytph1AKn83cbVdwGs40wV8lGCNfX
2TTp2xrn0QIXReqX11IjAUG+M0mQcDDZVWRa5h7rU10gXtyBVSntxuT51eUPXYLW
uEp3SFp1iV6fP87YrWOCDkKxfgBfz6vfig52Jm/AKG0A7EZkb6sye90DVh77BDDa
zHyjdp1zEtpY06XwZlX68uQSJQ6DETu16yKxnPnxcK9DgVZyHxGXaGO9/z2co5aC
k6GAkckag6Cc3lsJia5nhP734HGzcPcdBEpSz1aK+uv6srYywHRPS/hOgXtt4RxH
t9FaFhTgwjpflfYwEcyLVZu+1leGjrIrbfRK2H43jQbbhgsiAhXUj2wfuXgrhMkW
tFAE8bVrRvC2F5oxKpDnsC7aJ49827q+ac0+eodfDehWpeKmBjIYIWt7qFkNDwKJ
9XSr2ZDFujV7aZXt7A4QmMTnJC4cvDhneK3XdSb9o4fZIeP457zEigbyj3K6Ow+m
9sTVCZdmCGySXT78Rn4fbLiFmJjO+ZJPODQKoMHsdjzmx+CQ8qPKcOUD6BE3aUAn
ByZtm0ipqo32o6K2CRLQ3ojKJJdDSwaXW0ad1z85ku5ja4k5SoEbxd19Zm2dKeZE
iLPelbuGJ5TgCWelc7MB5j7V+Yuwh4epuwXvq+NPbEI1RN9cnH/ev706SREUqLvf
nexk9Cuf60faOPXRzIB5si9cxW2cIw+ZlgZPeBYOsxRwXkpUdHsYX5butE+0CXZL
UpOU3D5Jh341ZVQ69ROTokOQEfcJQdratl7jH6rbfD/2eg6z9mPKjXC6YIFLdSMS
pXRQmqQ/9t3hq56maDo95N/QLTaBt6dG6MalnFEMrE9pEsXI/gQ/W7bwpUKSkfLC
ewQPKv9kKAWSxXu2YSMMQwi8EvjVFG4bCQOAp3H+tawttOIbZjHvRh1fJ67h5LcI
m5MSsXMd+ZOQT289PILDknsFXH9/5TMioFRO55aidNkTwMdMzAVNhJN2fE5A3NsB
iEVaqyliZnbWLFAlOrXDd45ous4o5RPObTaKAU3pKDCjjg1FIHLDQBgMBm74pGYS
Z3mnFCHA3S6o2kueVVYTNYvlGtCu/fBal17h5MKWfQcz06FaJ1fCC9VqUQ76yGXD
J3hnHm8YujJkZ2f+gGxTSFhX2bTJmSvWNxdELesJmDrywGeZWE1QlhNATdWA3VGQ
nugoyX38cioIoJ53CFXGcVXOygBiiRz4nOky8WmU+ArCYh6xn6LQNgbqxgfv1Tbf
c4dxsm8zvSBwyCPwbSTHAo70rT9l2alx7OJgL5nf0IUibTuDQgrHU6sgfOE/JHH3
P3zXOGApzTcATMM4+bmUqRoVFUQ5cnyi3g7hrR4Qj1mTx6l5Vwtx0ueegYFWH/DL
dMKTcFGTlWmw4cyyS0EDAr7WlPaB763w/sQH0+Oon5L7nA9jr13+LKN09fhRySF5
WaAVa8gSOtgGQZ1hs8Oh2CRYL6YvwiVzr+ycVdjWZdRTl9jzpfoVMieyFM3w5lkL
Lq10qJLG7W8xpBtO7eCX3EHX4XJuSblMsuqbPHIu56n5ZFc0er3m3sZUQtSea4Jt
xbFZNxf6dly3JX3/DgowM2gGxZW/DMUdzq5+93n6EWv1KhZlbAWXcZE3OrmQ68kP
a0dQ+AJnsbxT1QjpGfWXu/IPr4l5DwB0ckJVsTBxWPEHCL2ml398qysPc4wAaBbD
i8FE1v3YQ+B5kGeL2Nx+QxDhlWUyr+FSgNQ2AEONfVahBeFAxg02Lw0bIAdWEPMG
L9LU3KOan5NsuEhThX6OKMxLbGU4JhRZQViPLXTNHKOTFLrcoBflXtnRbv/h3hiH
wp3N7ppc4xpUvM16/7agzXIFusQtY96CRljGJYXpy5eTWUg2h93fV64VrED8itbA
/RJAK2mh6aZ9XS+eeS72VA812cskqAt3kxPKlsyaTRJsXwymCCJ9frHO9mTlHj2i
NrAlJOCRZamVLCyTsfMo/l3mHt4DQyKt38oak2jmPMMKQQKtdjGCVZ8QYgEHRlAV
U5NOKigJDvmL+SSWC3v2p96KNJkgOeg9rG66VGCEgw/JuZA1F/DH/kKrWmQKoxT9
H4j5IOaFrLKERLQc/VTMnlITVDwIqUSGlH++5r16pc6nD2G1jJJbULnj48hvaXfo
XNVNGq0YUsIi0o2FYR6TaTakGtvWVAgSdiJtkRQ0gG2xj4gjgBNlwG2nubUNKUiW
xDiPRxm4i/wlQNonWq0vaWDKJrPHChjCFPOzHHe92vyEObjn6d+L2T1OGMqKd0+M
RDVcOKT2JCox4ZPqTvNTmW9gAJE+i20lqbgt+q/gKHoJZgA3Mc55i7ELvR7zRWe0
xkMd6g8m3SW+xKjqAH4aNg9oEPjIeziZ/wBNsSDn1K5sQ0mF1MwB4YSM7I5L1Gd+
MVCfq5DGtRraREyT8muwA2ID1OY/Bd+C3dYvmEME+SXq85cHX1M/b3iv5mvJjcQs
mmMtJcW6HNX3E0/+BYNBX5ppH8NIfF+pH0DGtvnT98ezHkhlS+KR2hQlGZ1skdb4
cCmRxHLeaso/52jfNdkzluRLlazQsbFSsBoUMhiUse5bfuF6DeFlFh4AGKI4X2uI
HF77pVW+6DDNfMjlf2NmKFpxOXSIs54H+jlmgPe9t3j36WEF5widc5cu8iAcRzde
Fszr9IjatnjeCEmOMpXL0iLXJI52ZWdmzanUzPtJVaD7HP6+BSlUp+Pm3HbObDqJ
NC1Wgb77EzqPJx0vu9csa14zJxepPhRTwFRQ3NQmQOFAnzLsmxZb1b7VNWHAP+ne
9q/C0ZyB6DSzEgxLRFxs9L9LwRD3QxtuohSYxCE/w4wRqTIamRa2oXuU44ObN0wJ
aXwbi55YPovNZCPkByfQorqGTXQav119i++1cNWkDpADThfTWm5ozBMM4w3Jrf3W
0RWw5xdjcxKVp3O/YRpqqIPtwAz+Vi0SSackLRXECsb5yXWS20m1P/iTm3J01+kY
2SckMk+1E5cL+zFwK7etmS/pVIN/9mFyMlvsWZeASbETE2GK9v08ZStt8tFVkuMk
CESaxh5lgEue0pZl1Ctm2ZxScNxZ73mSeLu5cDAv/ILxMBA8UfotHXUxArS6Fd6D
faBvxNWCdbZxYfSZaXgdyanY/fbAro4oYuEwUa5la2zQqGAa5t1zsxyJTH9YeLaK
CNafFuLONpZH4ktHPtVcThR5RRrXsoZeMOoTSMeWu3TMnS55v+8zgFOB6haICA2t
pWvEW/1DWRAmCQUoWTW4uQp/8vv9JPu3nL/XKkTWettXnNC5IjLjo6yz5Bn38QhW
mjFzjGf/j+o2nUICVO7IJUBkB1iPaelTcvV2APr25mEskOc6AEHIsOGq/j/Qh5P0
Etr2f1GwZmyVHzDMHx+Wy7iSXRNaLCYOMgJyzZb3bEou9o7tUQ6v1JIvmJqFk32M
xXphEzr34HJfnC96dqTv4rUYxG3pKeTRt5C5NpqfuYNrV6qVbVz6eIFsq9HSqe+E
G3ZWvKhdYWLf2iQebN4PvnA23/QMrDZhJHPMC5DqCmBNExdB41U58J77Cm/y3dyA
J8z2+OEwGVw8PPqnbqMBm40/QpY5Zh1zApzP/dVwHAgphFPY8nw+xop8xYpznOaM
XetR3kkYtI/q4vhwDJS3GEUdJ+o5IO6EbzU1430zofK5zlkQEpGgDTiHOwQPHHYW
mPZhuR/D4bgRhJoUilqP7HT1dxYonZZ9yjpZuarUXyEzqOzNk+p704OQrjEtxxEN
VMZI3dirlMY1K42enYCTf9Ti3yu19xNVG5IJyx4aoMuIjv47iQBXL4dqhGQQ5K3y
JBqLMjVCSbMXF/u6E3bQBQvSITMVaBZcnGU14RKWQdaWxrsnBXwe9iCxlwoFVMGH
wkuS0/9Do0sRssSpDWNYbZfmFsoeHcrYX/La68QQiHn4I8YdfUUMFEFVdnp8CaZt
vyeRphqPbgTrVAJO2AtibNtUAF1Cv1CgNqqGLrf054lnO/qi/E3lsM8DrSBKBcP7
XxJcE4P33/0u+242p8ogg6a5LhHBdf4f/8LbAuG0RdYSQ7nDjYf5zjdqrLUPPmE+
oj8tk2ijr2H27q3Si+M5T4yyF81TclSDZNw/MGkiuDDHgqfaUy0yF1NP8lnmGKdA
d7oNY57TG9HwmQnooZCGj0+Cln9dVV0Sf8tu+UVHMhioq9CwBhmagY8YgkBPBoIi
QzjRZFRHNMIAjnRpA5Il2+48M73DehAM0BcIggzQFQWNe6hNhxXbygxmaTOrp6XT
e7pEK26V3myu50I7tAlQGqDAEk21lIGhFqw4Uq+Xm+fTV+P6mxHrGPnoKQWUwrf7
SZfpUCm7FvVxKqpu7xxbMici1emtWs69+6z2J+OQ4ipXR7wWXG9IRb42LbKcfhkT
RcoSOCFxWHf0HWMMGA27m2dZ/LJUCX59YBLAohBrsXx18qm3IcUkN6nqRmuNqJGs
49+uwErgoNbcdMwLQtGuRjmYIPQeJ/F8f5Ztl0km6bXsie7pqRGVK7VPl0rgQZCK
Zg+Ob/mDHOMs5C4oKHBPzIrIl0YILCAAj3gYACx3tFp5WhEVJ8hmkbBGc6n0m4iE
FgXtR9ND/kEnhOXEqiw3W1DOlDEEg7Q6GT0mD0aEiWDRSWqaMW3/IgGaLkCf9e3N
35X94o08ruOPMGrRimpdYO0liCFocyRpbRidGWNReiAO8CUVaMJ3+scb9y+5bN+i
QmBztT9Mk1f1uaBBInMyClfR0HCMUhGCCs13rFX8RproL/cVDhIezF0O1ekqSXUe
wRQV6ge+11+oYrR5qtwoUYQPXXlvT+djWeRRhUCbMxDsVyPiJOf6hSsD7H9hGmXA
yzXP8VKbxSO7zsGsGz3IfeoXjCD8QB5R05pcqiltuLu56NZGA8863HHXNB1yqS8b
LNfnh3xUgfSNSupNrZOGTn/fsM+GD+T/zMyFHY6MK5vRJWdqNTdBu2sMMsFomLqM
puKMxSIJxvA/s7IMUvZaGuw5OPo91vIb/IHE9gkpQqmdGxGq6qyKwxXVTDE7/KXM
pwpEg55yV1NrQ6aH07or36fgpyWK4OyZxy8TKQa9n9yuKRdELohyKa5diocxDmkD
+pnhh9VQQpRBPQNpalnUxzDw+PaCjyVy7zTpIdNghPdbOH8O9hQh5qpxZQyHN0jl
taz26iz24BPZxruyuoLxi4zaCE5/x46OeZ5DSx4Htq5sGr550HP8CvOiNeYH9Bht
0JL42gF4rFjhwojUKA4sllCeK5T2lfQkNZzTIezW9lqlHnJqqwEhi/km9i2HLEJe
rACJOammda53bmcKh8oEmQ==
`protect END_PROTECTED
