`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YBojCb8fU8w+byW1KS2oXlJPG9oPZiB5/1FOheRb96SQVYAIcPDK9bHHSiK1MHqh
bLZuFl7662bsLhZ90SenkxTSA6qcJIlQkSk8vtwrFEyIJVzFQgdspP9wi5448zH/
6z3g6RUpRI+kNBchNMEQZY4mvpy3aAUXsW6W2G9SZYfRSCcMaPBGelyNQAhFBSK9
WP6UWKhQg6CgYNAIKl9+lWG3I2A5F4UjJV9abm/wQkHyXf3WjjJbW6yO3pL39AmX
TdfmysEsgbrqGE2FxotAsqOkmMv8DEkZsWNIvRb/wnRt1x9F3Pjnk8jbrgda5dNi
7XDfV6KDDqefagWdpQFttEGiChz5/iJvcTzjMyZTROCQiE27pwhpgBkbE00zGIDl
iJQ8C+wIDhpECHV2Z1ooe5vZXPFRqaNiv0ZHgNZ2Uf4AH5cYvNlC8gdxJdNpWRAP
YMNEfzLxeFHyl/XtUhdAFEgRaBX32wPkJKoDxRKCqm3+J3CaU+KuKSYgx59SH9ep
HjsRUSswZ4N0zjRLQW4+3Xz3JMvvRCm7zzLfps1SDHPLpRF4XjLQDy5Xfc8mIbFq
DSz7JY29C4DuQVzoQzs9Pm+Zr4Cn8Dgb7nv9lor4og6bp7oAQlbWSmBnG8/fMIkP
wZbSRM7NrdfDXYGFtUknZwQCrkqRvGpBrmpRAyZUF1Ky+trLo67nd7v/djQ/H1o2
LgZkcyC6eXjpGBb6wuuWe2zrpXVjLMmc7wg6akwGwxOvo213+6cwBcetZChhpPMP
BSsOqhS81NEZEnSw81xG/E4CNlCLldCy/1kIKdEU8fI=
`protect END_PROTECTED
