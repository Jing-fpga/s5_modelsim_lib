`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jLuOL+Fq0W/NobCdA4yOMZXX5GC+k/QiQnu7EvhtcD3BwRq+xXR8s+1S0S8yV0BN
peTfkoRMAM9UIk/P7TurvocYIQqxx/8kqvKgzYSYFsCwb3qcYDplQK8EDHLKSd0M
YoPspF3PzP3SBNSjsS3tzNgwCAPhfFc9rCA2cBTsT62YTLqGEfLNa3FVAcXFoZgc
6wAwgwRKuOwVnloiEG1yNzRD/Wv3xKDOW1TmrfY93RPwQm+N8bNDXxx2oRGNWlqg
dzWE1j5OKI/kdVgUzzR4C9ZVCOmPtwJpZ42qfvGLD4i5Dq4cyMc0CeE/vhas+Otc
lxwM+2bZyI284ZiOiW5aGZaOp2V0EDVR7zTJGJtN2k/VTWFXn3ejjTr1neNVBpip
DPiANqp3jjxKnrjVCkfvGZviUU0FR9UZ46Tl0iosfvsaLjklJ+PnqlxpjLnLZPke
4t1W2LZdj4z2D15ixU3NBKAFtvTdc2vg/9lPsR0qAmKKteHQQ/w2TS2YYuro+8LM
Bj3nriqtlQE8EfGlhhLWGz60M8/FsXuDKzOCXBtZ1j8GSHRD/+23S/ZF3nXgtk6d
lQYRn/oGUEUZx/uPu3nfYkN2id5kVFauRKkO4vB7I7eDmyczXVkJnFUc47gB8BBB
SqPUz+p61L1ALwgy8RQfKj19zxc/6feoJtGxxNM+wmoqE81KU5EclBBFgU0eQ7xq
dP3spEOIFFvwnFjJxPrVVzgJ2sMq1Jb9uoXhy41570hgDT+2/RKrtTk44I6CTidT
7p92oesyGDL4M0BVzo/YwY9FdnCjLp8x3WpLa3O+DwvNolHXzd9+CXdK6So+hqs6
e6rbWNe4xdu89Rm1FcSfC8Y7J8Zdtuywxk9BrhHh/4jZkPxzJ1CQpuFTTt47q0sT
1rnexD+vYGWMknAA3ObTBasJzUAvQNd98pyZUvkEe+9wdBbPdzxC5cc+zxrpL9D/
3Ji7/odh/xCBkJ9svawH9W5FnEKFsMIeMxhjorwpdfKXpUDm2GNOkM88yf0Hy+Lc
1zy7XcMZf9bOy68u81ud2ZpcycR1ome6IRD6Y3wl/2TTkqr5UlE2n/EW6WXJuqKV
dwC6/Aok9JtobMdn355Xv7wCScVB9vG2pdZxDxEmrlpTGy/berEspl6RPtDAfbfN
0Dk4NmPmW71diSvuiYlPiWrlh1mluVmequhV7ITwHyTUrt8jFGwCoJLUCGFvvnKj
4x+ea+2o16At8gLYiwki+hXcjEY2Cw+4oZ4/gTIzPd4/kqud70WIY+6txhqQVh32
4acSxotgTxyg0/IjDc2YKasHB3eqv7EZszIgMwFBgDAedOplSjfC3JYtVa3dLByL
h9+0shLdfc0ncqmWvaSSSnlFn5yqXFP1oZsMdjv1wU5dkhE15++lQgTrI6hMkzrT
qo+e+WYPd85hmRFvtWe2oFFXa3whVIWXw++NvJJ3R+XShVvOkDcVcHNe8me80Azk
8WRICeXAba5yFGhQ6itIKIDe+olDfuiXi0FFi2jJC23FM1nkCa2IZkGevtLnjTcO
iE2pBf4Om0vcM9VOMeju2X2duUbPVyUARCvRDZxiT0C74kP//SsIQk+gM0lWOKoh
CA4LEqLm0mnSRRlxXexyB+xZaOdAKjanTZHAm99EeN9oGLloIOwojGKEW7Mf1LKv
I5qCdDyhaJ3dXvAn2TkURXqi1U+lmKyNs3gYq171AWjOpYcYgUbWEKRsfmtjCWDe
QfUbEvJN4fEunHKkHryUW6xSH1Cyu7XXzVgMg4W08qooEUOJvWnBTr09mjRpbXB0
I2VJXqfgc3l9L2wPZM9XgUoK0qqJG6yFPOuzJG4v3ygCrIjMUaZVc4uzQI1bZ7DC
DW6w6KwRGpRcexVmSUxnh+YGZrvc4yjLuFYvhXRKlTonJ0QN+hfr8nMeoJemYRfZ
f59pSgEWUVNdY/WI7uJDC6uf4bxZjRbVWG/2EsmBh6mFR/ecnkur8Qw3K8ei7duK
IFM2kwWNwQ0UYZSHu6YLeU+pGu3IdVU/52mih9mdn/jxASlui3UgOapBoLRSiqbS
mPDHpohAFIRejtQpuuTEjgiL+OWOI44Euxk8BdwjBYMaoboAyXAvGXJTfl7fm2Xx
b/uf4SmPwPsK+jr3ASF166gvlpmT6ckcy4t7JgfrBpDPAwp2pIkSrnMRfALJ4bqQ
KdXue0erYy11mkHatJn/oWaOKp0iviCgHR575DCbLq5lqo+8JOUF2a5kw1kX8LBE
6xJT9Nwn8Dt7LOTbLkqNDTg4Y69USPXWMSoq5gI2WadmacEDmH9iSruXR8pgVkLa
0cnY/Nk/pKRp6dU9WcrLK5xDnCYYNPCFSk5jCUVTlD1tUT2gV0b0sBUoURUUSJkr
AyX+o/zXImm1wbj8pvplPgMON5Q2aXG+Teb9YFA3++uRJDmOmkHEa2h40JG2j390
Anwyx88jHj8NcxyoxqIh5XDOcVQ4rOiVN46aMHwRHTVGM2tTV1q1Sta4b9Kxk/Ag
8qsBJfvYCPv3HabA8u9rO0BEDnrgeLLcgKgD4BHfx+wC+Lbgtv/o02MBAPRgO92U
BJBuauDKNZlUeQSwQ2plem29GkH1+nmrsC/678gXnZn9RPVGF6SWnfZ/KwJ/Fwj9
p7d9rb0+JWWlVL0cfT+o5LOl7N9vH85wlPJzlHc9sk8mOM1Am1/Dw8PniECnqNMF
9P/VS/ZVdfe8vqI5fFsXs7vStvMedB+MJyJCNDOCZEbrMO3/dW7Ex22xe9MJ9bY/
EIFVMKkKBA+dB7pQfXSmxRtFVKakBESA4fiOBhMgnP5RuHVQfa0L9WDTP0Qikus1
cT9qZ2n2OWhbLUJv52Bq6tmRd7F7rQheCnwlFImrefQ=
`protect END_PROTECTED
