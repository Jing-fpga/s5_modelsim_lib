`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KE8GN384M395HvQaFSbHTP3D3G3hEaguze2glTs+DcC4kF1fRO2qxoklAJcMgxpS
O0NWnESi4SFbxHShWpf5TA+qgEFOWIPiCBpQMPhfS2PEdlfxVfppWM7nU2RNvcIq
v9ncs9ts7C+WIFyYM4t4zYqPPkC4u81rclc4PWxLIJbwkQqMsyczVssovjjE3Uxn
FrgZlDXCsp9pPHzUplUYPl0X7GlT6T5UtxXpQUaEQrAXlxK7ZPAKoX/EnA6CdzL9
N6rPL20AnlnLgcE2OXrYRNjcSH33tMlpBHUX/ylM4RHkBmz2uxBhxBKROk1WjCZ0
ReV6D6DhAsiR5uVJ4AvbxhzG+8VO9ExG3KvJ2lwi5WapG6my/BfatkGp/sr2YH0A
ar0pA0GZUxabMj8s0HQWosAJnmCIQwkiCjMfbQEdtELUPgoNZ3YE5jG8U3OEXx9w
ux5TVKfYv5aDhArbc80AGW28w+5PY1567NqpnRWpRKdttH3Dbd4HW7HZGdEE0jsD
d1qXgOkG13dKQjsN3dtCrRfcK62ouOsH8I4KhUcTiEbLWcMthhOiMZULBhBL1LiW
3O/uJ7dvuxFsiQJVromLRqlBtBrMWfYDPtAMbuJgh+wX73nDoQ3vMqfH9W7Dcob5
wdH5TEid2FEQdsmG7bf/f2foJIgA7SDdY+qmY/JYf6/ns2mzCfbL7RL9Zyy011Ub
o+tNC1H51gmtumnV+TFEQVBJqWzibSw/oTmOV8LmhiYfSjgB6Wr6IIgLY0cAsNcx
hISwQtnP5lp/IxbqvwLLhHHR433qSPp3pDowibjNTAY8X+np+fs8iTz01w9t14to
0g1zU4qBeElL2502u4GA4IeNTPqZROhtq8dHiqwDDPJyIHjXfxPSLSHjhMu4wHqf
jwJ2atgAgKblUM21V3cRtrg2dluXJ45/EycDUC73mrVbgn++nI0yx13KOtiH79kD
gcATsNq2msOSuaVT9QjUHX/pXBwh6eJ7oguwf1cB4h09bhNK01xVnanbBEC4/mU7
SODK2FDo8qrqYRLGlfu3MwFjISkNCWqRSiyAjoBq/9s1OwZAflfkPxu09ObStrh9
O7+fNdzvmAL/I/Kicw18dzXnYu8ZkflDElS7/vCWCLUVxc7KqKip/yeNzFS9w2Ho
aLhvGudE4gsG9qX1HYL82Wva7QjIthDF9WSRH8XpBXG/nea/5oujyd3eUd4j4vzJ
aaGdtB029aZ4jEJkmcTxnQ==
`protect END_PROTECTED
