`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oPTb+tYDx/ApDRGKOIULZoF0eCm1wh4VKTwvjcm425ZWERgEYcRExgUO9x2OS/aJ
TZl+HFwZOQOFmZBYDGsbhMNtib+iY0dd7wraSbe2sEak0WyGNlHFicB7b2EF46ye
XBOW+u7O9UZ+VvWtJUzGDkoBVfz9bzJrK1MZbNkAE3RyWXiKlq0ThatlQUVaT89b
BYWmxWCA5E1F98rHgl/XxS3OdjWnxQrIp8yglMvvVlHPfD3zt/bfwbEErQontz/d
5VpKqzwdbbEwx86ySnWR7creUUxTv+JUdFwVNAS+CMWbrl/PoZzwDS0Vg6GvRnUh
XgeTMMFndh4KKip+MEdPkv17DZC/1Hf15mU1AtMGY90f0g1z4j+QpTx27p0n6UeQ
xch65Z4bvTZLYMEvGd5mC6b3rMrB9y4FimjXQKnvnxpLrpNNl+PcPVwxHLaZw3Cd
rN7mlzpl9sbMQgujaS7TLWAGjgNZEhAfqsfKTV11iFvf0DazC4Jcb7SB0jwf5Jnp
Mqa7MhWA1/PT5mJ+tOmbXVart8OhgRf1mmUk3VaK9cT76XTwkLEUI98L6kaAJDJB
tfXblrafah1fFQvfzMFiJVa0RGemhaZmuU6dSq3Feaf6RBKVTtO0QL9hhLnp6Pky
tWA/i8VNkfvsK/iuSZJFEZs2XYYIW0FjWpwhJ9iPAVQWRXWdFZZEx1Mlm4w1bqIV
xTswHMmUBfc20ZHqYsSUPDLiggnKu41HfhkWIdA2kkJdMxOnEY0kfme+LiUK/jck
XUueqHPbyX16NQy1SszwYQgLIVAMcsDaz/V/aQ/sfEIXo+1889vFjsq6xieJCj+8
ZiGUNx4dKW/fjhcp7WawaXb77/IwcD5kwB9GjYezf9oifQKmhAPCumV9V8Fyl1fR
T7QDSEI5mWSqYBnPksK0kJpXG6jWluh4/JOu0tQuygdIVjNxBWGxbXI06KpapH51
4WHDOM+oQZSIqI5/j+gCJ+A2AxqMBhONMxBEXSP1WsCPb8gw01/BxXjeLisESvl6
8nAiYCY+ot5PGdkYoENeDVva9qgtTkNdHnuV6mL1RaRrppIjYoQQYNLcmpbiX2Na
tVMuE4QmrJbmR5ZLwSlPDw==
`protect END_PROTECTED
