`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bkeGrPUt+3pkcRnKaX+C3AwU+t2Zi5y8MVDubAkwhYykmaxltqP/x/CjO5Vq39x8
h/vMC2erdD/iJdvFKex4j8MmYX5hEZz7PG8VyeITGr9oxPcaGVYtM9wxqVEhdJAU
IoW9uP3imIGpyUkcB6lA312N1jwCN1V0hbDeJpRPnleLMCAym0GmuAaO+l6HAVzZ
g51E9jNoQCm1KvuLLO6qwika4EeZq/wKyLaiH4ZMH0fPky0o6UaxiyDnb95+1gAF
n2x1WcIVEoXGQZg/42WZ1okQNsLl7mBC1cZLByD0CqFoidRwkRz79Eqb08q919f3
IcfY0yewZsFgvuQgimBnGBgVX/S0e0KJwljUxQ9uutLM3k83VJM/xPHz667Lgdj8
IbYOrKJXb8faD/z2E//tNhPCcAZpOv1wZ9kww8tSAof3Qf3HzOD6CAThFb4CWhcd
J5Dd+hCPhJ0XLyhpur8oeirVsNbjUgexHlVsFCbUi6xM1DIoqub43Kj18l7kK5HR
J4+F9HkKasOtQwXj66/dIkd7mp6+7RpUlBdA/J34JJmMtpywLinN2PtGWtnMAdjB
gOtK/KoyiEqsjIdIVKmAxUkSjKiHkW3Hl3J/1e8xbo7Yywx+MinL/QJRQ+ONK8Fh
AvmU7LY/ZkYPHuwyTVPEq3EzrgzKRSNWYk9nBHKR9/CwPL/zro58JPO5J2iJ5VwS
IyPXvFB5NOx6QiKbJvXa5hb0X8OW9y0hlx1KIVL8xOJj3u3UxixqN68SsfXmh9zP
8GYlybpWZ3cCtkTLAH8IiZZxjAyB0AqaYAey0bZIaPpvoHJNSTMvQoEm0yIOABot
HzQKyzEMWnGOJqM/ivSAlFLXm/nXvlVu+Z9LNyFBivFF9MZd4c7qqqzeGP8Zgh1G
hYtO7QEOdL/SQBlJATUWh39skpddgx3XOVFCjSBMsIS5Wm2ql+ZdrJN7KHPSiqH0
64TcsDYjZ+A5M1GNKSU8HD2weuk5LM6UheLwXa5FETXoCdLbQ5JQvXkNoRpvKRQB
rs9YK+67gk/U5ks1uaXu1d8WJp3V43MYqPMNY8MEQwQ2uxPf+dl2VmNky1rHgvGG
DTiIy9PMYeqIjcCvBJKgAhca5aUjkMtbAM7kp3SaTfLlQkc3NZGz5OB8EYv1FzHi
fVARuJbMHI/almfYVJFdRxTCVczXgSUSga1FUmWHy1l+iIOF3n4xOb1cqHRGsLRR
VOELUf/N2hHd33ebD2XibHlscairhqsTd5IpOdab24IIgq87L2s8N/KJjlAqNQBT
`protect END_PROTECTED
