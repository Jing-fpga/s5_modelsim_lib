`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SIkJephVob7c2vj1CMJzW5rXXpC9Sj2fOnE5YkBNDWPssbTL2HbnncNFf4Ecff2V
t2rrsy75pjXoZw5i6wGAH9koaY9KODJ0bssLnEhaYG+9SxsN18nIrTFRoX3Zbka6
hzEzvDtAQ672qDN8CoMMjArEaTsZ9vphlQ3i3pDkklxw6BcpVH2YNGDCb08XRqCx
x5BAIYf2sq6kA4Z5pWQbP8bdWnYR1ZDv8p/iYEgsZ0aGar/4x0p2g8E68YEzsn7q
Gtzzb7+SRObsOtPaffpxUmHhicZ1yAghOkjGcxhPNjhodMqTAHlE9BWzwyZF3KJO
cwnE5i3bTUauy8zp41ZghrPJaQW3kzGeAhKBxxsRWYcgl6fm4wkXGintCZGegUAY
Too1bBu1g0qW3jkQZ9ooxTQtvWymnlU2Vf/smi/RIU0c3qkDL9NrBE8ArOPVmqyP
0pJ9xq+yrEA7w7+M89L+iiGHKaW9UqNwWpvey5vN2Q1bN6UojNwBAJYjK4/P7d0Q
K3mvxDih5vNAWhNfuRGfstT8Imm+NAT3TmL/yiGkg2Vc5Dn4vso4frls9Vm1CHXM
j05F3PWZI1HD+HJMnx5T8WSocggLE853hnrHBcxaIAJsUaLbaEl2LGrU02vkpaAp
fNU9EsFo68KWjv+LeuiWBkwpTmIx3IyIO9lO2wzMCC8+ZOjZG1yvaGFU8hy8myK9
xbG0YPUTCVD+9hJRpXmCG3EBty0C2XYRhHnlhNGnt1BTVxgavSdE6WCu3RWqHKmY
wS1c1C1Z3fPsbVwmdRPrw5095ZBzlXcAGjWYKtD1ejnryoVNwJ4Gb02DvQObVja0
WOlQf0hOSTJmT/vPg+oQ2YSiuPlj/THN+nLoARoD1jEvUxqU5fQY/FgtzP/Raoxb
dzTWACvqbRXNz+32cm091HuoblCLXCFWxIfM2kHYAoTt84kilfj2d5oC/cUpA67L
jWpiFjOROV+HYl9xsB2HbJkZVrUB5O+21ntTF32hBhmsZylcKzG7PdaggkgWWNBS
CcUwVvkpCTMIIl1On18Fk71GLC1tgG2osEVNdq76clK69wnSQKbU6/UYuYm5T64t
n3OIA2XYMt3G5vhL+C2UhaQARLER2SA3grOacZVd8Y+KE/HoZ43Rs6wapoMNP7kT
Pw3tV3DjsmOKeRE4wKBQq/Gzx0s/bbx3cIXnPzw6rqIG4h2Q9sBgXQdsc/czFkqd
/k6R1lr92Ffwk9T4Z48yrtHcnWfGihZJrw1ZEf7oX9IDvxLT8U1oaXwJTPJAPIv5
FPGikO/EUPq7UqD+pkDWZnFtPLeZ10V5PDKdwAlr1GBF3sxkZ1uquZXDpBbpFCxw
tYk6LvtpVV+M+byZt8PuzKYCv1kbLZYbIXfCTeBqFcVc3IH/3Ek3jEMbx8aM5VeV
6I3gkZxzPk/7qgJOkOgBXUyfHDizazLbEyHUALDwDWV06zs5S0ZxI5Wo49sySsow
OnWtlvW+nzxIO6gUAqcAGSO/9nLZWzmvlxgAJzn3008eaUPodoyWJXefmiAl8nCj
u1WQXktnwgvrpcVVV1GYV0GM7gZikfuaTJdDP8cEdE0FNqy3sWz+vH0gg6ukqBVl
8L921jPVpjsYn2FiEo8J1J+F6Hu0z4ROKzzUPXNu2ZjUsAL65/rxAwoBwBTP5AMA
1sjYll8Nlq+x6L+0ZXQtAiRm55TiGND6YxEzoPZSGSPri2Klf34pm3KmUipp/041
rJ0yI4XbuYPHJi1pTYqtVEdkZtHQLM163dLRjHSR5+Q=
`protect END_PROTECTED
