`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9o6VZB4+bUanViE6ub8dgNuu/BJOmB6N1598O/hY0xCIWzSgpn/NWBC9g3ipR/E2
lRyqt5Gm7Cqm0SEPY72dEoZXuoMGulJpI+evMGIpSHYDF97uROxqvb0bdam4m7s/
nlnCXOK1cLcASWYQqJ2jymFvQIIxroNpJOAtrvgD9xWvru6HT/xk4Bc83oapZ128
jMyLn13loYfc5NQ8KPKx6oNtZ1E6k9olhP8u6NN2KNZOoqCcX+mEgCPFOf7SdUUf
IVgCCfme3LYNBlQR2Utp5ssiF3nthgDQM4b/yjqMWLbUZXNrBpILqgC3B5ywpCxv
MRM0mCWa9nrTBRZzttxwCK7I7aKUNC2Zh48E4f0QPZx7UKkXai7T1kjoJQzIGDt9
TxdL38iGbwIs/0P/hPcCxyvogQGwoV/LdKEaC/Zo05HB+d+V0On9h5jNJJehI0Ry
r1BxyT0M7Yi9MmsePoRp9UCVFKxEmQxnm9dkWBEFU6RY9T5gN4zedmnb8HwNjpK4
rZF4ID+z1gB0a6zOEL+9+apyiK2X/XHcEwCHUVkN/O9gJXMM7hpxcglEPFE3phxo
Xbvwnz2SGHA/1cwOV88rLxUMufa1+8vw4Ly6YpTb0ayqYnk4rCVaaw8WyHbymatz
oW5WdiA2D6dly38VU+4YYqbsZbFGpWs9ufunXfrl7yhCbqFn8G2AYMrShLt8A8I9
ITvRcvkZiST1xDgZCgJfvZofotVJbxJQRAZdhgmvviTa8Pw784ormu0PxIj+H4Ic
rdFcLnAly55mNU4rGjnJLISm/9w2R6im6t9/ootqjAoJSH4uEh4yduUvdvlhSyDW
OGJ1xSdXXYKXjHhjWchvanmQRvUvrFiaylwQlGuO4pbh9bnWuGxj4ujZxfPXbTgt
cGFjJLzjzCN5uQFP8sFFnCrohc77OE6CBKozDOovaixtCjKYlBzY56m0cwQb9LAA
lA8Pf6LihpJy1y68qy/deQ/5Dqx4JyyPblux7HUt19E3Wfcd9hK0KDwzz8HObwSk
GsUSD2lXGPr/Q6g226Y48yya9vnrSuhRsLyp5zAoEzHDIHjLjqhOkr6cGlxh797i
tnr3LoLKAPHHLWW0/b+W2WxZpT1NKgiRvkMVXmfsPn+bZ2vJmBevHoHNrkPJOSIg
3yQq/sbN2bmjhyUQFSsN82a0jCqHmCw1A9b6p0/q0MQhEUplBN+dwxoww1Myo9Iq
ySKXTWOe8Pm+MN0bNhXSNMNvL8RTERKHvBjDEH+KojoZaw9xtgt3fxw6hZAx/4CK
n/rf4XOk3cgD0vBBHWRYiSbcjFqU9/YtsaGTKG3FJITAjgilNnXU23zZ1av4S+GS
fKFoCHQyGFfCxDyFKS++VdVGjQ59rWDFj9JyekUIWHP28gmdPJ4zZ35241PF9VMh
kVXsijPKCAI3xdGfDKBSKUha0imTJnv3hxNa1Ha20Nju6V3DkLjg2r4uhJTR2xFh
PaxjiCVREImxWwtev8mYNQ1di5B1McjtdIXrZcqCc1fnylHqyhPD3YXLcp0x3Xee
aWOzADBaNoKdFw9WPH1LR0mvtPJlc8o3ALCzR7gUKhiJQ37c/LWHOYOkf0ch/uBr
bWJRlC2Bz6e4VSMdKy/93gfr3+bt+cP+oSeNKudrsqVxrDLmOcKen5Mdut0AbBG7
UxVq+yRgC7WmZEUg8mw0twhdIF6JSlDgAe4uyCMzNaFHNak4jR/EcBj0Cpig8Zej
NCl381KYpK4ySdw246XDIydXpFwDXaT4upECAivpnZbiWKiMxDp5kr2iknKMujcj
jsi7jmKCfNVzVxpjWzU5dWvrgeZ4Lj1CLePVaDdHYaf0eaPAF+yATSLPZ6w4xLTl
o5vP7/pAuEg2o+bZJn4/boVywuTztt4qaJsTXJE1bFnMtS7h08iXVU0oYD4f6Ep5
Yu4Wosj1kHaiorJi6g/g9rV2ukYeYZ9GKjTTXLxf40FGZkKyqCiMbN7eNDAbqEp/
ibLDr2uM/yvOXxwzoLFqU5+PL5QpO6hm67RhIkalk6Jbc6vlSXLubamKVQB1vytx
49TPCmQoFxhDxIDHUx6CA42PMyvNumkQHbJwO8RyB8guhIeuL+ynxOA3d+652zI5
KTLRJ5vMIMRNhalkHVYWr9Eb16QfbKWXlhU5Pps7nZkwdWL6RixrmeUXws69re2v
QtPegL8TENxBNceMt4zAsA+KO7wNfnt4S6QCXRJ1WIdJz8tqFWX1TcYheZvajkjB
kpTw7itltBDUMrSN6basY2MwyR2ANHGfVkPZMpNsUThozmtaTDlXc4y0UEWXnIrW
EMTBzZGWIV8IpkzMWBUlhxFkDYa1lUKhsSfeQXAMbSSU383K/HF8pYSQcbng1XLU
G37vhEDAQRV0TarPQUgfyjiaI43XzPMZ78DWYqZ1qHKqwSuFTr1DuOquhv0Yre52
NYoKYloSnexVtf/4BGafyaplh0DJk0iZb7Bd4rsC6MCzGICGLZjYFGidNJFN3TEh
X5lwRAYqouakXvgqHm28qBhz1wU5iIAGqYoTzzWOCQskAJK9sQXLWdzJo3GTckl+
auUe2CkyH7PUmMWqZNSbgw/VOxbXfgH4aqkkj5RGCDcNeH0eWhVeJVTk+b++WnIs
RwZNfzQL3CupTuUW0OP5FaifkFyhuaHacaK7RfdS/Fa+Yr73Wfq5fWU+OHjRJjH6
OxoqFcMlQOIIKrKCzyS/JeolurowTtO1Xk2tl86OHpI+NEsRrLyNhhGMy8xqe949
36xfOu6jea4WEKFWPESxahWEVtJg9RUxubMQOciEJdKGdyA+t7jy6E8lUjdqhlbp
BiFyni88n8dAuF9wy+4Xz/IaveWN9N8yVyahFK9y7z+rV8VTCai1yQKOlwASvPAY
okXuevyCeIH/cEc6KlgeRh9FlGWvrz+uEbHMnPz5Tnyr86Wk3ptAORqWjoFizkoy
BxLrjGWg9OcaAWEYcUOLmpBaVJ3HAWFchCLSATeUl5IPEp5C9LxMmz1EgaRH6Obh
UE2P2GqkwSkZcNfJ276k0kViGPqdeVL21V2iYoi1XUKRXmUTqDkEyEraC8nWIJH/
8Nn8eUbd6wOq4KCsnE5dObDdksoNUGI4RyVEfhmFUpONgR3S9dKXJ/ENmVSbkLA4
Ziu1oipjLxwiMBu+kPKqKbtL2Z9Nix0eehaoNIrUJypZaqQhCg439sXFmeZyov5/
v5Ns3Isdw58dBjyPOVItxcm5vYcUhxXWMnZiX2T0V0Fhvaia8mZAck3svaxSTDOC
UnNxo4zTq8FafiBKI/1slcVN8fz0KqfxRc4IGTT2Gf+/AA2jCU8nzLf5SVC2aR2C
yUIRoWOJXkOHlgKRDKyopGwAEBIIHuJYvkqUhbPHySlBMUtOqtQ+eIJx09W3DDKK
cCKzygVV7BLyZCS/qoGcbtf7zhbb+dpTWRX55AnGN6syWfBlnzKAkKHwGwD3xzQO
c2kxWyl3AV1ixUeWGf94fLjiA91/sMc43SXQ3wavvYZPXR6ITdyxWWBzaVIJao/Q
ZGeLBL9Rk9aJQGQLkmxrZSp8XnAqxeEbIg2smWXKRjkdSoqTmBS6shrOf0jCFVBQ
UYMo9xVFfv7XPck4IbrbmE2y+ipGvdWy6c+ooMXOv7mSQpaiuNqfNhu4Dh+nILzi
L34j9T/rUtg+FApwk6l9/pXNnanbZIb0y6ok/D7spfj7sb5WFUNIWFYUMgcelRpH
VOLqNuP5k+XGq4F2HxzhWljCGx7iTKy2NugaSmy4pNspVQ5O6KfRI0tUqoh1pa4i
oLAELG+bNF6esLQphz3w/J6Y1xNrqyDUPR8zZDNe4NgBbZFvkGtPHVfBxLTwzM3d
A6EBOufmVaAMwhDcUXfnkOBHR3a7loKKaX6IMZSSLD0EOcdEXnYAGe5Wtj7y0yi0
Z291Y+LSLNOgDVTINwF9B1XRSRoANEcKs1gqCSDPam2+fHuPgDsZ2FYmz+FkbnT6
EHNinCBl64/G07uQ0YWtLuU5U8TPRKWdjhi8vhGlr0nFJKEqacyfpW4oWu95AisJ
sJb5sFOpjfHUJpiv9zJBA3RNeFJhILXPHyvD/4UI1kkQjOdBdXKo6XqFfzJQPLf3
XBo+GbKQLb3nWZcLGrAr/Eymo6bOiyCWKeHzJPZmx04R7EMnn/6DPTQx3zXmJHtl
pwCsmPyCQm5nfKQbkhYFfxpz0TpPuiwvMRAKLUddGs+kc1UZ/pH0TmvXNXDzdGw1
GRrkzCtzX8xzLWkXn5U6HPy5aP8YRywOcuXPF0GoZuIm/rbjRd5hVkVm2DhZaCM+
LvD8CsyhbsRAHsSAC/UDjlLokB1Ms4Rv+uJsB5TQePfBuR89DSBAaU22RBjKyZCC
Nd4e5VRW7exZ2bFlvXxwvyfhejvexRfHVc2T/aiC7vPAGgbpB6hsYQp4z8XjVuoc
loWwPgafLgh9vf/0Q5rJxZHczxE/7Q3U01UfpK2/9rEEw7MFQUV/LtwsWCViCbbR
RO5S6Y/FTfO2jDiO/V7txxJ4v2dxURivey/PIc5VwNdVIeMGdNVdVA1K9EBzYd++
cADKcU3bGtRt7v4h7gIh1ieH4GYQfxGPVDsJ3LJFOLbg+/a4cw7PS4i/lJM6LqMS
ZfPjCJXTHSMYApVZw1a7bm9JWla2tT7lFOAvgpgp3/YEAwr/h+8N9EgSFuNFgkdn
K575V4kLr6effprDc0v1mv2ts68NocUB5fGfs00w8iaAwMcqWCgpj2bi4CEn+yFO
aK/NnI4L/+I7IOHUIP5nq5+ybHeW3EsjfsJWg7HkdgzubCZHXZwBKv0+bFz2vZhA
ARD6FOM1pI28JeSN4e8IdwM9YiAfRj009rxXXZkgy2x9gBgPiRloypT1AB5oq9jL
7t9IGl44gyEd/lbYFmGyZdBKw5zKptgqFJAZKn/6ErK5p7ymejDsywCoiAc9y+eQ
T9vI568Quwncq+RhYy/U4TwxLHku8jgiGmxL1Kn58bec7HZ+a96oEiVrZtabLlX/
nzblURThazXOdthbqnGO46UJywtkjnGce2gwNps5UsiiVlXyeUCvIHE/LZW0PC7m
kWyCBUNfN+Axo23QuLxW9elOmzr+Nh3sDiNDtnxuQhN+pKqxeWZTijQRxday7M0f
X7Af07Xc383zhG5Dj76QehccslgDV7i8pyDzV9wjUbOtrim65av6J0KtKqE4643H
lV51tWf6gGY1Dy1vp5u20C1wSZ+LjpMYXD3ZK3cAYTSxWUHIciUsbe/gQkaVwfQ2
PMKEE3urstgj4Big51OpJbVNiBgNoZYWBPgJ31qS4KgYe0ai7xNd7hwyB7V2yLWR
jTSTfFUln0kSHaW6L5nbjULDzxGrUKOlLZdyfKHs7ENECjDT4SoaHNo+RjsuvNsz
ayqAa5kRc403SO1GIjGqdoPPDi3z0MuxIdpNlsBlqhc4rcSTIT4yqWusbQ2XgFhx
6/jkUu/wXx2zxiWhShNvPvtu5fU983eE6869mD3/cjkvbt2xrLF9Wp9afbRbqtTM
rrNA0WDAUeeMu+Neyddn171sUSbTuw60XgdS5nsfA4luDxllIFNNYZjJMfrb7tYS
U1VTw8CuY0kykIBMHorS4Wq6G5IQ6kF4E1Tts9wtBlEhKzSgmFGwgwstWN5JI/Em
A4NhYlyOYUAQPDTsJBLbyw8NsKi0sUAJ9ooP0N1vRTua9P3Agipd1cFX4a8s4Wm4
8sdY+nDlX7rcfOUhrQAFOcM0rEEX1NfZW7Ao+ppGkVMRwdYFi+6wod5uPm/Rd9SZ
AlXQKobvlTLuO1Ac1H4yAY53FK+Xt7r/RN/56vTQVxmNB4GxhKs5cG7JWpfkVEic
Ob4TehcCnukPg6dbpe1f32Ge37pgs24K6PfnRaBz4tkgAxRTt/86v8YzQie7yP+0
nZqn8cB9SWJykKRDGukHB3j/9m1A1mA2Iw/aFCUsv/dINLnF/XJhMymoOHKtsCuZ
fVfWbYNyKnRXWlRrjYnpoxdEPSj3xe0lDzUkydVKylaWIAMgdJzAMnoIe1n3jO0G
SDE6TB22LiofXAqXbobQA1VsRq9tYsvJqRZhBaZ9+D/p08xyjGJTHIVHIn22ceVd
jov3OJ1waIyrNWX4MQPwSf8cEOddXV6lhDw81vruoGlT9O9Ux+r5X4TTMCm0twiR
XgnGIZk2g2gS8aYof2OdA5jA730UZyWBBgdGsHInWfR2tVxHEmhiuoLP+7odh/vH
2WTelNFUThuOQTRreZ2fyQJhZrHKSR+KQC6iYuIb3uk19DLHGmYT21EzR8f4B0aq
0ore2SOebYenRs577PRAFhRH1VufdOwhWisE/ihv1mDHxchZBthmJ8aqaMOgijtG
x3UD6+UdaT567ZBfUNejtUdxRRvdzQLeecy/TkEOhaJop7mPzbtyD0TXOtjZtvoN
4f3Nrawn/TajaU0816xY/Gl9kzIUXzSTOkx1+2RWLoFT9TYYqUr54q58UV4n6b4z
O4RnQTJsrwCW1i+LmuVolf2R/7+SrI77Fjngj6oujALYqaXKLsZEVxQYBGrk2D6B
9y5O9YO8ZdE84MnTwnV1Trdnq0r9cniY6PPX21tz2BGN4w19OXt75dTt1o6NIs6X
NzXBrLlElUqzKP1juPSm0NHgBnqRBW8op86Igtl9vlrsWZgxmy43m5E/VPpq5lwb
e07jiifqxDl+3mqiXH8sh90BwwEAmRSYKqBCDwfIOl/N3Tv6dAg95r9kVvnrv4ZG
o0sTaS2k/rVmPSn9ELDQHee6DRF6HTe2L4BG199khm+2Gwba4nZnAD5vURqNHq9C
J89qv2mRhQSDVLsINXt9j9G7bCElV4d3N3pHzElJcry1gYATbJLfWnxe95wIxrMk
cCx9LbK75Bzdd2ot63YYUcD9r+67iyH9aYDirN4Hw2tYNY7sztteS4ngtSCUWvTG
WiPkvtQe0zxOQXoIGdF+iuSKWlh7aAEce2jrEEbh8QFs8lZ8kl1zGRZC3dLA/AhR
gUxTMH2kfy2IRauF5wiO7TravXnnri6CHXZI2mXismMGORFVQ6clewswwfZ9f3DY
pW+8B55z+9F0bK8sDFSvgVFrcbni7JDArTTrLoGzw666CffZ5d8W7rqz/P/k3vFr
ap9HUSC9kk8KqFd9AeaJRtVvYWHV328mG9ln5QmbRWpse/vPMlj8ALOPQ6AMHfbt
62dBTWR1Wf8fvvFUR6xlw0rY8833oKdwjaHoAE34Dcmfd0NZrN36kzVDoRVcrUIa
ydvDNqj03Mm3jPo+l6JrtYmKZZZEVRu69tSigtwpsXlFnRjGCz60ACpLdlzYAIaM
CS92Dn2EREDPUGvKDQMhmf/IOaGKXn8J5nWEWHJAtJDZ706brQ7t3UfdNIGHYxoO
UC6Lt7PYXzq1K7cK79+cvtv/dhE/XsL6oK0b7JD0AH+aeD1MDxakvFZu+U+NZxPo
3Hl27ppP+svGfx3CmZXRWuUl9G/T32I5Hn/JbnQhs6IODC1jvPxn0BaX+utURHqb
SMdofN51GL/6cDgYSM4Ih7UWDy6zkcbAlSUMW+nAdGs1hRj2p/bIuDi4KLwtHRe5
TC66XvUwpFmet6NIR4auRME8dW8ziVOJNqYezPjuEkpzOUCL29JC6Yr78MNy8+BB
EUwZkRawLkDYuZunyC//4frWx3nLPEnCdo65MTCo/maB8thIkhQHP8JeeeRLwvGL
+f5NZWdZHYG+D+KN64yA3Bq5q33q4r01T3a/Pv2SbfJQokw37ozuMXpCW6+JHlo+
OZ+ysjKDMlls8n3z4lIAIakTYUD5Z3ODB+5oZ598mkwwqoPL5WJxL5yZ6q3meF3r
erligvdVsBoghbNJxAoV0BGoUNtoB6Oe8mdtLtJXFnZxir0Rv0bGMm2dAmnWppNI
uQBCgpggLCZYwwfznEK4O8ot7FxI1AjzboxqvGC9NwOwFXrc/YP6EJP6IoYN+vcC
m2X/gZWXF0OHzBm+PXbKzaaBWczsW6NnSMF6PGCe98Hz94EpDwwGTnnA9k3Ai+QK
`protect END_PROTECTED
