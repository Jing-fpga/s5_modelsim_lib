`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TJ0HcDcbFH5diQsYBaQ6DETisyZfslhwFfMFLx+NsppmjLBTvxP6npKx2Lb2nW3c
wMbMVHr27nZL39o0RqQIpKN1C/TWjKCegAsgbBe4iqKV7SKLPJFQFtCZKj0aKiYi
IfRl92effLBi7nxjOcDYtVjjN5dw9rJ0g/txVqwp3qE6f2OwcoeXisnf8a4HvbAK
`protect END_PROTECTED
