`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ZPG+S7V+6QchMQkwk5GaGkFX1TjNFjHRb4YhIUKCASq2N0uG6HTM3iFxYDvJvfg
6rbF4JCw5+HAeOdYQ+/XzL9Ygv5q6xbOwB8uwAJyqG69/OaWxnaK57fzwqCGHXrl
CEkTuNaAtXZNBV4uMV7UTEOpfNlU9IQWU6fwIphrP+UbPYH4vEo9EN/zqiuzu7U3
zyn/BF2OVwG6JBVfwcQ3qEfdK554vopizxXKtOGdaufDEfx/zw2OmhrMLIFEtGuU
mkIqL8P/t+qu/kHFDzrzXQljBlpGViHKfXiJCZOCeNu0p63ZxJQ9V9tGomJPKbhE
5OQQIREzMgP5B7p/T8MEnUMhiRZknby6nczNefcKgZ/hKQHnTKMtZy5KxgRxoHou
XBOqdKSlH6AfG05OIjBX9ZYOIkyER2Ti5K7jeWG4hRx3ForA5dF+uaW9AdXvFG6V
lafIzsmBQi1gfEweDgYrMXKTAmiBF/DyfTgLvHLWq6M1dWe4jMe2ub5mufb/Thj7
`protect END_PROTECTED
