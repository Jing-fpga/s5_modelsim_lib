`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WianaCtML7gPcQeWsnbLCHvoNwfndzAxjloGPD73IaupT37bWR+r6ycg9o7L17AD
ItqIhK0W6HCxdTk0RKR5BJ1bTnk/50D5LUcF6OCbPOu7cLYECYR5+C9dhhMW+ve+
YjqEJH5s9lexbynrjBBn63M+IyXWpiMzNpDr5Pi1qZgKhPKCHm+IGKzy1gZEe7v2
hwk9txJXNCE90IjDrZ0rXVOIJsauHLZLti93rf2Dt0FEcuTla2Yg1sek9rNA827f
Up83qM7BQwGoSuyNcgdBLF81U9sHzfYKG0bo5e/P2CQJ/hHyYQalx3wvgDPgLHx5
rk7ay/Y98xHCrfxjAFUxBgu3zwsbKsa9Krzu1HzlsHfdr63POQea22uc6UBljYxQ
4HQI0iQURtogyoTBae3Dv7jgvNjJ1iFL1cLVv05dUEkGz//DVTu3/lQqESTa/fl9
RlZm70X8kbQf31gwO23ZkxgEGmWyt6uwPVd5rh4eXIPSEwJjT0EzBTsBIqEaiiWR
K1JKnap/4hze8SpvJJGcTdmWo6mdVI0LP2IF72UnzwDxvVr8SKwAZZ/UnKXMNy5E
C1rxyupAyFMWYi4wGrHBachNit7mD+Y+gffU0zII/oaczg0dnLrInc9aw+Ne/D4a
1V66DVOx4qMN6w/dUlEjLMCm5ngqrSfaRZUXTKECV38MXO5Ew2C3EPw5FSo8d/Tc
sbLG3iBdrvVv/AGB5ehosA==
`protect END_PROTECTED
