`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9X6Y2NjTx9Oa+F9USMepT3pFMEtGexFL7NNpvKngYE+65NfzneGFGMrb+qZOHbMw
S9s6CoItshWg3P/atPQ4AyD9xLNe7JiJbx/MYm1F+vmDPwdpewSEGu8NJzOfj4QB
745lsdCgkIRvcmII87xfbANhCwAGkK0l+REIguYbMfKd0fQwgWyYZnCWJ65QkfO/
tWhmha+3lH0YxoRfAfHmcGwO7fDdQjplAVdioYI0tAZY8HXdzeDe3iRflPOrY+GM
Af+Lx4uZWjidXWcPSa4zCs6xFbqEYcgu5itJb4tJurixFPhs6WeIiGiFw/vp5nlD
LGF04IreOLCmbrAbxdwS7quI9BlHYHhQsOSXDwXBEZc1IXrS1WMN0hXQCJALAxX7
ikQhswk0zvUiFRt8L2MUk2lB5Nh3ZXtFJjCEIjHYEOJtuS/oIqFmw+I/kRQR4LlV
2UZEag86CQhq8KkMDXYKcT8V7SsGloG6IgFCoaofCBCjHQjPoqZjoIc+S3xpgwgV
lVKcJ7rIa8oJ52y9z/ye2En6vQMARDQddx9Dnw8UwNO+z1E6BAhWepuMnSukj5Sq
kjYbrbkmDiwFWRYY5LivIk90m/dw9CAJ3CcCbgApw/j1i0rRIGqtXmwE824YH+Ir
Zv9sIdNB2/BuGs6lKqdNucSH/AMEVWFcuwzJrvOtXJcroR47eixsRU+jPqOEGMNF
kevRqFJ7teV0ESv9jlOjC4GGvNz4v5TSxs8A/YpMNUU+w4D04pT5ZP27MgcmM8Ep
XMHDuw5y/bXgH6SKqwbxStSxPLXjE+QgBqZa/s0izg2B+Fq0YCGKJc/H3SAy2kY8
TeiGmOP0A+gMxu4UHWKLWKB2ojSFo88616vx5nbJWh0raMN4DeWjw+rGLFt9BMYe
LC7UhdxeTwOJyU5eVa3Cy641fTvZ5N01PpFMcy5V7WBJtnDKDlubWPF+Jb5AiOBK
UZw9BfiYWNK1sbiwnmkGRCK18tS+avA+0b37SUiVPXX7c6ELS0sT89y/1T9gF7c3
Ghr+AojLHO2l8MNjw2ucnv12an3TWtGtD7y2vkCWqk5R17xFwFnYIajir6R+atNW
K9+UusQY2FjQ4f9hPUefHGkNmNzObdPru9e1PRL/pggEAZRXslQrRljRByGHsv0B
N5fDUz1xUuM3bhdwhT99mqGlb1dTz0By3JxCy8lnwy6yARyNYPoke/C7JEjBy1iz
GyCu/ENGNlGGqZjnGv3/Sq7uuJZem1v/o0caPgGw+8q0HQ9RqkrZJKsoy45ijACj
+ci5aAZ6WjbWzVCxMYd+7MIHtePYQPf58uKe3drB9Bb0IUIgZdcC87EByr8Q5AiC
AfK5DpWgtuI0O+9dN4loCMvUf08/lvPblPg7M8z6scLhjBzBAnM7pvZEUnuVx7eL
3yuoWVuNqrrb+9jwLXZc9O0f/gtakdteo4AmzHC6SxmjODxUACff7KgpDvts9Elu
VvN4D3vgaGUrIJLc7aUAbv79y/B67y69Xax5OJjdKgVjO9YDYg7O0xFWK6sgSCnb
/7x2ZjkNTn0juecck10CBOX9aV2rpMPV7PPixNuyr0ItMv5AR0D3cNpa2uB0Xy77
ASD/O5RPqGgsFZvgwMx4Ullz2G/dw1SR+zp8TGcm1utPkQltY7AIoDPkEkcLaRQo
mlXYjDligv2iqsTkFDmIKrSAbNFAYxRdOtZNvtHhHh5EL0ANuKBuJoK2Gm20EnHy
Bp3NcYVBnegPmP7SsXwQd9qQ7BbGH48WLw8P56qj93VT+LAJ+sRW0G/DVg2OMboO
ASrbukDNdH/tBzBafU4Fq11k1+bXQvDlhHSUqKI2xqyedXlPBHEwLq50Me0ZqzKe
62rqPf7meV6PNDOdgnmccOrBNU1oexAQtg93SkXD0SrO4wKnHstWwJaQ5Oy5LPuL
rscuSv3FEsARiVnbezSD1spFhQ0bT6SquSuzbj1/FLU=
`protect END_PROTECTED
