`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6aokBpKaRAg7/OxuyZmn/6TBldNx9a8mh4i4PC9CXtlMIEYe9qJuY8beujW4EMTb
qNDJSVoVkIAFCtuLyRrprvB2Ed2jMs7HwMs0z2KoA6NMbnzdJPGFx95pJjSu7hpO
fghkP07vAS01kO9R/qqORHqBnbsxkVlOlKxx6T6C/hntiijagFAq0SPVHH5IXxiN
ghs0zJ6uP0JoZhpTIEs8wxokM1mDT268OQonPWeyaMAYu3QDwHS/Kb605vBdFK9/
qfCA7CQzgRlkMat/jSVNvB+olbm5H/fSSzJAGRycQXE8pndUF3sqCvjP+Uwmhsrr
xnU2XLTVIvub853E5sA3uQUINZ9kAglu9zBMVcEOkvvmejgmKYHhzpP/JXok3k6j
8TUImF9hoDTlWG2F4aOdPun7eZiiMnpI5VbTFuR+IhZJzaniqzRrvwap4alIKRks
m+hfTdWS2qZuA258LxaJ9trO+8KHAnzx60zwvXa3S7vC/KwViBpVXVjxl+rq3j23
J/nJUAQUnNOGUSwNpOxXQe6ogi3FZ7shOAygxvt+rOWXe8UV6kVhdIbpkS8PFflU
NvuZ6s0JnNwstD9q4RSP/lNvgdezL4+B+E1t0TUPOdplxOLJjPXDBHB4zjC2D50z
zKeSYZ4e3HeQ7ii9VM846nvOzTvzCISByQpDfXbkGmprIoZ5pJoSP9cm/HRbedy6
YnVuV3g9ljLdbPt93xQIJTCl2CfEiLhTQxKjBkW31knt3JWiRCHxQTlRbmoQV8Vr
2efmNyDQD9CqlZWXTLhJGGbaVx+PHQGkPF4Yb/aG8mCwRPtP6q/bW4VcTDVbiY4q
qWEkP01zKuUN7Nvloki70tgNhPj4EiP/Lth20hBRspLMlAykOjzPxMzSkbwIJBA5
6Vde26r+HS+ZsJ5AfgeupGO1HHzqDIQVsiIS0ULPzfaLd+8CvHweS7XWPFN0MuCf
xBziOj8EasLi/MbMO28N7ouDY/yPRrQ4NjAy70XMRJBxpg6dWsZW/Btpd85xlfaD
qPSzrrQgqEpXCJzFWNXE4lMUGl5RK2UHHBv+2R/XBL+PtGbA8voMCBDcWrVE4pmZ
5/xyNLEH6zEtMz+oVClCwh+2rZRxGYz3ZQpaoSuq6/j0nfpOz5QYM8bBQbHT27dP
LF7Ttmo0gMZbZ7MopMpUPgbQ6iMeDwYulA44xBBHCpvB2273WRzQTIkTlIINmEId
e3sqDiEMyFczoIWuCkLgCfgEtOdi6J+MrlCL7mXX+iBPIxyUtNrjXYsqs/Z7QNFN
lpax1f1hR3xsCylJeLdIrMD6J0lMdqG+neCmknsHrQuGzPbFku6IzG1mBSXYOmmy
2d4MfTTeW9L8MsUlwRycvDE7ceQ6FsOc7b/bab6AZXUzhJnffhCuQmwWqK7empxs
9DlrLXv7+eUh2us3+bgw7XMUBNmVjwNdfTk24ZLDbXdCxQyI8AhfpsNTQ/SshVZt
qrPI8KXw9arP3KmmwGYLSQrehP6mhO/eRcvVr4+zRrGioG9ddK/gBvw+y2ViD5mo
645QccWsB8j+kMkMd3bmBB7JyS8odtPwheMyVjZwFkQt+R+YRpDTwFo/aWI9eKUe
9zUjYQ96161euGip6Oy52DhfC+LivoDEwsUcWuU4vOLa7QBmxG7OfAN/B9L9NRf/
uWZ88pNePK4XQwQaJuikbE08DPG3CI7IX4GQJxp+jF2MJVAOwZe7dVh3NTjccez3
KAZL5ZPNupZ4o0W9hSqo6KzzouBiJheTIK2FmiEaLVqcgYMBYboIMm8q7KIjbHh4
xRV6LChuplt2lqt6uBuPYd3OTn5OI+IkH7VxiI2VUYSjPcU2D6+MrMzR/K+wzFQU
u7P02cuBsIG4ch3pNMlnSAsVzyRFTIA0r9c3801FN8iSIF8atSY2v2t9Kil+1VhJ
GHU1m/1riI9o1EIAYoF5noRdiPe0HLYyz9YAw4In1vhjokvwG7LCVI5I3+3OI/18
tgGaSFg6Lkoy8H0nMZXkkHcRykZ4DlWZoc2hYgwkNXvmp66O3YO5NrcHlHYyh+8l
CTbgppswfEh053ma+kOHfxpndAuvRHY1Mm+ApK350/YxkbH8RzalKDFcflZSU7f4
6fKMJz29DFvlUWh3X7djhjykFh0jmSVT70K3LeQkPjeqNbb7Z3KNwknusSmNYu6F
ZOTN1TepChEBRGr8CTHrUrHUWdjNfIBBUGPCdV6MvY/bCiOZz0KZontWafzV9JY7
Cn5xyYFXFqSMFTkJ/KS0sW4OS7JfaB7dRoooYbjrv9O5T7wjDIHJSufTYDgSfggM
/Za53fAZHR0S1fw+bpPIgNZanNc3wePGI4AdXf28GLAuvOXRgLg81E04iTuqSpav
Y02zz46lTfCdL1akBRpz3SyLj8zc9LTTSYUQrkcEeL2/qRcC6FZXMaUJXfSIlaeq
wd5K5BqsA15Px/sG/A6O5ZSkepCmDmuZO8Z9SqC/bZ+KszOquRyzN7lpmrxLpK0f
PbgOhRSR7NPoNUuoELghd/Nb8X1QLF/8tgup9yQSiTu3k7VMqfb+X4FCy4+g+723
VW6DP5+3GW21OBKYX1UMP1Pdv0vChC8IfooHYXZHZvyh0UBbUjLFmJfMuf841ufY
iOFWidbLtoGCxbLQydHqBsP2tUqnmmdLD2rXMoWbAydNCZsu+iB4061Qhkbho9hH
8eIghWDXwGRo5wcOErTcI4jLhSI0xVDuLnTiMUP/NtlCLAmAbDYuqMLHIdYU1cEZ
jFq8+69yEA1ya/Zdam1qbFvf71E2rcyjgwSAOSe8s2wJ18BSLg/KHadyJPuNffHH
g1GGlKx9G3V8kd//tYg38oj8rhKTk/L5gMLa3DbST0vy9r/MUAt7KsyqXgXb9tYP
1KjT4DrETnvoyeNTvQNqlNoxnk6/ktAKJfOic8wt4RTjH9fqkyO69iBpaTnozzRS
jUQhK1BWLR4koEFwH0p44D1AC+7+21pqsLKKtLXyqCJN1/XgWJvKK9LtLsVHViK3
Ko2Ep/Ekrz9JlweAXZ3ypUgMO3DheXWcJNedYnvqEEacOjcSZQjlWK2qfwTGek+g
gn4QO7P/Q54PcPjdNvgtsAdqjuMyrMDKKdDMLVVfES6Gc/IH7acwthvVQPPMXmad
yvwqs2+ZvHwZfGDkObTxx38G9c6HGqfcc30ZS2Sn2xA40Qux+uYzm2ukB2TMMhJj
jPaft93X01ieVh2oW8adrIRuAxRKXJTdkNRsNMhDEUfa+KMOCCobBFEWRzLQDHH9
G4CZypbbVT4FTCjWjzc4NCFFGwCqguYMeh7og1RPwQoVcjRKn+D4/8SzYHHtmzY3
UEMqVj5GeNUyRm5e8Q2kvq6TFDvY6LHaBGAP/XhK/ErGw+m5xs2BjHoLol+ZleVT
XsJHPh3mmtN7bod5PDUV19IFqnNraMBSGKc50fdN3RAOuHzAEARmNrxuX8Zxc4tH
9rYvzTCS9oPqxiskjN2PgL51ieSHYn65x18HmIcb+QCMGK2SoAfV8wjTQw4+bayb
v20VONlkvTT87ICE1VmqHpUKv3jGh0yd10aYNywCfK9nBaCEtX+3osEnKwnZStul
qd1+t0+tV+J4AXH1y1ae339FzZxo09iZdJnFcspGjTkT+QdgFW4Az76YEaGjq4it
Qd9SsrWUcLWG0ry6EY9Wpqchd49M24WWY6VCbn+AlVyM83qhrcNQ2fC0PxFkXIsQ
VWcSCUBJLHqgeiunI5Eu1X2Ki2qs9MSfqEiRjdyLb+z3QHDqVVuqgDCbTsbmhkFf
wvTI5G+5Kk9Ho6wGpSeb5D8u45oNnTFIqXoYc/SGX/pUdhmeuMFWP0I3MfZSdWLs
Asry8D/s9rL5s7P1U6/fgikMPj3i/zfoY6dCt+DJJI8OO3sLV3WhvCS+dTXVb5lq
DfR/2MXHw96MwOmuG+BP3j0fRwPqzYLm/okvKpQn1yLHXu3GD1lu/TomuW2dPTGI
7YA89S/5xBQPZWIRA6pJjANaEs9/Aq644IbSoHMc20Bj3zHq6BqtOV9/IaA2sBZQ
5MLlC3wnH7yfbbKgqfrbj10t6rSsnygh3YhOug6IUBYAlEdXWU0EQx3w4uvNPcH9
ky8juHwbmMz5otrv9CWL5O9y/AB8r/CNCEEUe8ZmxbGPq02GZ5LyA3Gtgrj3M8Bn
SXTfSaAX1p5GrbZ6xCOkwMgBoBfcdJ07mCgryN9CHakxqsvJ+jWYEU/CWyplCfn1
rJHZXeTfAw0klJvpKBUlhZWovkX5fwTMGLbtLyZuH4HdF3E0AkYUYh6m1tq2O/cY
bj3k4CkliKd0BQB7ujEqF61YcqSAHqIq9QdIgH9fjMkjVORUuNkb5b5Au1s0I2g/
PYzrImHxOvV7TjJWkL39OKR6fjETublGKzEs324EtEujzbn37nX/kpSs6OP7xFc5
C0WUSAVWdBGfSdfv1GOl6iEloTltmTT3L9RTtn+8TBQTzwsIakISNv0vIfvquZ9U
h9TlbseqTdciqKifIPMttKjJAYZEQG7PLsvh5y9skvazfcZdld80qOljOBisbP/C
8Mrb+CJXjMqEdX7ZgD19CKbAhE9vmrSvXz/fMM5cLVo/YC6x6PPR3QIaXCkEFMbJ
RwcG6asX4MXwFOP5kfQoABVsZmTr1d8ghL7dXTwN4+W7nh6uxOmCNukZmJ+uoYQi
MK9KuzGPOcZpSwF+++FwDcEguP5y0sX+kHzIvcyxpdoj2foc90x3SwwbTUYLMQdR
u/r8gYBSlZnhSfmpSqb+sdBbP4CsFc9ZhuXY53VKoW7wyGC43v0KfUy6l7hCi90T
GApkhVrA6uN1beqWEBDIYdm1PmAzdZvTwdqVwNgvHjV135kG6fbz5tkA3u15k6cd
n+Vob/akJb0WVdwkTcEfcj2IXLvpLNGRoShBeBbTrKdvj69zxlBclvAZVRfHk1o1
oDTvT3lsPdTUFvZDd4TFiS+5ptX2w2TA+eeoXDwJiojDSnGATUv58p3eecNgcuM3
967eCyLUz7gv+zeUOhu1zR3sj12TSdvwKST2l81a9FBlAs2pOuQwt3cjXeXNoR5Q
R7RpZGG9tg+3BL3nxCCgwTIPfVs47orfvqEuN4ssgr+OQEXLOGukM1sq7x+2nlmH
RXvN3o2mvw6jGLli6YU4EU0CCaecfSOMwUC3GMH45F+z4SZW4bgIKiKY1MwqN+BI
gsePf9EGA2ijyfH3MrntjzdBD/WDB1nHSWHHT9CmMyEfNfGtWwQPVGuCIGN+woQU
gbknwUFbFhuXOOu2b1w67bpPFXeHy9CI4kEp+gkkYZ7c4fUnMR5uHixsMmOC+7n6
t97K0O0bKtB9eZ1d+Gy5ELCVyPINakGkYd7YkpYeykY4WxNwg62t+pYjYoSxn4KU
R6hmH7/0LTFRxylR2wxkkWjr+zRKNUSamvZ05gsySww51I9TD0yIC4AGIz9FRSxs
FoBzGBly2tvncMXPoPR+6LS2s9S66xlKo/g9lq4Q9KxE6dkuCUcaRbkdj/cBusJ3
0FUgEDmdUtdqWvBwAnwgBsPcQPvEi6oRGTpksPPi/VdaIbvOqbDy5YLrxcPUe1LF
bRzUbo4tnaCeKaqDsAxkpyD57Q6gNaXQ/0mptJ6zFaOmLDbXqFFZZ43iNtHvVwQc
Yowf2YQ0DAz39zdIuVcoQomDnabKrVzDlA60DU7Ps64RLdOLk4kHChLRsfVz0tLZ
kxwqMQLS9aUrhNG6eolRzrQ4L1zSUcgzOJtkg5945p8lCQgGVI0o79hZLZQWhlqq
OlV7PvWawfWab1zwryOQtZ07ysh9oG/sSBegue27nUu87akoer/dEyX7ohta0jHu
AXYnx4Vk8be+xH5QG2cxbP7d5+vDvwlDO50kHV1JAXyW1vKDliAtmoh+pd9F6E9F
vq+w7jq2B6jos+mBfOHn7sh23c/25SJM+C8Ad8cszNiB+67ZDECmoPFsgMGzASBY
0z3+pAhtusNIPrsCVYnxn/rjR6HPuZba0KQwasM5TT1hOddYDyQwZamUciXVPNF5
YSj+D5/AHKvsd9CocZvigDJ8e/QA9trOJAnR5tCUeNyC1WH49YdCV20NwAux3/do
scG+PW2KoUEuQxnfRbNm26fG07VnlMnTS2wDpgcxTa1zoxa8lfLV3FHfFQhAsrSi
HFUBxwQUSum1SiAHVgqcc+oUrMHmX1I9NrsAsT5Gxz/ua51FdBPhtXPbrH/2ZzD3
BSX6013PsaBWjimLUeAh2o4OKWyYp1TCEiyfELajIDT4H3V1S8x2aqmXKUf5epjQ
F71vjvWL/ydm7CxINBCM0UH7t+RcXu8h6qooc+VWaojrAZpCsNlSgj/7gyixo/bC
x76PBcV48CzM138WB6y3tRZo+oHysFFZ+kZHOBLVctvr0iz9qmqhg8rbEs8S4dnN
9bKgn6pE8HRw9YjEFgAsUyMa31QAI/xCDoXrlczLBqOVHRb4hpbIjxuv6OzgPiB+
JFW/q1XK887CnD/CxE+R7nvakzJOlzfvvu9u98eCPOcJvTODObV/Z4RaoWW6yt+p
ZEBKVxjc8+gIZpNyWObS844hw6XguOKN4nvatpU6KjKB0U+nNHh4jhypWvJyCHq8
I5piFRJ8PoBky/SdwkU0uZL/gDaZFT+ZEv33IZZVSRNXUa1DPGw5aqxaD8j2YOSt
v9rkKu7JSdJsWNW2Egh1QX802vJlfadjAylM0Z7XOMRx7pqcKe9lZPbOuUruNnEJ
cVO9Dksyl7aiz3E/h/mJGlTC1Wq4dtEGEH1iLWgJ1i5CaCVmm2itmaCdnMKyFL+h
MXej9ZqBeMrx020WHB+Z8oAKbdBhnZd6bOWPOkAa2/OXvV3HZsOzk6qDZSMxG3Wo
G7LlLgIP5hM5b5F8uOTNtov8V7EuwRSlYG+zyxAypMosLJhlu+7dvDsYOBrQWfD8
sCqJ+cPldxgLDyxo75np50U1wDu3PO0DSU/1lentdX9QHPGLLHwrKoRVF9bMat5U
ungFTdbQ+7uK/nEfg2Nrj6VC+zZmGJ8yS1Vr9aHpW65LFjOpL/lhkLTeMVm2DWYo
VSrIqsOTMLfFtRZYFotoqhiHw3hFa6lLnny3cfnh5yqHeU/44fqrrzp2I5hsIIn2
78ksNL/t/Qwx5Bk2XjJOirrAV64ja/okCauJPqWfgsS/NDliJT4WkfLoQyA5H1uW
/3qr2BTfaHFCOrVCzmzoG4CD3Yj+w10MPgpGdbkABkptJ3CKWWs+Mepto+V6VZ02
HbBJjPAM6H2BcWWDSVgW37GXmtlVkasxl7rHKRS7Xe/OMWb12h4RB14COIsftd6E
MGiG3dc8x2M1Iu+73T4CXSnRJr1WHz9rt5JgPGqIEWbwDFtiPHxspObRzZeZuc/q
i1YqB209GNtnj5vd900b59UL/OJINXRs51GPRbZ08ut9BGNtyKEaexFiwOmZn05V
e089gdRygk3BtNMYeTG0t6itvziJV8c0kKkoClKzYQRun/LEH5tbd6FszIb+khGC
SA73WArE1huF8IwFsVVzji/2e4vpAltytNZP8gwqs9csvX6vR87jWvzVONtDoPFE
SIxo42BaSj5/1htf5yhjp2sOAvFM2sM3oIewWVTiBJZEv2kV3OAt5dwEzcOfaEkP
oNW9BUVibexAoUCCZlbYpg==
`protect END_PROTECTED
