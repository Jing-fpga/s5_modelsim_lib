`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eYLjB5vwpo6eCZWF7FDJHmyUJCU+hBEeN4ru1Yr9bZEjRSxVoHprtUsw5CjXwkTs
7t5lZIZW4wxerAkYcJfWbQXCjWkuzHPV2uAXsc/eQZ47QM/m1PsiFG52VRGVFJ4S
0J2aPqFBT0Jg378vqVyNkniQTSp+dvPC0yuhLMqnmr9fDctitFN9Dgt/ZPkjdVRE
6y3W407/ZSTKhubZEiYk35h/jo4kNb26sFBdGeNsGmjNchq3905uGgX82a2nuRg6
nNFcRAOLgJVOnRs5CQZlASB5mRz/15dj44ON4LdZEOFoth4I2W+EC0jNCv+9UweP
kUzcu+xDYCHDbFJGmdqmMFLSWKgPl2xJF26Sf7qVMraZNRZa59Qax3ADTmWtlJ5L
Yjlt7NSq/YHt69nTdoakvMIhoEPnBtU6PngmT3aRyxxUbRu9OflyZGgPQnpMBJlW
5hBZCECVnL6sneZAfeVhBz1qDTMXDuivYul64zzKVf+71j4M9sZr9qdugzwj9eKA
8l4pSLAfY2TJf4y+By7xLstQDg09kAV5Kz29BzjLCwA5vRq1u9cD5h6crPsK5vUF
QLCMKbkC9pIISSuq5dMQU+Zy8C3w1llHqpRwbB7OjBt8tqVSeq4XQ8k6peZMNTN/
LsyEtUnCydPL2UCHfj0MqUqeWjbrbSFnZyPhnUVlzr9kS1RVN/71u7zENMzw5/NT
8+r2hWIFkDgaYivGUosLNzPYBX+khmiv2vDx1Sp36TwmYtyLyUEOqtA41v6TDvta
mAfoxFBgh4eDE6pI1autOOaTPgVZh+Tf3LTGNeAdVSR9ACXLOSXAkVopXDecamGa
AO/tIZd9cSwKhCikYLNA5H5s1ZLIp4eaHt4ddSTXMSBdUHw2XQxN+TFiEIxiTMEA
W4H/qMSmnYBUfQ+SuA5BrRlndafrlMhARMxKsXAjI2aN9JM9WsjjuuV/CWaWSKZU
KMCwzKHUY8v74jo92ngzf3HMFMcNdPwhXSHsyzjHZCAl6nL8C6BUqil6Y6exsDQF
HgiAKELllBj0DWVKNP5Wa38IKxNrKLnrXpPcg8dmZM9GRLGpghRiHR//05IEi0/+
r5aLLXIgva44GYCQ77u9UoppoPmevht5ecUm2xolb3E+G8EbYNuDNGTXUCdJ9Xk0
kY1sfbARi+Hzi7pq0F/aGobnCzrgg4DfgSWQQhxbaeaBetNjJe/o55FXYG7sTzje
dBro3YNy9g2dAuo9T/EB5yNrCLU1OU6eaInyvm6nqJ16fvWKqSu95NBM7OPCdauK
7nMRvmJRsZSBW1HZZwx834nupFAgPrAppVIew11P1eI5upZsEkkt0WXgjkkLfz+y
mRIzubtvnEuHBYTcO1McIUlyZoj8iJ/XHt6jr810+1meQCvVLqQi8QAnJz+Y8/UB
BkF5/GvO5bsb/DppkOnZbdgvw8bCXkHJ7S9JTeDm0hdB+oQFbxlcTxBlTd/CtbSe
teboaqn+lJPQIP9CV6ECTTM0fjXjuK142vpCQORVbUpBNWd5F6TcHjWFsMzUzQlK
Qtg7cpBoDQ4cXpyVtnJGM5GICIR4MuEnGU0Xr63k4xe6ISe0e3Ke+1GxQdoa/iLM
5iOKqr1eRVzYPBU1slhX2YTRtNNthfCQ4Cf9Gz/V5dkvXsMIOlSykI1+YIS2Ndcr
G4JQZ7jN+8EC4h50wg+c/7evoe/UUil6MLn4R9lTPI97aAqEDTlCdb6dZopbv+PR
abnzJloV5uEe6NzoUSZaMkvM69/GPiu4/QCbfM2/2mOxRZKEsTizxtJXB/R/LlsH
kyPVDYKjppX0LxZljIJyJ7h9Bvn2b7vM/N/+kRQ6zdZyGsUswVrO6QwOs3Ta/Mm0
fLCAqR3xAWze3HEluaOyNq4T7kshZiDQzLl9+Sr2dkMkySEfFYBBd4fca1/zCr1Z
25ugtSfptEs5OzkadWggi5VMxC04rJ/XII7NZv4mq3ZUp+BAvSlcSxrb0ErhoWnl
QXFRMmP4hrKiCS06wdQH9mOFNpnf3DMxUkjmLY2a3yUCVFLhAr3fdsvU7wjmKEy7
4PJbb7P3EAMZCq6yQo7a2PDjHD+eYktM0EydlYEGKm5qM9yhxMqAQovoe8gjXQu2
lS8gfSTXxIUNyCwh5XbnYNT1SZkKwK1+k23SoY47hfgVVpOGdfbF3CaM9X8PTchf
bqkq3i2UkQofWkAS7DUxWJKESgKwCp2QpolMFpdWsdapPZvYOwK/v4EOqg+0QK4M
HXWGcK/wjq8Rq/mHiiwsDeHuNk+WITu2444PB2b9JSaV9ZmeQYp9UbTdZSjQOY3w
RHALWcPOA11c2udUTxerwjJOisrZ7hq8oJPWB0DMNPY2fCLGRft2+X9wZBpv/ZR6
pk1HTRnQbrSzcMOp04I2BzGCpeCLsPv2IwPBVaXCeeHZasg2YamhoNaDgrxsXqYB
m2la0q+rEq8jQC0BeDGS0aawS/Ca+wklZL6S4332anvRVtZ/+W1E9qwnXnN30Y0i
uI52Ukt8qUDPGSpv43Ip1QFgR7gjrfHp8H/4fjOvrJif2Lx8qc2XB/z2E1tM7pfN
qD0qE31u/10v2BtqtDV+56iCNq3+Y90bHAC1laGbLIg3xjta7u1OP43M3hoOTs8M
XtXtZwRUaYw/fS8lvOwdFr3IB0KdY0Rpz7Up6xo4/UbgqbzRw9liy9ZQ67peCjXJ
mRs9V2AZQTyJIBaw5kxEHLFSa9aMiGzWkTUNNxz3Y9MkulFloIp3FhVWCxJJwDyo
DNst/ckwKmwrKQ4ymdvbRddXN05ypMDda20d6Fcpi/2hjnZ5Ra+pzy9Ycki5Cv7D
Wq+rrQoA3A8CMiuK/xMDbVuXXjuOoQ/YSQAWWd/sYuKKDEQiFQK6V7XPadKWoaLc
1W6gqJ/yKlBQ1SKpr4iFWbq23D9OWN63/QZbi7zIVkgiycCUIL5cfY7+bPYDtWpm
zggod0G5HqUS9dKQRs6qr89hZ4/hBcz91CrzKBhxo2LRkS9g+Pol1nK/jLQSn6+y
NVqRkYhR9ryN6xWBKnzw76TjTFDHmqyHakGiaHBlK9z9lT+VxTcIjZxD+9qbNEc+
ootuEZdkv/ijZ6rCuqWumeKzxKFZUx+T4ymC6camB80zEvbW93gzwmuQHs2Ke0XP
hk8rJN0rXZruYnwRFMJoILa+GwH5a+jevBonMr43wavSNifdutCtvWpiEaXN2qmZ
vjrPUTHoSlPv0tcs8bgO8NmVwt74XiQumlS3l/0DwCJehe0C55jYA1ROGMfCSlMT
jLpUtE9QBrclZ4GDRMtxLYuj87d4h3fSd4wlinvC7WuyGzKc1u9IE2NtR3zt9JiF
ZVzxt/pjuYRwrxdCUYKgjMc6CAt4Tx6/K25Ukt8GxhmnDdPzHK+lY8O4QOxQ03/l
bTl15ZSJKpb1wKHgNN0EQZYrA103lh5WjmesWJXfISNgYig/1X1KhujyyOod5o/M
wkE1STuGbqXxFOVAhSTws/b0h0E/0YBBuNuy6v1AAC1MMpNu7T6UyO2bOVe3FbKt
GXwu2BzN2d3+4SMERWEydwPT0Vw3KPKNJ4vh7P7woraoKA2Gi0a99x84kEb8ooDq
aGc3G+CtJlMMG0kzDdqCyNS+NlNFVSfuh0DIIDAcFThPNCN5X/U+UZ8dk+USqyFA
JSGPHmhiH2uQ9AApaZVhUDaFVAZeuFGdg3wt8SDwBl50tAdGMmkEnNQlqyr7THJn
MoA66PKMv/0LtMoyi567wsNipVhRKMVfwypiEUOvy7qyJ4cdsH3ZCncuXfnXUAhA
r31yn20CAfkyDGqa197jq+0olLbbjDNafJJ7UBoruDMjYYvXKOcAR6ajyh0q9Cuj
FLdMErFYWSVLT8hCvLOODfS1nbcfp89wUhWnU3DtAGSSVvvsOZNAIY724VgmYfy0
2o9h95DYRXIplfsZovD6J/A5hPFbiy6EwIyaO2qhVq4ph/CZfMKPdjNwY65Xt2KI
MqTJlbfCjTuMqJ6T5y3UX7sIP79tj8CwqiRRW1n6rw5+QqU2EPmaC9zi+LNLNKh1
KjCGhrod8iOil84BcoM63kxLHr8WpU6UmXp82s6sKmTNnREa3c6QAZkl83nSfCmy
2WGlaIrG0xq2TwfQxksG87nJYVoBS/pnybCQpAOMi9pEg3o/+ba9ZxKUsKSc4MLO
R05gfZaVxNmyqbJA3jOjhePge+Nnq/CqJfLIcYEbHMP552f7kTrWCTvnMzCqheWn
V6FX8WcUkNfAQOpdonLEMKBGGFhaVBSrfb74jhanPSZFzShnd/mNnQuUp7uf5bn9
s4o9ypuScKLsJejiRo2tU6ssbESInwvZtcFa1dh65SGD29SSxKM/de264m1NHwpW
OGa8bHLCbfMLdrI/J0TcmoAQxnl7cEYzLgtG0+MqaPPb0lc7vPns9YqTiQdtcn6l
22zwdZ3NZJ312hLhUlWY1608Kyk1jH2TF+eUuehO2toNOxmLUfkevGW+Y/OCuY9a
6Je7xY04Cp3WwfqU/sB64bx86FvhxQWmPA9/3WmUeKJO6EzhRdjCKewKt5yB2bGU
aT1fsduXMwqonNFna1/xCpjaYx4Cv1gjIyb4YRRwtHtISUh+39PPTXhVCiMmXPq6
BtBsJnXgvL6y+VIDEqy4oYNd+v1cr88InNSuANo2ke9Xtky1LlyoYFZZRGhRBAaa
5QxFPFcQR1hqbIhleI2yL4av5hoP92pYMB6N09e5GurRlaplvsDPSr5maaqh+pkR
l7G8rGDzL47C/rM0bdv1FZyax+se2qzN9gpp1h00q5b272UD967t8cCeyOlPZD7S
IKgZitNLfTAilW1gzdZ3xZZL/osWlb+REQ1xZq+2idFLLSf4PMMK6n3BpxFFQV37
XfAbXomiUVzHoXZcZC6QTIjeWkcel/8IzfyZNuA6vqaVRi1NEJB0rcPcI+zC9v3T
+txRlKgd8YNUfNJX6y9yl7Kbauf/ucDu7O5bpLwHM9Ik45qsKYvcdfV97EvhVv4r
F8jzwh5ey1Q0VUGwSACB04OCqoCnqx4E7TLxSRMM03slt0tA1g8vqDjHau6bi2eJ
ryDxylxApf7uqoxugpoyfl4rKVd7lFlxDKqvdtixe5Z0FhnZUnTAz5XBg6gAq/GI
0cZoHvx3d1gH0Ew8oGO14YYgQxO0yRHb5zt5CepilJlC3CQStu7wv+VAjKdd531h
rWuSIafyHnBgrdkjbrEvs4Xv8lP4GLRZulrZUUpFrFZOu9YAf7hRK7zoEffcwewP
77N8gVyCf9hS9NvEKE6c3hof46myXvVLs0U3suFXcqP91wKpAUWF6xrZKL5irC8F
Rw5RGkKbE2d654PtQHLt16i7xVllWGg2wd5NkwGFvm/9WX8KK7pqOvZhYqfs57WB
eredD6RAynbH7+j8fAZvsRtIoOP3jjCm0YGgPjWe0YlRotZbJP32JcopjwP6UQPl
/VMgt/tdrLyHDZpC0wajg3Lhm2PPxUwsEMcCTxUVetqtkMy/mPAVwxTMjX3PowBm
fU7p18+CzL+YMMMUO1DwfDPZJMuGwxO++dC7AQr7Am26j1jN+P6M4W5hg/wAxtZ3
OmemazDtTfk6M9eYpjCMUEKwBEEa75nhR16ZzoGMPaGBhZmAMSK73OWFEjTz6NoG
UorUHKGv/aYwJUqo+nMUdsbZcduPhSv6F/o7Amx3v6Z5alwNtZ41JGS8QvmLO8b2
sA32q6qxg9GO//P1BEtoXO+Q66TyENer5p+NEkE2140G21RFHkHFUSCxaEkzxwVv
/V/GzjXFgsuXvT1wD1rzLbIu6XlKlpqBRFDAwVIOePKCJTEU+lx1Pd7v60ksQJ9p
egvRo2En9JwsrIntVN4MrPYQaCwGO6T/Le6dZzi+rh3WObh/0std+q1Du0WS3DfU
4Ia1LRDnDvUdKvtOvO/IvWeYQf4K0S77CWlwCRiBZWP5Mc2BsA7zQlJhTApcM7Mu
yh+FpZQEgRFpvLT0w01tQab7aR6z1BEe00zeniZsX6Nzl/yQvCTjSiZE2ehobxK6
9SIAgR+ZuLtfppR8+ttRUPP0qbgWiCahoTnn1q/ngYNqnWYSvuS0Xp5qFiJ+i2xX
Y257PReCek1YWYx4+oWh5KDrgZRGPbz2a3VpF/3Z5zPM6sueQKMcN0KTljMvVVCq
hx2SeEZ8GCIIfPZfiYYpCzCUVyTv9eg6r7fevtjClPxGX6V9OQVPuLg2HW8llOY1
LQRH18CfUrpsXx1pKaQEtmKPEOH+4peGZrFe0zl0K7ZGGhqQF0ZORjlxpppMN0Z8
++fQ7rCQmhxfYNLEIMR0cEC8IL4jM3wXCBgv6/ct0BZwsG/BExyUDFng8xVGBpNm
UhDJicasCSX/NV26CIbVKK6ADh5/SVy/vSH7XJJa15VHQRaXwPL9jrCpN1qkVJYJ
rll1NOnigYjyVmBMGkbI4BvYS4Th3UsEtEoaHeWiGLjoDMhojZlDNRktBuDytfDI
pi+tkvjEALBiqbSQqSpO0HJBXwhrTBqDIPW/86ATAD6yGpsWaMg4Ej0OIQ7Kv7pp
pt2r85V9o8St4+Y0exwneTPvxrdByHezi9p2UNyp0NVIj9il8ZN4SuktuiK24HED
UG6kHPzG7fdUK9hCJTPxVJNM3AfcezLIC5U1j00hKPFGLnPdiJBhoQk+H94KtvQI
ejPzCmpciKY7l5S40wHXeV4ITQBkc9oc6SeMdITRwwjuljXxOVIZvUXbpoYFCg7D
DE5SIbCMEY9/FPCcPpBp9eNawRxfsaO130dOmstU1chRwxJb1nzbXnGb/Rl6p/Jn
9xZMQk1p3obwmnEjNsp3PrMrBhE1rOYHo5CUHhIZzD8F5Efmeh4PN4ObmMxP27ML
Zu2vdBvFgj7jDKWwr9pqkmFpUTpQdKLo4RC9ETt669AU+h98FHhDGC2SDsmJl1ch
vUaxD4WCCudXyRl93dwdB0T7mujFnkNd268FX6CnLutDWV6IxMaLPRw3gpuQoxgu
jeX2jLDA2u/I6BOvzpPFeb/l69yOF1K7SxcTWxfF/VWs++d5ZbvvOgk9m8E5SpvR
xz4GRgkqrHRXgzATfhcvuunIwZfWG+jAi4Qh2hjOJgD67d33xzV5RnbrLXk0Q4aJ
BPL9X7L3Pc7VUZGHriDYpmPxEwS8hUkGWrXAjs5TBXIBeAIFi25ChLVevnkUCE+j
FofnN82RpEWIbFyxQBhfFyhp64FuwTk2nctNqhSEzNPalfgCx3G/3JXgdWPS4k47
/8wByPlf9O48Qlc1P2ETFlr9Kye6Px0fMtLzvCeJBPYx6kRud2XUi4nwFV5iwapU
N7N91qJQQZu/Qdihr1ogaq9h0Dm/RBkjyku4eiJne8LozFksF/pnT01/wq+KmUGt
zTrKG1YZDvaLhBl2VuiXJlo8zug0TjfjMem527fMwtNjbYdhnSkMoKYwo3tHTlhh
ARryRx9yGnxbFwrvxFKj1tjRM19TL3//tm5M8Wn/CgT6eWvOdvZRWJLEvI4mOTJD
k/9zlsg+Ue7lbGyE4ZzpmoDjZgwd6pdHK0LJTMJSsEAvVR9rmdLEf1vZ4O9o/bol
l1fTSavYgXes7/EyxNImte2TPJClNR/EMohV3A7xxIUVKSUpQIXFmDF2saFu3A56
FQqYbQeNTYtD5XOoehe1Ztg/mS4+gPzHizlECJY7b9JKR1BP6OqUZglqpMtWNLnz
7UnVYgphkrNZYwL/uVQWhHoHocYsEgfUDtpJWIsyfujM8JzQm6+jc/qkDl8VOim9
ilLOboaWqZneGoq5RsAsLmZgEp3m0OtUs9YmN1RMTnwzRIOgaSqKE+X4iH/ne4Fu
P2gtX6N2kwMa8pxum+wIPxJhsHbmnvNfC5NhUvKuv7x76jVAxcvNdoJWLygWYbVf
pXVUdS3qL+rYDTiUJI0Rm1fdEo2j/F06cQPZCJQDxWHUtyq5Amq0pZzRaiSB6ecG
qo0m9VeVkYvgunBegrX+1tDF9rqzVBwU2LdOPcXwGMsu25MnhQrKOeU0PgBxQnJw
1oe8Z/LLomjGn7HC04mqSDisPuht4Vdr6DhnkU+i/9ScnNGpQFv0BIYG7OolIRJo
ImqS/ViQNmMtOy16U9vryk6slNCU1H/hoNeDFTQLiSU4akhBoXJUhnM7WwTIHf2m
OykqYXdCS06vzptGeNevAl9QYI+7Fk83RDc8jKK+9SKvUozG255SUR/261CxmNgI
C86WNc/D36odIl7DxhEj/eni8rCukqLh8KhL2KQ8Xxn5+DYnkqYc+Dqyy/xwWg3r
t6//oc7wIA4cBN+wxzKYL6WDGR+26SaJ3pawlvm+pqsArMqQgbBFZil1jELo9il5
/H4LTFJIaPVpyfO4/+RYKxb2n639eL053x1eWhTtDaT8KpHkfkQgyiPY44WCFCjZ
1fxVLO7bqMSX+wam0tVwhLmIu+BYjw1HjCVuERbNfDF6FcZd9+m5rtksIacamXNZ
tSi+cK7u3UpmkNGKmsPMZBezNeIbhnNVCqfeKVchn8hc/ZQq66AeHScQ5+VC2BdL
JeVxhf94Zi0Wm7h+qKwEoipSJpLKG6TCkjnVvZPqQUrKGBKMEP9YzdyLC188CriT
nCEG0phJJ3H0v+PasqomZzBlOcy8Z0LOVafifShf6P1MCMBJRS4bRp37nCc/5K5v
tVzRNFpPi1uCZVRznCHS+DxTMS7YuZzg7p8xtOXFCAnCeIZHFOhI15tbu1+bOs3f
h7et3ky/jrCbgzICm0WPVKTy+2VNyZHNy+0dwv3uKkfx7BGqJFuPCoECK1AOb441
bew8ZLsAGytIsvihMXbGolQLFMrZ+uVADJUg5mVqhsZvUByoUHr5T0NKbfsXBYHh
HMt9Knb1MUmfJZnjJ4OY/5yFLRg8CNVwFbS411U8V3MCO/mYZpIFPj45gERcItLd
JQG1z3k3ZMvyJyFCuj4ITKid6jc+XGHdsfH1f7SNib1t2dWhuK9WiK02xTZf1O7W
KsbGsToVkd8HAhnDLEtmFAIOHvuip6hM0KR0NjJ1P4NPC18GbiSIbKekDnTrTSl2
FoHqBuIEH6cuDyYY5PlvzGCYoTq7UvRevJlsJ6qYA/ijSVRFGgp+xAgPwUnSRUW7
rtmjX40YCZLnbf+V9nclPNdkAvYQ4fxa4wFKvjU453K12TB0pJ0X3Sw9ZEpWO/PT
volMty2C52xyQmUlNshQBKpIlg/yd6tYcXIrCTxUJYukCmOehNRsftWvYWKCmFCo
q3hSdP/KmfHaYhukzUfPElRczQL9LdEbO0UJFXMR/lzryIVAznxg0d7vaJ+MdHnA
gn3NL24hHjrDfzTYb1vLzQyLqtQog3jSI6mh6EHGpEcPOohEOu+9cAhGXLtKW5rf
qhx9qO9JWlVY/0TbUv6myjlTcwXgkjHA1Zot5M21xWk4P9mZfVTJ1cM/xDhCPTAx
28hSl5dyDOWz9owfSxsUFl07sfxVSoazTg9tChSA1UtOJRe6c0yKroRQM0vZtSUa
MmNgwDWXv4K16MbG/7DXZ9atDa2+SfQLUdqAm956LyyI8/aqnjs02BVZBRyqIOD5
5Rajv8leZ7PsFuKZfSw0uwgcDVrEjrr1nkHEqkL8S1JAd3FowZZ8GQlgT6tV4P7q
9+X4uTRrO0o1XVohifzFavpSPZAhVskIfePAzd9xweqDFDS6uECaCRqT3YO8DPUb
Vo3GdYIXMTxUmkjLgOOrB2V0ghU4fVQzUCPW32JgvNia+eT/xuqpQEA6Vs5IpkD0
nm1qtC1lKfn0kweY/h1pB8PRqNnCm0fbh0xW+NHT92bYAgp4EtxXF2lZsF3G8vh7
ghljbTs11VgZktGfyMkPyd2ZZ/Un1N9PCcf0WIC8smzOyhmfZHxfAXCplLOignvq
39lebJWSUSBhpBQrd71xuGO1B1+qMh2PY3Ml9YV2Y0hkHnkvuSVZQYl4RQubUSCx
w34IwvoVSqGBoyoNSB7W+84DpqSftTAQhLRarEBsvmydE+1A2KovXx5R+GKmcjze
lJG8ONWrEFh2ALtdnbOgeLx/ZC/3VzqGKjwnQ991cDwU+ekH4EQQmIC2AjAh6s8Q
O2zBCByc1+SGGCLDIqPHQ+EuXeUf9WqNV0wLe3Gzmku4o1PPz2LsFS522FpTmiUX
vq0/aKxn7eng4tC2Vkal6EFvdd/tmaAvfM7MOAbytEAdC4KxAIDGr5xDsjwab7ex
Wz1YR830u2wLfJLgfe088MAg4xDVrk/dqSsLuv+8wmlQ0lp+SfYEFvsUzaWAyPCK
4+6SHmC/PLIbUkw7k5rTkH2hlqdSF2nDWzt0XjF04lTEu5PyUX3Bjzyo887a8Wte
9UWG88C3hGDYZYr6fXH9Jn0d+vMzGvvIeKFAgFy9p7CdaQ55wbHHmUrrXmHwM08k
HFEh+huzSfopygjdrvx8oeTdHrC/PbXO3/Ow7Ikxw/bEBnFAtZwwfp+3qHXxscaS
RwiBSL4dMHWDrur0jYD3DAhNFk0DRaFDmdQUzE5Sr7ovsf9Pjqaxch8gThgqeY5D
RD5hvpoQmZ4nMp1N+usDnmx8SyEPCHnLJBcivTEQsVraPuLK+lOWom+qImZyBNOI
x9OSDyrd0DwCnZZ5nu4U7gaH4lgi4J2mEs8EFOEge80i+KiLwOlK9yrsQEe4WVHD
TQua1p1JtmzysbcOAxER1J4Iu0UATWMW+8vSNv7RhLtYv01rU9srsgxAtHzy1ZOH
/HKNlsmEBx37clz9PnGt2iAnDG6bScjR6m4SiU3/xvXJZcHKwofRU5e6rAdBmPJy
YjjTXX6QQhII+WR4JdphWB5Hxq2+k1ibKcRpic3PZbrriUAf9wvhrhdaT1IE03gm
7cE59TQJDA2uJ+u1ce46VXf0Xmwg54CBGpy36UIsXvbEJYjc5zta25TzB24W+QCn
+vTEQ3ROuY3tgyHdvqJVmK1TdwfKceq6Os5WYNOTKZKaddKjBKR6L9NAbJfqV1ga
PJ7g4KsVpFvUjawocJ44pZG2lSpsAhCWH2guaAZ4tg3+ISMX6WlohObS9ufq4dqQ
jQFaLhC88kfVEc61ZyxvcsxXNzhnyBSKLbAm89BTsYI0Ms7B2jH4xaOCZKsDFUd9
y3j9MEKK9HdUNsgXKgPBdHjrygZmI9k0cQn4DF/P2wJqveHVa+yEWeYFJJ9W9j9z
DenaeSUTqN/1wD5fDe9x4+KtPBOeOCWzYfAkT+sONUsqQEnjtY0p/5uw7TuWSO0q
/5MSTX9XVqM0NrBNoiyMA/cJCGWSgAcr/e2jz/NXu8t1zE+mOJZYF4owmn+xQ+Sn
5Pl+gbsjA349DgOTn1+b8sm7NISh6AraS0qelIckNVOI02xG1L39BVGZm68dTEqC
LPvZTochMD0Gkc0q55YUbV1Ea90fjr/+5G3DefW30+R+UWVGD3vZ2W9d3quh5eYI
XLPWc5LGz8KuK+NpgtRCkt6dY5g3a57gDs0AO+LAXwUZ2RvjqvVJdy652YnKO9C9
6wajiCKJHB+UbNem7kbuP9oC+qtbasyuEm2Mc1zyYgZq8FYwkfjT5MDYOIliPhuc
sa/2ojXcIOpGIte4anbzECanos6pzLpjNb75HzQ1MRG4NT/2ASXg5YMZjP8/t3Rb
oz9VKSM1WUuR1vI1l0+1ayKcU8wFXGiT1D9iwLHp5pVoHZT7IKgaf4u2E77om980
IoWg+gIoAQyitZTFOI75W1v99sjrVh0TqMlv3KRSQj/mjtVLaI0Hk57M/Md1xjvX
IDre25iFnwDqCGFLbcBEPbmUvEW2pr/tD6YAxjREPN2+QYacgSFkEq7a3QGM+rs4
SdSPZDik4ssyxmsubiaqLo/ae5HATC3IV5CgvlcueQaY/E3PDQHGXwSy20DE0o9E
yARd/t5oz/APE17ZcztPM/ttYumtuyeKruGHLaa18hxoxfmkieS1HPhXDsiBRW96
bmhmghxOvL4sTS/ut8m6/zeVFyHd7K+imppnJJlW30TEaZt5MQ0oPePGXC3xxQiQ
jwmqBcW+4PcV7ui94C9UVzieDnVFV6eymPIxBNMw4iJJgWAilDatx/ghGDIH54C4
ztCsVuyPKB/C8lMeJyj+pwvsSbwTRQIZv/eSiX0YPYK6RhYaUUkcGrIAWR6LExEk
fidczIyr0q6AIVw0QKkQK5TX+S6OAdUiBHUIaV3w90W2SqWxTevnlXB/9eMtLLBZ
AQ57dEB2HlG2Zk3KRO5tVjAVK0uS3IGACeEmQ+TGiAUVejCoLm1KroXpL32GGZQf
E1sy501YQTJdLJ4SYQ5bC78QaJxsFwFQjwFvl/axviNrF5cSQ8xFmAxZRczqVwYw
RvxuFLL6KksAZsOa9EGCnGG+0x8jzHBZe5CYm3VFK9k5E6tnfkpRKwC6hX1O/NEQ
RU+fJBQqR7JO8NXgknNzwyApHD30KmEYjPkhnT+WpzbN7/Pc+Dvw0CS6uyWEgRRA
SoF5nEzPsoN5JLw2YfbU5dMOtSgNjweWj8yLAe3xydQKDh9dPHmD5sbEepYNsQcN
0eFWG7Q2WsLZb3EF70qpa8n9X0t/cn6UGVwugpBVvK1G6Od5DEm2D/YP0TS7cMPa
EuDYPcwZGrBxJrAxPuqpwXzzbhsvGg6+bmVJ1lZuNFHuZUQKWMeB+wOZKrhtFNyl
cua0HWY+71YxxSjb2I8a8OoYcVTHuOcm0vR+wSMKqcKZCqXreGw+9YJPSGY+gKG5
g4AjekksDXYBG3aXmSgty8Zm6f6Va8Q8FAL3VOXKLZWoLI/nbNWuBiDMpnXb1oU2
4YlL4LTZA+JHOmLLRD3ceLlwmlJ7B4MkCf3d+UoECH0xCjKvjxpi4gVzTmexz3RM
7rOFrvZvO28fgMKfsr9upEs8Sm8ZLoCzbzjpKV3vwcIFB9IlFq35e51KiRtjiwbV
1Czc9gmXjC9vF7dk2balG8y3LcP/vXD1QHbXWmdkUrleaMj3kVEfSO0QYixUu5IH
kw+6lSTk9OgyPqk0ovdffUsOATKDXLJUcfzeX8sKXx8LRbqB7EEmumqpWPKRJwC8
jCq9kZ8fmdldgpjw5U9/eR1fQYol4f/8Jn9GT6U2MKoKR2d+yhr6CXSPB3DrmkjY
O8kUsMzR2Nq3+n3pv1HriuKKhnbR4hW4egonIrQud6EpmRHol/EpI5iXanCyIarV
zvr7mNPHybjmjakMmDNNXTuaeTfcufeDWLyoKUehZ4KufCdIndIot1LHmMqEuE/2
tSA19C7HamAIZOZELFzilIo0RDPVvDcGA0FpfWOaKbK2x4PP4qs/N8JuDNynFV6i
Xt4z7O5J6Wkk9oQeVRlyOubTJK/+fWP+2gr7KrzcU7XDwy8Tf+9Ey7fxslJLxY0b
ngFJdBpTeFiTpJfaToN+N9Pzj6Ka8kHlDXT+3s0ACagMQYmk+f0RYpM47K1XUeEo
kFvZk27EO2G5BM8yoF1LdbA4GCNeukvnVY973bqQvBBc1JUHK9kC8CenSjlRRhQa
h94WCzz5aoER4V0FQ78E2P+DldEhyLsfnSHwrWEjZMFwBQJ7ciA/wWuA2NJydsx+
TpPkbLdYFfwARjsoSLw6Sdfyan8ZUINx3jvFbX3CwN432lssih25pCTQ7xVmdbAl
y9WQOqW9yN+tWRu0RH81o0S6ypoEH6kEQSyCa6459aiBcjFPE2Ssf5Kg0F8O/47B
JTH8VKp3zKhaJCtBZsbRhuwYMlQmt6JmKGGUF/GqIvIdZ4CzwYBSY7Qabg7jfG38
/vN44QaiUxuKXKzya0MTyHtW0exYCa9HUIJ/qnt12UP2LL0t/Egr5hvByOVvJ3lh
0PxXQdjko++TDWLHG8tfEH/k4DCAPA7W4dSKMLrminQn43cttNyvEsAZ1MUv2tEK
R+qQb558uCZ9vO1QClX1O49X7MZRtJVtGCei1GQ02yikUvxHxlHlimo7wKe0Wo4d
c7/OCjSA0Ky7PDwagMtsp5hEPvRIG/DlgumX1dopF8KvnaQ+ryX6GcUxJ61F+PB7
cIc96iDjx6v7A5vY5QlLnwPOlxFquZfFyQ7CNBZSk2IKlltgUNX2JPlhdBZFJB+r
rWT+Aa+8+pe/F1nNQy9fg9QWFKu4jbUI1SaMS1lvcH+5Ua9wg/+tpvNa37WPQA4O
dXhZ2B6WR0FoMEqEWFNsu+BzoioxoZGYH76N6mrvwO8ViRnghzKhT5XgsBA9Ihhh
aDLXh6xxARaqBErJviGe2W0lR0tXVu6ygqExVFs3nA9owiNdEYSvN/V2IAKaxja9
tthDcF/05U+bd0AYvhBBILtBB2FqfffvL2kSWj2WQLhEZY5VVWihtXOzPDbQkb5J
8jlg1Sn0WOSOdGs2ikkpoWnqEHmftcrAikshWqlwhdcfjHzNvgVz32sWVTNRjAmd
tied/jHRS5s+TwWP+0wyDGedDh4U9xjyHYEMC75hOZ6H5sZ7Crf8yYk5QKWGGhID
ACpEbugWrhqhGq1EjnlhH0wWrl4XsJcE9QuCVxII8PvOKxS/KwTJN4QneQQ8rGMb
ztopP5jICGgTzODHDK+lPbiEZ4NDdsmsag2ZNYZX4bT4F8gkaJTHFFwY3wCfk7z7
DqUR/nJujqoMLOhWv/aULgra1ytTM5D5pnjrbAjcye1UTUrRrT6IOr3i3ZOmAmbY
rsN8TxVi4qwdoBSYpKClV6lIatC4KHHPk6AWUJ0Tk0Wpn3rXhnIbh4nJQ+9sAviI
YNIp+AMC9dwyVoeeh+KtT/ahR3Aba6E0mPUHxzviSlIMxoTdqk8SjpV+SppmatsN
k/sTslfeZwh917zt0yp21WoER0OwYE5bmejAAycPUxrHWvaImtpiifN24NqUQI+5
Z3tMPf6ithb3Z5o9QRifOvOH9gUQtkOrNOLhOBR+kDv1mQFHFhWezP7JyQ+DGhIE
EqU3LPsjeeFDd8cuJmntDBUjbknL7vXbalWGPaliM/3AhQz9ajDK9ZMKM/wNxeiD
c2oHwxMwyc+RiDYK7YSyXq0HL5hAhjcNxnsr/SMM/3Itoja5cXWv7MKk52mb05BE
tAccrGfsM+t2U4ShUeNQfdfnf853sqsAvuu8IiswZUe5U8PfAuI0TGFW8uOD74Ve
ullZNl/8v7Asx4ggj98WvI2deSdAlnzDXqmLDJyTzfQ=
`protect END_PROTECTED
