`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
waSInq8NyXwE9odWsuKqiEp1PQqP8tnEfVLxEIkvC3+UJ0VtYLW25wA/2YVYkj4+
8IaxgrQvEeUqI9ImyyEl6Ps6UQSmMsIUlfH2Zd99FymBZZKUuYDAIdCUdI0TyL5Q
/TPa4VkqsBTsGsyTEk4WDUCErDvf7AjfNnX/WkJ/TsCKUHl9f8sKY4ZZZF0Gz5cm
PywBtFxzMdzxuw9kvTSPVPB0wnjUZxadT/728vZaGUuGuqGhP97k/diGFlSMrsl/
ZWjWm1lygN3VvgroXyCPHcpeSi4l0FYmwQXSmuLB1SmkwXPpk2MiqVmwFPJozCvj
/UR1XPRjXrUkG+baT4FgrqKb9vw3+Pe/wYG7AdZ5UMJQfgP7nI+t3MRNuVNe+D/Q
NnK5wwyo5NM1H9236htxgXDyLGjXnSEK+0T20BejiaLCg08zixo5p1dHhXtzf1OH
S45rNwzd7O3xTSMc5CzYTdjQgWNPsPhOKM7GAqUy3xqToHRrUV4Ac60JiO6pmV3C
/kc8mDPR2VEFgJJNO9oFil9/+xkXYQcoaR50Vo7QSnF85oawXM4asex5nxIwhW1E
z9IpAsylhswDzSYa1hN2pi0wM1r5qSjehFi1Y862/6tVzwj0wKCj4WPbL7KcuYca
HlRuW218dhWr9iTsR+AFawT/8i5kyavMK7DAo0/zrzpN0mxJTFsuJQD7aLC6JwOr
BWElNvTG40BqahxpqQIVoxOttuLxyZwSX1gG1UgYyM2uUqUXqump1L/Nu2Y5KTwG
prSjZDGn7gnbpLPy1VzGbH0tE/ul1Ttv6UHQKGBPDYwCwfGz9VsBm5wFNFoFvzQo
/XrAYiqvmWG/OyMCRxyMSd97MoDR12VOGEMqVu8Quc4SIvijn4usPfvb7w10FMif
shaaeIL7TrhQ29i8Rl3hYHGt5xfZYInvNvIVycPVovWBHHDcx+zIZWObPg85FQ4P
5YK57JTRJXz9c9C+UXZSt5NKc9Gn9oY6pQpKMq0nQWyXbKMjRfqfPkb4LI94sJHB
wpAscgqrEA1f+rAzLGz05/7428jXZCle/h2F5JXX+ksu7M4GXr+vR0lL9fxMsYAT
H9JDaFVCgR8gnB/7N1YNjsM2xom+tiS58Ey58NPLVyeQ9Vc/Oivqxv6WTJgpEgoA
N3A1i9HBOf0Tcu22Fnfjc0HcTUGwQ9UaB8s4TNL7k5zAb8NFgB+T6iEXOVZ1wKPr
dKbe1lYQXhXCQl6/rLt4DFtYNgZMOLObnZmJhAqxobDaVwoJ5z14c1Q3f+mWNkYk
I+YucQqNh5pWGXnWBVveW6UadVFBCISDDLS9Yh9gnUQlGDSEpI3rwBhOcmEhHJ1B
PRAtLcyEPLbBJQrh4gkwv2MsXhrmNmcjknsOjuPhfCmbEnAleeMfn45iOF032Wjh
3+saRxNmaFf9Pgd/dGsOLKdv/NHr3ETG3OT2GurMSgB8J8WadQqLCyVJF/NKCH4b
RN0c5qImnut1n1CkhFC5tQR2RKZlQTj7MEBRQWkPADfuGARd4NOYsMwyBu1yX7ez
KH9y8ITR347C4wTOrZx84pfrSP/Be0baBTwnJI5faMFaOVG/lYeB66RWe2jXCzPw
sPoszkUSk7uRQ9GX9tXmFMXLJyzIEQUshaoZhrxIMV7MJPQikZ6gHGMd74xfxKxT
V9/DTNMQ4aW9oO5DkQGSefEJQN4vzhWsGCQbag4z3BkDc6LqjNRqihYxtzB77mMa
ezetZ/u9smw+BHkqKWUzzm6Nuih6sFzZks+yiyEKfwi/eMoJcnURdo6jyDhkxAvC
8tTuynwgxxwVk6tG5UO4er8yFfGohCZ8teiR0zXCN+Sb2EONPzNnYsTW2opZlQIt
/AVcR+6pvrRDYSHV7HZaZAA2TI5b4gpEznm6+vBbWLg+G96aw+x01fSMakmayJJh
UsiPLo4CLEPXA/T84iemKQoraqoPBv5HEhtpLXtDqVsjemkkd5QOGE+sncgxf2+/
rheteRjvq7sBpM0WMnSkw5G2nt+O/JPIq2OD0+7z6PDwaLHlv8cQ2EFVIRMZH3PK
nq8E51mUmBu645fqwvzoCtwur6BhZK+QqcvSk9KDtETW4Pi3JPTbNBobKJtZvs6o
v7rv3BLIU6Wi/+IllqGGY3YosBLlmzEFD3szzfaBJ+95lgSHIkbCgHhvbytRAV52
vOa5i1SqGW5OTcC9gYeta4g/UioGYf8IfosVsxMsaDy8LMBs4UH7xFGPT4LBWY4p
E+Ks0NsMbo3bOlO1ETvPvF4NSa6JBTSLWEmAxTLl57mUzqZIoVycunVC4uVb316Q
fsFEmCwXGOj2z+jFWYsBcXmrUeZuSceIWzeVNLfxFxUlKDG9+FtqnXdYNorpxMmJ
iE0/8weCCvXsrnXJTdA/hI4ZqKJyRQDn3z6G5nSBsRV0x21BaMQ06AVFbV7L05/W
tJXp8qdXjXbCle0A6bHDvrdCxlwAVbfjLhp9x12wIZagj+yuq/sR/sVM+Foc4f64
SchrTCAOX3VYv0nAs6muL/2lcaGxScHHhQ/+ly5sHRsq7fbPa8hbCWzlZft/nO5g
wgavLDKewXpFtc2sPg/Zq78eSANSeaG9GQtYBOirygk8bIUSFLxKCFDwUUzLvnjp
f4S7KmikpPxvUViC9don0Kxu1/HcdfRQauDAT3YbrpSKdQHuD3ac/sVZLKD5GDBQ
+JSCcm1joPMo+zX8YAxdbH6tX7F3d+KhjfmtNVkSAk6T0OhkCSKj1EuQ2x/hAN6z
AB4MJvT+/UjQUAmAI4aZZIaa1+nV1+L7BQK5OecYD0zGeu7TZRKyWN8RjGtpc9zH
Plhxwh0QFlnHHcgP42pN64fgYFssGzN0nPEnolY1mqYBxEMo3EhcvO881jq+5oZa
jrxnBJhWHbscGKdD8c+UKZwsqTgrDnEcF08FbkwA9qmvZ/beuyZkNfEQ8GtI0KJq
IsXEuTeoTS2WQgwabQza1aF+nt4yEV9SDb8cVmkja1Q97wzP6HwYmprv1hTLaqut
elM2FfUf9glh/3dSj5pnp2L4B4DH69UT6/vdE3zKVnA0z2dGe0enRq1EC9GNNNP3
VitKTXZ2amQF4LERiSuIi2I3D8jf8f6KfInfHPMiDTbNs6Okkfxq67Ykj8d/VYZE
N5nDAWkRlyXKNqRV3UOgmVBkSTmMjRRNb1VA1825JJcE+LatYW1Vx4IXnZPAFQnA
4XRu+Q9wDNH/V23Y1H2E0fEDP296K4VqJVJMfLykeJIw/651tL/jdc6fwS09oSRf
ZJ/697eGD1MsV1KDILlM765/ZHFYphdMlk2jsDRiAUJRQ48lf/ryz1vNf83na2Be
SBcD+rz8Qj2ymcgEpfCjoFexTojtrskO6AsJwjhhvbM9RoMl15gqltBIiUzt34XM
prEyhDzeyljwobq+K6ehEZ/FwT/6xdF8t83eS3t6FYRVoNBXre7JDoVJWEpXttnD
GmAx2SGOi2nyhRAX/l8CjkQ7HQPuYIyfTTSds4zaiEJuvh4vAU863hwxiEcoWnP5
eC6G8hVu7ZaB5xHBy7PS4jK3Xp9w+Rf5MVne6IgpfLZFbOn9+l5Q6uCFoVHsxoki
a7snd701Ng6Al6n4X6sE+RiMWan9+tZv/to2L9KbEE28CzLUtKL/aZ0ULfN5k/XR
a0JKWRj9scXHN/qvXMRF9URsFWLH2yk1xO6B29DpxBnFehXBPa8s9iyOR6mA+Yt1
22eJ6RDVZnH8YxoIAxgaK2YySpqSXHXaeEVruPbHQx5rP7acvd3IZ2mBq89IZj1T
lhTsvW5qDF9YvAzH2TuE/SjZFKB64Mjw3ZCqiN/WKVsMPdDofj7xJRyKkfsWmtF5
+q91mmE/MgefmO6jYALNfqXj4M7KlbT+uXSb8qDdH9imkNEkaMpqXPzIbWmJzVpe
Qk92SP0BCPnA10Tt3tYjg1GGH5+XZFi07dV62UMVXshF0da9cue1SWuR+RMk3BK/
A5DTt6P5xlwEs+36ucN8necNyEW2tPe7vyjlB3Q9vwHM60BOP1HNglrnSLS/XJtT
wpyVk/ubnx0Ug2HbA6Q6FRj2mPFU8GU76eoqTtIpuGU=
`protect END_PROTECTED
