`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FaHqsV3fulRMkDC9666kWO9xN0oY9vm342+j1EPwsQMtoOIUgyuPbday7HJ5jJSM
vHS1J5xI95t9TNuXIIUSSEumn207f4JJB4GviczGS/GO55cxNbxaXkYD9EIVHthB
C52WXXhGNpKGqaZbxAeAqW1o8bgR0xn0+WTJrDjaiwJznWkHBXIksH/S15Di2699
cZUlYjsZWRD8WLDvbdcxO0fh8p5vMknnfIvwq955yDPd4Je9VpqwmW4PvX9gYhq8
87/lBaQ5+25FeCy/IH7BJcX8fFip1OVR7OWIL0F2prO2ZLahFYhOM89TJ9WdsBGT
auXLKChxjPzReWXXLCuCylZfGaZfbitzLzZW18/JqBgAuSle9gEm68XtEUJZh9ns
1vHb9+6I4jweGgYpcBnwXuptHWxzbwaYeuW2YfjyJkaHFrK0R26j/xb+gM6bQDAI
rGGzpE7pcKSwA3EHJRpGG6GvxFcPCE9ejCYyqIjaowWgH7C+SmEwK8gTwNNFUa7S
YR4pjeWB8fiHeYViRkJu7OBSLWeSDU+VglNbBQt8NR2PchnAn+aOLmcUtpgx2Jg+
vAjQwTg4notOKkjAIxr0lH2J8oH9dSYwlgxqQee80GLnRzA8oSgjNkPRyJ6YJzeC
HrywarNjv3cAWyEbUPQpGA1Wbtf1xjmdS525IT7xMK6u5hdXV6ZFEAzFw+JRjSWa
jAeILihc8F7AVfR/JSztaofRHX2PK7DEhYA585BH85fHTY2ihALPo8G1m7J8O9Fa
MKY0IEF98v01lp3Z81YZtkxThwccXAq+WEk3Cc6MPIacVmngDx/6Z8RexjcNQHd/
0ycdIX6UHN+sYdci/zKl2dDiDTx5jQCKdQpnhwSRyDqHrqccKXUgHPRbXg8JtNmq
rHYHOBpdNPHpKLrvIS+CliL7n+ZUQz9PqBEtbwFCODSd4K2Q6ZykURTWpP1OUDLF
wLQ718Z1fMf+Bh7MC6rMMcIZyIoxVdmnwtfn83aQv+bN+vlFVxA3FKvUb0mjCUGC
19IcqkBqdBRRNaCYKnGljQ2lJ+B9ak9KqH3NzL5knBcU4Jz6vswl/+F+OZgWg9k9
FF1qWTR1JPdmKns3KHEdJwcsQhDdFAmW0YGRDaPjwgFt9qllGTLPSTg1CF6+IwZ7
+LCJT0qa4or8R17544WE77vJSPEjifqZ/n9oEKkWL1essazaOixtZ4Be8O7qU94g
jGIJYMlsXXqH2fx4kkAHicml+BfC/ZhL0QXU01Xnrr38BIiePvDS+hVtLDZ24aR4
TF+OeDvait9SZvJ1pQowVRdBJDbEaBpsZ8hhlxcnkTKyFGzucQDxBU04DR4GqyMM
yVsrjdcNWVfNYnuQ0aJ3SCjpdLjM6l03xd8WzYDfYIdlvBCnBlCRAmu/XLAJNKyl
/XwR6M3t/DwT3g2CB8RiX4fMw/9PGTHE9r0Tg2/OEQw+xHBPX0O7td8j5aIcw2ft
rSSw5kLHvsSCGGAbNq9Jhg6V/m2rDC8H0VYNBfUaHfpW6QftXsAw71/KOc01FvDq
p7HaaQsvQReVT/B3aS967qreWL0H53x2T1eZIE9p5yO0IIADDXkrMro9oS+dQ5E9
5SoSU/fXd6OkQegUYTHV7ExIXazGWt5uzH8nYGC1v1jt0bRT62Amb3KORtrG7rqK
HDq8y7PeFH1lbUwhSeKyYGhC5cUjrl597oSAEo3y7nPc0kihX3veTn3GhQEHjD0l
vm+5ITdDYacPIbq4jpVwvkwuKW0htAr5sIlzxSzmzSuR9pgjDDCyMlWC1e717adH
ANtkntag6/EWBl82S55A7JYruxGvqio8R0kNm4otQsrTf0uPZELaEUnLCi2+QRgU
cQEpuvNhJQdDFRnBeGqn2juNUrs16kbmzGMWlIGT6KI+dmmGzwlKycoDTpbwhr/j
VR7EpBw8PI2yvO6YQbX55UYRfG10eU+OlZFYaNT7vvXrFWlTzyo95W1at78xZDyK
if+ZnV28ORb6wU3ZkuP6EOmOotlD5noUNSmEqMhoNDun4JFpq40M/JzKN80nfSqf
MtndtEZum+wohnNjNrpyQNWZ+jT36FOIyaB9d0ja8Cmhf15a/QiL5BOY0tQ3olxI
kBF1hpng6l71J+WBkQBe9Ow42LCtNi0m0D3Om1vE5YY=
`protect END_PROTECTED
