`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vQVqnh1Lu+KtPUnUaPwN3kGgWqR85dLW+LNUoyDXAw4eEhJ/HaHfIODyDlThgZi6
Wcmzsd/Jkul9BywTfbYUzGXLz2MiaFInFBuLmwW+5WXAfagUxZBGBRd6M/WC+3XA
vs26pRytMMOy9p+WvEBprbNCvNepg9gKjziqhAftaI9qGBYtSHBYG90v/9c9W8zj
Giy+gQAwBGgxmOMAC7+hXQ9zw6LaEMf8hnft67MnURVlwUpfzC6SuTjRkjWuhNA3
PXOanZ3iOr9BRgI3hg8MHvN0XhHBKppkmC42KOGe39vtJDL8GhdUGbB7QK0RlECH
MeL8E8VJDiMGnD3aKSyCJ6s1/diy6oytIAuM1gpVc9wnfaJ8rOO2B3oLZDw2wVZs
U/6jjYPN6V6Eni2qdV04sKUXElp7sAJ9k3KPmOonkmIReC7gqJG9i5KsZhtaIlp3
mnm2y3mp9pYKSxDvLdloOnL73QNFvxQkJK2u4znxkGzNgp2AqvGXLvtWA/q2jDLV
U69M/3vCV9EQqzcNkHZA2FQ47+ALqiYZzaURPz/8FnMiKVZajgZtDO62D8mbQhoK
/ljy8Y/fq+OMEadLRLlBB2HLYJENY02mVlaV2dQe+OtONCbUSHKq4LQRBnypZcy8
0lq3DsdI75DFno2o/dRtJq/u+XlMwAfIkf6xI21iOK6v/MTwRT+kEVW0fHECuYay
Gw4jqqOFIsAaGeNAWXJTml7pJTpRpPOIwaA5WaTwIvLf12VJtP99D1QU/8vpR+G7
6ZxiO/Bncz8jZc0H18DTH7jb9ra2fR1HcTv8sTFRoIrhUbJmn99lelXewxzHQxZY
0ZvHrANC0r/fOmtNtHzIYEyy8BjP/rgj39KI/Z3rqv71biOC8EYoAVVTBsgL3yvo
jBkn2XP96MkfGca/HNA2w+rYW9CuHzU+pmeHGIlGqvOq3AA1FZZSNcO4HE0butH4
sNa8Rl6Gnbpxh3VYXbc8vRvS+KSWHV/ta+HrVudy/d1UoMDiLbvnmbhzTgd7fVWQ
GjZe4w7ARygSybUnRShgQshwbTIskHxokS3yn/0wWtmG/P8cxv++WSszoKHWeE7d
bnNQX9vHCJst1fnxcKSAKPl5sYHhCb2ZNRf7XgDMxwm2nYuOYtyr7DgDv91ImGDZ
7Q9WCTBhvT3zhXRip5rsv8AFHFpwqBBGmjreEbPqU+v6F500sjBqJCKPVzDC0eVb
OiBhx99zIqIV9YlpNMvRM6o1iN2LURYjh+sjQ7BQF6HqCh/t6r4FLEFNi0Sebf4P
uMWelbD8MsR1UuA+zK8GfSwBBTteF4sE1TXTZD2lCey7hz0b7UiBu3bYcC4Lj4kb
cj4LczqXp6SUzl9wLqffsH2O2NnTj3OdiPZhq498WuY7op8Sw0p50Gxdc63uawjZ
+C5sNP5nay8KZyftDYAue19UEUAQYFu2bfFdiH4A29EbS3Ms7r+U44NQHrksxYqY
DMD1PnCiYYSWxv++vgL7/+7WQuzHMvtmb9UdJNRIIbWYu3zdd2CBV8d/5Xs9xk8M
M/19TRKVC9/wskK0UbASpBHX+o5znn34jseG/20dduyk54bDhW7GnjhbijHU5s5y
sBKrxQjnBD39fqQvOY31e9X/TgkziOJDiP/+VyG0TmRBJ0AEspIYmuf0lfEcjWTt
LQMGZmgx7hnMtw6jlG9DAyXs5OqqHx1ok/akb+Jz99h6ZE6Y35CohAIMnpg3zly7
KPmy3/7+4EcIKs1zFdTkuLWHHZIlGVE9SSEStDnw+XSec2hyZFZHpR+HswTBQkqP
PAi0pvrMPjYT06XFaeHFektXwnIYAWPP6R2VWQZtGesxt0hmFvCyomNAO73cFkEv
s/GEMdOQke87WtQ5Ln4Tj0YC4jWcJT0oqD2oXbuPb/9bthFyED9GeRiVHHrPQnJb
eLacHIeOhLSBZwGe9wqrrSrSvBlYX4BfpSFqc8kfpTGqzknIDNNmrFTN62X1l7Yz
pPgONS66Z9y65sgFUAQpbJlYhX+BV3l1ZH1rExgoSGF37lX30K289lgNC0qFb7YS
NfHl0O1nMIS7dOBsyinchVrBPbPgbsJN7qeVDfq4dd9/PZo6oFc4n9u2omRDu8Ef
hliMBlumLr11bqHGpHp7pIF+HOoD3ocWgUH149Vf3ordknwYpVhwre54NDn1rIAz
cYJALLK3hoqMC9WdzweLGUWJ2O0nWBX7X+mFiySyUbOZ0whZJeWU8QDVBCJ9OcO/
iIlYydFTNaZ1OHrB2LlFdwZkBQ6RpGUezT3OZODvsX5fVfXnRYqi0/zs3qYEO+hK
FR/IcjVoWf3bvdjKgr9ui/+5hiRi9l2SegwNi4Z5WOBQv4NVHR6wFu8g32E6oTkw
Hz64v1FCCU3sBACeb//2JVitxSHUyUvWtBGJbmgLEn0Q8lQrUeOTIo1yUPdkCLL+
OXAWRQqHBDHEZhYfpFPeZQF+5gxwdKKoGv8+llii9b9Y5nAkayUDDdSBxzoTIHfq
S3Z4aOT5si39qdf4ms0sshnfGMniBQx4z3LTFgQS9HE30+uEM7bRJVcdT3VPDwk8
tcq5KWBRUgcZJdUSsRyhdfLU7Jkmt4XA6CWaZ54NRSlsyBsM0w9ZedGM0UqIzAvD
twGrQf97yXV09ng/zsXp9qiZbEPPgurzdVkJ5ec38qKMbQfW6AHcAxJuagd/iwW7
L3gAejxPWY9O8VwlBWIhOlya2NmMr9paUvPNziyW+HmHaMfjJsgdfa5LwQcGtOs4
w12a7wlKXBXFTZBu3Q/rMnaY9Khw+VS6QBOIGWbOTN31SUwNbimJmchD84xpAM86
bNmzdGITvat9z9RuM/lR1k449R/uMenAaJ6/daRH1Wg=
`protect END_PROTECTED
