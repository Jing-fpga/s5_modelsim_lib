`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K/N8d1UIc1rZ8ucptmpkqp8KU5AkUP02p+rAGw08BuIVdTHRSIvPajYxKAlAbVE/
RPyJrscvNNDsYjwU219oMPHhdTH8B2p3xRyx9rChfsbe6bIQka91F2uoa2Pd0GJ6
wvqWU+9x//SQZd1ZDhxj9HzEeGF1ArpwQU51IxEKD1Jx3rrh1ScgtEf09EijuWzx
p7XFpZzigxV5Ug/LySXyPyQT0cK/OcZM7CVAt3bIWQwvtF1rSa7usQlnJY7ByX4E
QXor4ea4SncTTwH8+uoRYVcGwHNXThG3+aKY3CpOi1YFjvmbb4flvOhoAB2fFWCD
UeyHW3ByJkRQOAo33zudgDC8/jpMXo6AEDCyTWL25rW2Y60NjrPbVTBJCRt89eLP
C9vpqeFeCowqxGBfAkUPjg==
`protect END_PROTECTED
