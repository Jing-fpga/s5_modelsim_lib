`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KyUCjceOnxhfD2golNpFJpv1RURrkKCSUIAfKLwuxshqkYK5FXbtfoELbQEq3Nrs
e3bkVqVQXMzill3xfc00eOjbfbhP5GNZdXRPwSyFRv3dO97++xH1EO5bOT2lKq16
24oiobC0iXNBqej9uW+PqQgogzfT44n2UWxC0AAjqNUPjZJwLzLcvciBpWA0T1bm
pyrC7XA2i21oQiVPvn6uomJe3mYC26A1gw6lP+OF+bw8QhPuyyRoqwKeALEV2yi6
qVqeO0qVTVY+k9oDE3Z3daHutLo95vox2WApQSfStQBImi+qPRsMZqOq6MLtUXyb
YBBki724p9j1QPXWCRdkg8bZuVCnN8pdFRQNzRncBpwcWelU1Sfrr6RudNQIHI/0
huiw2/593Sy+NWSgUBElbgYgGJ3lYNrcymuP5oBCD6V6J99Kqq7ozBObHn68IcVH
gLvjPKNxuw3dcGO2RQzUhcxKnMxEe6Y0CurTkFClgGx6G2ejdKlmdt33W63AMGUn
ztY5NUEG+Virtoa2fBW7VYQa4RR/T3/b37KVcoVNjG0EiWMtYNJvQr1h6ei4nf3l
4m4LkUGeXi0YlDCzrz9aUIidi0u5EUEWsQPJ99lEEIQir0JmfpUCJOhZ6Gp0m5FJ
7KCJfE4yL+YwP6fj6LbgHPsiPTPPqgX/Ah633FDARkyJQ3WhI810J9Rs5WBNO95V
XBxKxmut+/5iWGio3R26yYSVtq9HAu/Cn+4J3v+jj1y+CGHPTTME4Ys9dGz6bnBu
PCquFxi6uky3na+WqvyNSZA2/POacT7ytO7iR2fiMFQOnKA1nEIgXlwl1Bnl4dlN
iqtguEU4sT/GJVS5vgA3Ipj1e9I6EpyUKy1yaqotZOPm/Efc5dKDdKCHCUqgnGag
3TcuMt+TtaK3dxu1ynL6PokNW3D466zvDWXQMcTA2pHXgdlLisdP+YYmmELvwsA0
5xyCmtYVBACr/pgGgozMkdKafYYOCeOiwPwz011gFzjSdSyZLkMLhh2sMJDnzii7
bgQuGvWODfWQ5QvBcYgp3zrswWuqRTvvem/UjGfVVVqSDvGrWe7FqqP+LwjWqcm+
UMa9hF9RwMeW1maAeZpjM81G3Bo8YHTUCNfNUUabAGRAWjSBlt1apfpUz9Mssgxu
QHy/dWszUwSXCVcyf1Bt07/+EXLCWwgx1Wa5Puih/9MNotqO+SmDEsgIoNKhyqOK
kzZB6uobaqYFYaH4gAsx2gzA/yEq8BI+IgLDU+v6x3nOkdDWq1QCBsnvtD+F0vj5
E275MrdOklwH1NVhf/1UCilaIJVsHw4R+MjSp1exiXZQ4RzbTTbL/OqWoNhvVsnx
Gj2hH3w8dSGkzKgMYzpSClipnzQqltuAL9qE5JKPDQc+2t5la0TMDfA+J/MnKAFu
q4tgbz0pPFGFDWSO1ecr8uQJniAQE42Gt7sbBYO5XI+3IXFl5vja6MGSUTTBSP1z
`protect END_PROTECTED
