`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YZYyQ4kJ6MNqww7w7Od9r2nXSnCoyvWiFsDgQRkbA9jzOFgsLhxBlgsNGFL4KutN
UjTwB/pyvBG6NOiociJmqVT/hqXr5k2RTR8knQIouqWh8w8HfX01oUzp7McCtPLJ
z/WdBI1it3YVamqKm7SOND7nxyqpdRgPef7yquMRgAFvTExLlwhwsRPIsgCxYKrc
KIByxl/+SPhF+uiTc3FZwQeBsFh4QOjNHKRvnlMilfE7pb/uOwxUomaa9jUBxKdl
KOLVm8/Sv8wqX9AVw9eNcpj+2p2kzvJY4Noy1FXugjg2EgzNEcU7blROMgbTaTME
GPKSy4XjH1uD/9hRsjs1558QMJ7RfRMryPLgNzyadEkwIqoo5Q23YLIS3h59RQul
hwrzOs9oCyXmplPSoQ7+PE1HoYruJ/JtlJBntWqQdB3CG4VGJ5QhVFzWnHREH31p
+K1DxgpSqCFYH9Rjb/9ODnFz7ix/3kzrjJOFXrToq1VeFA1gzd/DK0GvJbAHJQ2p
L78MMA13YPsOavxeKgAuRDofKSV5/TTXhdAudbaCGEDlvt4gYHk5QhBUYzgTJbus
bHTsyyBvGEmVNyRRffJdf7uRDeralXXe9BfT9V8lj+GXt/XcQN57iNVFwss0kZX6
xFNxGpst8zjo+WCzVlnJHyaWaZep2kfrnuClWvwjZ42iBDc1gh8yefxMT2n/Wnjt
XaDOylU0ZmwzDAvXR+UU4/b/KPAkKWCcsZFNJwuRAtXpgnPG//BXmceHBR4YkqVu
y7pUSAVGuG5eb4ZW/6c0BNnd1FQB4qRyw3TkXsKURYvK3Y4i72xQ4vK+VIgHbMiA
T+L23RhEZpHC2djboF3QC8WPlFXoGgw8UJuhcNgMa7tx0xb3HGJlaWFZjy08CjR0
XAx7Je6t8miT5ttL+geI1XzwyFYkNS2SLc7VRSZVhGNNIHNUmtFhE5BrtRGe9oXH
2G8ka3UhhYsvcJ9pCy7QKxyRWHE9Jm8CmYJaBHWtUnnoGI3AUTYRzfRJZ3kgwH68
yc8w0Yp0lyXAuBgieulxJesagO3297oxUzSdR+6NDir+xgaNN7AAg2/lpPW8nyk2
+U+p4dKHL3S91XVsNzNtfYJBY6diKdkXkhYnqJXI1Q6xd9CXxbW/o6foSm34r8pL
VjGqeUI9KwU83nzXNett/YofSdrFFsb09bJAFtkiOUSVHBtCudFIj6gLa8mAek82
6XM9lhDfZxQgKLJWpfkEETQQWrF+DJX4PQA9QzTG0J3ZuG6AS5dAMJSgukwDHBwC
p3wuzaepLZgnD5iBJp0ZVqN65r0b8ZRktTKgtHoE2767KR5g+Mu0A7tqRYSDXOqZ
+F9crxE5z6gvzPcQ1fq7puVHTBJdTaqlQxpjfjYFqqn+XSEVOKCzxIR82caLIbpp
YLBGHekhrmO1reOCRYst6kE0DkjLIOmge2U5zPJfhRErGeRJqH2scMEruuSOh3Fx
0aXbHP7XfLLmYnP5n4lW3GyIf4a0qQRhwOVTYX0OAZZRFwOUefDqwY6HavqgxiAA
7cUoKYIKSR6l8SAdWOu6D4VDkJhmtu68rzjcsYf7146Dl+P5OU1qCz7T4fzfZS6y
V5U+skYqlV5YbAVkj8rCsBTZ1KvikAAeiT22IoYUckH9+ZW2c3B1rEsn4DPwJM+r
kfREB+qdB15wNnLv/YsCdh2/1FxnzBPg3nciXjVYmVrk6y41zddSBr2F4GWl8jE8
sXQh5s5Zi9hIYxWQQG36ydwsI0o5SkLEjrw6SUTBXiG11tP8H9hwg1YgwDur+zVi
SpGZb98hR8GIVW8DHP7lPXrkVVaMBf/mJqlRvALFD6T/dFZFEHBl9rRs5qNL54Sk
rj5vCsqCoBU7XdSajJmZvSqSJmaPpSkr+dq1qdTidCzCFeKXKWYDpDLLMahOakSk
++MEuEgyBJj2hTVu53Zd/YdAOeUqTWN8NsuGgyJJJOEy4BI3MFMayK5LGi6wX/4P
zTb3UB9gyJVx98D9VqmDLcssQGzet47g3Vp7dMKqO0GHX0qpC8U+t12BTEcxZ6Wb
9pMEK+OsfCGwuEatQbEPuwAi0ics1me5p7uYciJtmzTz7KZ16h6w/hTw2Ux6faRj
TIdJDd3fSxIVQYUH8Wu+/VAR1tUYfpZ/sWpBEmP48d5W06yExebqEYd/6J0Al5i8
b37Egf0Jl1Sx+cPC7PKBgecSxcRTRLelWkZSfbmjEZjYH2fv3mHBkkje1spFlXvh
MmdfWJTwGvlEaNUJ7xrIZDjZYtG264KMOprD9S6A0qv82jtIy1DVONJazWYHMcO1
5WzmgybAcSA5TltirpTOzk9sUScEC+4tRCbGe6wxUBJrA7PL5Iv1LUIDGT/TBPUn
+BSbC+mXBdXGewFDTFY+iBgCIPy8kVRi8N714KrNTOts7HfZXOoEykgBB6k79mvK
ckLAhp0AD7XwZKMT0p3KH6D3BOe+GQmCie+au4QUTT7LwM4L2yA2cTQZ81aPs3ul
j1Gc0Gc+XVYiw5P9zTjYmeY8xDqFoNroENJfbxY7SLgQh4DrTaNihiicKnwsUnPY
mKgOMnqclLGFFwAmKQ7JEW12SAddRcrvNl8rZm/PbIUz2GtDwt44e+H8M7kuEvI2
wGmezc4bsLEhjNcD2cULoKvhPdl1nFUEeCby2e82X2BaDR14AUB+oKbCixO5FUWd
KDfmuIrFrh18+0nzbFHAVGvg870+0rAGQTy8cbSyhwoThVfwnir95wRVNRQ54pkn
2LiC7+TMC1R76++pcDlhQ7Af46iPoMAg6L5kkO74U1e2/xsDX1J0PNu/DHXDcfU8
PA5+K+2RTD4w9LNb5nI8vK0VqpSONPvT/o9yQC4Gl/ZrGdN5ub0Qs5otinYspuoO
dr7hu7VYS1FnVB+SmoMiR7ZOiPSiiVL7vbbz1KKe3n7wtFhiV5eVFnh3eJ2WVeFf
`protect END_PROTECTED
