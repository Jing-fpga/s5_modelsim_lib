`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OqY0sHSxjLKN2/WMjJraGMnwssJ/+GFMnzXIg/fP8p8evLcQVGjDbj3mb/oj2z9h
NjZ2DK+WVO0KFXEZPFVea91Z7vKMOw9N4bx0+FB/ywVnzYBZd0an/dwNg7zBeOJJ
0Z68v2NIzRecsOhyBMKrzQNG8sPSRbV3Tt6VOWheo1uBqDi3KSPjlzk42HZKO6ui
cCyXvA2QFwgteFDsaJ9hya1+1UzevWPmz58Iu/VWy6OCXtmmbZL0ctxRP9maA1X5
buyWBHJCssE9msNFACiY4J+UZQZvJZHAprsLcRji1o1EBrrImpuBDYcaVh1jOW8T
wmSk1SORXkGc+QYOcet0zjjr7AKVP7vqLL81Fcji8qVfELNMEoolOXmYWt085jNg
cVhHyhLTa2H2BjLihgB7gSZ5AFaxSIMtapxpA5qN+YtO+jzuSwWb2yAH35+PRBVR
o4L5MQekT/thFWjwIx6NBg==
`protect END_PROTECTED
