`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SuSvdy4cMpZ4rH2onK6CUkZBeboXfwWfUiFQzqtC3Lzn5gI5GR+5WbFCExux0jhq
VA1FAgRBuuQw4QEhuQW3ex9ulfje7+PgIhqnw5Ik21D1UVvJMIffHH5Q/1YpebeY
lYtVj+nZl83XyAuL5yTAlVRkISa25BaSxNIDTJWIgjy7oPL98/wGWxiO0wbXgr2f
rMDG6dfYaNgM0JFm/6V+iy+3kADL/4YCCk+mVjfJsyc6psQ4bFshtQRRv+4CwgdO
QIuX/Tw8jcK91Pttf1M5oPGhLK6GDtXMebDrm2RY1SUCMiiWYgnr+Qxyx2wB4Ytg
2ZQn0MQyPdQeKzDY5gyG2DxnQIVPBzZ3w0bpO82iW+XLPxlISfGaP8XiS1vES7zD
yUlKyQ2icfXiFbj53Nw7ZlhH7hu51qDBVRXWNna7q27eFm1VM9d8pQIMOY+HSxUn
P3xnw+DtPLDpq/fCImRHjY+dltepgEBITk13mofVG5UT04NlAFqDMgIsriejVqbE
hesWOJVVfNdWLG5Oga6i35yZoYq7j0u0B1vvJl/HQfMVaZFdkzWTBlHW0/vF2hbP
ns8Q0I+kesMlfnjWMiaUWd8GqSO90rHH5Lw4lvCfATyVkiPr/QpKYc2AMBoVK4wz
eg7VD0vmzNuuaheVMk8APEoe/xLpL1GlOQbkh8QixjKtYRmUNc7KHomcWhLlcaf5
wFj1B6xZSx/FE/yOwdw3Oj8c54v4zURURwOPdMaShOUkKo6VBYhRLvvzpNQydS40
BL1omcp2EHErOUP6gf7wbrFBDTt7hqFR5bLI1FBxhpPyWwXduCV1HyOXaZsaLuN4
UUGpsA1G0vtxi2zJmLWhIRVsdg7GztlvItfgpLabQFwPnJU9A+4Dq8uxmfRXtvsD
IZh0cPrRipgQCDDh2CKrks7PmBYb2jylIcwrvSYPck5iW9GfEG6XAZhsdz7gFSui
KQtEIUGGIJdvqghi6jBGGotfnFJa6Y3XcKn40WnbpLgm2yPoI8icU+f414gKwekL
PX6NHqn2qmqpNzTC2D+G8YuJreDpz8/+evtWHQD6Im780783L1ccp90WAZuZCpEa
01almuYb7D8HKDa6WAapKhkzK1/y3BsnqwK5Mc9KiHGRffY4wc4lUwqt1CQ0Qu/L
RlVMMKieQ2/SBFCL1cQX3lTDYPcFLYsZ8XdHLUo+oxdBtXvmGBkv6relKckDHW8b
d9IinK0Lbk/ull2hdRw4IfkX9oWziqNzx6q9it9a1mTLMU0+HF041jZPi/VHWRM6
eSlWRCeTOC4fSVOQjy9hHqiYuEA/2sRODCVlBFmwb63cmckJ/IGxipo+mTyDXw7u
zdMiovHj4c959bzd7eTSYRRG0j6Uibp/NEpmJ4HvVmgy1X1CvklVMABy1j0Ek6iF
BQYjVo6rFacXdZqxkw3MeOeoEnLQm9PT5lyZDr5HzDXSSglq36UadNz3GzrpCVwt
qeO7XknfizBoiQhYaX7XhpV7YV+ZGBLxy3x9+QmmWYfjJ0xUZIytMfWEnC7fvny/
f868nZprkTutD8aSVDcrFAC3rV/X560KNqDFglVdGmor6waWYkvsgxJKgfWFfnYI
aHYDlfTFTQ5iYiemkYAhgS583ThD7YvL1X62wVuORKU8WOL3hjS+qJlbRXkBcZ56
dVoEPSy2IG/Q2NCTVaTupytQBsKIwtGHn9XRxs8K3RXbGumEcTcO695Hc71qJdp/
xC+BmVcL9rFEhm13gP7nHVSdSlLmUQ++xISsBGQGV2N3EHbqjcCQTVlDAgnmObua
zQaufbxvBNTedFp0naF3CjNK+prrFauqiut7Wej9c8dYvZKUsdQ5TzfYzT0fvgVf
CG2B89Ign6PszdaXdd8cH9XrEYYb5ieNwQyaj/xDckvDypPRQEhKntjlOv4nK1uY
NQbjQU2x8QEQ5Jq7AlTFsiEXmcruBoSKujqSBMbvqErcJ83gtBe7JrdsdM1Zvqya
nXKN5IOmqRmxE8E2VGtwggUBXvxZg4bSKn6PTrBwT5QERwGnnFl5lB+Uhtzk1Wie
ixvvRbMilKOwyWbwTF4loD+x9ihc/lzsyiWlmeX1FNo+8BmR8y+c0jgLdBOTzO5L
4ku953muzvFD1fkvNwEsIGLlHtCGcy10td3UPih3yImDAD7NTGME258ydhRDz4nu
Vlf2Jrf7OzpicJ8DS1xKdoEYcgnaqerRkJAuu16enOsB/OIxQWoJ66XMnd/L1jw2
TQieWN0JEb9E0uukEKhX0jIKPBvxroKW43WcwlhUhW9pYr7PW+vUXHE13TCZR8AD
L+oi9GZ94O6rhug01yrAntTYmHMRPUvAyZl+LHda3rd4AA3xk1iqUtm6gSfGsUnJ
gtrH69hkT28Q9/MHn0moqh2nxABijrS9N2O9raF78zS74hWhaEtfjGxAV/uMW9MZ
BQCKWm/5S7peX3M9Pyxqn4FZ1+ac7hiY0O+i94EZm/1f3GiAxhO1LyzK31bVt4K1
kwHnVTh5DsGxPd5aW6G4eXrArnaMxHBwK8UD+UR9Xp+nol8G0uR1VmAnF6xWeN0y
GqsXvP44AxzNXfg3C8SRFHT6Xk7IE3GyhEgCyIHpYav7NxleAFxb2hrPP9hpMrZV
uGy2Tu5nTkqyCgUvRygVqZMh/z0AXu+MKPBmGptCGbE3Jwv99DlQoi/WzP7nwQtr
+OLcJ2RG5lP2KRDh85gDABe3e7Ss7nxS5FHTqzaEGhVfUSe8P0Gy92ve/lViMApS
0734N9rh656ecyxoUb0x5bP82byaC1F85EpqmrB/NXoVeVSHGYdOVMDoBF2vjO7d
HFldIoDU9HSknC7DDx5FxSm2oOfRQ/v5GDdN94r9jBSuevvueVnwHdYVp93zHlNU
LjdS+CNe1tYuFMuyvN7+wP2pGkxEZNOM+k5gLrglbcLzTSoQvLIHmc0o1mWK429F
za41eSsE6wu02lh0qVth5/3BcBsWqFSYZiOFwcDBpHonv8a1hOe8rOiQ+fhJt1wb
0k3t1u+MIRn/XoD3cZsQ+4UYQH96Z49IP9ISTcNerST+016Ip03FEugHT2Emvd9P
8lIZSq0ioaR45NgvgsdFG9eh2yFYpl73Q9m1iw8uxUoMp8T563ZXx669OmgLU9FO
`protect END_PROTECTED
