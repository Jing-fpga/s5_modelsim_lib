`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v4HhHLEfmYaF9n2/jOLn1ezVFU0coQbGFnX2kEH4cdXqdzeCJJ1dKTxxBZ1JddHG
HQp/02MhwpGW3PCaAe1Zw5LP6dHZ7QGB5qbVF4WnSndPjGofNuKdNXJ0auFizKpQ
re56qV3xsJkmizbKr9EPgAIggBQ8BQ3XKV7Nw4YMTfXuLzmX0e9ticf9zlgqaovf
Te3hHYmaQU54lQsK9Zfs1XetD7P5zuz62QS+/oBIxtAyXx6zmQtVXUzBxjqTPSYD
DajyWyTuKB2FKSVTOV7V9bmrN5gQVObWN8GlEiLlV+/9FbGepsbtn3+Y+M/wuL67
enbj08gs0zf8A49+e387o0nwrwNyeE+lT8NpQTvGzbOOQqsTdSwdmnnjCh/V5yBL
P1Od8yPtV3g8irofVTBqXYufR6nvDnBRd0SxPY8yy8MrvFFs6ibONxFRCnqGxpq0
HvbHB8KljzqML4OLRo8kM1VwkMP5pdIYxtksiAW5kxeNW9BI3E7rTuWEglWL+r6Q
aryVYdd9rbX9axMKN8ep7LT4QNmsHIfg0zZ5dfxm3rt6ZFmyt+URXbohp1RTkJr8
+sgXiSFWms5VYfcIveRzfg7DUI00jZhQUvEypNkB6zRf3tv3uy5VKTREYhEOMSej
DmkLUmIWn/p/96GkbZRDanx0XUh36hTAElp7MdBo1GoWVmQDziNbF8RNbEGo2Bpd
Ln7lFbJeYD4hZenj77/1ptb7xSkKOOqhQ4OpM1lOalzTQapCLiF776bewi+yspMC
JrK8mBY/Lcpo787SLDOF+AtzrdL6EkzJoD1bZSCJOwRRg2M8K9TVg/z+JcsH0wM+
/+fVpFtky176FD0O4dInR0njs2wY0V9R4Dk6TSiRLwnfDIeHFO+vUnc7dMAYQfCz
BqehfWX3ccnb4uwxJJW1WpBUZkPLe7BWPoz+RXwpRAJiicEDP+Yp0CxWM9b4skK0
`protect END_PROTECTED
