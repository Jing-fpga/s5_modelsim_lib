`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cFhBNaJMRm6SJyAS1lUIPLRUowhYa06BC2Nxpc1tddYIbABM57A2gZOFKxHI526t
kvyGK5d6Q57a0amCRihMTNfdlKaKL+KtmaCISXpUzlAiVyuiglkowY2zwsh175Qc
ymFjd2WI0rjwLyxt3oXE8grOvAW1XljZninJ67a6ZWyKdUiqhjMBRQEQLT1n7h0w
zuLqhRS0/GKo/Cb2DSyzstAitaJLtmm3wLa24mNPIQnAcZ4H966QulMJdp/C0LPI
NJcZSDgwwxQiayKcfd9MnPyvLm2O59/dFfD3gu0dy2HcrUaZsenZn/1GBLcLbhuZ
PNg6ZqOAk/p5fcRZ4eRxN/9FiPOFZr4cKW/4JwLqX67vdGBaZTEAiOcuKZjlyYwJ
Bz16p3zRJGc4xC4wOdP7AbOezGglhzDvoxWSW6PvaDMuFmWaAzpx4jJC6PUy99L/
+LlAVgy7BHHwjRXmEwa4IZ165YolfodTtpwqfZIieg9cbglQoef3eSXP1W9GqtPj
EU/QbGU6bRkOZk3rjUwISxe976RMH/ArRDucCPZc3LuAH1M2a7pRYaWVh8YvUW37
4GTBl12U3dZJswW1Gk/vWKAfXOCQcZJjLqbXuojsruAi06vb0jKvkaK+pSnhVsUb
VfD92RTJDgo/d/7iFNO5BcrEkkZEv61x7DEIGQOyKo0VF8jYY0+LkKoJEHq9FAEN
L/KNIHJ7v2iHsZ2yq/tZXxqjWkiyEyDPRDU1e2nxEnt73cgpJy5RHAjBj7b9ZhxT
WIlMEUxe0cErZZJ+LGl99T38EzB5DphXWVd1ymQC8UWt/1t9HPGbE8/p/FJakqze
KRh0s22tuXIHAZDU4a5/hXqGj7t+ulgxsZ5mXZMaOi12ao/SSgwQPftaHcu2muA0
OGFdHTkcfbg29VkIGAznviTjqdOabcQtOhkwQofijtB6f8+qfC2u7f89LaybsE+V
M4ncoHSZDtPD5AXQD6Rn2kCbUkJSLcz1PkusUsn7gohCHuXAF9eVUvIucLQH3Vnu
CjI7xqqVbeNRqaQqjkJ8YEJPkWnWwuAi7hdTi1BSrWnrq9mdaAXjCCEEWzFUZnGs
ZAKz+feiUqT/spyZwP9Mg8+aXhGTvHXgjee5SpRUu85a+HJjEk9AVhl9S9TaPwbM
wr/+11oG2MeTjl+UskcQCSuaJ9TJYYSAdcjU+jl1acE+oEjHGQEV67a9ku5ZQf1q
b8HFjxDDwVXCCNA5vKml27WwuWINZt3Nc9+b9hZ9OMvT9ef+ke9w7vWrwNKMOM9I
jZtmieS5AfBG7dcdbHpHtFbLKjPa40Y8ifGgmnPAqNKAHcE57jvcwGXizR3gTiz/
SfB1eiwOzfB6bMmIUb7FhPTrusVAFRbhlG0zs+dI3TitdVr6RlIlpr9CGjt0ZslE
6+tiDxYLNYTBhsgfQ2SnQpwfQ1Zx5N1ulRDGVSXkJdukSJmWEKqa2GMXzdHCIoqm
flERRBPGegBnDqZ391co6jRiIGr+Aig5vFADtmP3JX+FbVjWDG4mouO9UcEUEEYl
GOOcXGWbcHcHNJS84f1UjfpDaiRWjxXor1RXoYyn4hNZQanGnoBUt5G/nJbzWlBz
hVbjfGTvg76kG1bSpSbiik+KvebtUoUwdYZ4Z6GsSZKfaKcJmVK13Mkn84qRajP/
lUf4t7KuamYK+pecFNnmQTe1JD+wRKcbHMvicCYTJx+ocYtOKumQ9Z5ZJqCfftPn
emglC1xj2ju40P8kx7ar1GzLk8TdW92cv4QUKJ5KSAKFCD6sTkKIAkgE6O8EYNT3
uxo9xPbpCiKLskRbgLNzg/1JgqhfVzE0mxezrEgxnF3ao8zqxFQZwtoASnzivym1
edJO/k/QPil2iL/bzAAvm1OJeSQ/qwWIqcxsQWf+5ZQIgqD/oCtHh9RbwSi2sanD
vq8I5YQnvLZeyYmYrWphbDmjKWGDR3tIfCqIT54daxH1d7tcrxVUz22S81387PtB
RLhPXLTks/1lFnFweshkQ9SwaK1EbjiAMGAfG92t5xJ1n+GVv2KcVSr2mjb9AOEO
sfwC68cmvt2v3mLR6dY1EQUy++zKve+MpfNy+Bfk8iqz8XQ17A+6RvsTplNMfTC9
A0RvPnPEgj7yZ4NrUFrp/Cb/Zxpc7H+q+oxa7qA+mNdVmeJbUsZXbjvMtlT1iiXY
1uhXc44l8po8kT0UdglZ8HoLoUP6auXG+jdAL3obesCQacYZgUUSH/TnEd1VRinK
7qQd6pOb4WegTDgMt5LakF6ORkKe+sRlv7Dq+OHAs/qjDqOiYaEUaxIhqefpZP1d
tQZ42I+XSVBNH7zj6pvSb0geRbzxUOr9VIHPf+oc65qSwbmyNSP65T0We7KTpN6N
gMfmp61lbMpx2C40tHn18JWawJfJFgWuRZOXpwypWU/sIuqMb4sZh8/sjGCo/UuT
pdkaPgJuivnJtZqNe0jVTI4XLTE6QY/u0EuKEkt/yuttcQuOrWZuA4lftdkJPjZI
HNOX6PfIhPLfSxuC3fwwkrBfw8QctaKLxh8s4Iqvu1l6BjEhmMfBdJGiSnkJOqyE
NajBQgsv+sCSRXFIRm+WjykvhJ5rnpzpCK2cA1e7rJLGdAQGYKYfnieIeFrjjQBh
VpbGIbu11zk7ZUDJRBiKAyzR9ahs7QoPp7SIX2vsEPKIl1YEefnspSw69WSLo/JS
`protect END_PROTECTED
