`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BqtTdfcz+JCWIdXp83ZUniEBKkyb+1g0IXTNPunaS8yb1KAa3VPAxITuCsMU86xL
WF0MfN/1XuZxAY44H1NsV/poBW34dLMQNYiahWdQ2aasFIAJ696EHaMw0f1ERj7G
zSu92CYb68SDYjTleC+uDlmfrGyDsd4sfchkpBUyXSPuH6nmAmRw2UD8fX06q0Sa
eIAqRD3YAH/X8CV0PvyN9GO5VhCVPN3QbsQfSG7gV2qqVY9cE3Cwgmf+FYdx9wTf
mSUG7C3VRJPsSHAbZBIBH1Gb4zOhVWZC9P/0OP0x1TebB/yFSKH+qrDRULZ5PXgt
kvhtLDoS4YvluZ7HqO9rummzrrW9pURLLqLEoEouiFU98++EG4jt+gmTx1Mdg+gt
ztQ7xp6SQ9k3txT0g0vy2wS1wrexg/nI12PuDOqR0PoQNEp7czoy0b4LrHre6LBP
A7HDXaMVe/2Yzjb8bNh6diXo+mwb8jNzoeAvjhhXU0J/B7QM/wXo9yUVKTTZm/QL
vX0DAt+0yEL+1V7httQVjevLxZd/OZRXvZAK7ziz98z4czKfaBNRnhFPceIh8AO9
Zzbo1Ec5XDExjOz9uisYScobGfgl4jzyGPSXklS0Id69Xb78ra8ETvZITMTICqRV
XMvS7Dz+nrMR6bSQy49CTiDtVZRpipds1Os8YmCiqx2TOUVg7SeWm87TdIl3QNJK
ofo6w0yMZu0521aulPHroBSuI3v+ipxIm9OvOs8RXirZZktxc9v0CD8b6DlhMV9y
iRdsKjq8BDj+/U+WzNpqOmIt331HmxKPbwjhlTtEiQzM0cSdQhRBOGmH0yGfs//j
37JbZEdQxRAQklUKd+arS+zAkEYohJRmjIqJlpls/xVw12M9cKfAvzzFue422kpS
xqF+I7H7cnF72JiD7abOvO3z4ddq/Bgp553DL6w+o9cdaoflghKF+6wmN5D+EoOp
cefcYivMnp7pl+cU+E/XVv4IBDwtYermKQqT4QeMfs8WQzXAco7fY3FGjMHBs2oz
3q02wZMRV+s+HADI/gJ8h8bE1eclK9viViisVSZPSyjmTSCVRUhxa7SfLyAI0JGP
xpxS73JKTQUNgi00hj0e8AmMPwHZWXWk/GV/ehfFsbSufgcawxBtdBpJ4Ub9o2rm
FpuKGTB2VMCUjTvN6xVVNlAiR/sfH5WraaQXx6foL4QZVfVw3cY44KmA93JfIOlP
xZbM+H66NRX8cHLQwN+Kt86qi+XM3gLHjy+1tqo8fD1MTj+f+c+nvS0aXfTdJw84
rPhg0AK/1zQIPFoZEUTqlisN/K0KohOA5Z203Xt4VJA++gOu2F6WyUOfEAtNxPIE
I23rUqiM4wSrijDyYRuMjdRCVQ0QIPbIz0ELRyAo0iuYZANZ65/GXSS0CnGPNHrR
1U8m9qDnS3pCZakvsUh1Oea2+g8YBd0Bib9gloJ8yeVslZqzAtaW2BEIsbNxl532
T+W+1CuytDDE9Asni04xxRtyW7qe45022f+kyT1iKDW+A0SxV9e4A/l18TbUGe/I
h9aDNJEV+HARebYGnXfSUFlrC489/asvIsLQYXCu5dfN+s0ICBwFkppoRbg2uROz
4dFoyhSaRQeWyRRp8+6INU67wdKbxHOkstfQRkEseQnPHNRHrF9WZhr73ylSg833
nKxShhy1N+XiawuGMEP2h/DWXh8ZzuZjCX7Lf9yHpFvlSjIXu3opU64LtKpX7UsN
ly0N2jXuoPOK3UOiGNnG4OD+Aq9vLnH9G3J/irXpQKYtkINMs2BGoNMzonOsggH+
Mjhsi4kQ/5hgM4b3vKCjhwoXA20sH6uS8qk0PCsIlFqDy/pk5PJTA43pXdlS8Zgk
wggp5TspGimTjNmtThS59qATtU//iDxZTk44R2EPZ5oRJeaiIrYP4kUjeiOV2OeY
dvHKDnzDkNj/klvmXviaMKzp427k8s0/KMZ6cUeVuCLHpuMbWqlfYv5WDZLDhVCt
uXcjbkeINsbspSYe53SqU6ThQ4Wp/BsyXT6iPTLNpwAcFU0vGIP1csyGsS0DjoSF
dl4v7BTqnJq5pkOGybRt03Fq/dELtgG0ipm+zV/pijG8pcSSCc5m1uA/id5nShoJ
/Li/GHIPur2R9D9tu7ZDpCyPgs2z9CYO9ZHyYPqz5qguq87iOPs/tJHrja2aTguz
`protect END_PROTECTED
