`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ysachrfCCgS5RybPxHhU4Q6nvPxCuY7L4/X+h7I4aqiyxdYLUhLOrXQee7ClPOU9
jSZPv/wordkGx3Jq/dxfPWYOXZzdiFWKdz/abUE7lxpTwI7dPmTTqbHCHbdS7kOO
c4LNKV8See/OFktm6q2AZaFAez1HnmeIVWf5hWOVyo4Gn5faW9EnVDiQ6hhK+4J6
cpC2YFhCG4ItidtpOUj3HebH2V4rnwYrR77s+oGjoVjh39eDy7rnJomu8wsCupa8
txyZWyyS+4V01U47d+0wZtmYJNm1LTMJAZXYCXWV8uhMuJPICcz2FyvbtnSIsLTU
Mq4N1R2eej35MtVGlVfBlLXDIuoG5XY0fN+t0B5sdXEs0Xi79I+ImTUMoUvls3dI
UFRXK6kes8gmuxaZ/+GiNIOcDOlqr1KQRVREoH/9jDhH4mVGGxMU0JyVzzV/Y73D
e2sMnxQSX0WfRv2l6pOcsqDtZlLpV4jT1iEyTJoYAUhgHlBIcMJpNJ3NqhVtyZYg
Aodae82kNb8xZ24L8nUNKDJ1m7pfRT3KjKmSdB+bxjczNkRI6blBHi5jshah1B6G
4myNMaizZaP4v4GKGiK5NxKh4TZBryOjjsNCvfCMh7unMmqnOOh7HZJsFRNFjcxe
Ok44KfZHlQHUDtjqU5fuBL7qaw9kW5fGpHSWydTVXcY/RWY1McdnSIHOP25Uuq9w
3qny9zCbf/Gm/4rQ15k+YEkSnHvOvtVIzWt2MbZGk4lEnN8TlNheU739Y8tbe75Q
ERpJx8PuaiKqRNkpGxTgfIqD5B9z6In9ReHb6j6/EXlRn+XmBLjX/J0CAr4uTyXF
6w+Y2lVvEO7YWDXnTay8HUpyREhkw4BuPhr02F84k7gi27A8c1D1EXTdsJrXVnJT
6PVoSLECQFLN6Luu5pFuTIm/yp3dKIKdxnPobdFW8bTjGRBi7gTwDufy3TlJ2uvP
oZRtjpO4/IiXHmq6HPXDRXxA91DZw39SLA+mY7x9ulLegJxgMaTj5Q7ywZdXL8B/
2q49hrU4RrMe2fkV4klElHXEgkhytfj/GL3Z1iwN+KU0yQpjnMolXi9SfM/sfdJl
eC4g7AEmQB3C/vu6YnsPYCIBhp6+5KDpOkZPZNWAy9cgUuWI+idBrireqkjKJB01
h5mS2g1dvUO4lqZO2xT5EuI/eysmJT7SLPnOtpW3ZXOl6dqmuXev1oL7oONi3dDE
z1AJo/GLTWngQlQhZR2YftlcXz8XRNo0kW6pTgBt3BeGC5X+F3+bEnigd4CRuVaV
5B0KhlRFB616PEo/m89p3fFr0TM7zTe1NoMTxEfmbIPaYsTDIfy0rG3kRJ4tJlSY
0BNzFnAnGcRydlBORYrohu852wuppEN2f1KWrAVVLlXNiTXwWARqPXEUJBc6c6yL
9g1XZLVgmkh1LSIbC2ejp9pJlTQw3deEGDt+ANc01G1Z2LfDz3wtm/kyDS8h1zYo
A6Zj8PwTnu9z+I2Ng4TZoGK4mVZeP6LLIRxA1/eOKXSq02G7VFHF+0QoRVhi7TT6
PuLqlz+WM9vjFTdDBzbuNlX9lcRYFml9RG966dPp4ii/QK6I0w9sNSra/jeqxWYE
DH6Ex/Hls14WkvfmJnrvjiCzs8XPGe21mV7kadAy04/Cq2CeA5wIdRsA+IGr+qTO
z2fJIHw3o4vmEaJgDN/HqdF0exiXxdyBl4EAAwY9SRgzDWfimATIzxToQL/Ainbd
J1mbENHu3JCKuoJQC7s24tJhuTeK4Mp7QHoZFlhL/9xxJLWiOvsFz4y+XmQLVy2w
4OfWPm1FYU/uDXIkNfswnNxVPgVmSyJQEui8g3lgTDMO92d2DSn/p0PJyEOxaDZ4
l0e+Emhr+LU+FiVbsatkL0E5StzePKQkg+kI281rv/nlQFPgpu0n9dj9R6rMljPP
NSuG4Q8N3eUEjjTjueHRVChY0i1VvaWjldULE/JjRBAUD7qE8jPXE0YJ9pOVMXHJ
BJFYr0Sn9D2wh6WwQ42/Q3Q2MGTdJV9vLkGtSc2x/JUZqy4tG6C78HxzP8NTwrRZ
LNxW/1/v8uFOOaPKspRQW/CiN0536sP87ys4b3qlcs/sWZy5T38Wg5X6B+yI32BK
txNMN0ASydh05qBdkA5QxLV7Hr8M5QA0aXTqNWIUVzjj5rourY4FfXLLyMfCMXmY
CQRmVuGamE015Db9O9QUZQMh/tPQTrZkeOvp+3d59voVZfnvKj9MDHifs2bShM2p
bo+0WV3P3Gcesf0WzcDTwwJlmq9LOHtwfHv0Bl5p/wJ6YqEe+PWO2lM7Sj1VhiKp
uU0SrAuUjWCrgDee2qTbYIwL26gjmnl/UEbqNZE1/1hRpxyIpd+fC0j3er67iIeq
1YPvsdjB1FiqDT93qawWzQADDnACKY53qdxm5kQMd/xyFwpdAhjJTDKprOuQYLHA
rnrZVt2eUgky9333+DcBF4GIcK8fcjFA5c4UYr9pBOzdwDsXstJmaHU7Ikywa9Po
PlYvqWchcqmv3DMnTe5Q5viHuccuxgA8YbFXE7ngix80ihjyP7iNXrPQJ+bPCXqk
yoom5e1nnzO6o7on0r8IqSZp6/700111Dh+4E0XcwIYHoKA2cNsFGSTeKm6bITNT
sbit3yWBLnEIk35qMHR7NjUJjOVy7MGaSNs+eAnTV755m4juY46qiX6JVcFYUVtU
kFUsIzDhW1WDgNkGalM1za0bKmXQNakeXh9I+qnCnDuL4SCt3O9oHFiJN8fHdu3u
WE+F7L2OwQjs7JjzhhIovba7q1H0nVsL4VZbMT3DSUKYHjYgHkp+FtwYmR2777PC
ys/APY1fTlq5VgETu8rs3oiuzK4UVym57sXqHdoLwN+ELEqwu2VZ/EMSaF49nF6G
7sfo5DIWOxbqvoxGOtVWm++GcuH7ZzVDb6Xq7HH99mnFnGguBrrZrjZIbxOforHx
IKUtY49EaOvxnFmDvc7bAROWmlTJHxn8qMqhO7EC0vQYtatjYps1qmdJ9fAxVyP2
Qs7mxsV5+8EB+F+PYPbXKXyl3iGbACr5JeQxHONPnNgS/qZm/m7mCER9+jyMfoUY
W+4oLjldNSPXkheFOcSXVPYvls8PkEeHi2Bp4gclNmitGOs3eBG3+w/1OyVO7Eqy
7YmxjBVihWsHL74J3fMFqTA1piaQqVKePL6ko9FYrBofG0Asiiy0X96nkwpzL5HG
Hkwwi1+/MiGxFQUDd/XHYjtAui8ykR/rCytQ1PohFaBf3ECDy64qdVd+F0RKX8tw
/OT51CjQTfsyUFIQDOwBzX/GjhF3jjFXU8W00DPYPRkGw6koojyXiTTmdEClqM0A
v302Hc13ZmOceCZmo3q3jO896otkxzxPUltKP5dulhwb3TxYB8QvU+4OoBMURDo1
aHntELprqSlD85G1cI7KbIfZJBsv76vQL8fE34QETXPpCDgMAoFJQlvtIZQPvLre
U9Eh1j6/EDuSaaSAlkR291dDZpU+hQw9SFXuazyHLcXdL+U41ne2j8j8ruIi5wIR
9d7hy3b3q9LBMw8DHOVjrQgqWy8uufDw766X1BDkQ/y77c+zhQb+S1FXts94Oz2w
shztDPo/AY7Z/El+S+JGpm35sMAfDSgfsNullmOxoKynde0YftP0HDBm3Ug1NyLo
P0lC3+FlyjYcSGNcDanxWCGq8BvRRnjlpg44+cv1Bp1dTuJsjHQBmqcgkscDLSQU
RAlzioKugcn2SEUw/lr93r4fbVfej4ATuuhvdKRwO+tfILRaOhzW6vh37Vg3YbiI
C9XLE7GLUgafPzY359tTV9oGo9K1lyg7RtaQyq8k2Hjs+ZixSKs5+5j0D+wD9c95
SrXJF9XufsJlSjpYc+9uZZsMo6UacBJBimARpo1XWWyp1zWjChWwlD7EOsbM35AM
iMjJIA7r9QajQIFlwANY6tvxxPddmbbvZPh7QrrF9QA/hECpMUjdspYRvqjBoL5d
Rb6e/jMgVsC0tykjxEWwwYqyG7B1DyjnkQr5OrfzHNn7GhmycOmN8V7vDa8gNrRn
cdWg3s20tEYPX5+rLpG0Vx9WNqqPvR7xMicXqapY+z8nKZtMphi5Q44yRRBYKaho
Cc8qNXwbfAbrdUrs+a+Wzv3cmSyOqzmT44iQh8XdMvyJXm6enVdZZj1mtQEUrZrY
6r6Fdjd+eEWVX//zfEc4kVXNQ9MBTo6PArEa9/GWKNl8AB+EYg3B4k+g/XeG9itt
+ecqMTiGTlX5HZ/3k9guzOjDXwbdrXn4hsqPjpqdyNJIXi0UtDruJeNJVGtWZ0MM
sXoBK9uPKXjkxFxHMuMgjlQfAJEuy7+IlRuo21KB/Pd33aeLA1CpEvJI4twzAWrV
1sGrh3EdmmTklBRK+oTuXi59yLBqXDBr/n4acHQWyrJqfNoSfIfzegrCJzroIwRs
r9XV412q1cQDZ2nNPfgS2bIgv/T1g6erLOtt2GYBhbZzl6qy3hCZ3/dwbqA7NOnO
wXKQYFUPfXz3SHVw25ROUBa/evOxgoErSC4YuiCqYa5726UyPa0yL2UXxNupW9p7
k0D2JVxxjT5i/Mp5fcKT2OEoPjOSJtl9OXEfZWZ0Qei5zYkwbC0AH1L0oMdAKVzZ
PLYt/91YR7MLr6uYX0xWVmnjhDcV/39dV4QK3NTPf6GKKjDUHRpJJZ/4S9DxwIIA
Dp1RIYg30kscAHK7Vn5B7hmjQ3zNnPMKrEa7yY2LFlc4ZfDTzSDqdqtClzPp10vO
AnrJOXHFUDaygOIcgeN0cIhU6LICNr9vW57MQfYxoDBKQfj1CjkgYyLUQvFGLc/w
nUUrXZ0gcGLuDZqrSjD9hGhcQ3uAad4CbiRoghYCEyjU3yimse7pFZg3OXbsBQN6
Vo03Qk7hfwaGeWIiqSGY6BEpDXKo3mS6XZnCZbFODitUuo3JYG0mMDk2I1seGz5e
k01NuR95x9hgWqy0zUBlFZN6OsXVH0ABS55ILgfgvPoAVDA8TewqXPn6yWvrh9hU
J6VIijtcP5sGOOsvEu+zRzpo5GYLms8pkLY/CVsVG6oVR4oPLvMl4VtFda7UQjlO
bn4nRV1Au9Pz3UDk3Ug1Co58qAaWD9ISWOo0y/TySpjbp/h1oPJQsfMpsDneLqqA
6hHiQzcVW07NNiep48/zw+bgRrOOrxKuCLuM2XR0c+6N35owjE1KBKy4M6vhkMms
mEqmakUkfnJtR8qOxJlUN3Vh27QC+FzybL7u4+gu4HCDRUDuDi+8Vv3EUl+ukHAR
f3+KeMXvgudU02I3AU/RkJYkkXS/e+bYyzIci37oNrfBvoTzeJbS3PnIDAs/exZA
Qof8t7i+bNOoJsGPkrscmwZXk7MA2+dJiWvOZyihKVVpOnGrTzjjWQtfRgLeXMLN
2ezNkPUdBgYIQQvXjLcaL+MoAb/Y2u/tfyMYXqLLPZv22WfW4FHEYimBqz+1+/PN
++iwtv36H6Lw27KHGUoH53vOiashzwt4L5Wkta8DsVVaObndqWZQgjnlch7objIe
45rNW9MH71flYfXmv28KrbljuxdnOb2TDE3mz8d1JEO30faW1ihGXSlXnUkvQItM
mNlJlrm16ZKzZfILL/JlqnwAyTJVkATtoYeMaojsCkgs/+Lo0+EyUqERia6HzNjU
Ytu4OzxpWWS7JY5/r7FldIYP35m1e64004pt16bJDSNrMr8nmoiD+YfVGhLph/RJ
CAYMb4Uo/Noqry6Ag/4hEt4jgH+fZDFcNDPY3mJKEnWn81XQExkpB8M4MzWgW1QK
HyIBajuSvDsredicD6s5ZgeAyKlHhCsPfFrs3rNfQCp9kJ/A3LILA7JpA0q73RVc
ubMwVjBne2sniJBn3PKJ51ef7iOjJitEsITWaAt9JWupqffbVhGIPkEHxnmjjZhm
7nslAKiNDlfzQJ6OVxZ5+E4Xfhd3tFBDdUgoX7cuwM9Tn/cU+M6H3opUYRLjM6SJ
8aOHx5vrtSspXvKZkYqtNXyDVBdr3s28CbO0HENQ7hdiJD8nqhz26/oxANvmhi9w
Al1PZ0/fYNhNgNy1vj/zFY73+Rf5xE3Cfba4JtEHwtCrKt4PobZqB+VJHGphIFAc
Fq7nOfV3NmgGn9FOYj7Mr85BUTNPKj0EcQCjL9jFMyh9DHhrGyVXJgtWwrgT1P8e
At+Q4Fq6CgvMW3GduJlV+bT6odn+782B7Dpf7HbbtNn+vBW6oVkFN0Cw14oJ+OMS
AxbhqaZvVvRBgwWx3fPdWEjen3Iz68PJ8D34kiq3Lc8lV/XS8d2TtOn9xb2R/5+y
vj32Ml3AjPC26yZSV1qYDr62ji25CukJxkETO15rzE5qf9TpnyB3RXyLoLUnYs7S
zqzsfoubItBpIkhr2TPu35+i6/fi5IKj9a5Da3V738ERrF/asg9BUM18GRJMhg1X
xiCii4ccD1ZMczaYxsCUnnQ9tocKjiD/75ZObbIcVxvDUiTDCtLUADpqXPoONlAL
klj4d1MUSPp1loDmqmsmJqB1Iw9nO7+OnQF51UnKNbs7I6OVgpJfxNTkwwpJdjg1
V1RWSo/+nmV4kWUVcdPJXXydxlCl2ekKkHEHItuR3ox9kslrtqdDpEEIFLoFnf1w
h7zfEZ/MqKxgAmg078aCQvu7wGTxF4O+pvR6DBpGRZl58p/7R+JcgtM5oRX19MGC
ezSopF8EPK1dyxtnnFXSi1qIE9B/QGGNWYuh8fguCKfA284Cy6Qb6B2du9LqX84K
MIhsDG167E4keKiPi5+VV0GlhWikAbY+DD+voGebvNMWaDOkkjSO1H0wh+A8wuX1
sPieHGJ8yBSO6hGePyPb91Yl/ny/qQDHKtyWu/tmc9t71mC8eZ/ZoTMtTcKD6uQ8
Ba3jshiUSOYJ4rdhPGEJ0tC+i28yNubThr4Snzv2fGxBLkRwnkUbEIkK7XrpJmH4
xlzuKm1DcYCh3zE/sjsVIQUQKWDoH/WESUyZ+e57zzO3GBjiZMYRoEpecGqQ8bXY
cbdSHg4fwfPH5oj/ydllv/roFZ8nIk2HP6x23omPcAkqC7WtmlTJIEeEZmdbIMa6
2ctlKs1j/PfFVKfGIg6g76Vl/SRx4UDaNBCior0g3KtgaaDUhYPhqdoeA6etqB+h
aF3BgPDKMyNxb6PtuN0+GlXmyFa7Tz/PKugT5raVkYRg43T4z5fThUkdhEE4s9gh
7sph7CQaVXZnTfXbIjAR2PAxD3TQXAE7HkDWIiAxdsSdF/Kk9s3zfxdnYPH7OeLP
Iu87AyyisUmi56nSsUScjHDuYLxkMq7bkdVYw0YyP2RL8r2M2+dtsKGxi+IpVKLl
0dSFHpczuQ/Zu8hTXCBj4DJDMdfKIDbK79NBZQt4uXQ4lKOi3o+K69gfBujCZcKl
Ara/NGE7S+Tp4I3w14NhIIr0hjopyiDoT+rNJaaU65PsVSbvzMY5Gn/mKupLeMd9
i+/UkmGRwbZ84QbsQssIzZnoCz06xfHby2hLCKxRWmXuIkgw+J+QhvTjJCa3ECfh
U88qvHBA78hrsiEss0ZPrk8n+r18cfIHgPpzJZItw97YWqMg6eh7h3bCyH/5wmI1
jQxh756qxhHdWkYWqMIcgcCDlOtdrHJ2VDI40qC3BBMp3lj3gg0IbA7tOLZTH1Po
aR3Pny5banX7FproxL9wFHzCdgWYtfcgYgjiTEii7Ly5zFdwJRGEZYP0P49zbbNz
Wm0zNGK8yTFX1/J863nviPTeZ9YDsiTU6XNjqI90ilccQrWE0rTEkk7Bg2YoB/tY
Ls0h1AAqeh9EBQnmL99llsl6dXYDtsT+aePTXR9LVS/a70+FjUgAebvtB6YtsJF2
pm4fzYU+VhifuvZGjJAS8Rr4w0b1C56lVI3EhTM2PioGU87AN3qXh7UmDQUat9M2
+g67Fo6QtGV/CVraWyv/ihcX1fJW5FEKYBHfpexdEIoh0DM2qsvgJrIuMTk99UwM
4s3CssRyBZ/jjKTGrzypuyx1NhMGb+UJm5YKtH9QiBLKMqXlsxTi2A4f8zKo93nU
93CWK+ftahHkJvUxjX0Lxuxv9E98KYVRmWSI8tColeLdUTerjjsODU7FdGMc7Sda
m+zIxNETDg84fjQsuUIU/cqwWPun8bhN7Marx3dLdgV3JL3GQS1dW/Ct/ZfurC9v
CJhNX3S4ytNNOhOi3wNzBz8+x9Aig9vTfUNzOc52tlaJBdqUGT3iSykSspSHHeX8
Bbulqt+fDtaBSUruUhftOCTqVWg1CTb2aCILyyDsTPA/F/oIyTToviNuFk1xR7tY
nlmZa7u7JKizCQw3nDkENHpolwPvY0QqVp+NBWCFhvIzJKXX8kQKRLUkfVKwiXRA
Mu9HMfcTMVmgfrKJyi6N1K9p9NgysaulBU5Y9Wzbma/8B80ZxiZa5nvJRNXCwOsc
+1mdPaTe4LiYpj6k1j2SQTOW9YHTMSa+F1qRpLAxWJkRGJNBa7MlddbWyKwjaxLl
KMz1OVxoaTi7dtMGK8ywDtnapkSxwforXunkBloQKQ0TFKJKqpuE0UePXyAqF5Wg
07eu5HrGc0tmqVu5hi6YshKXxMn3Pm6X40SGJLD3LSGsVWwvK1d8zehLU/V2q4RQ
x8Anq80mOfi78ELJItISZvRjAaFErhHqh1/4WVrtrShh25UaT3YNRqxUplBbehyo
2Pgs69ZEIKu/UzbjtH5SybqBoTA5v2GvKelwXzoTL3xs7x9siUjlXzLoxwHXFmfR
69AFODLmDjNcaoU487FMgs9gyd0okPlcAJrukCTAbxCsAlPVr+iQegfLXVEb7hkH
dnUVHwpFfQhrDgX8F6/VC9LZi9tOmc8JP+ODwgxCBV9YVugGayEX4X4oGmTjAUmR
xbqamjUi569DG+AsFPOv1hV/V0dYo+Vkmcm5jIihT6pf+i7m5phSZPhsUL6om3aC
nW8ZYpfPZW+GRUiyqYP+cJkIFsxh8tD2RZg5ImaeKt24H090uNesre1IIm856q66
L83oDB6fytjZvzgJinQ6m1WEPp54o/hMBgymD13BCkE9is9ScF9e04xbyN4dCiv7
f6V4u+CVYik73DH5ZFs30en/IbjPugYguBd2aR6BDHSZqymM8LvPckwHfxim14tg
OeylEyfTmKGDQNdRrf4TtyrGwdplvw87qxD4i2Elx1oDdialZbAg3AZQpbAImbES
PlBccHx3PdhPUq2mjoNy+zSLvpaxANzoP1cPSVVBuHtN8OsPepF733XUbNSGd7Vt
rYMGy6iGps6H1NfU5SKMoWYFXb8E37tvHA+oF8fuQja2DByWlNGJgTN5vqBWlc9f
nBB1aT3uIPXaBxk2FkbzFTOtuvMu3/yTtqydEed7/oDZm90VqmIYqA2VyzGFoPXn
l+dYHbB5288nNFqQYovdAsSlm30iAZYy/R80Va4KY3s+U4sbRUehN3htaFdAg4v1
woorEYy2Ln65/lX20EyWtjkS179JFICYIekpgD7JiDILl70PM/Srt6nGgfWKE4g9
gjogEsVlH2wrcq0AK/0MTCvJ+ObtSk4Zx/KppKCcNgxxXA8TkuNicAETKezRnvdD
Fe2hafMq4VxvBYRdhAyZus3li03lUnyAnIfs60Ie5mzKID5OY6F7k9g/uDSH4Qk4
7ohRYS3WxQ2p0J/3/B0SOc+gyS6OCgsLfFKieTYgDyQhGAs5DMmfUBZp+6XC7se0
kSXp4h0DEH1egAlhRIlk6HtXnwIsSnqWEGTlcU5Hx4Vg5gXtc9lX8iafqvOqAXFi
2R9qc/Dx5aEqqYzC9vlABC7El+GgV+IR6HdFme3E0CKWJOPS/5kuaR1bYMbM812o
GpwFty22MTzhYnFKfDUbq2T81lxOdTFprjiIA5q8IxgFnphi1N8j+8UxHosh1mS8
5+GOjAdCRTAykpia23bcGVjDV6HqUXh7cmwdnbVUCmLD9BA25iDapPkY/TDrO0QZ
6QtTlG/kP9Qshh9Uo64qlw8f8HtyYxkHGBp3Nu/1o4BOPmlqXKKCW1aEq1fPY0O0
sSzSt77YLQoKNSxc363AxzoJNu/rBRtMP11SvS/gtl4c48aMzEtcqDNr8xeDW8YW
WQRqwd8XegSEbvAG4k+56izPHdwMoS9dICQpJ8JZbXb6AxABmJL8wgFsbRwF2DMK
6kJqo/lXh3csOI0uckSZCB/Zp8ARa6Nj0zmtEnQhSz4WAvxJOfJtny2mWYWQm7qB
T5TiAM11duP9mlLzkW+1uL8fiMlfzyDxZQuG1Sn2I3wWKcZiYSWPClkg11vhiNKd
Qg6/H/1zVWz5Aa9kkHwWSdFkxicqN9yE35nRUZbhyoPgJfHpBZq5vzWgdmvUBfJQ
QJGAVyAy2iMjyjIYyHg9kEFDjTFD6Jm9cTfRUm4GTG+AtS4nmtdaTrZzyd/1GBgg
WaKkPJKzhRLY2/6ZaiugRcAxjfdFDqh0iV6AFdWxUHdO5hluzBg/LpZ5PgTnWUQZ
VMRlhDiaBpXYhoSxqjBO0tb20PvlEhpgQfu6ECIFpqbcdgnPMR6eFoIcBCVk06lH
msBUp+tKrGUkfPDyrWEQ9TpvzkT+hk/Qj+HUo+H9ABY4qUCdsrR8DTp+qiSTtcln
JWetOAPIyYiDb4ok+jUZAg+23KA0pjhS4Uo+BYvz35P7UEHrg/92DuR9Fb25uE5r
OaEKGnSYkv+YXY9pmnFq4m5FPtGqATvw33LVaqTjynRAjU6RfXG462G4WEgbhG17
X74tNUyS5Ep1GiZHJMVVqPxIACHCzrJRsPwKIPUHB+7Vf/IiGRoncJ+rHexnyItj
/xnNTIauHYG9Bqeu81gSKSPQ36saA1vO9EFdXjB5RTY=
`protect END_PROTECTED
