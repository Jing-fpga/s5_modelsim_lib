`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lag6yK0PrKSVdxrUKjTdpYhM8WdJDm1uuRTIwtCTCw+Ns4nTQYJmIlVpK/Kagr8x
a9/ElVbpUZdZLjBL/F8ZbSde3/X+ItIstMhrAC4MIPipUWXAA5usnkUCNhJl7iB1
g248YqteXeCDQcMiVlkdz2KyhSzhk58DC5KkdJ1DseWgf+2ADFhIzMt6jTUe6WHy
8JGjBoSYggGU10qx94CtK14SVE8kF8jNLCzqcU2bO5tr+XU3FoOHmfMEI5cWlLWn
TfJR5Z5x/+G2RWOW65bNJPy2vuCXheURW7aA8OUlX8s5T+tAA5IpGnoRDDcWs14J
Gh+REC73AM8GPnp5Jbdxw7sr41chC7RCeC1d/MEtZbCkWDcLLLl3VqBZopJRXm1z
Cl+OhjY6EIlNOnwqLp5xK0S3nKG4p2S0A1NeCWG1wKOBuzSutzdD+kz8PrstK1EU
4l/IztaBt34OLJwQ83mutU0rBbIHE9Qhuwa2USQ0lWB48Ifo0nDbAf6W0JTqprrv
AUD9FyHbXXmsElz4pl4a7AQAAkvQ1hcb+iESq0pxfelzuMnnIiewhA4o2PzQ9/oV
w+p4Oi5JZQ4PXHcy5j1TGsqeqbevrSe5IW8YCIYV/ETViyEUuVjboZkWUfUihiE3
mLds6q4f5Qp0JqCsP3Nd2SjGQIW54ceRWz7TunAo1WnRRQyCBsYJQfwD5+GYFO1b
glq3vTsfYbxZesGWU1/e+Rxv4dPuU+Yf6DfklkyG+SL1w1xhVktwJYwioTbIe2Z3
oErsGInwC1g2Bb2FmZ0+i9PsNowM78HupEyd1RWfU9b5S6HclhShop/SOup3qTL1
4gi/yWitWe4H+vf1SsZ1kiURIXw5h7UfuNBH0/oEB1xOKCSsxcO/DRzv1ul2JvPi
pXSH6mxamDptTOgCup9lsynT00b9V165tPvu57Bq43nm5ZloNP1r7QN3kQzL57rp
g6EBPKmpGeiWU6W8oZIB/EAg3T4X4TAuwUiI5mb+Y550Ijau+dqwB4zEwHlLTReq
5tZCICMp3fgmn4pPBai3UAZXfS54MRKiT5PzP66RNA6EOBOoleza+zHlIT2SFWuU
0PW2nmbfjUYztGAQi5TkmzmR1LeuBSlA39QS2I7Ts6QmJw+xcHgP/zuYXtpcW0BD
u1qozxXE9HWyiwd41tITcVhlg5Q2vxw6CF4SwBHZDa3MP0J+cj70Tdth5UvL6B/O
pbxa2U9YmktlwM7pLmtWEA9bej/3kEcIHtPQrcE30U5S7BzEixRO+eS7/eojQ925
xl3L6CaABGjxdj8Uz9OlImZSgzj4UpNiDRdlGV3t4OlCFjtmJR6bLEfeWRFYzRWC
bsmoyzHo9VD0h73AMOcvIRk8cnNZogp3RwHMJ+k+QsAjcm/H6aa62mg8hueccBzS
M9UXMM91ekefjs6kRHX9Xb1K3mwNWokiy6ExPFfc3V+0lKxb3EgbIkqiwBRPMzvI
u603skKfCdLXpSikr7QoKjfBC736tvO11BgUA5U2TCeMm6imhhVHDhQKBbGA/vSZ
t4/bIVh9hj7/qVCPBBvRo9rQFlIqddBn5oNrgs2LUsvssMb4LhKV16qF4Daf+nby
oNyXhLjQLw3KHeksLpYwhRdTngPBZKhXICLEzJLGPsUY6i6qQsj7FWytCjjl9AX9
kewvmrhvIUczSrEaauX6kQFNFa6FvbbFwRMhi+ovBWaStaNvOtuuEyYXnVw16MLX
eLGJjqLeQHqXJXKVKg26eY6dUn2MkY4ZRJbdzucXcaQLqn79LRYGyFVGm9QN1bz+
sRd/gDwwtsO635I/fwaDj7XuTcCM6XmkEN65Tiy7xwMmSvAnWDYpJYAiLXco1HE0
ehQe3CSmeEiZGvaJfPohlVSKUYRnTgfB2Ofof7Z1fkYTtxkN7hf4OWaL8KxdEHhs
rutEAhgX19vS3In91yyfWkvmgbBzV46nk+d8x05hK+HoVce5kQFzcMHT8nsP1BO3
6F2b3/oS7MafH/HKOJ94doAzxu3pP3w4fQX9T0whYUNeUlvDW8LTTl9vm2AN6yDR
cmJRomw5J4PHpTa8O27/8dIgcJczJsb8sMefUgLsY3tlgCVUosoBgS42/DKDzRbp
I/FkYdVQg+C3WgiX/CjQEgGYaOFz9shTD7lA5jawi+JGQuQ1aje+PMTggXpEQkir
WPTGmNl0cA+tJKS/10HK1G95Pky5C7sCkr/iPKAWcbQp7VFx6HSxCk9MyCs+Z4V5
BcUWUZK5JgYOXDwtRSEKBsF0FJtmK9YnTsX99/M7YUtOvc+Bggj91pvw7SpbjXh5
G6X/05SxtjfTlcbx0iUy8cbGBWR0FRwMvyns2l9OPBCABLCdloKnG51Jq9+Ize8Y
2wufrLG4pRGWeJgZQZQQq7hXQSWtMntUxtRe3bps516mpEMlVmREWHDWo1r1XTcP
rhU77w89F6oq6LCPt+isRcceUtn8jRKGtPz9c7mTt/dlu5CUR7l6sj3iO8oAQWqa
YkPP6isQsKRxr0jFWVj0MaXc6LHF//dwTG21feuTCjY9RxKvlqopn04ao36F2FhT
cXtXCIj9sjvXmMcsTbgt4Q0K+HhgTl3kQNoirAnKh2KeBWOqZI9WzW6wx3wgZ+KO
KP3f3C0V+fyXDfJvrjS6db2eD4KHNj6p8cXiWFAbZpo9QSxIbSTDoeGlzwHqOhRL
faEetvBouEgpgnyXVM81r/sVtTb55rA8t/kMNUICltqOBeHWKT0s7BhJtdcaIHLS
JEk2a/39IoUaCIVAHkMEiW1RFJq6WFJk94fpMo9Nu98q13deZ87ifE85i2vD6glU
+ZXhOxTtmzZdHpxIkMjlyoYq/9+0ufc0U3QGTSqNyXQZSRBL9E+ADauwvNh6mBnD
3XQE0yQwg2KNcSY304SLYRMAMcxuzG0Q/g2hM9YzmP3XlcxCidDHSULGZyeZTe4u
vt1Ghd+mEYD+qHpGavtXoVhREnsjLmu3iLwqp+4tE7WHh5QgTmbJA9IJdc65UdjV
kc7IjsBa/9OCVoiWvRUUYkAteZ5omygapqhFjywM7Gnp5WgEkhWnl9TCvYeNxfg8
JFLY98Doa8aGVXG5YUTx3P3HUbBV9BdDjfAWQsg9lstocqEaxQG2+fMNgNeueiiX
BEtx3t6Gfb1VUKvNI0CfnvOKk4BJ58JghZwd188ujkH7TOimLp2kSZq3N51hN5QE
10LtNo7rpffjGw6VNSbXz9F3koc2mmr1Nd+n1Xm4yL1k0OACplZdjX3vkswwx5Hm
+z5K5WXEzy0z5yFeD2GOAvZq7DJo1aWaVF17xm1wQhi+bSYjAyYM9tVfvnVZ0PSB
edmAE5FFxEHbi2o/rvupR96HJkJvaM0okNHWFTwYV+jenM98/DgByUeEzGPaPBjQ
+YAnNwXww1mgrGE5gXQzcM0jnWsBN4Kn3rMzOoVchey8g3RPcMwgekRyEPQ2nnq9
2P3w6agvGyXs1ys48y95BQNpb73n9jJZcaD4Bs/r0ICfYeEd1PMKm0OMDBJ3WVQB
2AIEbXz7/ec9E+OgvEMWPakm1ENsKYthmwLmZNFVcvIfftB/Yt0+5NyrmKgqtGtu
Z2p1F7L2jaOD42zMvwISENAKlmYw+I6U3mXcoJWDcTZh01qIZ5QGW+oV3A7ddTzy
Ff6vYCLw6iGw5jOVMiMzFqZEOpN+znMPC9BbQFl2XVgixdTIumnijGKH4HKPPuNO
EeSJEzsylG76xh0CYVs+s9x5ycIkfHkC+8zm1a23XfRvRGwMH3CtNCmL0E0j/BGP
/vyJARSnINBl1WTno18CQWBI68QriV3KFqfrO9LdcoO9FkA7vky0MaO85aqTSoq6
YjOfBLDFsR57l2jN/8fjw6b07BSkcedJ7c/1LIyr4/4JTC8W+5YbOoeN/9oS13di
WNbQhdJjb5LjlaFCnEPL93XANtag2unJ/SHKjabldMaVDeD3lcACEcqJC1W9VVsn
PrkXShS3Ohtgzw43CoerHheJNTbupYRZFCKI/1OZLP04kLC7BLdpgQBsdfKYvRjy
O+c75feCANzSDTkmbEnKrYwvvCDao1qSgAJQ6EZG3DChlHUZq3mM3oaYjXt9h9zD
XQKI7JC4AVJfadM/pXWFOEcunztK8y7+YTE8IsSwesg0oqSPQZrBqaKc+aYrKobE
QfQDe6bdz56dniffUgBJH77pkg44IHUJN7RR2Q1mBstBQZ8j+BEEAorIw/2QtN4x
F+IaHk9yqfertc09ABH9Wot9dgZ9Un2d+o0SpuxNba0mM4m5u0VNveFmYLyLmDed
HpRAMbOLay6dkkQw7SAHO+y8pwFRms+P17prSs2Y1pudL6yHUpmGom42o8RehbHH
IzE/HQsRa9aAar9/KipjpeSx1rYfHzyrEpUgrx5JRs1yh0p2GiObRFWrjEo+pNzC
9+pQ658Rq3OMg7Rqhbz7++6quSBJTR34HLAYZxJqvTI/kcxQPshUQExI2dw7jKkp
U9to9fzvxAU9vYGDYJ56dOFKDyuwV+igDlDV7DfnetJXngC+t7l+5+m+D0hOvZ9T
oU+51FqlVNwtzGaYJfn6b4OpegsvMMedJUtrA9nLltf99wjVpSM/tppdbq7sUmUJ
gPoFssI4Sjmvwaloukgw9E19dB4fHYgiiAnsYg4DWR1W8nmnwdGPdIaV7KuWJm7A
wf9cpO/ON1KhA3anpu64yqwQgkqOYITnVvOl+2gyTJr5ERRfZA6O3Uj067+e0pAC
r8NgdCOd7e+FIZiTMKPnITWl+Hp3POe9o2nxnKCTp/KHB9XzQQOJOdQr+7tWa/sF
WQcWk1PuRMg4I2e9PCPKm+W+PyG2fitd5vYSUGnVhc9Y56TNp7o3YXt9VEYOsHf0
bB89Le7jK8G3OsUqknEvgQ7rEFDZDIAxwCjwBBtLMclrlKkt8l9bvOyXQj/Ih/kS
1isLCG+2sCCilyBFjW6PK9FIWaF6cIKuQNw1F6VKRf2y08jmL6gEDw7IeEUyETky
RDiiAafs7oGzAUo+5uaOmOMFZAfeKEeEDyCT0xRfndFEuLlWk7JtfsHjPXQ4RW7W
tj+Th+S83t1ACeoc7g8QvOmD8SCJGf1dGTt9pQC/JKMQTFPsxla+ZJL8sWOcup62
HOmnodW4c6H+Ml+AvqxQB0TfU+Mu7Hs1OFqeIYE0o4nbEgHrsKa3G+vN6Wg0o6H+
wwP4GRqsl8uX8rY0GeyVbI+8n1uq4b0etEtvWkPEWuUPOJxGtD9xg9rX9Y7P0Sp4
MiHrwHjA0bW5jTQdEBUCj5HODoL0BlZR64AxiMRX+NnW6ubAfBfeQ6fgdj/lT5Sg
UFr+EDUQOqDBjSKVfWyzLQAhkMQFTusqFm6r6N7C4JbUtOaosSk0aKeSBOWf9f0h
ZRRRSFA43g3EfwWBPcUav/QxMbcOyxPYOGKw1g4hEkHmRTcZJEYT88kUXbjpTj+M
QCQHSDjr9lcykivihQ2Q/SDhiJwj6sRpygWQtUI+8oOQyioS9TSfHkDD4UEwQiG6
6toKMhyopoJdIEaOKxlqMSZ+YcFWGY/VoiAF9ZB+8o6g16u4W6b87R3nd8soxbxF
B8Fca8ksdyntmnvpcGG8QdIS6Oyv0BxtoHud52BE4p5delogm+jgFW51pQOdLb40
sSQtUt0otcK8I7WpU2yPYkb/E96EZJP/+i2qIk1adi7Iujw0htM6+cajsS3sxHhT
9imfC0UCjStA2WlPiIqwmD119AzX/LqL5Kc2mNp+n4z3TeKW50jD0BNYvxiEyJG+
d4UGTMPLNLUhvkZUYcLW4xJtMdkuIYLfP6kkBsVeRzkBCoti7QshKG7TqyFi7d1Y
f8hLEsu44dWNmBU6VADUElAhoEdDtsSxazGFuUF0SKuBosu+txHLeHNH72RVDhc+
hvFnYvRKfz1yohAn1Vw0WA1Emek7rO0+jBLszCucYm36cb7W4nZ5wTBk7trE8q7p
5IgQPiPbVmzL81M1WIO6rnyIJ8xYul6K1ho8LU/ChsunO4W56YAW4P5uAzKMe0hN
gmguNugV+dET6ZPZWwoMQ5BQmNsQb3lpcBc9yshDLR2xrckU89bsaX/4gI9+mL3B
`protect END_PROTECTED
