`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jx35ggCFztIDIj9AsBmfSkuemIa043ZWSOVxXXBtTqf4hnAg9kbdoNKaImsjLtt/
fpmbIO4uEVBjjoPgfeU9mJU9Ena145jH6zMqnQVJZl3wvhrOLH29CW5uhyPUBHCl
ebv9fJiQV+lTaBWf+LkX0Xs8o9qi2bMMXbkBMpzV/pEvU40+kC2YX/7vvRryVhxy
1zJ0Pms0IfcLkpk8YJJVpZDDOW9HazIxnKoiRz5/GrofH09PWdEkhNm/crsK7y+d
YDgn88dudu6yYXDeE2er3MolOvcoLsSDN7Byivei4Rdgo2yHXlwLsWKZIYYgJxeQ
QkXsT+6Dp867+IRHSAYBXke83857dQVwUKypL/XsUF0uSQEivWZZqxOU0ReI7spV
qpBW5yXQgaEDawh8PxcniOuhrWqwep6acxjas6uZKyR6kCx7jRBDpwYemkvQ3Pgu
ool/86uIM3cBY4z9pI7q7XBFWgVwv1VXM2LDqqKZRWwFnP1NAYYiB5VkMauUu9xj
mrMeKhAejlRdew7EqnH7pj8Au3dWtyeTss7jDXubSpBv3MXTzr9d1OVckKy7ndXJ
WmKpOWSipVjLqadR+bJkDa0afbSNtMbaKOZBPEZjsBM2AFKswqEPFWWH4tbzLx/n
vNfoXu93Fycd/Kb6f3jINZYJF+dcIG8bibEXVccO8xW+yXdmSybPoPkCNVKtUglf
VXvS5jBsrHk8U1g2VOyYEKytBoNOkuS6PODiAeIqejvX6xLzI+EWCMqehIoQl03Q
B783TScEGAtM/G8HlFN0o3wJLx+LqxN7S1DqdHMY39LQ8RANUJcBBAq+rOhW50gs
sHYldvIeJYpdEil3NJy4VIcFElvG2CKGlOjVhclulYjZzT6OxaMIn3fYtKrZHW75
niilDzSBPJD355cRWh8bCicGeLJUisH8veyJjSBEyfIQc+VjPXr+QgfjzlUIljAm
iv+GlgBfwcUtRryO02GN+dGAjf3oV/6kIOr3p8uLVUT8sWbburMDjvdNOTfpszjv
VOBmw77lilJTLfF+Ke7wLqVRQPwYLzkwwgI10jXlVGL0NgoDt7Ob5VxryQBmu/t6
j+/VdtLsYD5jhcCLQpG5qLcgSRB7Tj0lWsdsNEfkpW+BxziZxH4Nh3id0pEH9upG
Y0GwQys2wQS2+6IpGK8fObDxpdyGVMY7DZ6XoY4lQW7WhJrMvUfr7wLLP1YUadVT
/1pnG09k0INO/QbADtL2QWfSGAvK21BGRofU6jKyMh6Fz8E/xmzspRlO3MU+Rcbu
4+OnucS41QQ/CRR6CqKSw9SvRz5HJO8F+8YvQA4xFhP2IUnHIx6rTTpR5s9nRTV5
AeRNKDR8Cw4FPM823h1CyIni9XL3gLHV/CmYdD0K4bGmMqdMe8xGfunGRjPrWSbC
lkglwjkBReYmccRKOpI4MzfXRBpyjj1vh+JlUO0mSrnL/OuKkfRVaGZfgGWqJpE2
LYtrNWF2jttGwBuOj4jyEpm59ZnNiolcYp2QGCQy1jLWxAQJ1Vzv8iWTyoQvDKgF
oECdZABvN+LklUEvkIq8WG2nLiQn9okA6UGmSe9fUm/f0xUdHG5rd3JHtxP1/eaI
2H2t/hS6PhFF42ymMqjRwB8At5SGbG72t3lAQu0GGGeQKD5fjo5y655+RoryVJVZ
ulgNr8LNAWA+PHOsRCUIdSyB6dqU774pjA8UHj98UhsPyj0POQ7f+MlTZAPDrj5e
6QMeAG4HAe2jNglCSelqHqWbl+CvBRqO3s+C4qNC3dFamK7QOoSJAhQdcquMBqYk
LMEjI4LX8ac10QaNoAO74qpROz1AsGm2D/p3gWPoKFWINNlUP4iQrTBayc5fimEN
`protect END_PROTECTED
