`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nc+Ln8UUJQBo7S1BZeHqkG5L9Ud513M5Znq5EYQcuuTfGmn30ki9Zz5GcVWphYb8
yUl2xp/hWvumyRlOpU5vWE66vJ7QAii0ces5RCvn4Zy+I+7WyIn1qRbDhSf0zMda
pTF/Qi3HQrx4lB4msoIFNf6DDKbelaI/EG74EOydtTrs9+9txgme3eGc5cHW7+XV
AouSq84GotMJu8txxBCy3REm6am+5ktPUpY450OyK8A+vVk57IbZ9UdR6JZsZZLh
3Rl/y6MddO5hiYkGIYmSlBP+F5unX4bn0FYTqFVM+NcN4j6V+emvbBdwTx87vr7w
O9JNvLWBuaQzxRGnpRrylLnNDANqO6hDgybKYurEFL1OpdAYqrHz+Bvj//uiwlOS
eQ1gRbQ0sKZBgydYJnPXDZol0uJiv67J//xDk0V9+agIa+CpUTF3uHp+m4vyDoeE
ecamqFaxbv+qyKEqxDLJTi9qR7RdAaQE/v7Rt1hJsQjsies2S3CWyiGXwlTfg9ap
Ty1XON6KFVELVtCt4BgevPZdfiH+RW7Ias31lANhAJjX6HwvNTKLJn3Kv7IUqCmm
AkF7BVl1lHe7xy2s45AbJPf9jiBGZ11OJS83VXqKPaZJJmt/DZyQ1Q0yz+hwLSrU
h83oDMP9DtEq/8pvNcyMQ3D7oYZL6dBYYHHUle/DhNI9/ItpJXqic9F6sFZ1KVWb
7tlE2415gMChqBW3Ms8hz7+kcUiCGzgEgOPVafCeSpTotU2mgvmK5u5jnoSRUYA3
90VGoCbmruYBlnbMe09Wkq8BRjWuMMmh9R5VHi8/DNeYH0SsIhnATIm4pYKN5VS3
szYg2/Ylx+gXEq7laHehlghRR2h7lkI36viGexcw+QRC545xpTFNn5kLqGIqH/gS
tvw7NikIaF2MbKnalKkpAXTlmfG3JRULo8INosxzUc4bttl8vR9rpfJMSUfTkirA
oQAdbyEXaGVir2t/JmaG1zB746FQG8cFdKLOGhAn17yt0z6gsF6DNwI0yrhuj+tc
r4wlMzKHwJbMuo5bISKPSG7P3XhKtDVoteFvZSI378QDLK8n5MywJijVFC4Ci4Em
mFlQfNKCKZZKB7n2mW9DbOfO1d1qf6+LTaoZC/a5sxhg6mUS6bHxHU9yO8R6EaFm
oSNCiYhlA+tVSlDaWx2Au91I13rZAev4+vXh9P2IsaiMueDoSmI0PyKPFeQcQ7/0
sXF3JNg1Cxom/xCwLxV632OPcIU/fgz/26GFPcbEEiIxyMdFuR//jPgJZXyTndKA
iiliXRGAiN5InyCeIhEl07WEMgd/2IDbNenyAG7P9mdCQusBmlYb3OSeLr9Zw2EF
kBhggzAQp7TZ6XZ0/IE11FC+6lMSjiVlXzhG24+P2VeHoRstVNgMS8KMDNQM+5nN
5QYAKATe3meDGeIBgrvb+iBiuAUO+dD5WqlAZlQ7tCiHeiwiD8HU/xDY/jNMZ61Y
tIdgZjTmO1AMg3g8JL0aqfy5WhtHMguGqmZhT3SKB/Iw6cbQwIWL86LR11EZgvm7
Xs0byjMg6uiDXGleRvOh0nPIE1F1i7yXOYn/YH8hvu4BFVXA1ysnWKgiradiff3F
O2tB9y/tBnu3Ab6gvE7a2hK9b1YtT5vNsxdJkM6/jz8gWDLuMLRsc5BQW2SVzH0B
Rt6yZDVN34R8E5DxzrQgAKImP0ZBuvkzWe8f2YCgYzkWh3tVP9oxQeMoxXm8irmz
DrpZJf8aq3gtNh1WxgWrUTDcrBbwLw3WA1+hlnO9kUYFmMAMZbnOkceqrLhbEa+6
8v4KzTO55PvDDp2JXrhRLHGoejKPh/txA55S8UCG4ZKIQ5LDfXOaEv0WNzDzSJGl
Wb9FEyQuI5Hr77+t1G9TSDahbDfXs7M5DOUPSfR6efNuRlg5X/KTXed/+2+ImZSf
fJVdjApu3sKDnYLJvELoPkXzaui/SN3htQSTLWktZFWivi7Jd9CBk+WxRhIkLAaT
+o1V7aiCUi9EAiEH+OTvZeLpy1A+P74aIsxIxHdDheSAslk6teUPivw5hzJwjvWJ
+FjCi/V1IyKEmthd99/Hum4FuWcT7D/eXBo4D3s7Q420lIaB5aCm8JR2T0MLzYwD
2MKqDDWsjPZ7HJw/Bq8G7aLxlO9C/FroLniXDekko26QemxpooW2HoeZh18kwPPl
1ydpkBTk8Jsyc9nK9L1uf/8wWJUkbG/1t6ylnbvJXz0uoRs/bEJFJcCNfeTqLOHv
NzGDzfQhWdFthbUr5nZvO4SuLplAGa0w6O/fxroibSSYJtoVSZqprfP5BHHawGul
FhGOfMVWkzHiLBH0Oh5d0dGrzMR6xbS439Nf8m706Criw7g1CywJdKWsbBm9Zkqt
3xVc5whS/YysF/46Vj5I76+PPknopLAcN/djDqV46DAnzZpq1p9N6/dfULnc5x8U
9v3EvgVZjhQzHbpTun7tnkMXZ+jOHbhwPl4L5z1769WQM5u7VZ2U553vU7qWrflu
FIgK7t7PvWvK7LyuPYHDlsfEHWT0eASwdaV6Lp/F6LmpNoDOiv/apGW1iCAxkvef
YASK7sgNOXLXObc9sk206O0c7lQnOedMFuihmX8NCZQh1NG5VsP5zYAAiEr0ODZ/
hsn5RxX84pR8KDpkksbeC+bncrIr+6NfHSExhDcNaQexu+DsiUIevGbwuw2FPn3L
d7heBEPoF2+gP5z+5SWBNfSaLTzTd6RlEq91xtbbZdQM5HCGHrUK2GlyZo+AHo2m
s4GJ3dH4u2C8S6Y4Bl6TfL9rSnRHWjlXAou0MsYl7Tbd9oRI7H/18Nm06m+6T5QC
JFMeJF7MN1HNRsrjIkOKax+yeVk8aVd8vQBgZzVJqC5JhccojaP20pa2V0tBusMn
MTcc2neVLGHh3f5IvEyf/3KRCeK/cE0XVaHK8XExZiZjScBwjSNwPAdt3C3r81Lr
n3xLvd5cP9KkflUl+Bw/DbsZ+LOjEf1qCN9Vo2bP3AtxvK2JPkIOp9X4PTa230uA
sgxM4DUxxWr5P1Bq/ch5w6d+F+783gvS5ZhDbWIPTD6bEd4zxaBiCE1TNQt3Qe63
TEWYO7kBhycJ5D8/QBP880CB3mr0Hx58RDoSogsS1UeMXl61lKr5Rc3yA43sKFnF
9vK8T16b/O1CJaKn+s/lvmsQp119EaqyiX9uO2P3DJWwnu3PpSasBMRvjijwfrg9
h5cv3mezWhDgsbBTpWgijAyfCLncuJWE7lJDA3GtaTdHQsQn+ZJjBSudwjpkngSN
m9WvtIyKOIabKm/RTwjKuw==
`protect END_PROTECTED
