`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8GHZMC6cylVT1ATQc775s7LYHcixYYK5zVei5JmyGiEvRGwVPLEleY1ud/8k3KR5
WAKKJPFqacOy4R7MfllIl9ttCwzjbn9KBe0KvXaWZu2CB8lqy6fyN8g+nvGboVZi
ci9iA4TlZRxti1D+mYnIANFjqpFFeUnPUK9NCLpPZTvil0tHHXmhh++r4OvsEyHq
Emjuv562QyEBQaaLa5f8yfP+Fht/0CkemJuQfDnszK4XErgkdwxyn2SZ64X5kneu
K4Z/FebefP5/WRjjCCdUYBHUd4fn1fEouJ57J9Fl5zAf/0qXIlf8MrchGE5KXoaV
u1+iR870jj/wGC4IbXLzImr0tUjgyGde9O0NwaRq4NjsT9nGEOq4N1rg2VYasIUd
GFkUa78i+QngvLFszsoaLThfFhWHeeM22RFWAEe/0MMq6T7e27An8IB7ao9DMRPk
J1O/oSXKVg1i638qxNrjE88kUA3MLWSLj1pj8hHyAFZYiHh2VJfEi04HAcQ9+hjQ
h/PjHe3fBCbxv9liLQce3xXK+23QOJQjAkU/+mVlJ1haaDl9aFld+2iRECuT3S4u
59Vhqcifi1ffm9RrO/jK/9/g/LS737vhZevV3PqWurAbQnBqOCK8bsZ1cPSdtKCH
tRrnt6kidcKSwOOfCTJ7x5rfToESJBHK8jogZ2r3p8ljpacqb6sG71y1B/sXeJDI
sXm8++JopASPFXk10APCaJJXh4IdCY6jpRIScnByfQyfkt06ynJYgfppz0+PL3tp
8W0trS2YbJYTsD6HK1WQvEN7eQlUBgUci1409lF4T/hHrPfVXuM5eJUW5VlkreY7
qas/NPQJWYiIRK+Ivk9xPgLj52xEh2YRRkke3jzwddpWIhoF2oBAt8EKhCQezYrO
pgyzntheomXQHV1oZ1NaHRFug/nEOmEZfLeC2ng/NGtU5Q3bqV2b8htcXLEhv4+y
pPZKYk5lSM4Di1c0upwDr/bD2rfkdE7U0V3jFA+xxiWLkE1mjOrDUNeMWKEG/GqP
k5GsA24valvEqNfpugBMraIWpD50TC99SiTnfoDeC0cynjwwmVU3rIAduMSwiL8F
kXw3ANaY8cfpgRSW1SzJMfx7zpQr9/nJ7Y84EoOXykMxglwuemwa7tStQNGQIOtY
DaBfd84UCjDXYhhRTGO7c4EdBuHDNMQpalNqpgo9bxcZNMUpdV0oB6PkIkPOiGSL
kMhlzoxdqFmlY+62eVnpM9jgx++Q7n1DDSniAp6n+T44X2iW+VU0hYTRBkCgSe/z
pohQxAnN2rnq+aroTqtViwJubcmQLIRKpRE9xCfyxP6HLoPepfyHYiMvPgBpO2io
+YpoMPc8LYla3Fkz3QX9DlYvpP0YW61YnUfzEzcRDxu1UYKYxBrYtfPHSpoBBBDc
RnPLLHzpc7+ApRLFRQ59obnNmsi0JRadKLOiKcWtIGshmvahHXtHRCOuOmGsL3XZ
P7E1k0SFMzCJ3SqSZusQfA==
`protect END_PROTECTED
