`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yasmaV9lbAiD6zf0cFxTI1A72v+CTXs/+sjszoOMkYZjEqq6LM0H7su2GUreYPQM
ulJmIi0lTvHUmt+On18u58bg2IXGZ4QCVc7FgPHxNPYByu1LE1QCg4HkUbyuecul
Dsbd2uNGp7jgaclqX36a9WaGO86grKbGHoSd5V32CpLt3D+HSzDfALbHc6QWIC1B
BdgOdffKy3V+CF3KIEF62efTlsZLrtW3CXyFL24tL5SNkSakpuxaLOcxAGujXmjU
dlt7Oxe+O1JRH3wIieYpN5OKwUZg94tLLLRKHjIeJy1xGxkCFCz8RG6qOeuQmiZf
9mCEzy97ERe2n70Wkjc+hXP8Z0zNXQiJNmWEyvAV5EUt130xYnCt81vkcr7LY6Qz
qOr12sOQK3NabL9fNEACJELFzWH+7oxfxwDHkEoXouzaITBVrc1Klmhc7VoUCd3d
8VPj/zpohLNoKuWcozuBsw9H+9q4KSheQ+ggUFe1b7Iz1C01BC8Sjqgh6SRW9sLa
Cxfqt41s8gu9LgAgy1F9d1A6sgjll7IwnQIemzO3ZPCa9RmSWF6l6lpS1+qj+iNT
kPQg/4zJhjDQBvMny0Dqo8r9YGhfu6fCljWxTCguaM+pAXVZO4muhAAVqzytGN7h
RkS526lnE0AICG1OL4ZCUnTIdWSnCHDQxVgVsLDElDULz3+4P+HggFM0VrOqNFiv
uB4Mxmw/syL7w2xIUW/5h29R6ZAE0RIvjpXqXFaQTepaBkZ4dPkoDZPs0KSwEyXx
+Om+roHfHUAunnnBQ8+4jQlDRjkXiGkZWi9mezJAuT3yXdu1TYSkyjicO66Vz6+a
uNzcYa4VblhkLfofruiIi8Z9lgJcOqawMKfMuaurgnkl7Rm7eBVGDOAG+81obzE7
dGDREHX1fJOJzABqZxH9/zBBdep4aGx0JDOBSNuYPLTtPlvTtW8m8PYEt8oaT32W
pL8eq1u6gx1u8bo8VSBHY76qqnudTNmp+i/+LrLUGPmpLegPE1QY1/k+chCFH4F2
p+b8H+tO8T4J3CUskEWkOaf15jGCfruRjkI3ZGEPLU0U9OyZ6VEGpsmbN2PiucJi
khC+8XqOCJSH3IWMH4inwNrKY+v/tsTf6qKdh2jk8QeqC8nb8vn8GQyFVsr/QUwh
fl0+6hS3I9/5Y2v4Aeg6OWMBzvbrpojNKPXA7jKreIGOK2HRzCM2ZNByRra3aGrZ
Rrz16zKYyD6k1j369qvOxrEZd04cxnzjHRqo/VWs5fMxxLN15rKTmQSO0TAw3P+4
9m5V2Jxo3M5hiir+szEe/Z3Defu1eTWev8swvmWaoqjYrpcjZrMruUIMxpLbkqA4
wMAl3Db/Yyj0I8Jrnbu/F0zbqrzr6q75peYE3fch2K9DK/PECo6uMdttwCLS7ilf
4BpJxqfErcvta/QhljMFYUUUbZvqNZBoBVz9f2hLh9JnlOol3tmVYzThZ2kofOsA
euKvBaw4oGT09UQ455t2JCSq0yM3OVpalFQZPg68ecJf75yhPWe+IPAL+CcRV219
aVI0YKzX8Skw7cxy0lV3IHg3Hi5xLtyJ9WfsaBseYGW2/mP5RjwEixta9nUwzmHH
UoLYdzOHmeY7h5OCDe+V7s6I7U8HhOVuRbpmFMfi856anot5md2pz5gDdkNkl978
l4ENpqnbj5otX04E+OwOaIsddaZafHrkf43h1xFy9qGYZZiypCneH3CqnF597YXA
JGcOJMvNdjoWyJoxk9i/khQ924e04/TtErwx/yqQrZEc8YoFOoLFQth+YbXq9YK0
2hmai3+bgbNMjOVgPZJ3se4dCX1r98L8a94SsN6yMlq9H14motyCi+2fx/K92MLz
6u2GKKyzCX+zdxTneuTOOHZlmzcidycEL2HH3waNjYFZI/37ZO4c6i/XKAhQojff
/GsfKdPPn5erwfGhZCwLngyOk7Tkr5jJz3K9IbmcLFlvpJuOEuvARlQ0TcXe19bn
WCbNnzPEVbj4vV4zlYbj/UEugvr86a8qzSwQI4kflgibElgFLt0Bh52mIeX6IE96
cZbaSQkM/aP9MPibcKD3A07LThPU9NbvSQArejRelRZfZvEUKfJ9tklJMzNLq8kn
8t67QJ3sq31IcC1KSIWRccPfj2Hq11trKenVVEvpsudo2kwcPAZtUdrQ8YYGXEDe
KeHrIXYMpcVBarM86Y5mqHkFhLooi7j+288DaEZuWx7r8OcIYv5neJXYSGft1hpN
K5ucE2LoDXmsaj+N2G68ZXTZWQAUvX6xyam63T0TEghBELf/RCLq2ZL6XGJ3lWv3
CQTm7xFb5FaXRg85aUTDmaoyjUfeg3GzAeyWMrJggXSXT7Oyqgare10xGCH3cswm
HlEIZceuN9OPaeBbBH7MV1WdC8IHfbY5v36MiOJq1yCIxqWHVdFByH6Wqkx1w6QG
kh/cAD5g5bGNRzNPiijDjGz7tCjBnDaFHTcUQkG4YvZKRdSyVdvw22zhpzV9OPBq
eme/h4yYPXqB0ZVJgRdk0g1cduY77HFV6BZ6ERx6rW/p3pv9WPirocl/dop1W5fR
xc/H19/X7qnorpmNh7n9JtNgyLLYSFD/RgC2WBEMJEL8wI9qDI/chbgD1W6Wec5P
P+Sfjck5bKT9a2XOK0XCuQ5UpncpknsVh5awrJ9zznPVmWKI2FlNo5b0irYKM25p
3WtIVnjNKeC+hEBLjjU5JkLUs1wr/LmIPFEnd2ieARo=
`protect END_PROTECTED
