`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xtgxAqUUlr+FBjhjz0hlvUF+v/BRINoCl77lDEDFWP0zTBFnJN5fmeRjp11NfISr
TzKVeeAgOLPnr04HkgbeaN0wWe2Bh746aQggET818B6Cock6/OGx8B3nEnajofov
avqmWrc0vV9JDe2xGkIr4kU3G0b9aL1f1d9BpKQhs+K/BYUMJoWy6mUuz1aRjN6L
Uug8tmZb2wREQ3/ZtfIxcMm2JRrWNgTI3MVb7/S/37PnvS9RDla2d9fqC1Sin0iv
EUEho/SA/ZWwK9SuytXMYOAyu4zNM4HaRmDCPmV191idY+UQfNMo44+TeLZH2Bol
Vjn9phSrM9nxmHWyHKzqWGRY5HHmZ4FYiEUqDA8E+Car/y/UwcIjNu5wMBfW4Hoz
Z047U9MWGm0cJUI7mYnCpVXBNNeGwQ1dOShMy3/fGvg+hFZ4gGxsorKCvqPeWx9y
VILI5LbLIp/l1uSWCgtZY5puZbnAQcVxB+S1PCLWpTc4b8oXkOeMGC6/cQgBtQyu
ERCG0Clj5Zp6a7vF5Ud3/KzBHhmPXCWUNsRPaxBajAz2gH2miDtHKdc9zY5TVtQK
96wo2Xel+CXFGVVjGhwsqExkXEUzZWnpkiiGQo101x8Zg1tXg9RViQ0Stkd5mskR
gjt9uKWnFzxMkH0alTVyvg==
`protect END_PROTECTED
