`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OaonvW3yrApjHGhxBE+vgqt3KSo7Oms4Mi0IJ59wkR16OGe4j4iI5evJZmQAUNDE
9VxjsVe+mICu2VWI5/9Z7zymlLC6Xb05TZZtjOeO2EdHbGoRIeSh9BCuF+75s9yc
n2nRM+sAbrVjEadfAhKpmG2c2x9tCeXX/lh8XHxOG0qPI7EAFem/MyYEaC9oN3TM
zD0cjuvqHbX6EjKrmURMB534+8pJHgW+NANfMpFqJOxQNxXuaW7ftDFuJA744gn/
7T2EcpRPHFXO9zswLV8bG7yu8fwrdM375cPBgiIcYmSCVGoGIey1HkQ082pPluPv
rgPOr4T4aj3aW0hbKbrElvLUcybZcgoPTFEotvhN3JBN4+kK/l4wOZUI5CSc/WCM
8TDD6z4lI/NXIoTApSbHf7gFBJGL4Bsq5lP/TI/Xq55MQdTxi+5LvuIf40Bd/bVr
7xVW59xXkSojtIzl1nsrzGqAyazKA6l73LAtvefeTTLCKrP+cxr76QmhtpwRb68X
ic4ua1Kh/rtNj99oYXRXoa4/ofkDXaS8LKIzgt1JQol5u4uZSnTExQ8KbRVlLJ9i
G6JLl7N4IxPSTiUJRF53AOPM+cWCqR1Lb5hQV7Lp9Dao9dcu8g64XYCHybFrHKm7
ZBiYPBJNGSAvzYlo3z9GpE4V/Le9I1IbNDhc3UZRXNrUUakoScel4Id34RPJ3Ey9
y24PC2FwKPuwZvHmX51o/5Soa/eN1GQbZw9+eJNluknz9kodP/AU3or3v5hQRhte
DfC8F1mlr+xT2jq8kOeHRA7KOZ6Y+JGnTxSXkcUYSijAv0EmpWVso4QiUDwnZgua
Z8pyLmhgAUSCzoLQRYgXkrsNpHfzKcNPurCg3txJfbdJGATxY2/3K56wDNHL9OpR
XS49vYjhZSuJU7Uq75a+dQ==
`protect END_PROTECTED
