`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WhEPxJPIXoTGIQ0gqmR2wKkjlahvVVds3jUcYwA2pjvo2MCzm1eLFwhNwtR2uvwS
FH9L/y/bPrh7AJ3fSk+yo82rfMMMSFFGjrml3tdC7u8tFbg3FNn5XC1tz38arIle
CKKhP56wZ0SLBeB80UY8zkyZNtfWev9EF2iKGlVNugaL3f1T2QkVUWNiRGzwugMR
TW3sx60w+66oT8+t0fe5M7u+MHPS+UqKK9c+ckmbJ6C/0O3azc2wzZynW3KkpUtP
HO1sXswC9y/xp6jiRphoEu/DJzWqVt+FtXvAXLgG267Pla9rFbcJL8lPrrNa7enf
cwIjmIYz8vao1+4ON0YvcDkpHNy8i7UmPlGEopAfMu45JrccIsqqGwVYifbYrqKQ
Q4n0XS25c9+zUx6TlOKRZhlrbhDB9hHL01eg2xw5QVLMO+SJXVLpn1gJh35CQGOD
MhxShQod9sJZ75aUe25YNPTr4oKc3TYaPhVYfIcdoztXRu+vawV5A7SVKxN86EW5
E2aiIUQE6on+kHdzHeAWYfVITivnfZb+S4HTBtkP7iPgyKsE4U5O1VE2jX7HW8Sv
md/aNTB2dHII3hOhAghymwg2l1iEvFz1XFs7QkJEUcYCDE742aUNyuvsBwI/bWKW
VkxO5YbE1yQFwdoqKVygzA==
`protect END_PROTECTED
