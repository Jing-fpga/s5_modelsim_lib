`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zhJpAoxN7L/AgrZxcTQ10ddqRC9vOnSUJMPtrRs+2Fg3rO3WHQp8InS+lZw5qDYP
0Yym8nGS1D5vLfiaqufxoohy+qaJY9vjgwuW1RbzI5T2LG3YTtHouk35+E1je5vN
1P/4+sONkAFuSakLzdQNMjkMyBCwgifkpDmAoZabfTj4n4y7AIigkclRvEroC6P8
YngRBu5DrpS9z53OWo6noGn2dmOQwZANZpq9U+Sp4YeWkveyKBGrCAUgLVcQLdJD
OwYlB4P4+qRpoMWZ0cUylFlPvRV6xEMLG8L55g7+Uoe6037XtpBkuGfQbWM+zdu9
jGDLiADd7yCGt1Nfm2zOP6h1Pl1blw+g2RBCcWgkRgjh6nqXiNoyYZXR77ea8GIv
piKT+qpyRpSDPmANugPw7UOk2Y1gRKLX8eE+RLI4SHkJN/+axHsltXj1tKuQ1oEa
28lXia2PMfR1+bKnrkQpFf0o4nc7Tmh1VXQKvoKeVtxYwI+uF1i4PSNx6KkWx12S
YevtFFvC92Bpgkfbiwg5rfOKFZt809x3Nn9RB5F5Wet2M2RryqQ11o9C5L+/GUCY
r3AOXM3usJAs7TqotkHxQf0XrSnETxi6tpoe4Pdz5GDezpigLEFnybQIMRC1Ana7
nRaJYnvESXG+BpCmrzmpXb/lR0APlg4ebvyXlzL54Gv5YyAJplkzcy1tjoNkT4IH
e/PD1OTP0LBGkhoZHvQDY3+Lld1eHvS2rd0jsFHX9BH79ASE+YC6Yv46RC3odR8u
sShN1NDcICw5igm7/f803wb+dp0zQ9cZAYNTUb8wauO0UwOtvnJixViVIr3Ygh1f
qNihXatrSUFN9M+6dfVkIZgovd759Cr9dAw9M2MXfIoyutBJNNV88GwH4Mjj1+/p
GSfodl1Q3/2rfbZ2/WjUxpQUesloCO6SN83xHpygk6fyfK2VB2P6B53QOeY0Gael
XQfW9YEdsam+T0v2a/Dmrk79R19Inp9bKHGgj1HtN7sN16XiUdeWEzzKUAt2/V0Z
AspbWahj4cwIzhKcItVZ+H5J7CpjNRo7Ey/X+GiyQn+TtKNV/L2RSlaNj5EZD8QN
hKfudV+C+OQhOAII1J/w+SSMxX3tn/8GQO+HzWJjcOXzXPQEKHg4Ey4faWrR2i21
CPYB8mVEXBAgkuWP6oS0ch8OW/fL9YHQjU1tIebQFGmvYULelBj3OfXzCjNA2jl2
Z0j2tLpmU3jd3SrI2b8OzNwRLz8SAabFjAND75YMzm+j0jxbJXld2Abs6GgOIgPX
HPCrDccjN8ozMZFAj+Arz6Y5N1k9S/KCaJWgUSSbm4nmDGMLqU0kaY0t3dCXH25g
HSQp/32WoeaDNg49/IoAg6H82RiRpyYm1tcKBjtV4tVDezIlKv4vCgSxKac969Lp
mIx6fgFfY48B5cDRefSeBq69mdnXcVmSwW2cuMaVOUEkYlB/w4lcCK6UNElOWv8e
9IXtIOD8LO4/EzEhhIHBumWVIIEf0NSTaauxclpctYdM9+istd2YajLx+D5/lrLQ
smVQnJgOFIb9dt5TRRG3sdSu0CkGRuO2gW0gdnHKhgipqadNh+/lm4TOD96DCTdF
jOMpDYYxaVUmBgkp3n1qYJt8Qh3iZWsMH/AemwZdciw2M4gp9wo10R1BpDcipciX
B4xYjx1U+hME02ttzAih8j/oY7iOD/G0vZCb8SJdDXPHh42hyST7LAMbgC/WawDm
lq6haRhjUaLGeImyei41yYE5kqJD9xLdyVXscw9sIhC3k6AKSd4Xkei/Cd/s/Cos
kcXZsikDFtf4yvZanIk1oBChOSYwm6HjlG4A7Q0zct/hfT5t5M2l67v+ECSVlwsl
oUbg8VSAQGnA/DFEFKjMryl//nfe/8WblEqUlAihmkKrRmsiZ+RcRy6y2hUWzKQC
M2LFUpw5gHOoGsk2fR9Y8CizIindbNDLx4JgArOLpjJt3J2uoDTnhSXvNnSaylge
aqDBjrciaxkgKw21e8P2hWiJOHaGUo6ndraUG78v82zqyS79tZN7/zpiVGXxYa+8
OjWU5Ab+2IIsU2+bkoTNT6DP4NiFv0ZPzUomyWuzUL6MDekJv66DlwCrBEOdhwMa
v/XTZFQGNSF34tgtnYpeEgCIRdv8IkzmcaPsW5ZGO7yhaIahnIrrURRPr1tSvRr0
OV+teYzK4OaLy4wYxxOFZkglFmgggCrKc+CYbPPbqt22awHQgJvZtV3Nbe7YK8xr
fY2P79PV8bamr4P5UlX2zDuGVOKouiA81qVsYBHv7FRqCa0lsZrOdlH4xNrs1eOx
z1FbFAgGuG2615ypJFTNfnIjLAJw/sNIt7hRpH0m/Zk0WFzK2nGI2/shmyOZtEUk
+BLsbpdhPk6dWaO33t4rMCAv9B3fTsXvV/FOi1Fu0kWJ2NvyQtFJYyOr3yhWv6/k
/JAj28P35NtG3buORzapYXq8ReVD/tarCRjyl6HwuHQBoa15bEbXnt0gbT5gfxFM
tQ1WLnejH/ATO4oxqMy9yXTG0B8WlGjYucOwiTxQposQGsrOUDVP8/3WXs4rly0p
aRFEiQiVH8zcxBGgXqZ+8u7iENP2fa9vMWJ2+ZqG073T3WRynZkDcf4Ywrb9wVXH
7rUO6srbNTFkKEm6m7Bgewl/LTEGUBiE0w16KKgE/HWa/tIAMlfrvEFwXC42Kp6R
d78wmzieSudBhqngkA7hyeXme7WILWLqWFeOL8q6UFOq2MQA46Y0rPV9dJwdmP1s
pCg5Bf55LeFDg41nzLRxFBmGsHtmHXMxscMl/pA94Y9PtsHuf0Cjd6bVI+VfBi5a
xGLN45pQmSz18mn9OM3O3naYBSaytOgaQiw7gWqD6jYalNgfO7iwLP8gDrK8IRpi
7f3Zo8hOVn5uulglV9qxX3bGgJkx8Mx4fj/wWzrZi/iF5hfYFkQQseoo1lxP7CcO
J9bkos+9IpRgFWjRHeYk3zA+5UZD2EpYs4h5CWueKEyvdvIoT4Sj2eAzAZfaeexC
E+/IFiJDadlHIM8G6P4U3V9drPPYE5OKMRaz3LkpphBfsotDYU8Gk7jfidy+kzVJ
By9STjm4GJrzr27xdngIeMzwZx9n813rTZnUaRM9Vm3VRmrOOguQgFSuJI9LcueL
Tg1e11jDWnkFWU65bT7uMCS+OknYtxFtWL/NchuAr6WtF4UynyoVnGm5kI7i7H0y
43PUEfJqkLbM4ADxBLBdtA==
`protect END_PROTECTED
