`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2r9hcUclQAY3WAuBTf6AbqqqRZmQuJhX5gz5EvR3Ux9RIRzPecSUofqqnuh+QA3x
FtgwNUSGrqiCWlCqG+BTmz/tOE/JGtQQiTbwihjffCLm5CvWh9Fg94eia+wlgm7b
/kzw67ZEegVlNeKsbyCbgY1Zti2YGVhkJ4z2GSxfq7hkwoQunPoU82T2b4wQe7R+
861DJr4VAnggbF5rIY4CBVaVtrX+WvTDpPaRM8mnY7jm4T9NLGpPu9i8TH+RZ9o1
rXUwPLp9ngEPtNZGB0qdZ0LsjwZfnmtbmooCS8HT15aRdexza4v3wRiZC/oOkMkr
7LEHIBg5hkSJ7D+2mvS2eFBlpSJw4Q1cfYmP3whvIE8eQSyC9YpsCK6qqTab/UmJ
TBgeNEc1o4yb/b41jAkFQBRuKN8lBMx2UWxeaOZCbKRbhi5ZC4p8c9mTbT+cGcdT
rO1JLFcy9czh+JhCW5b3lg0L6FmnBF04RaYEgHKqPO+ARtyxe7sCyLORu9ct9Q2z
Uk445xQ+AXkBgpNrWSpz2O3hnARtnk0ALJTcSAs3SW0aWs38k60JOUyFUhfkUzWw
Nv+hJ80J2W7CSa4zHso+PU0VQZ9qzl7QMgKA+gmVda4JCsVHlMX/Uktc6cs/agmA
MqDquRrlKA8oVAETcTH/sy+ouR/RolNjB8jSVpQkawSJlHwHwedQ8A+wBkjzlOvZ
YY4nkEV2Ttwxc7+W03TJsw0KxW/HgBBQRyA13AyxaxQYimSOHxwnTYKVYTRZnnSX
KXVHFQkYEzPgbiQ2xOsdR1V9FBnLBqwOLHKC/qrxhKy5foutDKuvsxgSdINyXKc+
ZCguQOClgqsmD9J1j1YkH+vN9Mdg619rvcRhFinv4bX8zWisVckx0LgxY+6J1LXL
pUBMBnNfEMnpnAacrxizWAsqpQMjShQc5SuHQJOOcGlFAHyt9skzYIvH8gmEfvLD
GtThzUjCU1pGJrI5edfsPwYH4ZJil0++E65kx8KquW8hKXQHL10vveQGR5+c7rg3
B1liVqejvee7AcNbvZkzqWO+7s3E3beS/lMH6XrIXBErxqao+8lNThBjeYfLMdWH
Aww7GmLx4ntRMj2AHLPUBX+jB9rRypq8RzMiF1Ajf9jHZRWnT3Uo2k8kaMk/L96z
7ROlBY0xXgUp9URviKM2XhmxWLpHBtrhRsC4czzCyBxMX9nNP1K+kW+S4klaAvGl
qmPU0xTqqMhJk1RUc/aHubOXh2F6/bAWgsYXYHSz82nxtmnwxwDJBjjRGZ4k/8fS
SeebFjjtZw8cr0Ff+/rd8sieOQwstO05ESrU861gAasm13mR2jgifWgGhhwYQn6m
`protect END_PROTECTED
