`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6+BUvIF8FQFSIZEWLcP7EPWnwrMUn0l6LiwAH25v+H51A51Kf79/sD/i5Ps+mCe2
2iqiheS2ByTguNuvKhFzbGsXz6OQgfhoVWcmRE+7k8dfxLIlWjry/a1sQrzwWLNi
qwAj+IqddlFDM5tifC4SfK6ow1ntyZ2zSHWWoz6e6PEm70oxmCBAkaYFo2glZYX9
iptR21C4dTbiL1IG3Q9Di4EeALG8EKFYdnAi0UFsE1Zr6lUInv+xS0/cTbu7hyUa
LK+klXh7lP3IO0RTFjEd9czGBtVBVVWcTOxT0GjDme0JzHsRP50TAER8ZzCcU5QC
OBQcqImTZ787Ck/Lr8+ZG0Sw81wPZnyqzhd/aF+L+nIn3ufiCXeeedSCD7cvpReN
NRNPe1NygY4/+RKxR/En4QMy3cLaTSbHaIwwufjdvO22UPUPBK6m8LVZix/ZUwvX
9USkS3jNHgHLeGkmfPHRG9kS/NxI+Op7hpmm8hGPEE/9cyoTdf53qi1pnDbIVLG5
obGeIr/BGmX57ymbx4FT3pSEUWt077RcAOo2iulline5bRrTMgmVrh3ZsqEAZVBB
Fb7MkyBgPSQ1Z6ydTToQYKoDqFsM2BbxvXD6TUEB5lpy4LTkmcHvNvL2pssO7z02
kZa/D4HEGii31388A+i/C8MOG+bMreBgmebtfYtX+pdDVMYbLJNKvANwYzSiYvfI
XWOEUO1CnTO9lFXycGu4dMbWn8ucXAOL0T/7RSXVqFyfFxDRqTDcm6q0gGYluABf
auaMYmsbtr0XTYwpM71ZLqDWQvl/dkZ0oMaueVdIPj55EUKfFdYNnqH7S4O1k0os
nOO6j6fnn3tl+2iMOLYpoftJ34a0m/HCIw6XVw/gXMrpuW3MGVMegM/ksJITAWtv
SrzYXifB0RVhZMDFoiqAWJ+ZsNawljteZecOkEJnVPfQUkgoWCNwO9A8aJBSCDKz
UPYWYKaKXO/TaYetEUz33TuQtyD53kZ42GEx/SOIeTJLCDpUwx5xAOaXOzn+Z6ia
jkjk7QUviWu0K7eMEiwIuQeIV9G+iQWWxbbSuP6V1LMOe2At2t7CoC9DeasWyOJn
aNomnNRtZQJpi8UUqFoonM3EuYhw+Pej9fHqdPqYKqZOSI58JdZM8llD7jOs5co0
7b5Idia0U9KiOUYppXa2SgeRMbJWf9g32yr1KaFOCasfJwT0e7w6pfcQrtrn6Zmx
6CF5At3m0PxJRSdpBPZA1fXysPN/ctg9NPJfy18jtELxeiA6xhQd9hpc9oaOqyen
XeOnXwpEZCEoJhoPCvirRkEFhJBzFNKcczcXRqRZ79tBn57ILEeTzYBqDod62qmM
KdTHaLtiJJx8Xtx6vtUidcL3St9B7XqNgmypXWa/e5MdHNiJiFC0ZXB23QS/KuC4
CgtQagLS6blzNQyazIDNZcDFAMiO5rXAAxcaq/Z0KMjbssJBlgO858VQqmDCDrVU
iV7RQs6a9RkS3ME2w3N15ogX0coKzKdoyUXe4BwUqSqJY2fouzxdXgncvCJyW1L1
yy0c9c9KLHS/HRjBOSrZDMCPIhB5sPmqXrBsBUNXlx46v49uaNvGgO4O3u6//5WE
RiYNt8XVgKJJctlBd6YxSk0YK9R52hYLSmoOG6M8a6JezBTramsJMDF8sNElFm2V
zw0nNN42Q1yeVZZLnfokGQAFHXQm3xhanDuq4rOboOHDHzS8IESB51mlYWeHZiPU
8M/iHcHX0eqF+OIIkdN7kUvxd0M8lrar//+jUubxTIFhQxnKBGgtP49Y7V38V/rz
FbjK/d8JPOkgG+RfmS7tiPjXp9A7wrE5SWlmrps4ECKn64Sv1OwcUpgLOPAppdB0
`protect END_PROTECTED
