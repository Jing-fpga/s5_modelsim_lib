`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
evK0TsQTKoM5K+V4jf8QmYj4yAsI2heloOdM88xGG3sNuSbVMI0zKJ/tPZDZnWJR
UOFvUJdJc5K/9/+VDpPEz2vyKhY5W7QPHppEPWJEk9R7NrwzbwyCNlA8pvVPKaEQ
aHGzHTr+fhWXyILU5dJNjD/EF56X/8w+uHHQzOvJNZHCERA8yywQ6TQJH71pSVYW
g5GRrbivIJtmIGXJAzu36sx5zfQD6q9OG9bT0HsvDAylhLHwIV4Td8MZnUcyxxXJ
WdKNeOLl8snDb9gqSkzHCA76iE9PkcdcgUjAfWrr/oev3BTavGTxlngbnIxDDF43
HYLvR/y0AhYGt93gcwNBh8sedNuXiTLvrHIyPNzbPspf778slNuTsJpQwBrCd0b4
/tUvaJWDQpWuIltNWSE+LOpc3Cnpo+gPj0Pll9/2P4VEcDkNsNA+HPywgQLxe5TK
vftUI96XjdE5AT+Vw/Q7jYRliwE7QETraZKB1Z7ws7VCz5BQW74MADerwrS3FpS6
sDWyj5nXX8k0KTW3yLP2yRsIceTZa74wv/kTH5k+nxwhvsdzSvE/sp9IStT3vfnu
tL+SqRPRfW2VViCbYHmSQ1GuI21izBlm+eUttq1FmcTDCEYJ7ekInEK5/OlcRL79
Tia/OAMZdF9ARHuT8IGv9+Gb+Zy/Y4B4qcvJwh1Dqq92JNSYjYiyHPexPb5A9XWU
VZKX/EnVIh2l6MZxaTkXGs4RjPHL2IJz90uQ+8xtdk5Ci0akzCnobZ53S3H3Uorf
EpTTINoeMzdQaqpAkYMaucT/Qz3/aMd0sOg41UsslImXI3+xOCbNesoIZ/tYqTgl
X8Q+o1QUzKn7CFt/GWyDgUw6vwGOscbFvr4UgbhSyChWplweCuyfqOC3lEi+I/E/
vvghNCCXSnQBvpM5u/0PAjyMvDDrO128Sm+aiEGJHPoYdh323Ip2txj5lLsbASFj
5+a79q5oEmiyUg7vMnM4Wmisrspb5nBr5SJp/DL1Ug+/jPNqyxmorq0hW0Gqjyn6
gKUsgak7TL6ZFt5YVS+JiIJVmsXFV8Pd51rJmAOiUZZML74jvzxroeFN4x+nmFub
w59ScYxGldnVNdPr/FpJJNiJoLipjaPUK19XLsaudoS4vfa8Cn/oznyYAX1sizrM
+4+mDEUkaG4ICpTzWmfFZ6mldVuahXEI91WJCbYDLaWSM3U+qmvcbZx6/fSJLn1A
3kykCw+3Pte0Ak9/z1n7UIk9oLSZh2jgXU76GERvzRxWMAPasPeXUWv7T7NZ2bwL
Y3qFyZz1TY5m1N4hM7/C2ynmzbIp0F7fQTmdmyJydc7firR0RXvIaR0VazyCbJMs
dmp7zVOLSOZHTU+v6PKzC/WaMszPT0nsCWD94oMwIiNcGC7FrnIUPMjjHYjVjXC4
amBTbOpcEXI/wtgm+qD4li0mqwT7qyOJquHbZgCVqAhd5kyMJvjDNRWp+f98EDZ6
846xIZF40KIYS5Weu2BjbhJnaAb1sQZjDiHL5PEBQjS3DawjPPGIk/oWlZ52Kr89
dmr+/y+tl9Fu8ucLSyQwTGyZm+J73fw0df6uPBdIaFS44zPK/cylE3rfC5TGFlmo
z/voqWFcNIwSVqvAUrWhqLqkGQMsvwvAMFwdodsoVu7V6tt55uBHesR93x1EivtI
6ySCgrGKXu8jk+vThE3OOWJjrYjpiAkMonGjutdBCfUuY40cMoLDYnkFYgmbAvdI
DKPJT4ct3rGFvR3202qDXP9NQBkcAlSEiXKamklLNAHIMwGWgAsXVxiN8LmrwjPi
UvEVmJ6okY7ubbR+2N56pa+0KFR6PWnSA/4N9nFaIJ549UsXk702tps1sIF59pVx
rO13yqTte2gnaLOk8qdJOSGQE6bX4jtGKrKwTGBFQZqcDmfaOyZ6fUkl8oHfuVxb
8QcQDgcJlFp8BtXbESfhTQDYEGv5H9VSjeXCe//kX54ReONNUTL3SAFkqN7M32gK
TNJ4SM/FcRm3buuGkfOtkW1L66sfhIVXAIu27T5uP0e2sOY99LVnS3IoCbu6tMs6
Uet+SaF8jUcx33xWNyJRuKrt9y5yFgvHMxX2/F/q25ylsp5M+KKffagEg8m+06iJ
I6QCfNI3Sii+JYv7QY1NLBldbOAI3A6fFsIE2t3LsrMMpNDe/Kyp2Y4uQag9Dl2y
Ww7QUiAoiHfnKTqbLFrdxyV0Dug9zjP6wcGPFMYpcOJgaZ++oO5PEniRU8LI2QHi
NYoZID5zAL+cJInZMekiUrLkOyQNomHk+GO4fYlnP8pRGNQT9+6ca+UFwM8/cwEi
xAYxpY82oHYRP781c+YU6pTvwObnKNa0YcoJsp8d2VBf696HnVt5hwwgIkJmS/T/
xzb8R97fjCFwpLfESew2NBRMeoh+hKYmqBsdxzhDBX5KlpLjbCfxUtKoocL6DQ0T
DKRixX6h3brBwgrjFEidjhFgO55cIVio6z1M2ouB/r+Yq7LYyzfUQHWyy6I0OQcT
EqdO5nDrH41WgrAKha17SN7LPOnjN1QTKDkwJMULRXE9K9KgphFYJtUMYCtbzT/A
P937ncZD2/pdUIPN0RVEjGn3Q4g9S78uVVKMpYv4EMUqBPSswCXDtQibHplU/b2X
ozB+jl578eORst1LhLqUVEg5uZEnJREoKv+Thfc4gQtHtY/LgMZCerbSUk01dVge
8pIY9V0qTjewwui1Ul2lq5aAmWnYIrD73VrtRDg0FYLZe5/PepluAXZhAgagOdJs
Rwl+h0GNqn6U6lKHcS4kBw95p5xxICb0UpPDtUzWD8TD+J2A39KFDSWOTQE4reLd
7dDN55yWc7Vjcmw/WJdKDQETs0eORJzU7g7fcEqJQIA37//aHYJj/p3+JimH03kX
pq8k/79eq/4nsZsZb+0BbFsYgL3qsulozCmC9a+rSQHwGVCAh4yLz/hIlkj1AzBU
b57hO55JIWYcOCqd3S6cLd4gJfDLrVqCfnz6ypwOY33EhKDM/EFkXQl+DIvuzmT9
Kq8BJs+2NO7OSlNw7GaSQHOhpvmdJKGLEKQBjhtX2p+v39WUexGTlQRbEmCS4zPZ
JUumKdhi4nKWrqTfZdGAzLzbyt2o9bts5fG7CH99Fay8QEy1vd7yoNLuJOKpfEEv
dN47WIlpxClOHiu+jD9jHkGUs4/APP9W+rnZoh/sri1Lm+9xiJYkGWd6cD7d8W6Q
vKP9FWuq8vcmcyoPiQltgWeR5TM1ivGdCP+i5KnXRtIh23RBq3hAHfPloOLJN6OV
cqBBIyDV4LgFrMtue4OvQ4uIMlfQcEOfoxiJbMPw0kdU0PB8qqMIAael/+WvE3k6
mqP2NM/umblq5D9gKT3fTrRPE0u5J8y4llSnB6Gf95WsVKHihzj4wuXnL0P/afXv
254t5H1Czb/aF4C0OeDnSUQ5ccvxbOyYThHTO6n1ip98nTD9lLkRhK6/LIHP/hqX
wiQYcSOgoAHW+/npGAU5z1H3fvyj5VJdYDrkxaPQJujILEJOYhJcfy9uU3F2P3vd
fZjJiIiN54djecD7k37jO131yempaJvV3B1Vpj6XMyhRnNu9xSm14Not4DWMorL5
BnR37doYsiOX74tHN5Ep7VynyQ53s/unCpH65SSyTv8awPBe40OjyghAlSsSlbIW
1rz71UTTMv6X7AC20JT7oSLSl3vXw1sS6HD96jaDQuILQBHjj1984/ygrPp0xKw6
H0Etbjab9YUdcu5o1MBs5Xgjb/TUIEyVo9zyeXyvSP9fkHtiHs9d44TV1SPSKNIg
NJUCM+Ax4OvLL4TWdnj//ovqwldYKzjY8LNNaUDaehydNaNE6mMRJQXzznabNc1z
RmS4eE/cu2fXvysqKCMTjkvaePvQ+iGbHz8pUcFz0bX/5ojuzHvq4TGkBiy/ECyp
kyY02vhjszDaoUiEeZHUUIigfiTzgVTCPFlEtMYUxxV0w2Bm6YL36DU43UBB85uE
KU5v2EGnGWidSgIsigQosmkB1xMjWH1+H/KXW5CBNWdsofOfF/vwXziwNRM6y2/U
XovTIlKfK5Kbs/f9AOh68qUgM1Qp1opczE63nCz4oeu9Y0/O0AtBAuggd27Ms6ig
wF39lVqDoUBo8qe8fdGDSfkzmvc18+M7PvdW7mVhYhDXz3AYv0NS7uzyv2uN7TYZ
Vz4zLA1727QrE9pMHbU1SMZViPrVVayf1HxovVCkOfxo/zr8Jed/hYI9W13TRKHz
YfaZs0DQEqNlko+8nchSDkhK5zZlrmb7ZGWy/umK3Y8=
`protect END_PROTECTED
