`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i6kJYeLk+NMJu+6o93ZM46YSPrXehXPLubpAN0DThKwfwO3ptcVN2tw1ounjvwFY
C6jL46eWKJm1CN4SGWhdGkV4NqH3LhItRb4pgRutnC8r/2hvMWjzRRn9+16fMb7B
WB2WwnRhJcI2R0DjS75+k7/lB9Z1wtDcOfD2MQft85V+tgpw84rAvFAE5KJQTipN
piC8eGePACTPz2p/Xhoha5kAH/yuLLyo4Ez8IL0AHTy1cc5w9RUVxZqI3avpVNMd
FspICPOH8FxWoO+E98c/i2KBVjNkR+dN2Ax1pIO3V5rLn1ktDyoP4k+4bWqXKtKw
cC8CuembvMPichoJjMf59OVBmMPGIxsN3sXChfM+aMkXqkH1JfboL1624fXqwvW2
qf03VvzI39uZnEkxucLYK7W5OJA3vB1aYu8XOW0VYVrcmattbw+jW/fhSrS92h63
awIEMo8Hj4Lcw8arDoGSsMdWcpBkiA547ng3JVBn6D3afT8YCoJ91dhquM0HHDXr
QI5f3LzKroxAtBXkyfUi/G83+ApsFrV63lfTb1Rp0ybsyq3hABQg+8H4txBwJWOU
v2tbyd01un2wtxZd9v+I08Qgx7L5nhpxaaXzQ9cnUZ0EVS78J8+6fh2gMEDIJLiC
EKeU0mDVGFzoCHlWa7NEpE4YL+bGVDWEeD98IptDrNE80WsAS8jUmRRWjz7fUSjL
VugKpr1HDc3el5r7JxdHUzvSiA1NRV7M0v0GPy3O2wOStnFu11ekoG5n06QVSu0J
hmnq5bTidHRwnHDhDMWCbMO3qxBkgHXahEGk8ycNAIK1HOeWnBqSNszTqD0S0/LO
HwoS9tiKK2Rpi6W/1oShMehHNCfuv2N3Cws2ZbJKpAOoGjkMuOT7CEuft8lkeEMS
ymRdSuhfEvEdfFS9u4YZ3+2S7opH8LZOd60zVCgEv26V2vr7mEBefTwysy5dGbaU
kjGlRxySiHks98roO5J2UDG4MJ4y7qyEvSCfIp3AG6NMKSSCD35wb8uxQJYUBqTI
nIurltCGVaqwRZc61npjhoqi3rM21iric1jM0VkjlWebuz5yAzM7cKzsFbrOynTm
sqzyyi6+Tz++kdVaEl8OXDiAK4+Kvt2pJWZAxBZrZPsjfctS8Quj89A9loZ9B/Pc
8K77INeQ5sntAtcJcFd3nOws/d83r462Ithhc2Ohcf441/59C7YG1frqXPFQv9cI
LShsM/ujnm2tt/KPW8oyc1HCfjW/RCEiSLzRvMAuFexLM4/5ua5c1SxS0MzjecGr
eAPY0rmyxIOPaFZD3jzBGk9lauIMJrYyzRjYbgFkX9Pv04PCeCj6Orqk5Re0QD/H
zFHHRoSLtvl3fTQpnPVJIyI5jfxpGzDiXQit3t2sx3bFev+jQMycsV0DdqfbXpTt
7prcWDT1nGrcRMM1zVePHzUlC0kVR5C1a4cB5Tcg9cAGGeRf9qWpOfX2Q2lS6yGg
NdYwC3/d21/opmRJA2X5MJ1M/VagPyvkWmkK/Ajp2cVze6ZD5bPK0GqZkk/V87jo
vnVlsdVfs5z76B1KgZc9O0GHQBHK4z79eZ/fS9pzPbH/UXL6jwJgqvaKz5DpzaOZ
FdfwTZOt+UVDp9Usj0IEUJmULKkkLRgnNgCyXjPRAbkmZ/8jP8CL4nPqAGL24SHJ
jnVjuwA0tiY31OMXfwn0t7h8Kz+fLjW26vNLuqLOBcrTinQiIaFNu4fdD0CYHIne
AUA2Y7H0Bp4ZT7Xd8WG1nfpBdtcyBrQNjO5M0eyf4HQW4RY499XAMz9HqYoD4YPl
M5VUgp9w9R+7rZ+rtgH+M2fQPd6HeCfqe/y8MNi7q2P1fvK6pYpBNuGA9Nkc6+/u
NzL6l5qwoSBT/H8j2q5mQcdmy1C2y0jgUZ4VHKx9dgORMCAlPhP3ppWPBCsdzmo6
WkfMu/4cu56CA7zl5PN5wez6FSuvwKvOPQwyOXL8Saj3s8jtCOagOA3UCkCUOs4y
WPoSf8kEemW+P4kBq4tRSwEoXShEKkEXuW7OWBwvLSuB9fLA3L5oB796jW7ayhQc
R3hLG6ciiqiFNOt2ObxnuNASsPy1/bjLvWLCpnro0NU4V5T2NI/YLA2PSJo3jDs8
DTT/Zd7LV5+waSMv7UTyrBbcd3HrOjy9GAUhOw8mCb1olkUOTsuw69qOsVNlb5su
AtTm6SVXBsf4Cxc9bzHrisJmei2bM/kW0bU9R/qmsgLcd9VEh5JXTXbDZIgMtVwT
7Mmc4Q6FJ+iM4DZDNf7AMGY309HqbByJr5kUQ0ufwO/cCuXGf5M659bG4o7wvjT4
OL4xOzw9GxitEro4ix4gbV5Xl0piZqZtNL9rB6xiWouCP2NX9s/GYKaBKgCYZHAx
aYkFjeIiGcCl17Fz8n6va67TyHtRoqu+ryMUcOGMWW/qfYSzlzOJS22/s5jkeKDs
x4NAlmZ4pRPBXeivKRuFouaWVpJ3hZHrv5pfScxxYL5xs3tg2HGmaBBRub30pJIs
kdIY1MwX/yC6WlmkKCJ5oqx1t3JORNI7pD8YuNxDlXaEQSz8zmevLU0gP/FSU8Cg
X95XZQ7K6nITvb+S8TRdcOvYZb1PBtmbw0bCDQSQkMbIZ6FB1SSgNHcNcM9tun7N
LdWdvILof/6gWp7SF7JNlbpGxa6JJSaQap+qC/IiTzzSTSeWvvpTN0QdyuMMpC85
rpXRiznhn/IXTwNaRWPcdPmR7/lXt22yrx5wo3x0vL0s558z9mDk5rW9VrkuEhEw
qqRZW/AeVaap9IPaIoD3zLH/dNbk/MKB+myCMhg1Jtg0oYrPbiWzTI6tFS7/q4KI
BQaxQ+jrhLrQgFfVuzPQRpxQjrx87jsTX7nD3A2I6gI8VhqO2Yh5w1OcZoReGhZg
CZRBfOeaXvCB/hXfkq7A0wiPQBtslcgqsdZ5ZPqyOLX511juAzEEgkfAz93la3j6
C2kfkBPjFB/POcaL1fMOPumC+iMi3KeKQStYds3/QzZhFgryCmixw3WrxPA39w/s
wDFPpCfl93D9LObATeJ6yNO4qARJg7z60rS2/iOMxeieSoF3sqMCczw1GsruvauS
zFBV94eDQ7tRAJdDgdwOvLNga/HGsRFK+byE75fUu6Eee77eld+bh7LUPnrLQBzU
/LTrF2Sc5BuLRIWDBvoiErVJgaxoba2wc8wZLiI4qvjV1Jhef274G99nCDTLuBHv
B4tch3F19hnG4eYtGmr2+jheFfxn5Gn5JzJbBwqTsq2qwKdgfL7UsPVMny8rYWEP
`protect END_PROTECTED
