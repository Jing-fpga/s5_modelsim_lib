`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9R+2PNG75oQY4sdywoZq9uzU3+qMqGtYiMZY33vQrHdFn/OoIslPqIuHCqjvZCRb
rS8RAlAcKYdPKQl8qGpb28VpHB7cceh6Omros76dvyC4xaQu2eZcv+bJ0JXnAq7p
WO6LCTzSbyBBMM3gsxERv3YOV1gWDiWQvn88uiZz3g00AfPdFaB0qFumX3hSSFqV
on4IIYBD4aC2whYy0ifZ5ZhxCZsPK6B/YZi35qStnXaci6pqywnJ3JXTj60bhnsI
QKYZsyL+MuMICWj4NS7bW47N/Pf8kqN6t3qkvMS9167919kU4JXxCXRMGBWP/jSi
jQe3LrqvV+Dd5qiY0s8b0kmErWE69/PoxXK9KMuqeFyYkn71JZH/He13Y6Uf+ZxX
uCMQd3v6IhPNu7tAWlVq6Sx1wsg96jcca38fNEpRXaZY1VbHfcKEg92+2mR1fXes
mVVF0JkoKQIvzpa1BJU+wFfRKvQMsXWAGgnJsG273kSoYDLAERExZj6JF8/kLf/l
N+j2ogliNJjIouNYds4cXYlDe2Q5itgG9ewvMaLjEIHP4m0tneq+4xf5voSr3GZ4
ZNhYrVxDQdD3XzjzWaK7Q+nuGzSJXCZrfpxPISOU/whe6YvGywI4Z0ozVOuNg1w/
r7fzSFurfhy/H92RQ+9giG69h4xhiZyGe+Z/NSueYbXat5cW1I6rUc9nzofKfTIv
KHzsEaR2XiRfJ5qMOy3uMhQzniDUo/Zp0VjJQTZ9jToMR2GGB8bztC2dikJan3k3
ySNU4TAKaZQnXKAH3OEa18l2FMZh1zp9GKkpKaM8eJM/pHjL6KWNUc2yWPh2u6HN
E84IUYVtqrs8AKNJqZIlytAEDSp6czpHNgtHaS6q8tm3HM2An4HPrnrTYQ/wD+CN
9bKmsXCMpTCbZfE+M1iUlZZeKAMDxzo45MRUcV5+YF312CVWEjKIFIBTB5VB7loL
POsgAieA1AAPY2aIFtPRBGbLX+A+F94AaaDrOAw8wk2Hz0805LzF8UTYnEZp40zB
2dcErP+Kuywgm1vLpztJx7AXYVvIvCLtq7lss9qAYmNFSt09jdtbphlEt0QhCD5f
cQVpkj5wCWeRzLJCQO6zgATXLlfVVhvxnn7Ua9s4MHi5DhwO/tcWKR+9EjeXC/zF
2dpQlISY7GxLl4ebfbutLs+A3LiRomduJvfmjISGnk58qArPDQoSowRB/fs+j8pP
GodRqtT08+gLNQxmFV5n2Ab4ISvvQGCMsyLRC4ldJ+XroKp55U1VhnOooZyXmf/5
P6o2dkhYMNzFnOt8jE84evJoIwIAprF1nRtC7pSZcPKlUgt6MyyXOax3Q/2hh97d
4geo8KS9nQXc0OYiMQjgsTfNXX9zNKFNCMtIxi0X5yR1ZS30CSVZlt7YslkLEvv3
K7SFCoa+tuDQDxT3VbYIDXVE7LovtePQl+fB5M05pcvMmSrJ25twTpvjyDlnKfjB
BohJOcH3F+Ah56w7GzACxJ3N2JuPmucXyjjXlFd1sOhn3QVjs6fwXzkO6sJ1uEQD
XNVPHQqDNm4wQgnKJtOsc23KZhXkg6KRbJRl9iVyHfOElv3xU+qMssLJZ/YGmkFu
`protect END_PROTECTED
