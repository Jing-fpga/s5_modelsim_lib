`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FUVkVe4GkO5UJtWLhzfCgcLtOqNb1zKqjLwGjsLIwlHPCt1Z8RPBL07sHeyn7qYP
OZA27gvAPDsV+9j0gi9b0HriGm4QQPgnOQsQ26lx+LPeW0fOnCQn3X2B87o349Md
IsvtvNDtoM/YXi0WxMduU98zNc4NaQhFlPMIFgaFjKPplfwGiD2L3qfP1AERxdE0
eqJ4FmbKJdNQzEzPbas3feDDHYWXl47o/s6+QUg625QahGNgVOfgj5EhlH82Pn3B
oXdtdgkfekl0Gj7+TedxZGX44crw0WLSQ7j3r4G6BQBbbjARM1OAxFcCM5R01q14
dIiKU9/+sZEr85VKwXaFZVIgfc89gFmhRcaCKwBh5cbC4Tx7emZdDjJU0nkrM4/U
GCqfZpuJ+oA1qN6z9YnLALe8tBkp7HYKSPFeEQ1tUmxyjW+l6JDTbFQhL+pHjRfd
tHOncEl/tkE97zu5N1RyTFFqEdsEoTqSiWCqn+MzDOJuFF4r1zPwg1to9Xq/S4Yc
LkpQBY8dx1yCrjnGQMuSgOJE+t7/hPH39iRumJs7CN+D9xoGRcWvKU2dzjbZ8HzD
zHxwv/Dp/6F3Kx+jD4h8SOkBRlEI1/0Zz2jfY/skSt7i+FdNLWBOQ56vJFm7+cXn
EmG8jtIxwKxuwYr4lD4/xs6Kw84eE/Z/GY2vMwGQHVpSpijLwEW1zrjfhw/zxHR7
uFl9cCzL1jtL3PwPMaPAsE+23fcRoLUOyx8vKOkQe6uHe/IvC4zpVwvQqM0zG0RQ
cRyg1eJmeWlg4QUOEPWBuPkhLPE0w3JdnzEcKv7gFA2h0wx3WoFC6wo8+CcA6wWi
WAAxHSk1caizsoe9H/Qase9Y7T4cN+Y329okPkPzIH2qB9eM+RrvSJJfYa48eA6j
4XWJeWjBc/dYxD1ViIU5TCDgnLL7c18/nhSE9JMFIt9toxLFIOdwdaErUHHuoHGB
We78UDCe4mjJmKHuYZTIzfhpc3k1EMwNnG1Wq/OFpsZdlCW10+YyLCdug/jDVBPE
Muu+ngn59MTdpLy8fdMxVtP9ETv3fDkEa99reIr5tFaHvAuuZHoTuBTTxvtdofTM
ggVDYRcT1lZquRA9KaIZt3VZqEWRbxz3++pnzzHnbvYO9LcuAuVhKsQez0ylHhyC
B3jsqzFQd+iLnrJ+A0OnBcPGxDHCQ2XDyolly3+ravsL3qZOQMVXMWNsQ20JTGS2
jB1xqhGzQKUPWz1Jjy0pqL/yDNfRWh48rM7tdBVBvpO7QnvQQfdynb6ffBNRggPh
vNDanYUiHZx8NULrQMO57ufhW5rYbsSGBZlPMM7hVggSU6UJzrpQr6wE8zTRC1ay
ZfqiOC9zeoxIt7JFLfPgTOm+QG5a9qTCtaAs+QRIqIzKifJZiBoWxX/9L3mYtyDO
1/bMPVcTkNYgbwuMx6hqA97YQdhgFzo3dvsftt3rL234mvkWEmp/FwTk09NzOtg8
jyf1yKKxzpRvsDxVdlFQvgigcrgXt+lXEm2jsKQ2jqvPAqcqw+/yRBhO6hy7Hw4M
yzIddUBz+4uisNiwgTVb1WvFUR5Wd2CD4xLYnrX1qCAJys+CcqX3LUwHkby4/csp
7qvd8dv+pruobKyYKS/jSjDOW1vkaSJdi7YeqZGofu+gHWr6HPES5GXNNRPpaks7
aAQHhhr71OuCsV0sjzFTHQkUP+Uhej/0pSs1lEXdMkwHZP96t6Yd47LOcs7d9OpH
7qByAefzQsYse9ukz4W6ng+4EXgviuNEAOoQ2Gp3xRnnlMg7j/Y6UX6v4YyXteqq
zLPoNrtKU5e4lDUHMUP42Dy2QIlTz3L5YVvi+T/U/JobJp6Tx3b9vTFmwx5Ib3e/
UNmyB7BcgpTYTIcS86hnrYOcJYvVgOqLEx4Gxja/J+GxcSIm30CuF9aSYmjdkCLt
u7KG5F2ozNdALEPOW9u/BD667gbw7ozK8IZYrNMFZFpyKsWBzOImzlm37DMeDKyw
TUlMv7i0vhCqwxBCgjoUcz2R1osJUd/M47un16nVkz+DsjuyVz3n07NnkO7P73hY
9Ay4r9Fkx1OWFjxfZkrCSOBDcgEnd02Wz7oJLdusLCnG9HmZHchAu7vnUMub7DqT
78rsHn9boaxtXXe5va9hLe+fEfZShAMO8ZsM8xaNo+VjdvksiFktmiBjv6LYM4nx
iIRDWbaA1Zo6kvcdTAFhGpo7fhI3YKOlXCjPq9XT6LuxEensKCYzzc3NzaBEuHZ3
R/g53YOFX4Z6NhgRLh/kh4e946fJFQAcUjsgsIcX2EvrZEDJ3VVynjTxYGmMxv/z
FfVoK9Pwf0STLXMrE40+j+Z9YAZq7IMeifqMXWNyUl7nA9jrw0yZN/yb4O1OaF8m
53mY0hnJZp1Tt0PYa8lDxz+2RZLN+UeDhXwFXpy/Xq2WkEWjz0QFsHXkkGqbWLWg
DDdJS/+pQRdtifmQvYuAeUo4stYfp4mLBj4OtZ81Yibb92CWAuvhlOv1jo9+rE3T
pkrhoDedSvg5S1cAuxDE3apIxKj7Zbs5YBzVx5PNE114Zlsnoa/6DwasXFS9kR40
jiBQ3GUus5qUzLlywVB7AghZ4qPWXu/H1j0KeWTFpKNh8zBtYqL/A3rqtc+xAF3p
YxgrGUAUpzcHX2j6AYdDbBKe39AdxQ7wXNG+Vb6EISG6y3Y4/DCy4/muLl0CQ1To
v8UKGNbWJ2+UK1h5wJqt6R6sSq2olE38I/9fsd8Y9UKkQAFPbK0Y1FR/qdIp5Qdb
jF8uXH8ss9JPCbKDez2ObYTY5b2QNVPXcmqVM7f0mwHSHLbl2VqNC5y+KvIzvPm7
K0HxKlufSca1PxgI85XWSuj22y5vHduGX5mZJAij9oVg33g5//0/EBQ+J6X8sPc+
ZXykBTq9ZzcWvFExkezp7jOv2AeAiYJObzOgSMOTXXbrqHNQGuA7rENoQ+Bp3Ngk
+YGxrMYi1LlX2OYDLIBsFJcpGL5zuFNrojW0ezcKwd/vi9WzVxUfC3RnBhKPmYjT
CprJf8vAv75QVZKoTtS1qJYbvikbPLFi/ZGPMsDI5vo6/jdWZvrGcqMjsE+qJSIV
JGwddDtBE6l0Z9kQZFbkzvRAcDcPYCO/sjOvLTokNuoRKDRe4qwK+DMDQ8KWOkVC
ZWjPz6kNZIt6CoqbK1JXcdjrjGSrDLY+uCEW7vTbhn4HlKHaBXhNe6uROxzGidxz
agAUuQtikngBMQWwzEmwzQJUSkH2D6w+RGFcfSr803M5eT7Pop8gCenbJiU7tLDR
xQ6fok5pU1e5XAHT2JdLdj6CKb2sS11G2II5L87CsbPmPtC8o5ONfjmvtUDxLd8h
`protect END_PROTECTED
