`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wv8MlJ5mdj+JafjLd5WM6T8P6mSmfT9f1WffJRW9JQHP0jjmb84m53h17LbTppFU
schcOHAXQ5423ooYNQwoBKt8WZQTxOskDaImzSXjSkwrDBuUBLL8dV4E9J1DJBsA
xPjEAeWce9UReJ37gypCeXcP5xGUkaf85eel4fpok0b/AFATZaogI3lDhLwxecFD
kRiNYYhHSgTGPfrUBX6GXr4+wfKFk+ebz4x0IgZopZywR8xexeaeTUmaLjXigVBM
QutGlt/N9XdauJtAvopKBFz0h/PkR2SweJcFZONpbKr3KZX8Qg/ilH9Z5C3zXlud
O/wn42RKXt3GT5y6OeWuQp42GI47Y+SPhDIqu1jCorQ62KW7BkY3QD10vPfWFIoQ
KzTBE+kxo7Fi83smYAvSNAOPSrHLpdVV9A8dt8U8QY0q69m5OR4WH3u4L3+/2GxZ
2HjUHr6SwCWzUshbgZhhKN5KxlF/fisUoXnKn391t8wkFi3CAwBZE2KrNwomSACs
atKEzJvvsDF4efrE1xWGUv7QWZMP8fq7hFUKxZbvuLJhAPr5K4QK22qMxzvrv9ux
XTFO4oGYghPRG3+S6Uh0CPerHY5Kpj/oW/YnwYM8yZNOE2dkuiXB6VHSe8nAT67T
NszMdqKL50Yl6wAmISJryZzpZ2Wos4nce/A/2oggxae6EFlxew5vkS5VbAASeQ38
JGdpWPEOlitDIL9UR8xttqpGQ5Ggc5ZxumzzyyCl0mAMhApIgLxVmSu4dLxG9EoB
9v48g+auT8tz6dsyVCySzGh41klnMTnF6UGF8R/Itmf1SRl/DtZX6Nj7QMeySH7Y
WlTG4iXzN3chAjAMhkdMDSV6UGFj7DBny1ffZofRX9ynD+5J6f1caOcULUAVaq5K
agdrV5vA0SSR9vltkdHt1Ug1yvIRs/oGmOycwLqy3v5NB5SIH8d1opJBv4LBjeDK
bS0ivKNmAZxW+Ux3cmbRhfWQRnC0djz1HaNtpoBKVZgUhulMVA2LDDnUKezRUVU5
t8SZDFMlHvVr1+rkeydqWunql/FHBTP1QYJx3Sg+dAmCQGtLZNBDQoV1v3JdIPXk
Gl9tnQFzq5eqWz9kbFjEreNmhSxTHkLQps8DcDFK5lozYvawSu0i2O5kTwpdL7OA
nKXihezmWvWugQsWB/ikgUOMYJn+gnGohozSU6HJ4hweEabeNnQi2f84tTNVe30Y
mnsq7bKvhhdLdyslWn9HeINou/fA8hCvUw4pNykoQYvwaLE+sFNK7E4M/b900yLD
TA9+js+jivnI+xO2fqZqPS6u7T8vr/e40XC2mtsFEQ2WdVrkqlZC1kSgvWBAFNFD
jheKPQzSnYDKHkYOVTr+eARpIcF5vtCmWxMZclPoT07vhDZNZji8YTrsjgnrVMsF
QN4sjsmUAvQ6ezH7y0MmaAYKUosx557QiZlVg46qyZCZ8Bm1Ao/I73EeULX9c/8P
1Bm8QMgAi5QNmZfu3ch3GTqZw7h5C5HgDI6V5ObIdXq2gGs+GQOU4D2IoJY45gjf
bZIHRegQP2fDHIwnC9jDI70OmmABV5t/1cEf+/J+Zs8AA4nqKBMTFy28PeN8oohP
eVAtp91XIoVKsLcmcwccMg00gexfPoYyHrXBTnxgeHMSlh75tLwH6zWn0s415q82
g9Wn3PtRJ/Ej1ZGY+1RMVlHdx/rGvip2j+kV8ctONy5vggZsDtFQGcJPE7F09+l/
jPqbEexmvgfoy03kbi+X47Vc/LwpsTuHjy6Tr7iRIBMrPToE3XHl/T7KGXlvsGsE
wYzIRPd0fSBAb5viPmkLVu1y13iASbO6bSSC1eO0SeaDf8iFwFr0C2RGlFZ63YdN
DTI/Wb8lc82QAemqMipAAejcft0540AZqALilxDW/fOQr0iA328R7mrTXcXl3kcJ
ZUXU8qDg8nu5Sw/sNzDLuu5nlGkaJtN6b45qS2W92HJ2jBGoCsUYZT7NSKU2ogo8
vqU3PzGxInUNHdKJtTUEMsKjxtXL8Swj/dUfcBzTvgt1meNDBO05z57cAyBwiwZA
8vvthObJeJLLskk1A+q6XXe4AwcPaPxWIzQFPZ1gFi6cmhiXwkaA0B76tcLEg7vT
l7T3UyhVvVq93g/ABfQ0dbkoyE/Iq1F1CElnsNSkiAXMVH6frSyG9WDKrECKey5b
aBH8K7dJqrwZul+GfSWTZ/qDXhN8H4ciDkETBK6mwT3ebughzG7mXKnVodCH4yXR
a9ZrTGPSUDYsLXWCIEv0En4OjecZwCLKcJKKg/KsOG7ahZSjzIueC87/g2HXajqq
MJPxe+n4XjVzQBT0BMT+BcJ3hVU3KIVAM4LeEIeXcar+lVxMVpclKDWl+ew/UEh4
LdHmoU3eJwQQEgI+EH4JkLeSeNIzw1chGdcp8m4x15JqaXAUjXVvDqafrVEZZm6l
/Kcj/3cijxnReWJIf/mzMkyx9rdVIpmjTl46/SkZnCg8tl0f4aIGfFCljwASsg9Z
F3mt4uQJLeEaIvZ4Yk8ooUUZDxRs7j3YV7BMeGrgXICAVa+KDKxtZMRyPvWyG6Yi
bazsi08WhAHFO88ze/+nG4phgNwFQSnM19JmyP2KZcUKzYsw4w+llXxBqJJzEEmb
gZGmYW3f8RgbgEM6jwpUrESkaVFZDCmufIoNl4JJ1pdAvYPkZZpSHV4Blafpq4Xm
2hugHhiw04cby934+9KgiZTlAYwK31uEbzrA6EgbfIsxe1ZCn4lQ8JIEvrj1/IBz
oB8bI3PkC1vvdsjEPBfVrB7kea6+5nm0E2/hwTbmN9bFo2jNYK4eWZPI9/f1qezS
7Cjb8pKTs6nhwHQuedO8ZbMWT+TB/S+fmXZdv0UvkvZjOxCXw0pghNmwijb1NjfQ
gJJN1SaEfMjKddXHoV7QepGwKPZKNEnxiYni3pA/oUUzHy8kDSiX6I9uXb8Vgv2U
l6XYnv9Abw9E5IR3h7KuXzIIEjvn90kkw6/rH6WJQbpACpF5gUOmIbVKMD0EH67G
MEySvA3/teQpKzlSK1x3bceSbugUAVSQjcbiUNsi7UBWGRM59qbe3VlC92BZDq+Q
NisSK2bf5RK8Qa38CjoMXjMyaFhkEP7WNKuctYuOwhHb17rLSOOuIKkUbtc2xeaQ
sRGsBhxqq/U/7Msy38CE4uP9pa3ZfmFrfC8Vr34cUx9Ns7r8sNs19gSUeL9t7U9/
Ii5lTTZ5vukBZdeILOoCvIgFElx060MMQFH0RxHdu39LLRnyiYMLC6gNApg2yvyN
wvErBEybGqpXL9Yx+K1vIrvuNCeeBSVDwxAilowE0v21uHM6VVw2MVacbl0ZbJQy
Y0SkyggkP6IMdcGd8ElKcaARixrsJq49rT3u/pHGb2CRRNzBmlBr8iI0Da6OxoPK
bxg7YHwSbZX7hIpvUHygb38MaF9Fs6/es8ICvKhwq8vKar9ZYfX0gy/PsKeAIA5w
hwSBlGhUDKHGrQw5OlToAvSLi5qhK3XBZLtzV2tPPSZsQ7PiwHrywAQuV3Gh1jNe
XXjLkL23YOrFWpDyO6V+6c4AgU88H0mMNhF4FWqrUzeeN6H/qgebOD/B1GNetWGs
QtpIeb8UNMXwcyOjBmWAvfMrtG8C6rDvFl3Dl40ZoGLL+h4yV4m8cDcxNQhTm6Kp
lYatjo7iGBSXVK2B+SuuoV+OBG9Ubz9qltdEPDqGQRyM4H+2AimXlQ2oYUEdoXHc
XOJQMsyvBUTXEwQ5pPu0UmGstn7NwuDhWPZEhwsq0QG330FQ8u9S7Llh/0VVPP+T
GgeQxTaSprQC8f2TpK0CwsQODAGkBl9OVR5hfJyyUSiQJKl4y9Y5ueEYuturAr9T
cLQzJOK4c7G6lsC6qSeZWJRGo4knuyVevaoxLMstfP/d5iV5qs4BV1j+VuGblvpV
W2u+k3S/O1MmU9uFRxGd6b/1N7idMwD8pSD78jTbCyjZHDCm9ltce1HG1c7e04Pa
pkWyGYTbEatFMtDZjJDJuBkKTvES2Q6vhfgfTTHyu1E9uG+ffOpY/K5kJwhHITgl
YrOJcNJJKxoTgjuh4eq/AITqmw9Lde3Id9PyK9bjKZE+Be9g+Iwb6u2ISoGgEM1c
zD5ZfRA3n2CP46pq7/twifyDMOu0jvm6eH8eOHG++gaoSfoiu5hS+Xm2/tOpy3kr
SzYkzIDdiTCCrloKHo4UXhlkGikzFc7BnPl6ghDaskDGKf78kMB415k7qiL3nRB9
7PZFSZRvS7Qo9v007Dm+0WELxCDBBbGn+ZTaa1h8IlHNysAV4kiPtWkkvfZmh8Ka
+4SBlG62azrDgzn/6GLHJ8icQEolL2pqeyIE8XuNgrPjVsjMrnnp+Z1XOiPQKJaa
69xkjyZ6gpdj0J9BkNIUOPOEtxjc+I/Jdd1bWpUfB8IM7qkz/0lmmfv/dGym+OwY
oiwXUTlrEF6GqMK2kWSFBjFBK4uOfOIXO6bSTX/OjCrQ9reyosoHHII0jUfhLtOZ
+Dhd9oDQe84vafaddcqq26JKqSLngASVhdLNi/vmNbpmd2MT4u1+8ARqJzNYzead
Zw6Ol3VVlXin+kSHtQsaB5npifilGrvpi3LAKncOmsQA+qXwvNNRKDu/OOmuT5es
TrmwbcnZ0uHTm3hxjPwU9YdC7v2HZlbHdoFwfOvkGY3ru5D0eq01vGhkll7tlr6I
xvwtAfwvi96cvOqXxKp/xRc41fOPEIXY5fCYkkYtgi0QcoUc2k9yhgGHK4LOQCo4
Z6g0Cfvq+qQ+X2hxZN/7e03nmlirJfWVulyCqvcN3TqKRaCh8HCi0Pt1fklFBc2J
DXjuUGMKNyMRkRSYPwx9Z/lXHilvAyI2Zq5HVbr2MUHx7OIKV1kxGP5eClNF6b8r
knjInhrzuXLu0TwlnriqcTZzoNnOkgnhEC6+Phni11ttDjq9qobzIwJGfhPXjScr
t7IOPsDNRoxWgfjng62hBnVz641/sjunLJSSvHz2wvr92ZQnmSUMjIhjGa/v8C0y
QR6cSI4daLKxozUtnqDaxrO3Zmj7BiddQXEegnyGMEEWbAfoxu4MP714GR4bnOUy
lFoUpuo4AnSF4ivGjwJW0uuwVzRFPEv10zzpsZR65dANNnJElt7lUsammTM7aX0X
Vo8bqqYMhbfd64ug2oUJV8W7oVaggv/UwrhjL67HVtSD+Mz2suoGlPSgPNaF+bSK
JKRYRnZGF+K/QxbWQrUNVTfpa3X6DqnWqsBe3IhOXL9xXmD3sVMhEpT/wqEip/TT
ONE6CE2DXIoECms0gM/ohy2RWJBkWEJuzNWeDFkhx/wj0oey0jJhJXIv0EOsMAHd
x+BSawbfRnauty/vMZTj5w4WN2+TTFGo47dMY96r3bizDRE5PjIUKanvgxfb2HSw
Sa5EjnLh0dOXIjvFEaQZpp9xnbTLc3s1FIofy+RnUuLJyO5WF1L6Cj9pTbW8pEHu
bjP31BaNz1OgNP02I2bt3YLCe6rB3Gikhlomx8/fdaTGcMm7ae9f7FA4RFlTrC8T
cghy3GupD4XWAOAbQqWuNVT3MW3IqValpi8TIUwKdaw46ihTKhuZH24OTG+17al3
ePHlofUgSY1e6J8FdUeBtqYeKR2K4r8vB4riS9BDuHgrN6kNqrBumjwzmU6eg4Dw
z6/Ps9AfY27kpi3XvT3BWT4oLyvOATyhPPCckNuyBmdjMwiYObcPAOHL+4xccb/c
q1QUiKhum+2ojlmH13F2jA==
`protect END_PROTECTED
