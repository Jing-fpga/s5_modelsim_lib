`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W2WSRuV5MXw7+Ps9aA80tC5VdRdysQhkgAfGJ/n00TljLop+GaS3htpq1FKvLJag
ZhID95NzmvBN7Jt/GE85/TnzSIfUH+FNuy5vmyonb1QUB+v6/ENdOoJbcXoPE53W
hErrqEqvIFOOAlRYELccNnLS3CSYWzMxXCmYfs98+YHvqFsn0HIm94HczILgrlYv
ys9axV804Ol0vD40vhspBeOv4PETZ+UnXu6TgLGobZHj7CAz2KKam3CXww1nlb3Q
uDWlW2VEijRIrLI3ECUROWis0EapDRTJHdEiyS7CzlwhAF9LsA/aGKvYEMKidyIy
j5I3HELddR5IhM+IN2QeNPnfLAqFvGvItBbcmqzwpOi3jGpxO+vxAMUqtvUJg2od
Cn+ahSb7yz6UpflpBrhyLwaOV/N2MSpz8GqZKRKwmzRjGiaAK7AbiRGd4AJM36vw
CuPI2BJr6W6YBjmXBOOfBdj5VY4sdp6DTkvJ43hvrLD5JiHG7z7G65lY4vUfnxlm
lONowREbnYbvZ7J2MOe1AHeKNykGmQ7Sw4r0MTkK4LK4QRSitq7NKWwzL3oCXY8B
hieZav2OPIbBzrwJBqgXctM9Mps77rGABSGwPE9QesLuoBv+jOAqVfB2tjYUtsdJ
`protect END_PROTECTED
