`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JohzjafN9jP1gIBHAYZehuPXbV4/RMyl8kHCihp7d76BT25YA7gSOG1OIVyGEbiS
nBmR0+wFT3EpMZjmetn8mMXpJUK47f+iDP8mbbK62LZG086M4Slh8/GDa8QBEVcI
CkKMaesjZd5n6xLy6C89Rv8B50XmQV9A8PhCoiDyNEPEJ8F9h77izyu+ivHkz7MD
NYRkFaKDXu9ZRpT3fJ5knLHODor31n0/S9Cv283RcBOJ1oTdn3C6C7x+loj0jEpn
2PXN4JQea8wD2KEU4g5Lre5lX+NWwqU5qQGgCiAcgE4+w9U3gpGdqn1JLn/PkpC6
J4xaetFw4XBHtCOi1NsEZWrJ6ZKOHX+ElWtA84Tb5mmpi9xKnmdtMJuB3IGR+7mn
vduRyeddJOoTUIdgeqzkjDw8A9b6cSGZ7ZR3YqSd+w+4S4i6qmMy6ZAwM7ut4PSD
6geJ+yMDuHahbFKfx4raUuG4mgIl3uOETZe0XNW8bUSGYp+OZwqwGB+XNwwG3qtv
bNjI+G6IEaSi1mjdktKnk9in4fvAQUWMtvSuE36HJFzOthPqvb+Rb3k7dWQGz6ZI
w8QpPurNFyK8Q89G8lZIqFKdjTzg80Gqz2M0wlwVHEA=
`protect END_PROTECTED
