`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tLjffU+o2VMCDgx8nEO1jRWmeaDMhMxNqWPp6Qy9D/MirK+a1v9uBV6tcbBMabB4
NNPbOC0XalMqBQQE7/6mzmF/Ga/ZOuLmzAZnvWfaKgb7ugndg6MncqKNCr4ELyWV
tzq5FLWEGIyG9VucABBaYPj/G6W7v8NJ/Li8mlUv5pZacmTux0icYjY7H/UxDCKG
Os2PxVsTBHeHcQMaPoZ4JywtJ0akS9JP3TO+7krUxxofwNMAnmgtQNj/gh7DWwHg
NIR4l8tCtRFvDw3eEBFFt36yIrpJB/6f3oxyifK7OazYhcu/FDcSAq4lRCFLWf5O
H55TOML02ZbCK8by/jgy8p4h7MbzTD6XQLUqUaXhJOw=
`protect END_PROTECTED
