`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tklsF1l8wo2wbNA0oQPKpwN2BkfLXKjglf+F6UFz5AjwYCNe1CXDowo1zDRpxknN
y9rG4svU+LKYJxOlKwa/68Mw0xc1P/404gt2FTQXYazEKfl0xYpxdt6gKK8M5cvi
akcX2VxewwQRzxWK2DQ7/yiWwBYaTYoFuw3TihyduhCg6aN9oK9OSnspdfhTcfn2
Ijx0Pj/kifAu8vOd3i2UWPwvej0UKLVKPSlD+pILFvEUXoRRSd7HrqctuZkkjAKQ
N+9ABP3qlMp6nlKdQmfk62aDEbMUvQZEBQJSrs7b5lxUpRY5+7aSQ38G/UQj36oQ
q7Ky5pHxuqw1JQwh3IfwOCHbbTOB7BPSUme19tuu2sOeDgG77dGF6h32K7puhGsP
tD+d5RVm+H20ClfMZxQC+Yh7nL98loYqHMmhZ1knYif6PJa3Cu4WkL4H232GDF1P
ESPHvQVI2FoAvvEyv6fEWEwZoymEGG6rp3NgCC+DZvY75sUvPZxOd3qYA454+vmJ
CikhCAyagOIPUY52J4uVT8bzjE+HLbWabXt6N0JGnR196ndGt4tHZvTMmsL77D4u
leHZbMg0UEpJ7iWFDxOLvBJhXSc+k5t12roqQk4UJWtglVk+wgEsVE4x3UVtwzyh
xKhsk/Jn5sZg7LVutZ/osA7v3hhmqsUUhtqV6qUmz6aNv+fyjojClCcewPmc2ohi
CddL0GeCbjvMBGW8tH94In7DzPctu8J+LlObEWYuDYRWtRd+yKYBdbkECy1F98bT
b2B+l7frNjatKyC9toGEVI54me8kNRpsRS+ilubpAKT01QZaoivEc+UvysbA6wqJ
1UL56aPDK5npVq67jNQBc+WIAv3mQ9sGt8ka0btL6mEBxymjtglusyQunVRr6UOY
f0icWqCZiYnE0bjT3+u/hZOBkt2veeIQjQznB1LdAAgDk5WDsMF+Xma29fu9crLm
+a5Y9XR/3ol6yuFzSYMC5RhYltr/8Zw1xXaOL+k8kn13r0tTys0aoJBQNFX4NxnO
g61GIEhDBvqsZighXINS6ObPBp9e/mLtL8DkPswCVlQuwiwp/KXGm35mf9xScD4Z
shYJXzfGWQb7AQXz7NDvFiCX4xOF6vLX0i9+yD7SBvxALHDLkNxinAwB9TFbx+Hf
edS5Ov8RRH0joKKNH3ztfbadvN4IppGE7u5XLViHUmjnZxAZHhmnfR5WJb2takEG
YrE73ifuW8URMWibHidLJL4NkR1riDa0acVblRA18vrEIWo09ABoEQA/zI0u5b7o
GSCobYTtDRtBbc7TLxFG405XnLRVIg2Wd/VIIv/lRZY7ApRrTGoIGo+UZi7vvJAF
kHQ7hQ1yDFqGp5jZskloBEcCJHHu/g2KIQjIAnc92Q10Ft2at11+xu6JImzy7iH+
A2RO1pnwctyZz6ivznDhNqzW68UUbDX8rXNgFmaOk66FppGfx+nRujyxH3iEAIHu
vbvBmC1/JQh/Bt97yO+Rt2aVRKPE8HrXtkewUNa49Fq3vDV9eqAz7nloSiXCK7V5
Q8B6iLUOF+ytOewKFiIOW+BLLSZhtA8u1bEZOfgbmvP/t9HOMpWZg5qy/l/cPLKr
ywWI2+ngSMwnkGIqGw2foM9YrI9pN+8CQMwS/uvONqnjiYbd5iD8cvTuC7Ngu2+V
U13/UGJXVyjkFhI3t2CuPFLspqinSQPOtaouqDVAexnFbsTJAtZCg2tNx6pf9pS0
fPAzmKmLcjWo4PDCXqd00+3pgoujJnw4389zJm7YdgR4Tr1ElN70Yp7or2C+QsKQ
bIE6WRFwgPX3kVKdFqFil606VpPJq4Y5KXH3fYV/XHESuhUw3mov95bOTbhXsYZ/
LrtRZeG/dSu5yRgnmAbYb1uJPPF/aeU0gMYRgjV4wcwsVAMp9ARGThCMhkTvXPXH
c7GjRDvuTs5C4KKjS76pv+vTnJeiennxy5daOS7AvF/C5iAlnqNBjQK56hh8uzfc
WGV649xNPmd/Jo3a49aJNWMQUDzDEnS3NqtomTtNyN9smJnLMygFdrRnYf+elWWS
4SJigJimsf5hXMD6mjc4c11IZGfS4BhCiYitppnVQ3wGuRxNucjOGGu03NVtKRUu
dH6z88gPN6OqN4zSyLRJGl12NXNNMHkzeOGd/5AH0ljY26o1oltYz7gJCREuj0bs
tledVZgXwEbARhdImbJyv1BV2TRDHON4ZE/Yk2D4dJRsrg5XL5M1cX7/x0MikVlZ
0uOW8+0Ga62zel7qVLje/3NqUQLgqHusUhtnun1duFkir6cU3rDoWAC5GPZL1/5A
9WRl4Ck9Y6OE50hOAIQPpy5+nmd2iEpqqamrNDe6o9fbe+5RsAa0D55qrIiXtYll
NZAvh6laFqBMpa1CjqjqFwaxNJxCOvRMRdBYV89tyTivWpFnVNmm99weOaDSUhex
OgUD3pcNqQE3AyNjIRRz+psCtt1brkyr0nL66b+47nhsgieTOjB31J+8jXRTMHMl
mL57PJJ95dOgzskqVP6z+yK2Vh7aPWBZKzMAR9vFiZ7+U2wrgw1y19H3ERHsfO4l
r3DBI4S9NgSHlF4VImydKJXHMxKqMDVee34dL8EBh2NR5jp49Wu45RFpK7pSiNF4
7++G1Cyuh+wEPpFqrxOwMFkM2+II8T8qsxrOa6mdO7kQlhAukMD2JdnvwzwF/8Wz
i0OHWNgP23pdtxNaOYLbHHz9x8KF7CBgBNRDLiU4NvImM+7Ul7LO3dBu5KnUU0TO
RZasxEz/C4pQ37e3R0y0G/njHtDOMx6eBthNj+8FlvwS6qslpzmT4ikCWQETXFmk
Xbtuyqn8W39q5qydZXQNHsY/k6omSEKWXBQ1/4D1OU+N15kj0J4wGsgjXn7bv/D9
RD2DfcpkDpG1HO91NYotjTKQSLobMnL4UM5L6Y9OzpzkseX2zxzmiy1rh8LD9ndx
8aeQCy0wvVNWr3v7bdBAp5fbhYMRZmaR9qaRKrYtyFg9Ou4n9eSoshf+r7MkBH+f
qk41RZbMfeCDFXRMbkNTMB/9we+9nsmpWmJ4Z7aGM9oj8PlKq7Kz5TR58BHGu9Em
p1tOn3PsaiduR+NIjcKJFF1/IE68O72HoKZJvq2PW5bQ1EmYfw4puxdknycFVRXJ
pr6jYlkygWaoycVJlmZeHdsLCifODUOup1n8vU9XCTyLi2tUAmNoolhuKeqvdze5
jSJM9bU71CIOUr1vELfu+dctvgVjKjUw7PBH0HW24Rn9BxlnaPlbefDcGRIY/LcV
aiei4N63nIoioxbQwuubclN13voMkHfE/pqKQDrWFb8ws7yz+zZ/DT71lOA2Bp9u
WEDHaKVu69l+gjKYHLMr14I9+6Bo6xCYX4h6YbvrppERXr0eMP9AQKCLzhidcOWx
F6rdeawK20vklnfgU3dbJXDrtRwKq6T9he7eNo6GBJk=
`protect END_PROTECTED
