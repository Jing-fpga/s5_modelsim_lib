`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YEJwzUceq9UH070NXUDJ8kLldIW1i23RBnwiqm6xvPHXUF5nNg1R6fBe11TWyJJp
FrS0MzJyztW/b7jFtbSBjrjLGUNJI2awW0GdzDFLuaXp5fkw+1M0BWCT6MUso+/Y
3edT3rwOTCt+vCwmtbvVYNV5UzLsln9KDei136Bp7CrfyMmizmKXyCMLYPPeECT1
E+uSlrFiVow/sZ9nYVSOZ4OliaE+gFrR6eu/sTIWNuvgM7dAhrjLHGBA6k1uD9Zj
WSCN/Jz8qcs0Oi/4qtsrq3kYEM/tpEuuc30xoFYzJLjSvmxC33uG4W+Hiizv/IrJ
EdkNKmEFVWT79eqSwfaMeeHVgNzfn1bIOvMOiwe8GW4Z8lj9XbzVhrWkc+xn1yxm
bfVyKtXF/sM6bRH/54Pw8cvyPeYCcaOo2MxudFrA4lvMAij9cgfaiCjIAuem/Bkq
lm384UFtPDUuk1+ncSNTLHlD/xtwGSGE8NR4hz9RM65cLm+erFi2evEeM+WFcWfG
h0HRVNNVtA2s+4G9E7+0p78X+bGX/+LIgxUgLLVdLth2SXQNgkXjiAGoHQFcAb4C
IB0uLbPjswDwKFyl2IGmwVe/ksbk82sSAmysIfuEYzIi0dH1cwiwEIkQy96/c2dM
t0c7lUpP1ot9HgOSOO821eswo+5sLb5G/bW/abShUSxtuY3G/5Aoj94whHv96hyv
3LMSO2LaIl+KcZOu1jIlX7GWFtcs4JF1Jr8b5PGE9A+hZEXCe+jECRnc8XdPXbed
tlLwdRI7FFvKOHignBhCJaI7peehPodVtiMn7Qa8xlS4p2B5yyHChmXneqnPMOTd
oYMAJ66sQd1CMy1Kml+8YHSZj7SwQopBuqSMJkOGQuurUWKI9JRQy2OZadaOzv66
dn/H1+OKkPQAJQwVm5ueo+4TPPG5BbkQ/h5CWYsV7uLIN0UYAF43eBA5kiVlLNuv
NcDddYunhb13FgS6RzF15hi9MH1+xX+BLBQN+ofgx4ooa6LfvN96D3lKX75/hTBX
CHhJadvY+cJifaX7xGY7Uk7M6UqV9r/NSp0K6ghyNumDaGwFpo6YnsMUZfP9xC6y
MDKZ/hNpsjE0RjpfRH+8+Fw/6pMNrOAMfI0FbCcTIpXYx2Gd96OZY9RsPsfyCXhV
8IBcYvnQXxguevRq2COagGCEr9ejZJeWN/29O/oM9xaq2WQYSZDJgjx9coj77GJW
m0+482oRvbllCHOKTKljlhEmzHxEG3qFtT7cU+eToqn4wTv0JoNyS4vWBd+7NnOc
t5elMIz2C3Z9YHaEiNoZ+rTsdk9ld7u5AQo6jfyKauM5lg2BrPeux+pPgCIOGc4R
ug5HoGWmOL8d2SDSXrM+Zo55QZcn+29KMH37jlejztU8bH9Tg93FUP+wMLVWeJ7N
6v2PE2dzS6aY0SG9RDHA0D5fSHpNX7P8CQotDxeq/FMsX3E01/gmVOxeW6NrPhM1
tE0tjl5JfELtQXRhuqSXmSsQ31e8epI+169jYP77XFlM87UdwlaHMkLDByQKXhtv
8ayKTaLxCgaDVp+4Lnmm8iTF+NLu3bw+bnE72j6ZDNCAhqku3wNL62Z9+pIdWt4N
0bFui705krek3uPX/YVdbV/P3He5zsfs1btOXpvlbmsz/GnIoLSJSdnbZ+ktanUn
QwTfOGS4Yl0sWgR0HvY/q1h/5yZf6sl1h9qiYrdCNAP9Gp9EySvUriOi3TmplMjM
MtqNy3pXoDoACDxhqECgEWbjCc7+YrPfjzuQ7sO4NuSxl7UDT0jyMV7ebUGb4ZtW
6sthxfJBriuNxA5temQI9fuP/5RMY/FYCsUU0nhPd9op2v9rdoneOHgzyQiG5rZB
377uqeoD8daHR/SNnCEeHKrB6xgtA644CZU2W7xESDEY7MHGBor93bpykve6K9hY
RTndiCx7MUGcH1Mh+OBjdIVRnEaY5+CReN5jGIQoOtW4XX5Tg661x3ySAHuSZj/D
VJcEW2M1nuHnTwckAYu2h5gvpUUYzdlz9REntwkzFWQsmZZKOpIKU0KbEa/L84uu
9d2sZvYCYmcbj4XKIsrgkU8piHhXjrlhmdE2QAVKjtL/39R9/Pbcjg8tPLcLPt2v
iXntP82Q81m60yXlBPLeg4Msw5MXOLfvF5KeiOaKW5cqKZ1Te9Do5P5UWotcEsyw
6TIiWCAu9+CyT2gTl0Eoa67cPNvBC1tEpWd9dOwt9yNih6XcV/68CEhHUKdtd6bi
s4rpl5mrAzc7rVN1mc/U6M4IbVVv7p1UzA+kn4Pv4T5k4xnYDkKCAJGhUAlMZHNt
GaZf15BYfP0xwgnqhpS2/AZ1bfgesdwYEgJdNAF5sUJ6+mFYWe9ejReEiQSTpJWv
5ZHu5z068diam/vl10VQ7w/2nso7vGqcQ3+Xlmv3u++Aqo9BYEZGv+uAmlJS04Up
gq2n5884aichQmQWhMmMoJ+IfKdab1ULq059FQrHjeF+cI1tnpAfuQoI9szi9Olx
2tCjzGRtCgTqEqfnbJfITuZgtqs+1bQrYwEi8bPbbFs4F+1ooFmRP5iOQoys5u4j
GkGzBsOHXSKz6tMmAtq1yWAvfY1g0kTzVkqKsL3RmwGEmD1bDQy7UJGhD0q0EtYi
pzlNVEDVyezXDPvUmV5NUPpawcAld3z0+4gXZTr4qRatcy+ywK8f7OTVR2BI8G18
XmPfGc4GI/fN1uhGV5cM5J14ekHvrp08F2MowPmjlSQT8NoMM/o59LghIPbh/+Ct
iC4FBkKTC+mL1e2iX75MTJO2bxYNyzfs9lOi/g9Wt9bMT1Rzsq56KrcmNCsVoj+i
guJ7cu2B3OgJkihkJrBU6UH57wwCD4C3/GbVpd1xry8W/EP9jeZtnYl0E+bQkta7
kDoUzcqNDnUCYemXhEEvoluYUMKg9f6mA36Bf3LAYVnJCee05tRLYeD+cI6LuQZ4
8CIV0SeRes6WINUgMhbNlKvwFv9hj7jR8cY+fjLd3PyOGAkEfANV+0BA8cNoF7GR
q+2vY15HpAEIwMJpHwB9asox8hgmB7Nlw3ygX2mO58nXMzW8TZGtJxgl6jF90fsn
mQ4ElkC/4bELssD6rMhdEmmpoGm6sRzUn15C9ze/fAsBymtrk5wdMo/XwLQXWczK
2oHalvZjqvWHMVaNhwfUcPYjYz/AdVlmAh+vYUJjTjtFlsFl48zhBCmg2u/AjmrQ
HRDs26NPair0Z3Pv+zR9PawOjVr8oIcOpaQmbUNOh3PS6y3XxA8D2Tg8A4Uz8z7Z
9JptbSJ4QFTPbwMyqOHwfnIhdUAcy1Ruc8xoqSZH9WCtTZHgoy+h6bsao/JtAiDQ
V4g6/SqvN8VIJhWAU3FXXQ1mybAIoguste4hs64SVgT6v5ebn9zp0hLEMqsYgcjK
2AOuDVt4JxCHQnqbVya7yU7N4iOXXKqsqDovmWPkmKMODgT10a+FgMg1fdBpzvs9
CBDPxOsm5A1PWQ4eIH4SyTIgYpZmSVvOulYnohfDKSXmKA/Lj3eC6gRWa/UIqvbS
QCZtS6qeX694hfBEg7Ahd72V+DyrmBy0FtmitGCgBfhBsUec3+rGijn+L2bHj2yo
W6WbN3YLLhKJONhSJKjhPj8pwttMWDle61IgkYB1Pv69F+AkP89eF9p88nSNsJYf
n030GtfoQGwlQop8w/X4RyNJMRgKACLP1bNQyF7gls82ZWYK4DslF63IA8hT0bVY
lFti+PBvH7ilZpGh/o/hI6AdeyN7KiBRBqFT8iDRykqZvggKrJkbMk6lCb8hawqD
5i0dCVjvWIae5050PXZGTx0D4Vst3D5ZRcamA6wLAyzcDjQlleLT/BqVqxQ885G2
X/5dITymST52IKyhOBnIQc8kgvJJwMx2f/WAIuRHYFmxbixUo7E+3crczE1nDsos
ifUqPcSYDrfLwy8UH+F/v0EGQ9z/BtECfPjfg1rg+ojHhnVrELDSC6rOFeZ/hx3n
2lSrMpcOHOMwxYQ/UAPHTHr9lkVeebBGFPdCBMVxbHcg4ck1fnUMrZwF7s3UMQQL
APNMPMcxgzV74ZmIjf0PPt5jNt1QRVeSFbqz3Dybby0gTQHx3hN3qixIfMiKvuvO
CUD1bFc4ZMzjUNOjh0u1wHS1wdomFzmbswdhdXjYsIvv/W/j4AKjvzEVceVg8x1C
JldThsL/r3jSBv1GpjHoENRYt2RyaJBn35nz/shP1e+IPrWB8UU6C3qSkIZuw9fl
z4x8yEbN5qz9RBm/j8qfdwfClwZcgFHAKHrJwnaz1EhZhjuVsfhbFkmInMgBtklG
/si0bHk4Z6wX7CE4VGMyplXZYMDrTCyrNmeydU52TiqANqwhKFltPSBh5+VLG72C
ZcRoAwr2/4xNd17yjZrREqaFGrhZJM/wYfOLozHmIb5wZA0En9CJ83Zi175S+Vi1
lKXGtTbh0PIicfkwDNzN10lFOeGI3wXkOyEIN9eZh1/ktaF4lpfiO81YJaUemSTN
4XsUKE8lRLV7SgaDgyWMAChpDxs3pde5vd3z2mDyQJ0mOt1dmnNbacpuulGNr7lc
qJA6lCmLL6UOeq4ciuNaCnkeJ2GItH0d6Em9U19DNe1LZe95De2MwFMP893RjxHl
u69YNSM6vEcpUCENl+F5b34GUMeTin+o0yc7G5VUdl6EDWiRsAm9aII+RHvLBofT
/c9SjSnCy3vmJEk4kHGqHEoWbjZcE1u6/gORdiqdqz7KSrSETZfZyfpypTnRFURz
bCzqJOzOdNbOqxjfw5O+/y7XdgE5+V4o+o2mtOcPh0bSXUmvDjWM124GDumN35L9
hA+uzrFG4EgFQRpxgWNInyff3ka6AxszKs8IbCMNmYfn52DBvaWY/4WjshMReRNo
DPYL4o9qcoQQpPGwKEMLDYCtc+WVksr5E0QzKgQYVAzTtXPMJfMSNtyoByOaS/L6
P9Q+pWGmlNla0vnrpgkAWSNR1UPo4LP7mGYIQBRLxBMEG7Ia0JGZNoWkCqRpPo3c
aD1PpoJB8RCXM/eReJOtJbmFdV8QNmU8N3jb+lsy7Gf5EXju3tSDI9G6NNFV5mUd
oornCE/PfE5355CYaTZXSRdPoMQcXwPZ3KVQ0Yp6y5q26KJNmr3LIDwsQd8VDFHO
qTgr4zeWvmRPqsBm9taOTqRAtUqDRg1TY4Llof1udtErQhPgOUAvzfvkrOBBkMmd
4X1BaGuw+jmsqjrR6+vQ6BMUIaiQ3kNfRABZhJfIj43Yh9LEXWmhOLARDmRDC7VE
OT8Qev6XUBEZB4hZKe0yqG9nUcQJJZ5N2yKIpZK7UF/FJIPCLu4eZRXKSZzE/4bv
4x4ezxG5z4rdBZ6Je7jF8uATNfvjJhwFsZTRVaZqSBXWznw3IjtapZwJkgSiLv/k
Dtk81Fa7k+XmvJG32vabtB8Ip3uKTdHVCABMPPI1xEC58Ygto1KW52ChbFkUIccs
eAtrjfqAg3RHILHdoqsXKWXEiuwhsuJYqchHPl+ZODgqNK7JC6VLq8yTn5TIJ3RU
waDKBV3CP6EyBPSO2iw0N1ebAuVG95cFQ5VQjjXZOoZ8NVmvIo3mq4NnV+edlIDc
hRmDmM+NOO/I6ZOd1ACJRJFWh4B7DGQ6sUasC9PtJYrmTRncom8Gr2MWBFDJ4aA+
47d4TnmVsVjBA/14pYC3k6O0/yfAynFe3bmLdzU1ePWFnzjVMKkUD+/nPZr61FCu
2aITGjvFQTb7U3RA/rp0lqn+WxITENUvVCwPO0HGRCTkeDzWOY4F+D6ta4w4RePQ
DWI3ZqbNyS9FPbxkPFYGXLy63fwZxwg2PZkx/PYl26qSf9NbnMR/fXakkRFN5CPT
ErMt2otpEQkTGkmnyY8MQAby97vNboSNke9dSYq9M8kCOSseMYoAz+Ya3p8J9x8/
bWgjK8tSVxIl0ab9CGmqtBkox577JiuN+oDfXxjXTt38NvFCwBy/pR4EFDh1GW1z
P52mzNKgY360KvUtpJKpc9uWVwCyVD/WsbFbizXjBwQU5yitmDZdezEJcXfqWu7V
lFatZleJ5w42HJnDMuTxh2EgRPDM2kfAJbMd1dcwzvv+ZzUunXYrtDJIiUXLoFkx
3Q9iz+BpR90GLHGarBFD4zwmjwzVxuginCiuL5k7Ezh870TPcDLx8y7pvMje8CD9
glcPqg+vw5iGh4hnbUYOgawSOCo1SeG5e03iE8kie+Q8a0t1a0W6RKKxTTVXpDai
6ZKyo2CwDKh5KSu8sHJXlcul62Ba2HWJvvjHbQKs8dr7Aagn658FFwMLHTwK+9eD
804rBI64LRFAAWaRuIuaIqYv3g5L3muuKjNK+JvioW/gl9S22wR7Qs/tJIQTEZHz
waKgraO0suAyufI1ojmUfEIl0W3895i5SM10swiuItbQNQDjtoSDlC0GlbZQ9b3Y
B6BSiO+dD+67yH3ra8KDknrM1lyQPdrjauL+gnhr7QESEzmINXz5XsLAYcRC3wZz
bDd3u6yEsdp7J/DOh4j34X3ZeGdDZ9OaKwz1HvPsOr9gT4wg0Ua01FTolu7puhUM
i/r5Ye2bUi2nmuKG2UTM5sjoXiVpg4DsufTkR162H/7zsQLhG//iBQR2gj5/M8zH
8YgSe4eHsI+0MF3VadAcZ65TdMzrRrvKOL2iC1gvt+xQaRrm2YEgDwAud8gkYWwK
kAJ5R0vq957AfVjn/MK+DrhkZxt+DqRs5drKiJWUz1eM2Cb+yH3FHZLV3ilBHaPV
e6qOAvrGittBcLekxyX+bwIDOW8MlPR5VOGZH7HbzvK0/qXFWLPFSVE7t010eUy2
g8aRPcLKzUOlf8pkKIaUy17kDaY1rR6pXjX3rVwYL0XASOLu6LqenG8kiWx09WHf
0A9wWWFa9yf1ds31Ifm/alHeRF46+3fWKH3HD96vBUH6a9zXZelmYHa93q5GZacl
7RqtDd3vnFg2sdJKDKf3LXsL+OeLr1odhDkQ3QcAqOS5S2JYppuMm6Wwrnl7JFE0
XYyb9Ib+vkbfPInS/hFtLDi2Uk13sHUX2NaJArB/Wj7UmOxxoVnVv2Bqr1XQvxcy
m9NbmxV5ArMhX3MEhg+CpEkKFOTTO8kUXvZuBP0013x+NcOBaO+Jqyny/3EJOWPO
vIdlCCejwLEGVepzbVU3C3qh7ce3D1m9aQ77foZ2bjkmnmq99iuBz2+BHrR1YPiM
XZVhzGQTUtoZnyPbZk60A2nYwyAl2iuyWAJ0tBMyIyQ6XpHauYOy8/F4P0OM555w
zMReHZ9jvBp9W8gkEREnta/EEpNTmZf5sfywoduoa4Q9MPysNmZuQT95mCjt4tj9
JC+RYjTFRReH+j9g+pA35aI3hpKyolFKwg6Q5r2vsKa33EWDEk0JGCJKWy7VpshE
9EEUX+gnEp0ASDh3F7QZ+68eSh6T/+LBpG2Ud2hcbq/qrFxm4zXhYqAGTL7V4XiU
gvmYxdtRBfiOz7RYTRes64vG2or7k8/OpmpoSnFCz0ujuxTd5mGha5tk2VhMbazN
Bm8kUclyn+K9VyTLt8+IZtBdFw2CCilLfzSbvdT12/+U1ZI79zEv7y0SwT43Uny5
335wChQC8PdlW/he6tfW4Pb/wO8n+I7fkT1SDGy/k6+9pyO7zuwOqFyvTjSl56oZ
rBvUz81S1IfiUpHDXlvUuf1qlGcN02G4Igm/n6B+gNMSfmp3Z2iGZUwL63BIyxb3
FFlHp6jtJpaXAU51Stu9F2KrVW+OgQCWiuS+6duU1LFAXB08XYWBTBRcsI8+OISO
WLptfbKxeVYGfR2ilulnWLGMmGYBP+Id6shiShr2vvN7ZADFBd2iJNSAV6dVCB9v
5aGi2hy80U7VE1D71fNGtC5E2oOt+R8nBk/XNfjaRR4LpnpQ5iVwSODjanc4sZU6
En4WV4mOkSvb6p5L0+mFj4RQP6eeS80rhBRJzibG54oZIAQtWBHv7Pz+PQd8Tb90
8KF7Jk1P0FOS1OM2w6DxifB0Epzdqw/5mvUAd4A+0frSlhyeQIQXG6CcBNHIj1vE
G5sx9b5TsGFXt5i9QTTt2Qad6OqklLJKhZEIjPq3MGb4D+GjBMMjUiyBivgVoWD1
hdSSLQF4BP+0rgITBSzs2eYCT7CSz1kgkGIOy5KLZ6AnGBL0kOyNey0+gaFNKnKN
8Hha87MF1zC8ldhCC9pjADbyDYaeeuk3a75w4kMb/AUS7XcPbDqp3XQ4qSFP/RTU
WKJOwUzYUUrxRNzd3OWgEEuAUZ3E2r2npKWwLHrT/9PyMVzHTIDksljj4Cp9A97L
x3nKmh+9knUWp8tiX0/0paDrpnYZWyYWEo+ndMwvj69I+IWk3n5ApU9/BTBpL4Xb
tT/Z4Wy63xMWDBJWgDCDLc12dfAFC0Lv2TkTguUi3KqBQu5nf36+SGrZcGaGBS0E
Yf8PmFeDwAsZ5/aPeGkzf6KgVlnc0vkgR4NfZWWduljjjqLJft1H3TgfFMH+Bswy
9BAFMmg1gkY/2Xn3dFVvBaKT9Oa6vRQJUII48J7gmEal05sSygrv8Mgg0tQmx3O8
9CtE3dZw+uCgt8E2vMGqkcHoIcuN4VaAlGu6lywLSNbNQPrW9MIdud8E1wMIjiIh
D1ZdfM5lvuE05a/CwOIoJVUmt3X6EBeXhD77atAu6NyMCM0GVWRRpSN4v/PmfAcY
HA98ujUMIFwRkeWWgfUYR57hCrBvVGsVWgXr/ioup3Wt0NTdpUuPb88tliGuyFum
Bz/ubUtRxhvqaJYxkgj6FpXaJakuyDe8vku6C8AsJtfK00oP+LOGyq1hQlK3C9Ce
XRpBlrNQ4ZHt+bHLwmPWQmOOSLHeQ0L5Drl5FrH1ZQSzKDWZF0AF2jLeeVzYzpkp
MTWr7Oov2ToNK1ucNwv9ShkwUh/AVuYdwL4XCWv9WDmzLrv1FRfHa8PUXsKHwPMS
ilUss7JkPpHqDO19LHTNbVOrnGUnMhH1y6WixSNZigjHHvg0A0h0raT+9QUK6Crw
BVHwk414gb7FN6kMKQShr7gOy32CnXuxCV8n1Ct3RmyVw8PWFq9rtcAaaDzjD29h
/8ZoFATu4sERDhgWMAJkBzFFOvW3s/KiPDLBkShhjDv7OVA84VQEQw0HLLVSPCcq
C5Zm66XyHdtiuhLCfkkGwcEwvBicv5Oi1L9nVR/WkD53tK6CIlgwYhXLnlXDUz9H
bXMWZ89eO7kH24n+wK/0Da0Xq5/y+QmGPsmmln1sUu4oYiOqY9kq1uwBTe+2gqX2
1tUflh8gkI7ptYV13aDKvnxefAsUviStMq+BZfqRdKo4Kt28Ff9QE6T+8DhIKKXX
Q1BICkPdpX0hnPIwdpIE/Lf+vVwAVmXGelfk0uY9nfnE2tp/Rvk5BQP2f9yycfs3
ZKimAYBtdn55uG835sSfhg5gQeeqnG7uOIPu+eI80qN6ga8M4z+4fZRZ/+PplqeL
DCOUm1qFSruhbhC9MzD6uIm/8T9x6bTQb7wUbPyzROJgHlFGhCrfFpocYJcZoHXh
kGMVEO4k8FF/piDhJvSWNq1eD+bo//vq4cyaeXPAW4k4+2M/aqPW1IUln9qWRTnf
dLXxq9vSlR6R0r34hCIMnkaKNF/RA73Te7UCBzXvXiVGNu7EAKGwUwOB/8Snlt3V
ygzILB3fWuTgzu1G4hot5zZyIDoa4kK8XLuKbNYsgM2FFt3podi+myAli5NhdDJZ
b30G41H5UgeiHLQz7uD1A3XW8gCaAJdZNRLn4lcRDw70PH49+9TK94VB+167C6jd
PSPNIc5NQmepGe6c3Q7QQJRvYC3NVtw81s78sLolcrGgC2PSruM9HSYsuIHFwM+u
UBqpe9Ie7nwFJlR0b91/9ubzkyq5LHL3waRh+bg9e9/whKKGUdjLZjslQVoKzJrc
eyNir9msv2KFbbuP1fq8aaui8ly3ZKxrBvxHJ71YZXrrUsHbC+yB01JJj5TB98UW
reqofmE7/HnOppjorp2yE097w4+GBV8dcTkAlmsf4j3/1j6hSVwzDYSFgLmpWehE
tK1MyCn9zuAKF44jVWIb7cR1Z1MGTU4C49QNNCVfuAD5YZt1dzzNkUS6ykSMPaRt
ouL8oBrGpsj/AanotCbnrUdTvfV0+aqXfa1AEjYW1VqLBMzEXLGVZYjCMSbfUfe3
tfYpLuKAHU7WIYdLtkCEg4NIPvJD972zrbkxAI/A7lYUHO794ANjBLjoflAblmo0
f9f8AoQQTj0B1KO0zOSRDVlKkfpK0XMxhxxKxY3hPJrEoBsM2GeiDTFjCTf3FFiP
yTLIgXPnUlMgT61BUt3qKmnMz+6TQHwngPqaBquyTMv6T3GfokJxrm4aFtRbEKU5
llH1MCjyFADJh54tnJSl5x6S/wdms49EidWpPlZfvVjW7p7FY6s8uVNjxELFl6sN
dztP9mhVlVXPqcPjYsFyMH0aldJj2z4kngpokzVm5ZpEjFZFVHzFRQ2T09ZZ0htU
ESJmSf0mq0jsu6dE/UZY+PVWkLkVyV/YG3q+/vTwdruNorgVcHQ/qeSSi4DFNn7n
Et1YDGYqnK3cu0Fv5fjrtgsf3ZM9+n4GvO2E9M4iY7nZ7Yeo4Yw5A167NiuEguJY
E64yOveX1K8GcatLcjnofvVBr9AMngK7V3szGZqAqKXIowLCjfgErxhidBnTM6uK
LLiP5FTXBsXW1JtR/kfMXZ55GcTflnnBRj9CZVVf1zLrOGgkSxLktecmmHXBE45k
CJaBAy7UcGszR3U/CiOXF7eZrXjjmt4wrFHbx7ubxENfi2YgrHmKwScSwSFkgBzp
BRX91W/F0agQDjTFbt+9APmy8itruh2s9APtBLv+4cmb05FWuJkUZ+jawv2CAajz
oLsa61UpM+clHZI99WfKSSo5epsF35+hN9kjn93hq4wvBQJkTeDKlq841rLxiw9x
Y65ZAqRIzLozX77FPHT1E8VastuC0b83B8N5wKUGfE0DHh2pGQ5IiypBu/iTjgKJ
RHChXCwFmHyNi7HAaKnIMpDQiXZpqPTT31DcKc1MpOyv+1D8EY/GzviKW5ekUaFT
cH8sNMlappknUAAHspRBGD/l55UgtooBUyZdqwBX9fbWnCAVaK21lUtTIdHjgmpu
XR6wf14C+gG0ULiP0YjqbdqWy7DV8Rb4h5gyaPciOpiZirUifHhL1FCwkbWeI1kY
UOG25U/LcXIhoJKhbBD+fAtIXWwsHNYU5MCdHaydFYL2JlZ1pqtZmIsp/orpDKt7
tMhnV7bW9KGctBJI5DQZ22B+r0tMhV6AoambdidreBBd+JyrJ1X9pSpD1EsCWJlC
gb6IPmfuP2RCI2NoHkhzF03FT8nfT1DTUGfX6NceTgQHlV0fGCvvXA7secoTSxLl
rd2NNNkIwM++mBkjenxtjHJIoW+jC97IUO75ThFRfmW/IzK7PRSRHu532pZSY3jI
WQOfcHkUOY4gn966WBroU2GI0moK6et0mnWabqr877TSKRe7b3Fs2BFC2L14v00x
hp8rBNkuspG1sJ3gAamx9w9rru0xdxQ5FTWvBlqR9Lf/Qvg8WlZSLdnzPgdFGwxW
cPk5H4Y1LXRcxeqmrAhiU/GIFUsBU17li5uTuaRJn6Cw9AFMI64ntXHEAA5ML/Ad
mlNv7sTBJUKhND35Jwr6rC4R+kKz+c3Pub+1+Q7t1MDRCN4RkC3u5cTT7HrQnwtW
zpSBZkLALDSSh+aaldXOWwADEDvmWE+jlmO/WP7CuiHJWLsqGK6iu0pmgQSdFLxd
Y1WRTfWEYpEXKx8buMPnqn+sdWJ3M5JdudFy9O90S7yys3BgQvJBv04tDVpArkJG
b1DMGPp9WfvNohL227//q0b3COf23YAyASMgs3sELqBNX7yosCtIW32DN+TrNEN/
xCzw9zjXY+Kg9VmAtAeDtFv+C7dJlrF2kfq0ViMQqq660FbWNZTS00ZfmV277wmG
N+5bX6VHJ/db3WBaQ+vwTd+1JWpF8AEkf3PM0iPZU3Z4D61/y7tn11zykGRs6EgW
DBu0BTDO+j/kUB0sOjFO4jiXsmceYymeB1d1mj5u6OyPGwd97N6A2m4T+WY/kHl3
1SCfnxllAqF/e6Q2QxcLdyNKALQp3fXoErakxQzmBa4tfeNQ1dmuI5Fwmm7bt6td
prKTRNa/qB7oCZaodpcx/BEgzhyQldMITQGqmE3Pbf1gmiL+gQ7mxqYQFQdfB94W
xQp/uB3mtnwDws0yTvfiO1VjyFsIavwH2E8ORZa9lwPbtrW1yv6QEjkxVUbYwxfc
1P3P6DDMuWCT7jyGMHPYoHvfWZoj+ZbCFbzzsMW1/B6rh6AAFHGRP/O1BzZ3Cu13
532c4ZLsG7tYZH4Bl4KAIHLFQfGzvzjekOZjcBwwi3qFNY6jPd85mY/adG7xEatq
/FwKXPV5MEK7ngK5O40vdfUnDMdjrBDNZNbxElSf2fdzpAAeB0PdLH8fPBqSbkKk
Z2jEcOjS0UlMfPiM2yX0UBrfl9lS/MePJyuKOoPY//9YN+M5YH5SCG7UCsuYY9co
daSeaOoNe9o3HF5hlT5Kfxrl0i6ZZyt7f5l+Pv8kslu0obEWZfEh0was+xWQfltW
O8XOl34Sl8d7fLtNHHngIETZf+PgYgKsxYWyKxOuqCrA8d03Iey3KNT4BCoQBWil
O67XUsIqeI3LgG7eQUXLIFXDfHB77EjvMzC2FsrdPCVYAwALDI4sfJuYIIH4QfNB
6qVZ88dazHpXjjnPyiMwdqOITFzYhNwN5ciDB+CLDLuRmanE58cCzTUziOqg1ffI
OjXTNt+/DkJn/KVbpKG/4JmBWZrFVH/ecQf1vR61JGMNJOPEgPeFnDnVFccDSMs8
nvFzUPhk0rJhEXFrR6LEIF9Q5+Qp2tE6aAjvrGmsC1I/doQMkOvvx4EHAvX87V3b
q6PyvgZGzHxTWdYV6aGQfKgEUISvbhgbtHyomB9eeeorWDmJqXB2uZ6qch8YJY0l
ugybuayORBcmrbZv/O9X+Oqji49jYL+a8QxSoLaYnVqG+4/Wj6OSIXTvbjAZcyLs
imDoJVbNtfNPvDJ7qZf0BgxYtP2lGmO4iaJafhND6mtif+TW9bwlrd1lJtunBDUu
GK5Qp1e2LqeiGRRyqlNbj3cWvNZLhHJ0Ehc5PbC6XClaOtD4xXmisHIXPk8qf+Eo
Ugg7eM0YpJmu2k/s4OxN6ZwYlXWiHvsy1EkgnFs8YrUcB210roevAOi8retv1YyZ
0BzDX6oDuHlZFgqcUp54TMaQ3pYDswPp89ofOv0B+XdLaV/Am9QiVpSfGyO5T0Bd
hj3q1Bl8Sbb9D59ZpprKeA4sJ8HbmvI/Turwo7wpjfJxFKjJCl0m1chaKq+yS6Wh
J6dRnLPywDLWNdWcNss4r7g2uw2057oXO47ZaMSyR5xsCDvlOcHLye43iCZutnWv
jK1gAt5UDrzj4FffcQLv/Zve6SfNgQpr7578R+UGdw4nRi7Ov2f1wkXSo3g6uQYh
S8LDd3VVeeuJIKINbjp27O/uGzr0mo3Pyl1oVYCMzbeD/a7ye5AwqMkWWvu2F6Ht
G/Vrz+ccnlpICNoJ80o+qY1wPqP2W4/ZuaBIjPwvGlxPh8tY+xzABI81Oe6dG9Mu
dYhVv/ST0CAL8gu8HBErCPY45i7JsfOt//6ACqcZa9MLq7u+VstjAuPz19NqPNzd
U9YdbEM80KFaUFcIrXdQedThqXi0U/GMNBtzbDgsoKy4V+HFHFxNIIUd1/AXJzFt
FSMcLd4RkjbeaW313koRdEQDdwzY2Nv9d6tRE1Ko18gtpTB9H6IKmJSrc3f27qh4
Yk/CjYvwv5SPOV3TdOTUJ8i0z07fl1umP4rZEqqKRxm6YEJ+k8l/RrHsfvTX6gVU
W+8Gno55zNUUwM6ebqEjSvBzkRmbU3W/T7Xso91K8lsfNQDmTptLQjKCREALYfUf
e9OnS0lnM3vMoDjXuLdwjTQ6e5Ip2Pzml5USgkTd+A43yG4S1XTHsiVucoeXzbuA
AjkmoZJK+9F4rHu2GcdIZEfTDuwiGlafYIE7T36wumEAduk8H/AhrkQcozh17Zcz
17QlAz5wDyGUktk5ZYK/SO4ROKNG6GuQygVDFr9P7DBqHq5mhHYDxlFM+fisgGmD
qH+erSkhm/KWwRIvm/18vOnSU6ktU/aKjf3XprmrsxT0g9lZF+ZAT0VRbBlDThm0
dW7Jya/xwAEWN/jmdd+nGDUk/NtzkKRp+26zpyNWqFs=
`protect END_PROTECTED
