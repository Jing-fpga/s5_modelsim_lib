`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D4RMZQe9uO/fFX6nHDKqFIHkDjO3giF3FI7IXlh2rj0HY6oxw4UFgN7sUznzEDhP
CHwIlAdMom/OUNe8ZpUmHgddRkeCgwpgf/EB3D1P4PlyGrON/DjCBBp2FkhzAJUn
z9bfpGoq/DyPtcSSXeYZ0W7jED5ph6VXVEJUnTcK2s6NGlE8j+FRkqGxM+hCwZDX
pOH8MxRRriw8aHe0Oo+3U8DxJG18t9PlO/Cph/YNVkAOLsrhXpsVKuXB7sV0o892
J1gisY0yF+UVWNE7Pf50FevbLqfykVCjB9BnplA3dIqNuDpkY8lQ6WvmD0iewziI
TLqGCg4v7YNi4gUQ6lqA1Bg/XMvuDr19tXLjSUbxopUcpju7pN6UWk3qGhFvIFIO
4SK4GpGsOOhIMUQXcye0rP7D7rCtW2g00zXAN0gOhdBpufAnQP/n2rA01dkKrerl
0LElVDIyQXRkpXd8nCDGs10LaUXGS0vVT/mdSrPsJ3d8Yyx7iSSvg5UiwUKMBUOa
1cTMwDjo8+Nf71d6gwPvxJXLnVL0GpFSZub/2HyfUrEY8eBOOrdZEJKQmmILCPuo
1wLWJR0WlOu4A++UjvFZqAsDmU60FCThhKtDXFwAZZUH+CqKdRTohxrC4HuKhCaK
fuawlLKgKBga0gvkv+bXgV8t0tdXcjvTbUeI+yFct2XGagUS9dm1OnDc5lJYqUTd
kopJ8UbV3p3pIeGpjSKZ2cNm8VWdfQf70XhXhQYYPH6ZqHmem3ze9tvcDM7FtQow
kG7Oh0FIqHzLNRq37rClXXq71Fwtnzb3sHFlI8kgLitCaD2dT5utP3SH1FiFnKFG
lnw/VRydLJdfJuNm0/qaFtfFiwwxHD920TQyb5hxFrwza8R8LLb2Ik0HJwgE3WhB
aIq8BLlGaWOcFZC++oKPghsCWx4SGfwgly76WxhArslUClvDYpLeFOz0sPp/ttDj
ImO60uHpP8htmnhnO8NDnkCcxrDjJ8z89XGSIOjtzBliwEZKlvmlL2PlLhDx62e9
oW51v4dkUFX3p32bF0B31TNkbK/Y0OvdnRvjkL19TGj5FNs3C6kXlU1MsagLr8yk
crQSoWPKwG8CWPJB4hIeDlFrzY7hUcKUdUwFEuq3kVObzP26yRqzKX8/3BIW7Qwz
SwQj2A4KKNEJCRTdd7wzpBe5pXHruxm4QU2erGjUfjvny6G/OKJvlDDTiZOXUyLX
8FFAXJfP2LfNGLOjV3i9E1ktOB9LCQMSPM3thKYPMZOTweU4K3XburStX6YXFVly
8HzYMp8M8lgkcp1glnLTwFOJCwL6SbDh9+ljdbYinkVO40G3Vjb72Y1OyNOQhELN
dxGx3BMbTJ+0j5lVwRIQA1svwYa8EMu+gF0mYfeLDt4U0/cQXJL39sx6zcOx8G1W
HgeZLzaC1tk7LodFzYeyufxbJ8Td9JMR+46Uu2sotd0EkdiNoiJZv/h0VJ5UYex5
li+N1B/65XvwZXkC3lOItdLK2nwVAaUAI34a66M43EeDPpBNNOjoXd0kf7oWfX3u
7mYZTqdtldVIKXytH35zCtR/MisfufubvrhoQqNfZPpHKcRyLnFzzcKSgG4XRC30
a7YPBO+YtRmnB5eN8bHOcfiuqESnnTwNtIy4toEbXs2AHp0YDede/U/fv4+/c0c4
6+ftQ6tvU/bxaHe5MpjoFvbuyjudpB4K59bH47VtuCCfEibJ/vUqvtRdFerZ9WbL
BiNOF1Uu4nfYNvUqAb7ZwvWcd1ZsRJWxa7CPl/rQxLMr5MK1KJ9lwJpDpQYQOe1s
`protect END_PROTECTED
