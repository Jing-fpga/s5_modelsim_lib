`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZiGj9NbYQz3+nIuPhHqSyW8IlxVrZzMrPtvEK46rYJMeXgA6KnsISskS5Dcipra0
2wfsGBPM9z16U6iNjL6HKvBEFxyWDZozCta7cQBXdR6lN5sP7H0i1gVtKkjOjHit
FDYiy2BNMBNMRZdUJ+G6JboDKjiir+g+oQgNPeoCRXcgr54FiZLnm76gWXWtXZwu
2tB2lYjxlRQWAu2Zg98va5wW7vhtUKJ1yOBwRdNvQfdzQvJAW/9aLJFm8AQI1et1
766Qs62Mg/LrcmEfUnatFTtkOZki+aJ9UAI9iU26iEVVkg5ukkCJv6Lt20KIbfas
3HAiuwo8+mMeIOvUYvOoBqfeKulDS4vxO27IrSs33omjXLewAEv9O/hCiqtqLgFq
l8XnbRu/96bhaJSQH91oZP0MuloBOdfEAILAqyWTHVo09wV1BXTr90TM7CMISGk9
0xtHjS4Hj+5zGnhFMZV4/apM9f6HCa6SlkromrmF5kRzTi3OINqNro2fzOmFY+9G
KQN7wgSFRbGDNWQyxN5OYXAIZCA39YA7nJW7ygNOaijKhimV/4MGbWxZSg3c7zOn
Q2AqbfUHWUarHQMKaB/qgmc/UrcV/XjP0sHxTJlzP5P/gOV7jNKMHa2GAtmnR4z0
O/bzGBnJsPiXHl8IaYt6jtWfGGbKTR3mRwXYb2uD6pDHL7rHWhmINjTAxp/qmwd7
CtiWPXY5EHY1BL5QD4LFX3uy5wZ/mMgl9k0YgLn2lhhNjeC2RoRBBXX2+ggXf16v
TSNcEXPNTjb2oEcwZZ9ApKUx7KlGvTZJZ72KNZzjuyOZZaIjiKKzvSMwQSot1Cob
EvOxCOGpTPCnuXUIeWZX5SKL2WjgxzvBV9HPkMj4braqCbz5UGr+lqgIsmRHxB6x
Gfqv2zC2Ya7HSlAuwL/6WNb0cJFgDyUaG1nOX2hXDFa6LiYV+AU0kRRwzrWc22/6
+MZ3rW4GaWILOnRSiGjsUH3zKWUhpqrTl/nKpf46QSdp84mcPIBwpHUBLn3vKZoG
CeE7jPO/IdDw2Zi2mYV174bmJrn1mZkhMQWJqQZq7W+vxYZg9OTWepXmtdqvgnHA
0OXw0tJ/j6kE944Vr8pCUuJKKcf9gLFjSec19nmIpFvIlSN6jrFK+VlG+fEA1oMo
A5x38mU/vywJAi9Wjl7uORMjonm4ER8xYgAzyf8jMnWyu8hVl4jgNoGwNIdjSWiO
NuEq79wGjm6Pfpeo8lnTk1WTQcKYXd5sKgwFlXJ3RX0Lsy09NTmxoAwEQoQoBSKq
CtFN3Wl8I5AdD1bwv8wEOh3QFajJGMrRqJXOKGmc8OMY8FkxPfCUqqrSHItIzGn1
yhmAF77OPvrkoXGJ1YhQSIymqs1gYFUP4TmumxzPhXrFpiI56+hFQqZ+Lx5hWE6q
x0Imn6XyetrDqxaRaFLcrnj5YtPpMN+DX9cza2GoLX90UcqIk9KFOb18k6tC7k1+
dUiLrLa92pMUlx6b+DB2a2JCJWzJR6pjixdtMwKy2/OSDDcbfQ5rPuVicmDJDRp0
lL6wPgtpWUnQBd3umpF4gu8ZCMcnGLyg01/sdMxkE6N6u6T3Um2NBGOll0InzyfD
2iIlErWACh6PDoBI+wmWtJjGMLGPhRMY7H8kGRjHlUqRWUe+j5GbF0SIUBXGNWPb
JdjXJ5lYITSfMofCtrgNyprjmF+rFhbj4YRpJK9iiLeBhoY60E+h8fIorKgDeGtJ
OvSSEx5yeL8njIyHeP+iqrYBcrukf35j7NYtU3W6b/DRFDDBSSMYFkqm3BlYZ4Vu
`protect END_PROTECTED
