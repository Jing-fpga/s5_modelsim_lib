`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i3ChXUyvqtuayPHb4T4Q7m74jQzG00v9xcwS1XmWk29uruqOxPWBPV6lBcz4AhDa
dPvIxEQtIvSTW3qArDPOlo19RPZPwCl8GAI1LTJZIIvyZHdYXmFknv4Y/J2mUGpL
l1w2uyWVf9SfeEEQQIRUEVoKBXj8cLDgIJuGgaYL/FqWsBAqLZlNZtxcyEIzvrA4
YW2XFzIsd/mEVKmCZY3J1n7xknZSJB0I213hVAEhKWyUtyWz5EXCn+KMAMz7abG1
emnZ0KOI8ZR95SenLxulnRZ0XfWqMqODQjDbc0NqQeHTJraVEbUJDdTV5fS59/zg
kxgUqRGi6l+/LARgufoKkNHZTn9eOldNJojQwsG6DIE734czes9JPSXMouzIUlko
Q4Rrya9HVl1YfCWSY6U0n3q4bSkbtuow0nGYLISGavZW/psIgDZgaWs/2sVq4SrL
7NeSaSIJkPr+ia57ZL6mK9JixzOKgqdJHCM5RpJMURunJTyr9Hctoa6ay7cvhlFj
VEc8tRXNthYeBZu7wzBWtHYFIyF50atfSuFf1u6j9fCSjigXemOXU3SUFD0eVIwU
+A5B4ez5YYKfibwOIrus/lWIZY2geb2YKQ1WvEKnOZzcu3K/KRg3TVJelCprLs/n
+aJV67CgSQ8u2vTDE43PyB+Jt0eOKpkqg1UiN2uotM+IJcNBoLDpYSVHnR0gi2Je
AJaHYfAM58vahy/uq9MS0UhcLHLUO17bWbo7Siwfe6mCZHJwszvsmsMHqLBLaU4e
1FCqlY53VZ32GL7F1id+la/VHwl81jVjzLlcfoY/M3ZcEQS/7EPgDWo0N4GA4SKV
RRK/mdxeDmgoWjeZz5cuwTtb9x6r0P9EWADNpMHCQS/lrNZHTLgMcYTOoBVryaP5
dFBMJbN/8aM7hUOKvR5CPTPzsANTagt1kKOOaGCD1VfMtxgoZitdUnWWnHWFkIen
v0IPkKWul44Wpn/fNWF89H1AlS4LO5PmnPfDLEd/t1ORRbu3uqP8OlESkGA+YIf3
l7vjV2k5T9dPNKaMFOkCJZYfgxA/+HFZbRtvxzjKqfizBYnHgq9QMDKoZD0Dicq4
luIJsBjEZ6bhx7YB6dn2AhkDSO9nk+TZUPObznt1HjKtGM3VnQnN3do6c0ESte7T
oseAOD69yAr69P2idlk4hfAyK6SaCm1SQzcfDFvpNG34Rt9sbf+MRsznK2UawRNP
kRHl775sh0YZk4fKqD7bgoPJIJqAlVDPAIZ0mQw1PI83i4D4R7EaYkrB9+g/o76E
he5l9rQCZrv+LfxETiwx6MW07YaBX8yBvTWiwViX6gLcL5BDSFq5hcHKsU1EU5N/
zrJYhhRi2OnY162pBPUT1gkbjxyXJwpRSo10mELHOe7uwZeGR3y356A1KDE1XuMy
pDnBVQvbmcRA5J5cV2EmJ2BqclEcFuo0IJbsAUzZsBgW/z1TaBCWxan98HnR/wxD
2oF5oUK/9fx6aedaZoe+3trNPfMIeZ1ZXOBc4MYcvtI=
`protect END_PROTECTED
