`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iokkkef2J4KA9ODq5fPKvMsY0xCByE5HXLsrpbOC021NAZTa+IiIonUcxfIY2fxe
KL35XTggLEAjVcJEWgX9f1C1l7+GlYBXaR+8XaJ8RobQ+rHrKBWvja10+4xTvPSI
2lknoIwYOU71uv4rntoVCLSfajSC2a/PMy6UPyfjkz0fWcDICbxLF0oSUn0DraIH
iGOKLNFoQQRiP/hzcx+tKy2SRCZWHJuToB0yL37285BNiP4kWZbm8P45kxRIcjTc
bykN8nvoL3EbJPLqGsCRBnCImQ/ANvRE8speZAOoXS6BEsrR35CeduvYDDrNfe4b
/3X3QXYBQNyocEl2aVIaJnfEB4Or05rmtoIr/AsLmAGbcrZwJIPCMfTbsDXrGV0+
7dcWK5UHWWXIM2FTh7XAHDVlj5YrIuI3v/Xt7PrA+O2Gvcf0yUOxoO1X1QTPY9T3
tkAb5ijSzJdaE+pkWxaqexDPLOAV2rzhtAyKkFCfk81nOy2IBqVm9LKkGCOodLll
LoKe+aPD1xIPZ/UlW/99f3Qn/W2SUkQN9THiyJoqFkBSA6wN4qa5COfqAQQTdjfS
egEt5S6Upgb4Mp4rcJ1XWHf8Aq0r6zxqk7YI6E3lr0BvtimvCVBQjK5R4Z7f1Xcq
3vWxO8vs9/LJwj6E7xBEpm2aV/iFEUKsbGtkCIqGGask63v47IMqLssHXtYCiCm+
`protect END_PROTECTED
