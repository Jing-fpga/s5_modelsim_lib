`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mAlkhAl6NuQS2SQaD5QcBXXCLolL/2bR3+ZsEH47qNSrMCUGAR/dj85DbfJEp8rM
wJu6ft2tD+KAVlv4X6/0kBqG//zZenVnGxAgcQ1yPGaXbCdWPkuOkG7zS8RT2LkM
qnCPCeD4skGT/B0u8EGyS5Xg0t18cstsZRKwo5QwFq430egRLoTWV43wX/FdbPuo
QuAqCOHTYucxy90Hm7aGfdzRdCjRRMY2N+REE4QW7mENYKjXkjoNvtWyfsEPBFbq
vdhn0TnhSYI1q99OeqGMoTKIlEoX23MBPvagcxC6WblOs1yFORXgNqZHJ1+DoEU/
qYPTS/sh/0gr7X6Lxe4ax9f1hq9expL6z8SdIO565rc=
`protect END_PROTECTED
