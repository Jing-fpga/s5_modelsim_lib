`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WWSl0CVIiV1fUEof0PUzA3vE8RemgmHmg6aBkF+OKGeZFLHo6gqBzn8gvjXLompe
1swhnYzxC/lZ9KPo99rm0130IIscm33vLif5FxKTRQ4jhQDjNxVlvY1KmBHCK3Ed
1BDPfIIC4o+5C+Yxyimsnqq3rQZDDfW1tl3kaqyN3Dp2LVJHMFEluUeGaBvM4cG3
g1VWIuUGAKZGTi/tlLgqSSvKEVTazgp9lQXoHK31PO25vcAuN8+1nY9O6BOqKf5S
LlR2VatSnT8/m8YDK8PEiTdz+bnQkKPcDNvvCziM4owx9DNyMsvJ2mEc8Ucmk/Zr
q3ASMmCHfTcfgj+hVVcfb1NKZxUgZuupK2QqerB5PXWVbSnly5SJpQf9St2n7Ckx
w9D3u162Ru9VtzyhY42T+JuoiEX+BdcrKgUL06SBoj0eIt/VfCZTzO4Grnw9SWIX
gnlt7hcKmFvdobyZ8Mhu8BVoN2jY77qpIAhUhw2QBUrV/naYKUTmLkwO0cvPK06F
5tTr6hqNWLLb10G+hlZTbAo89eTNuVy24oF1FuIOtKf09Ep4h/XRtJKVMCP/SYeL
NdF6vx5VGFyo7E2kJIwjD+1/0KGr5gdRr0J4waIEKMVLTHePLdRqpqpoIK1i7Of0
WD//fXB/GE5DUC4cVWU7EjtjkX2E40MBaKvf7NdxISaBHnaYseGUUBNCtRfRS3iY
9vOZRktI6wQiDaA9nyCGTB1L6cBzCXqbLT6rrYGI1mBR58vGey2Nw2odbYSdrETw
4RQbz84/rfTuBmvZNKeLFGLqso6EUwrS+IVPYjTvKgSLevZx8E/Wd0U34qeeGljp
017qfSYWzaLqrPLlmGpPPmzRlluczyBz7dAmMluUbDUnJ1Sgp9Qm1sIwJQq6joQY
ycivcOz7aDf1ZPHqxIwXg7chTAJMZM1JHxF4xNQAHR+pXgJ4nVgJfIRQ8QdywtB3
LZCh2qj2JUfni4ioXB4nygkKiRqII51nwhECoyJzDBUuVqZYuPN+I+1v1PjMtna1
hB8m70eeKkym0UWHoZzVXc4fj5hBbriYcrxQ4hZoWibfCCsWc0pxDaDuTPrxSjnP
6H0eOiNz9SVbqO/3R4gNdY0zJcgkrKxeNe9NOWcGE40uE4vXqBwYtEiBzU+cm1Vg
RAU7odVsdhO1MaGdPsec1RU71GyK7bqapkNnOa3gya+BDNVx4lTUHxqJe3aDAPeb
a7Jgedfmg2Q8fcOTcA5qFRHg8CxIEO54KcF0345O/e5i+yqJorLrwydY7NrEa1i+
RdPslkop5eTiIilkUFqia/h9PobWrcH78BWpB/4gNXyxgKj3UmFHcbB8f9Z8xGT/
0GA2lV2uWHQar+klWskd8ODaAmc4cqd92UHg9TaA66lv47ugPgpwH67sscBXHTmw
nvmVqXBk7Tb1p+0LddsMTod1TUy26UmOPQkc3BHsLxtyUwKK8+ILbwGjAdv2AzUX
4EqbHgZQqyPtvEX2vnDFiPmhbv2trJmaCOmHwpjS6VebTYKm/9SDUR9A/f1ypOtx
DVE+xRdsMsAKXsf/7r7w+O9q6UEoQ1sbEkZAqYfECwYRHl/vQmQ3nQZOcxDAHJIZ
Pb0TsI1XpHzBr+9Uff34S1XtDFm4et8pVPW1thh5rcSLx3KY+uCOY94+QohLKo0N
ccBirUqOeszvK//+25ogNujvDm8SeoR71zY4VthQ4Iak5w1IUF7ya41S2CHCotYP
UXyKRWC1gqjEbKzxxgks+oFmhDjxTx/kWDkT3BDNpvchUlUKymJRqKbU96D2W77M
8GMCsNVzBhcTrnFDIlHe/YgQfs0Y7Nf67yRwQZ/ZZ1lDzY+VWAxHlB8RB9Qkfx2l
VcVtMfqhr4tvqTnaO3SjkqkGQK0VTWhOJDrmeR3VB0HUwJYwyepw+fHlxWLlaf1R
DTTq0FFet2QRay8H0FULDCfBMLCJ49mCVY4LcNSp9rfVPPb1pIyWqUs1SeoW6XjN
tRwyE86F/Of3cL0eSF/m6Wd/zRmhp3U1Xgx0hxEvNgo1QB58RrkwG9gGYqdI7+eP
zkDJX+g4axnqRSdS4iNAGQbY8SfPv25gHbiCgvh5MXHw+1qOqCYbci56hIfOHhV4
Qq5lbEK3U1dSWpbRNyLiqgS8pjrTA/cNzDuP20kH8XKWR57ItY9ZBAm9mWZOc6xE
hUwMWSCw9D5lBtEj1g/gARn28jPGKwFzI/XBBed1KTvoJHBZStUuPtiDFI3FVdeR
wZIjwnwY4yGmOZ9ptO+9aAW47gEkdvRbpNFJjJfywJGopWuhrSTtdHaTP01LRNMn
wfXpP3lEH0voGBeMXKSUm42szoDnRVuTAK72FdaYbhQ78Muq5GmeS3uzBu00bPXF
+indPUWtd/zNaOL0LMnRq+tc/2BZ6L3f3ZsM9oKRlIPU/kJSxnJ7WOVyCH1Dh+f1
xqNJkdca6nmsH5NtRr4p8KfD6yKvNr5ffCcJCbNz3qD4/B15CLUVbcUR/9+kiS1m
SNHAzz4fa7k3CKUEFN82yDCX84fRc2Q1HqWmJUd71HVWlms4UXh+H9bAFf4w4/T9
9DSfUtkdBg7U5HLIcqwOzPKl13RaleghQJGHj+LCCNKCV0YZJxTCDo1Q81MCXN7l
Sia60PgTGRAu1cqYn7670v0uVXiJYzJU3TV2+HhoB8gIPgHbELp2b8jjn86NvIHi
`protect END_PROTECTED
