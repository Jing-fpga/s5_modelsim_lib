`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fl5BU6xJlnpLsmt252UuzZ+y8u7RVI3pVdvR192PPm/1b121Z1ohtgR4RJI830f7
4eVd77H/O4xaM1aqxKq9Qv7Adr1GPDK03sgI0nY6xqtUzICVn6SgOsvbW5Xr/KPs
7+DygFXrObGch751BpXFueYAm7XsWNbbai0G2+HZlStipxov5G7mYTkqdWDPHuNu
KxFBpmdVWCEzRWi+bh2DQ6IQkCIuKIfwFO6PB1FTXBbwR9uxsaMrjvx/RpxwhZTK
qd5GxBus5lDc7P3oFQhTZ55SP9ZDUpaVmfiWcmiByj/Vr7Bg7Rrm3DCgMAy2rNcf
Awn+UITGrL5wDgDUYYhDWI/PlLYP/8oUwBaQi4KoTs7MDHTloH+MT+qFfL5wCzI6
8+rIagE4eUYcSM7cwWcPrwGCvUsUYDIHotHW0zAFPYJh2G08rXwPv0RC0wWhG7ee
lXZyHHn789QqsfoZMOSI0SExZEPnOzq85IURXZlKy/mjA5BoTUe4iFje+azTKjVR
k5rjK1hVyAX9YYCMYLzFkcHXwGUdUZQZs+5VbuUsx7xm3rbImrh8C3AwFCLTCjqt
+EF9RHOzlsfrwSAOrYrOZylUjXeIj7D9afaY+XuyBBFmr0lnzkvIcgVEjPTk/qh0
T82LbeXONH6daQMRl5drL6cX9zHfhWkTSG2cO6twJsS5l2RVXJDBAQXrp3ax+2zP
WKJeMKA/xBHCtz6uiIMx4szfbTkTiFe9oZIjjqR/jKDr/pblS7MkmJ0Ki+o3Mmsf
zr84zKmDuMD61zgkHaQvkSMj75CBm+L1xMqR5O5gvpGFbsYOMUxcrFLTBDzpx3Zg
k4f5poKlPpQiKZuiMA70qnOMNhfo+6dLqiPNMlZkw1PhzJO1Nu4Jls/ypagYnrJ9
9qYRmvZKUPR6mh0MgogqzlGQ4qPnZwk6efIUZJWOQS75dTLokLNkurTm6Or2Mqp7
/w9a8zJw5UZ+xa9JvmvTg3nD6JpVy6DynuXznl5aHOGx2+49usmMd8UUVQwpichM
JKMl1sGsHxL/JDUOFv/Q0083eEi4+CDrtTBNl0TQnqm7qsoDlL8UC4tI3WKiE+bS
lFaZ+rxkgEws1WvygqAkv7YyhWsZup4EOkXLBGH6Vegl3unRySN1Fmgrh5zyXA/X
dRTj2aIi7Y7YLFOCJ2cPaU7Trnxvod0pkXRwbuLSIMRdKeOPsrQhaI3DxkwDa1KN
fA5AaTCqYZAOqnE25sXqtyGIQhrNeapmAb7tKaKIfZe+VAaa03K6eyvFKUWkJcWL
2Mv+G2/8Q0oWhZhTSphEUtS/H6lwI/7MAGuZd8H4TEsAJii6N6bRO9ylXm2odMZv
XxHLUGsQVNb4VxEX/y54dHui80eEbT77BAAPf0wgx3vglww8vk0jRilZ1cDXOcFy
QdBFPiujQHV3Up9hYcggoO6KU/MPve4whCRqcLFOM+rlQ1zJ7+Ru7Jx43++9oaJH
+tytROZqOok2snJU3vw1S/YGoY0Otb6h/iZFuo8bPBS0sNUEvtkSN7toUuysg6hC
vrKvKR3ImftYZFheYMWwhrI7F0ABH/2O6n+GxjvAWFKVjTdiQL1HcaE7bqlkhngT
Y0Q1vAYrSXV1vu5QNpmck4WFJiNMIUTn3zABz3nkt8YfZ5pAJsfUOARUso2HnEcJ
LhuzT+29kR/sIiBAPm+meWyfvBAkW18SnzF3+6zkn23mGWJ5RR1nDDa0XJBqSSok
5rGrukSIvQCqBqRPk+328D1Fno0fOD8ncmBFQ/ucaiek0SPNnjnL/FmQEjuvust0
NvJqMUG8u6pmBhGUYD+dOsRKD+bLacZc08VYoDj07KPeUzMpnscGFbvIhlrsUp08
DNp3/e6P0BAPjLz3J5wK9A==
`protect END_PROTECTED
