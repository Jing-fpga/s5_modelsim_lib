`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vZgIUkhcFI4Ph/VvBQ99z5LKLp9ujVxbmDQxYibkNpW/y2OO7V+jlpzZeOYrEgEC
RXxO83Z2U7cXS5HmOFVnMRD1T3+LOCGH0MTyjlJCiTpLBC/RU5xYx1FltJwgDGIm
U1Zd1P3RBCBrXJs8umXg4Ci3blyVdfqT2l4aN2/6FX1rHMlNgYSuTRDE0DgwotGT
gg0pW0d4jIDUvofreQQuGCsG2YENgrwcloXEUwnpVk7sMK0tTXnvzceK6ap2DAkl
R5JOfTU/bMacosdMXy3P6xveS4Cuup1IfYBPN0lScnq4YCYjXCy90p/sgPlcu2Z4
icj1oeyx5fBrTfYcOsf+y9yxHlw19Q1BDoAgRWr7uvvUqaDEyH7zYbfru9POWJpa
Wut6SR3KEUVSKCEC2iHmSTBr9wsEaVYWBKAf0URSbM6s+qm21+drF6/tNbVZen1h
0txXd2Uz/LaogOfa2RXzqeONh1sWK6uEZB3e5OQbwn4h4jRdzl8Bl+Ve21c6GbWh
V/r2beLklBQtaKPC8Hm90ynLRJcyEXawun0qAxxKV27yOMQv9wdHLH4tkkmr/AFE
oki6bjQn+invxe6q9yCthV2d3AK/iCr6+KdRlvHYeMRFBhVWwP7xXYG+kmE7tR5T
07GUba475xUCoaGfDBvnUZKq1XImBz8xVQ8OpbGusLalobVkG0QvurSgRXat6H2j
8HIhge+53A1m4eD0jbkBcJ7MzF5JtOgG69CGTlyUlep4Ic8UrgwwutYgNWOj8C09
dn2jLTZxUV7NNeXrvlM0avcdfpTGOENPrmM9suhzK4vC0cVr62YWtBObS6ADsQk7
EUl2Yf+TFS/FuIjVI01rqB1wqMzvfK/4K2qj345ix3rR6C2RoI245FvbDwLd+L05
0k/E7XQKBSWbnGt68wXl5fQZM+LCKPGW44XX1ilZ330=
`protect END_PROTECTED
