`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
agIFFvdpQ+c/CJlWfqsloObER+2SPf6xWdA3XJBV2PQ0QPVjjz8ColPPEvUQ++cX
V4OJwagSOx7O1qLMBKM3dlGbOdCmohNJcQ7SPaeEWsrthR2kuoDtX2uOPHTVtHLm
81KePiw05++PcqfcZLIEB95qaKttslbhGO8DbFz3DYFEt77LLh9ZPexHfBKjDfeZ
5DCANmzAQ/fNkqiqy3bT7RH01jeLCPjie220S5CuPFiMq2anzvVy/YaLbNMo7qDY
T/AnSDOZLCn2GcjHHAgIFLdDTs7tyZzSUaSjupGGtoqLIsms/POm2eb1mYRhjvkG
/6Ews23LEgak4iAjfsYIAJMzZElNpMK9vTxUB5Xx/bmaBukUm32TiKHbdyCcZvpg
vB+JVjzRU1EEjk9dWAdHOjxABwn8SXqUA1iSl1qXgGm/5pekuMzUn0X4Co+P8FDI
f5BfUmq2686Hx8MhJVWk7ABiu/Q60pbxDMyj8O1zDrfWXH0wQgEHofFDETRRLeDv
E83lzGvsMGGzkVJqnr/6UhEfVlsCNYvwIer5K0eUGjn52VPlnId8m86gSt45BxSa
C+WHIh1ulQo+5SBzEMi6kBdW0op+74zu5a2mp2T8Q/UTXsyyS/zA2eaHhhIpwkgs
R6x7TT6oxhrsl5jPlsqDbUQ1lfbaEpRdXNqZuyRVxP7BjK39UsfegUcOT9pwzLfA
DiZzfgtE5HYqDCrd9tL0onomA5HbICMWZ4liBXyG+Le3yCS7HtSFF7SBtBX4wORw
GGIaKkF0sqUM4YvnFbiZGIL1sjad3tae0PFVYNnValF5suhNyKRARDLJqs4OG5oU
BzTXKhknWquLAfrNEIioPTLiKLeM7lQDycamGLLwelc8hau33UIBeM6C2DNSpzrb
/EQ5wUqKyW2RBJe0dh7I4a1/8y42CB4pPZNQRIOhR0XPS3R/gwTyCJCve60JnOYO
CFKKFEQrY5viCapJjXue3mKdCNn/hKm41nig7qJ6m+jirzccQU5WjxVESoF2I/9t
acU+WFqfyD9A6VJd4EtUgLEdxagmRkF2KtH9Q+FEXcyX14sxxN+acMNVZKubCMn2
Q+MAIC1sYI5GB5//Q9Y+krLsiG9wnub5f5oZmqOhZVYK7uJCIzXmW89xYN01Ob4E
KmjcordxI12M5BOkivzNV+zPrUejtJSwnrLYg3Wm5pvwXMoOPTwBMCS2fIK2MdXa
Mp7yu4YQ5CfexokHCoHoxujp3cSsTkabm834vnYR/GA0DBksbt4djsddNQAm9P93
j40znctBj0c/7Iz+KyRqw2nfvr6TMqn70OLkJhxjZlG7c1oqmp9VaHagxvp3ZtLa
EYvPKMQJGkwtRQNjP0xviq+khM1T6xqK7a1lrB9Ll80+3oJXJ4Q3p6Ed24QNA/bp
9PbVpC2wOjQY52Wf7bKwFaOBoXJqe23txak8XFgt+hrPy2enZD2bo6z1TaRHiQ5c
zQYHj+/PhHKeGFU5TAlMrA4NavRubizb+H5say4RRE3ZQtByFvTCFbScT3tDBOXC
1wvw3OuHT4LLF2O5kc5zukNaNUMwmkMfCpq7Fiqdh8JoOuIT5BzvwfSAj3J0RaeX
z+vUUkx4HTvLBt7cnTkIyNn1GchVjUK9R+NGxqwWuwp4pmHIDTp+ftno91ma+1Uj
GVzBT+Aa3v43KB+xI+M93em9oY+9wxXuBw42NHsZ0Mio02Mu8rjtdRwNiTWgqYZ8
ZrGMbVHf02dgT6US/cC1VkcShvc2MP09tcBtEgzK2PefCfRRZkP/BCa+j5ppkVIu
58JqmH4I+RZ8VXyA10lRsUzrMUyuJQrXOzDKIv5IxyofTM+dBbQQu4o8zm6gtzpp
pOAZUxIvEvIlwjX0i9+Hl997fsWNCkcA6yJg5CDBKsdGk24JVzFxHeCbsGoTt1Ek
7FTJne6BzfKAtKy98Mksye0CF+yLb92F0nltQgi3MVa2QxHIg2SZ2vLq3WMF2QBJ
bkb/vlwl2HU8s7uD5H+4wMUAwPDktCkRBOMgAVawsVS+KSb51vwxLPLG4U2ntuZK
Wy/YnYwDSdmeGx9l0/pUsuX4E2lB1K4B+RPJDjZbMYG8Y+ZlAngL52ovtq3yR171
DGCr/0SffoZ92v9cwdkd3npLNmSUZivGvQPPD2dtWBZMN3Bx9EMbm/9m8o6lSVKS
JSlo+aS8l2OqIaIxc3moChMy3wY05meLfswCfrE2wYKciXU0ddQCzTQjn9tYfdaD
+g+etHFMMqvTIryNUpVwCus9n7fq81ZH2a+lmE9Xo9aGVM/+zAJb0OLi8eZm8Kn9
EA17QncbZ9+vDT9Q3dKhZFPhKWnq+wsJ3aFLuIL7UiwNoaWlMlTkj04ITtfo4sQ6
9ceFIm/Z/BZIjj+/Zc5Z/t3Od0JUB9rLYbkv7emuAPq9vMawjUbysebLaPZPZz57
C/M7ysYSTuk113ZOXoLSrEFOLwuas/WP6MTfe+VoGrccThc1J8SrhefN+veYp4sp
90qsxL78sr9uIw0oQdBamP6Fuw4nc5zPRoLH/KdmG7dyPmvPoqqnYZDAHHk9CrKu
6g/Mo5DXJf3o+IMQo1t/9wdkNaAzfVgB+mO0Wez19ugvM0wRpnwX6jHtaBrrFeDK
yRZA9ReQ7+H2+rNDBf7koeJxxvqggyHA7LPBbUcfCB7au4jVqQkCIEhN5YJorlxP
yA6PbLhnaFkCmVP6XToTE0M6rMo2uEra8oFUY0yZjnq0ziksKMd8W09MUyD0Qme+
OrRwzf6xzrlWvCGnQcFaxSXfyYOdrRbozjOdyy0db7asfihfrIzzz2gV3y4wkCqa
n/DbZ2NXmezPpVioa0TIwwUUtLk2yP6vrtcTm26lIkYTMUBKQzLaL6txq2eMrAlr
Ub2aCMXjVbhSgM1XUvq5DmWT3P1U7ieeNLlNlWYDwQptN+WAdSWOSzj1t/1kDdE4
sPd2x+glPjGitw9KTRlEGWo4OQN29CZyy/uwN+EM0UI4bAdnEXJr96GE3qfSHs6W
7nSiPiz4cLaHMXA1ekZHJymd4AqrDY9IuxwxNlGZqKTBWmhWVC9fLfbzDFAvaP3a
YR8i2qA/Y76fytz5H1kbBW9+vwPbeHHKlSwRelKDhsFUrUTQiAs9k/dARd7mwNV6
Ioe+zILmT8GFgLrX2ORViiKdf9y9eItMwOHAuUYeir2X8UxutHtgODfpv0Eg9F4v
GpxWmNlCY0CxY46APDt9iulZ7sFUojJ7mZpHKNx1JRjKb7oN2jPnQaJHyznoR28q
ql7RtetSzzvNS0W2rKcbPOYubk5XQfQlXuQGLkE5uzQmi12kZmrNbSAn5/lQyQ7o
9Cl0tMd7klWQRPlpqaeciu6jRxrL+uh1Dnh5+un+BkbXBUaBJhvpRwo5bk6FZL9q
p+JCCr8VTrZh3veSnKcAtLqKF4XiTjaE3Lenwh+D203Fad47JHM2xbf4ykXnHumQ
guQMCqlx98T0IIepU+H17w==
`protect END_PROTECTED
