`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HBYsQcJQEv2ikdvgdYWr+UXpChFglcENM6cZaeyJ/ibvETUVdg4IqJnhgRh2eM8b
CjTAIBiISmPMvOvLvE2IdQekYWGx/naoSMVE8T7J37xkubzf7utNCfcHCEuk5V5g
xtaWh1/KRhAXwcT50wGpWZK7q9/FAjPt4NkLu8/jc9g32QZEqUpe6MI9Sv61E0Eo
rI16n43sB3DblnBB/5c4IeU23n2oCkBjiRkOHyYdwaXJyvTEN8gimGKtv/AxMBaZ
14pjHs097JtSxKqrUoD50E2WahIgXSwL9EafEoNcBorXFXTJfYl/MkMnUErjuv/6
FTnDPJf+V+TzptIUWqsKsiA1p7nzwkyhC4xaQIucCFx/t3X3xLWL3GiumIVaUNA0
ofHmuEHQzaMQ0C7998CDw33fL/PESVhgeURiXtIvm94r3MZkh12nZaHo2CqZWIH8
BYIL3nonfClgIIlL8m3x7kHeORCyYMgLQr+b3d+bs1UrD+bn9XGaEt8b+T5WwKpv
ZY3ztbEtK8pv88OIRGrPCJG5yfuCkz9an8dQPwXascf/m37quvxO8W1HBT/kN345
YV4uIq7Sixj8Qa4BTO+lhzAXjOS9M73vwY9lHJJQ5waabLXgbhweoi5QnpiDkc8T
OL97YDWwKUTdznOTE4kwinFVcejj3dUkFM/Huy1feqaEIZExfI2bkSDYUx4GXEbz
`protect END_PROTECTED
