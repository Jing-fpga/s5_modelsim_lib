`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bSrPpOl1pq1mIXEItfJH1mhZiwCU6coG+uGjd1DFynCMNZMmhLK7GqOMPxnp6T+K
Q4tyVTolbgOy8uV741pnmUEJj9gryYcGWvKfVx8Bk6FUkzQjnNWxWBbIwxBIGjdT
TjHwNhjcgL1Xiyp963tp7iYv/4HpUDGyiUtLNuO8Eu/T+NwUY9s2usYylfjPDksk
/GZQaDix94f5zTc9VsCQr/7z1bZnP2VjJbJADtU5OQK8TUlguFc1FwqY0RgX8e84
XPz6SxDq5Y7TK4+WSDPbo+FzpGzKTVhzJkQNbU0MmcuDdip2rfDgum5EF28n2kXd
YV9WnIwVZgped2vkvsrYJQnpfEZdu5o/WP8wg1Afryq2X/RQEsA+B2FeTA3RVjEa
gEwFQpJofPIf/oaEjEb5zHMme55n3s6wAnMf2oJMk9GrCYPbxunamb8DyPgATlD0
EZMP1lshRT229rCUSCE3PAIoXpsOTnufiAyPzB7vBf79fhomD/y9CQQgyIxTmxML
u5d/EQpR6tdEvQGHpnXm08lfeIl4FY5rsHRdc4Y0ziwVMWcXjcoccjh7ojw/uW9j
DuTHo4N+DXrGVGiRwa83GsTHi9Kw2kGeXUjdKV2RGx0gw9ZmKUoQqspLQsdfEB92
/fTvg7AOyEVvgiGd6nQX1IuKhLjPmx6D6KcFAiWW/CZ+vb+5erNOj7bC88aEpdCo
RZlqkcr8Cq74lRqf2eleDeH1uulEq2al4YE2o9YBLt9M2UK7mD1FyQ+XyOZ9FG8w
Gi6UsoMQoR62DgmM5+CUj0zQZhtQMWYrlbOhpqhSbq1OYp3OEfwXizcZsoDNLgQK
LHx7itxoacG6ZXVKxeWW/Ic2diK49H/XFMxxA8Oe5vokJ0iYiHzkFIFsGQE7BlnQ
0kN7/rHPz1jbA6h/yI1LmN6UGwhq7YhVqsQ6WhYIGFepiwIm8XIPugEK1pa7OXSR
`protect END_PROTECTED
