`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AmShTim5CYD9oEbhxafh1tUtLmYAZk0zWaNYOAJhwD4cVfJSqMp0c0NrMo9wEZXy
lUG44OeEo7QW2j0WVrk+hUghTWDrOrt6PbzYsaX/SjSF9sJ+x54yVj/tPalQ3kgd
tole8Dj7LTzdo4Rher6cMQcsWSC85Xgfct7UCI4AuhGnx8Mrqg0fd2LBXlZDFxWi
pDYVAlxRe+kGRSkiPHR9cB3KRbEmGVVuUrLeafYqVcqGIQFpW2TFj7Wg3720Ah+x
rr0ESkMfdOpWsAazcw8sF//c1LxsrIiWtWIttRoQPEeZcEhgSi1NAaoxEfPwlxTV
o1LsrXS+lytHiOQGbGntQupYUQ9o9FXehL6genbpij2heG1Fg1tp8ajh+/nhczkI
x0fqTpCAIIxwmUsX4NcnfuppFOADZ9tp7bUZezT0ro8cf3rN6xtuT9/ifyMI0RWa
Vfwc+j/QoDyAexBISaHE08OUlBeufFsMJSkzg2va80h6asScdukjtZBWUnXsNg+F
0/HKBnTdHRstIsvDjiFtMNLrNs4qdtkOB4wntJblJ/AQMlcAbA27u8twpnjN8OgM
hCC0B0qwBOkKjvx6unYD3+3Urc7BBGaKCH9Q+lMDRi2C8NG863iqCD0ShXFJBxBE
Gcc6mckb5tCzDar7Tlc9GzkQTwBc7YRr63HNHDxsQDE+BhjeIqbQfOLIfcg8is/W
aA4LPm8/Wwg5LFRoelJE6mC9slmi/G6eqa6Tz49lxHKLmi42q7rHCneoJzf8LItf
Z6gF6sgMltMevb5bmRks2vwsk4ifcVaPWzj8RAjajByueyqoOEt/BB90DVY16cmz
GiS8B9BOKFNhgqTG5OAI2xGOhPTSD9Lcp7VaOnEIIrtzx3pCHUOiiyUbaK7MjOWl
mAfbf6CPUSjw7z4pV8I9mCTM+yHTdDrPHlqBnK6/n6gcwrfqIPg60Lm5ZjYWDC81
ub2JTGcxZ4BtodwxPKavbRhTSe1xGoY1aCbbl1bfEqzzU5WkwqoIFtA2b195v4cn
z2VX0AUT0YoyOHT8CKYgp/kpOlPpjt65tHGvFj+G2szqbWv4mgW1GjJoCD842s0L
iKgtGQ/z3GSd+Ca0kDvRpk5z5594rMl5rAryfKUYm+GR8M30JcLi3YVdkIYfgR59
QYn89Ui8vdZkOBdZ6q0j2fqoIPEMUFDBetVm3G+DlMGlsOVB71ar8pEacHXIl2QC
hsCI4cWYeaLv/bzmTwbiY3cFJayFRjXHFGN/BG7cIXiHsmESqxh1nGxUbRcdi2fL
6DpNVKFqk3Jz7dQ86BhsVyy5MJpDTe4pRurlXvlTxd7Kt6azH4SObNp/aPcS4OsR
2gLg1xunLBMNkDhmJTbkXev3dBOZEjM0xdROfoq+EN3CCboABA/2DF6uGAzLBuFH
Mt6zuJ4doMHr9oyEIouNCyqv2KxBAG+jg257czzElmSi2F8azUbKtQiTlNTs6+T1
n7coNZ8227yfcf0WTrgq3ZYN52WF9u0gyyNz05YQElNFCWNFEa2RyXi7wylZO0F8
jkUoKfNmzHql7eAwXqlPvnUkb4VXtShog3K7d9BZweDzsXhbKY0tUzXhCyxBwQmr
UGWsKcEOkw5c5kA70+uxbyeGC6z1C/Snn+2wVr2IH6d+Otq7u3Q98J5WHAy9kbz9
YkMO4TS9BH6I/xUvlSr9PRksqLADRzmVyNg3mCCnkaCN0gj/WONrDcq6hYCiMvGB
w/eqXAf6SKTut+lT0qc4o4fa3b6SMKWRK7FZIYi5Q5Ax2gpUj94sp1pAeAEI7oQk
o+R+0F5JyteF1LKaRcv1FhBBRp9+2py6RJ88J73OuJ89ZKsRviotM1z5sKgr6qQl
OubgBabH3WNh4sif/BwHDXahCTtl74GH3DoX5RfcNi1yD0+lluoacHqRsMniZ77O
ZQignNbpSpHU3eqHFlBVlp8rG+rr5XRvE9omwTkv0vs4wfHNKZIKZmm4lAnknS/t
OT/YP4xjbrVbwqZojzlyonqdQKUjnqMABbh4QpNHU3NIU3dVgNgdNvyvR24nvLg3
j+fz7BWHX7nRUrhrugDDEMVSLKdtcKet+s4XWgtNXjQlYaAWU5JpOS299DVCmUbE
yB4cUAXqY9NYJy+3AGs1KnyOdrpIloTiDVXHGjZKd5l7zA6MGYI+1AI2MAowbB6q
V0zWoRpHaQjqVum82OrF7bj4NgDR5YWGl/+EL9iN7tRMNYLSJhWf1F1IHsAHP59g
uglsQbKIv2ZJlFJquKRAlMRCBHSvZ2XfTdJUtxuPa2lxMATvUyEibLteh7ILRaJS
kjXqJm1g+t/8NAtbClj5bJKsAs6iCy/gxqmUIt0ii/dQ8rmM1SYMSKxDT8IrQDnw
t7ONAbr41fl2tsG/6hrYl3+60NY4h3ogJEu7xUotUfzrD1u+AsSq7wj/cEdgua+9
xG0Niy1SzwWO4OD1cqFkmXidQWwbLFo5WjUuXqRxKPrfrCHrTu30NZU5B9f0Ts+0
vhyr0evHcLkyjBdyYhCvPftfW1JCeuXpafknK7xXwmgWUcVQgRqi6TT0mN1rGpoX
vwoCDksx2GLpaUvMAiRoS1chm6F/mZRC+IzTnJhsDM3RHh20/blAd1vK4gL1b2NA
zcKr6oRD6ty5Sv5VyerwNxHUvlCNiOUClRSHXKEKEhX/PzzMoD2J+7PJXCaslZqh
mqNN783tz8gkyjXb0WxnMeNJWDtXEu7DdjO58q2Y0VoCq38DO6iQqcVnluAZlMjQ
7D5rF4JsyHaGYyAiO68NhSRVNEfKWjn7Di2eRZeKl5o+5DRamRpTUEg6ov9HNrtJ
tGMjXosIEQ0i0PZjpsKUCraccpjs4priXDX1dccN0aTNoUW5eclLlIlqP0F4oE0O
UEIJ1L4Bni1WljmR72hBWfKq+6WjDfQnYHFmA4s7JWw2/97CLiRp42aNmLe7LVQ/
hsNGe6bBblPc2cIDnlHI2Y1c9ELIeuHe0yfF1X7Cod8fvk94db6vl2BHbAPZ5QVN
dLGAYbvxJu5tfGc7Qb3p1oQSwjc2tqlz/KPNKOUMh9a7Qo+RS+3zNRFDqLqcdyQu
dLOyC5ScCmQXumTH/OLadAdh4VthzqIV488Y1RuBTn3LQg/00wJuJbhSgNEEzTgk
HeIOmBa4yUYHylMHsRoo726DOC/qqrao4IrFSTkUk3YWSuaYltTOfYENiPdAfVV7
sxC4WtecB7PjkiRUeW+GsbWHPtUJ7Buh//Pljg7mn5C1VR0IactlOd4CPHOJSTtF
wMhvmdW92JMFaQCf+9cl68ZHv1mLD7ZuTQlB6j5orhNORxbQgEpLFdDurbRTGjj5
fex3UwYDQSH58c/9nHnvaeIEyYkCP22LGAHipCk8qKGxowwOY5xkEFkB3D1+6rC8
kxm8a1B8MVLE8bmLlkWLcjg2jxKYz2pW9D1ILq97cdLrCdIm4X7EEO4vIKtm4VkV
/3NmwO9dtMooxOcjbKpF9A2BbNNnjP4/alD4HPpT7m5PFJwO7EDFFkI32qk55wEa
qlzR1LXAqPBTCKJ2Xx3xe2T6OtrKf7I9ZNa9o7PceCJcgqB3CjhbMGYU7yGMTcSp
491tgws5Oh4H7ssyG4nArJCZpWtrIb42oUCqN0KOjN/A+SXiVbIwY0O8ziWmPT55
CXCLfpdvkCgK7qAblyT7RY5JCNcvUn52I+Yw+6zOMV5ibkk8EYV8bafhLqnjmdUo
Ai1prexESLeYkPMNiGhKwAZQAPA+ZStYW33ZfURQc7lwfDH5y/jEOM23eM/PSzJJ
pg8LANModzIPLn6jMyjBTxjDjRO+Rc8rVgWRozUA9VymhPXTbEribGMR/SsnVBQc
ZeZhwMfP1MccsSY43ks6hZmjReoz4JeuVeGkjsskaaEs0iNjTpLcrf9ULVAXVMs2
zUkUYklw1c95w/plOEsa8YdwWlOUVQWPvSgNg/NJMvZdJKlr1yMFTOVOtO+EH8Gc
ZTRTZC3x46Ar9HuHCZ7XaUx4Qrq7JTGvW7kN9Cao8W9eyir4h4fwl8fTFc7oqFAw
INxXeqgU/4FDzZWPhVt6DG37/lKJNtEh7UAkz5bWMDlg+YrSIBrgccVDs84FZeZQ
ezpS8AuEM2sWJ8K7k7Yycvb4FazUSxH9H9uF4MKLMQys9v0pp9HSLzFFH4IA8yhN
WOxpq1tWDSkvrwXeZNdyh93TCXKgoYoTpyiv3WD9muhijAO9RitJgOnSP0zOh7a0
P0Sqoe7KH0YqF25+DX7B8bAnOaxQUyIC8dDpSiYDVuou6PYe6K/mMnmGR5YPOytd
p1C8NngcwNzE4qSP2MjL6lp0ivqEa/SsN1hhanYPvxCB9GcT8ESwdPZYWtEJGkWd
3Uzbhz2RmLWtY04G/PqRALriXQlfRVoFY/41NCKP3Hqqgr/oXdrKMdwSn2RA01JB
ZI0gitdZwpFai5+Ut0M23YoQVnBX7SCU/FcAbWIFvHMANKAB22UfwAuoJiFTGqM0
HOvqjKX4zNzgdWnPEwEeGlbLYREiapVZadm7ApTAsQ9wY5kectiV+p2FQBu42UX9
NYd2QBae8+arRqXNy2yLZnRaQYti+ivnsM30ouAaJ17L9L/jEUb0fHbWB0PuLAKu
y8UnAvoz6r5MTGS2r4vRx+73OZ7rxW32/oWhN82beqBwnf4cnjgsq9t3TBpk39Wl
27ODIvBDp6iU0E4pS0xM0Tue6Lf2gY5MnjXSU7CJ/6X6xO4ie07qWppxhJP8jW6/
yYOxNu5giPycQ5/pXFqktMenesZLKY58fG2mcTbIOol7vw365T6r/wYQIj9yPZiT
XH5cpfdbgKg73cleubnET+uKZfEVJwEodRM2KLppRsp+6FdEqh1+5+4YWD27kOUW
rz3IJs9jPGSMqqFVYesGh1t7svXLl0lt18m/RPQuJg9FhOwWCEoFESkIWx6juLn/
98WxVzYD3clCQAU8oiOm5Yxn8LblPsY6ZkL72iLYaU+yLr2jgh/x6jivxF/ZaZEX
soXv3UFsT2MH4UvNNiWSYnS2J8SveM/vVZNfdXest3g+3cQp4R21u+bj9JO7IhES
gQjQ2ltHIjfnpMXDZ+fYtsKl1O4d4nCS/BRJX/IWSJFZmII54oaOrmHK9Ark47m2
piNwoUAiS61l14DsMiOZfPpU8sWnf4TsX0ODx6LjPQQzZPb+rAnnsWz1h9VVWVoZ
CX8BWCQ9+qgu91cfOu52cuXq7KeF394m/LmKxrwAWfHKT4egwhTUGfyAxtsMRsJc
OhpcJjXDedj5JmMeNdc4QxU0OcF+jQR0BD/Yp8IQ9TYOdAmg5t5gMClcmaA+Xdav
KdBZ9cyKj5ZIghCGQN1j1OC4tWroPjxV99QhSpqVT462W/GcePsvic7ixLoXcUEQ
OLzlPQ+fU0yz5k2+mglAt7AcVh3yNg9h7eHEFCGFdJI8P7p113ohLx93AI3vf0kO
+yVS6NAliMPvg32+Vd09cLdXPLvGku4qbqx/zyF8vDHy0tDoyZeR4yrYhjwFQEmP
Ny5hzGUY9phS15iknaI9LPF6SPh1/jHxD/XDxY0DBo9g57BXibHzI5RtpTthdl27
/c5Xwk8KK6nMA2MONZ2rVvaN8dAKwlTPCEBHdeNcZBUMGhoq5BG7rw/Rp8qCRV9Y
+OriMJSRnpTcCBXl73GW3neQfGso3Y6oVJtmAhhdDyi6t2xqNEoifBhoRbFEs/wo
klghjE/5xm4f4Tas+7PllYljq1D+iIl+VoleN4B/xlkU2BVosNs1aQgEE3aAS5mq
7krqesF8AIeBKnKI7FeX5kpcJO+QqC2y1NJEAQdt/4LmB/b4mmzUULiQfUeU1OLv
o/A4F7e4/tvQG18Kk9eHNAA3TqoX3MXKKrU0nXlDviQ9lCK5IC2ycFRIo8W3T6id
z+GBAQii6oVjPY6XSx20O2xKXiCBEpzfw76cAiRRIv+u+EedcLVemT3a2VyAVIf7
blqIpEntJoHS1263Jyr9HwFoCXzSJC5wdudGfmwQhI++QH/71f4YeZVX1OP9epTQ
txH8QM7qMc9Y5iGGzf/QGeX3fYjZjVdMVM1Nkt3rWYfwAjyb+QZAMPN1VaE0XKJn
HC5VpS0Cil1J6EdawBcmTbcVduXJvtyovO9G4mjpfoKQcpFAJyeLSjR0YJUhi1C4
kRxP39xyEiS2a9jL9CpmdWaKCyCmxzF8TUIeHOaMx0xh/LzPpln+aWpzNlDT6SWM
+ynY3gyOhSTICOh4QUFXAOJF2XymkpJTZYhJmxxlPU3gYmMlOAFG7fuMDXUzV/Dc
LwIZE51rAuls4fQfFL+028NwfKiCtFfasFPZ5AO8Jwkcf47lQIMkcDQCPL/lo4vY
X/v4jq2GZw1VfsFm7kpQBD2oJjgap2PnDQ5HmPq/4TFGceFkBaXNRQjIwJangU7E
TXzx5Y9BqTVB7vIYaAjVVo6ZJ9ElZLtW7LQ3tQdlFxIKFE3f15vSS+GLQPr5QXLZ
akcpOgFRBWRcW2LGryGXdZhASFo0pmp3vhKr97o0dDQKw5quxcRB4YRh2S4773AJ
/y76iB8qa6Qm4bqBQPLrMg5/pz/s5KPb1N/RuCjc9nz9t9PWAlmq4AkO613JbzVQ
R/WJdxn/VlTjS1a9eRRaxllKzqhYiC9Q6bBGm5bl3w9ucfBfTr++xXf3bB15R14P
`protect END_PROTECTED
