library verilog;
use verilog.vl_types.all;
entity stratixv_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end stratixv_routing_wire;
