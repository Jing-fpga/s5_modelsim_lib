`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qUgiopoDUpb4IxlLOYDmgYC5f0hinFJvhX8OPHSyo0hfkaFpecjrQepjfQ5aQmDj
yJXigFJ0V5ZNU/c411mOnfHwoFP9jEnAmQg7s6IWVdJcArc0nxwSjTmMo+TVCDP9
PJn+SDJ3lgVTmcPDQZKlf6gG6vBYNWH1nCje8sJPUaF+EHFokae409AsdmOyUvJJ
zII+iLtDrP478WgWav0G6MF+is4Wy73+F2z8aThI9gvqmiKnDg+GQa3IBtTMr28b
x8J5WWx0gAu18g7UU4S2IdKvNntUxcqYqtWZHfQcrAyPhxLkMaU3UdxXq/zOhmXp
zEdQP0Mv/BhUA5hLTT+LGiLgGjmMmsomrBSrnxlsVlCBb+wTO0ziAjJJbS+C4dVN
niWAhL0c5/2wCuAkdx2jTNyNFRctvlvBwebF+biAyOAKmas8Kil6huS5skIg95Yi
/O0A8kdysF1Se+7oFg4IRR12wznSYb7MisHUB8BaBoqzD9HjtG+jvxTTBWFx3t4E
4Q4Cl4blKMPnY24QEoKG8IJxfbXrRc9YqVQskOP9AIYd1GhCrpquoK28NtKjPcbu
l45WqVvyG7jNmg1tIze5le30yh/BzF+99fHbSps1ubREaf5GuQS8fbfHQOSsaDIx
BXhQWvH5mGLveHmJoozRzRh3cEUTRxvZ+Q3V6Lpha1xU39/nNLUiPdX+XLCA0Sz2
bKVPYbmV6Jn+Fv6KF91f1iz1JXdnBpOx1tYD6tknWtE=
`protect END_PROTECTED
