`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jifT6XXDIn+p1mblTvYH6e4z2hzbqaBPA27h9N5eyTjbI5cuM0jLwBMbWZs7opmF
UJxlFQ7704hycsFai0YgI9H7jNWKNYlYf+osIlEs2c0EMUU3haQGw1d4WxOerX4C
32lXzbFUZPbll1e83Kb8guVGLl4wRqevYP4tPAsY1c9qkjMAwiXqTDMNvm8vP5aK
EnPNq+B2CuE803qKr4h50fZ7X2/m3OZW52we7+tPozjC/ItL/abTAuCQiTYTamIj
2MzvdXUaTi8wzz/rW4YLYRKDDrsRU8Cd+5uBqV/ZRfEbNmcf9e71HMD9E2pTO+f9
qw/1hy5hiEwa1ObDKkk27feq+r5xGXP/xW8pKlcZnv1GtUhXGp7f//NTftQsfoSW
ISGWFEUSzaJvnTbKSMNln5Xr5qa0p+4NatUGBRxPCv5Ez6BYd9aCgd3pN9obGVci
vQvIfmKCgXGhdTnT6N1c8ipYmELtEJmABnNLa4HunnYjd0TnCByM22fIWWcTK55r
U6EwuEsgUbV4Chewg6+8AsgauH0Sfo9nYa6I89HfbPZE+jwwVNE2JlQWxb9Ts/KO
h8TryvPptJSa79P5I6NDhvXnc8BdJrfZ93+OnU/kJ/iIsAm1p77tU4s+wMJdeCwr
F4WwjI1wHEgXdyzc0zwgfYYz+vqQNqZuJkGCvCsBtg1KdS/OZMmPfipkzz1DERFK
EJ41IF0g9fPsLB2/vmjpX0hUlsQXdH1AsdSK8hTgTxN2oHB6V35ZGyiDRvSPFA9Y
U3bkzDKzUrjasFZC0HnzsPj9LicR6BPvd2lDREgMrvCsG4uFqsszBJCRJ7AWSjuC
X+6vKSdBdbrWryWw/0nzqBk2LUNaJPeILhmb0GHAOvr0R0U+pKcej/H/VWG0KiWD
+udR5XceqyS0958D3dJFoh0R+59dTrbXnYL71qk4Dn98yV74VWsMbU7i/aaaM0Mb
shcQqk//oVMfDKGnHjSxuQgcJn6645kNkPhEBM6d8tIAOvEP9v9Mxd6EEpKxmqja
onUgvvCyhVuygbwcCAc8/mNYlfHVB5VGaceeYhLyUoEuNT8YqCLA/4FKUdJU44be
TMDcboKe90a+67/YK/xDtIOUTfeQB06geHZPauexue1NttPhE5qRPZxT0oMVFRv3
3nfhTwpq3jYeeEd1jqVl+StPXAkesOhBP0rCRnLs2KOfew8G5M7nFY7PYk3mrSoX
v+TzoSLYoyDF/+7cOO040KgBaw8KEPwI0190e1l0A03Qvc1aUIE7It7TpMgXHrE0
pFiIIdoE/hHALOYPR/hZy/et8zk665j7CAdKw14oz2QdCcNIuOSdmPsVqahCpjuZ
lrp8dBR9mykDKaxdGU3q1PpwgcDmpQKepuD/Dz0HOtk+eHrvf3TqQdx8coy/bXJj
q/FzMKE/6z7jqkW68aFun1EfCdM52dV7xuHYKu9Zj5jCyf/GGANWlT8YItWonHhm
Ih12OKdZFOtffdXYE/7YnA1hYaEJ39FcgdjVTbM+E81/3260v8aKVzS8BtE5obqn
rRsRHNTfCxkluHqRLyJmOdoWg13z2j5VGaCtxNsr4QVW57vW5QaqrdxfLTFqOlPU
3k87Bbo4TRpW2Vm1ovA72OLzsNpF4gZUNy76fQzzk3Dp22fTSxL99/HxQfBcsnNq
J52fTJmuqNcB3kw4cFWbpdqyKhNk/xYt/ERH3FDDTLIXb+v18h0xF3DHx7+VN5RA
KGKChJQ4g+mlqAWLQ1oppclnk71PwPGZ6jVMhJzqzBSB6WFsQB/4fJoRp7cS0XXM
I0648xBm5SidjBMmt2C1d0zeaDf8foLWm5KVBEHk/PA/YibgFd4SezJ3aEigGEK+
4ijjcBqbF75whwlRFoHu5BnRurywaPDszt4jjcdi5zoliNHJDSg4fu4IFiOUMH12
43RbJJITgrDBWB3KHYWyN3BNxM+Z7Ln3nPd4OfkRxojrMo+WP4AoZ3lgwyEIi7Nv
vQrNS7Obm1nWZ9p7zKz2eO2vzc+bK71dyaIL1/L9yGmLsfKBH9Wpcj1ItglIU/MY
pj0bkza9Zc/h+3oZNWvObebd8gShN61tpdDf04I2/6uClpy/k7nLcpZCA4PiKYxx
I5EOsmqGiNfQnq4m7EPqoPbIx3T86quWimB/1d2Ra+gsSF93u1MMHXMIL3GjVgMd
qlCz7IGKfvzEHcsResY93lvK/YhBashyd3HCPEluEg0yP8Fjzt8ZqXSinbpSfc7c
/PabgmqQ5aBXJ+AVoTS+fYvz7Pj8jyM095N71+WHchiBX/hdUJtlxp9UAoYTJIgh
AG1CG7cIAGflHlcsZDxm8w==
`protect END_PROTECTED
