`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eufvgQi9xhpNfTxygeq8lGybnGYztlna+Kv+I3fcxi2BfMeZWa8yQ683QT1jC71+
cDDqP+HQBs9q1kbzlOr/wZCN4C8RGqDi23GOYiXDfPst6bcVGwgxiEEptdMH9mkD
tPceO+1wiUekCeiWqY9E6Kl9iA6pzJZDnfGk33uDwjRQEQx42UUPRekNtQB49MBY
5TUCCu9ZWNY0Zi05Fc2eV+H4xCgouv5d/9sId/l/akbyP4w3iu441fWWVkMzYnKS
lHHIWMQiBlBlN4Rlfhzp5Pw6+DWeGCl7BpK8Gi86ruBPdAUOpaTmFDjY1yohljEa
MOAuB0N5yP8lwkuXKfN256UE1bdPsXHyi6KY+8ak8v8FvVjcaAknQJASD96i3Cuf
1n1TK98y6OCiEOJSemJYWLtQ3vFDtAU0UUZLAOQ4J20jmzZnfDKEzKk1Hu+XKY0I
gDO6VrZaC5ZwqKiaJJJnZUgoD7ylf1QoR/GB6bHI/vuQydf6BpGbLO6HT7jvE6k+
nwZixEkOWiIHSLCL6N1CkO3cFuithFRBre07eIavwpALxscTA2lxR55ZBhYcrpF6
FuPZQD8LxH1oWESZy93fdhcrrYnVPgR2Xb5AJG0oHGsVAfH31otJcDZan4Ftj2Rm
XTu6jeKOSD9fGSJbRb+ZGF5b0/J+WqarHuYbQ8r5F54D+jOlL39RVDows8vSGFn+
Hqv/7pLFRp6Es43apKF1/nt0VZlvw2iZoPdPG+bX62tHWa+131qLtqkmpUZhTQO5
FkdMGZ6fFJHkFayTC4/57cHIgCnGJSbVZUAxV/capG2RgU9dvQNDQeBCd0GFZtUg
MJJAnPXfQnWXzi4/WOYCUtWkQq20VVjs9NlZGmiPqsD56xRLzlQfekeHfMX6ZpDW
R+sd5bUxz9VH6QIoKo/PclnWC6sVPyYe/4Y6lXPCbcttY0Ou+4jjdz7QDWqY+9WU
NY9+ILMY/cNaq9FjFQgucZfGVQGFv7hR85CEzgmgM93qCL6jwTySHoxyMZpawSSF
59LVk2dJvbUGP4k22emM2uxa39cPf5g4VZHlsW5XkwbThg6+qpchMlSc5SMy+OaC
/Am5yQ/stEZveXvquQVT+2jg34pEXtEGWu9hZU1Sdh+KwtsWtuhTYcMe6r7NziVZ
m08L3cACljd4djAYIhHwYqxwfUt9MhaS2kIhhfepIHkTHX4waT7U/e5qStcmurGG
eVdhNRxeMR17pQKYGUZFORRdpQ6zsIoIUbrZpvI3KDnt3aCZOK4ZMF/4tpRItZGS
mM69wl71+O4JceAm+l55fLviEtJnJNC9RgOF33rySf6RwXkxv9+d6A+7/Hyl1cV+
p89QJ11NFVgCXOKhb7b8YU6ZkVOuxIvUDX+1SXCKvf+2XcBH9NdR14MgW3MjwJN2
6cZ6kdWJZ+zvHNg3kin2xmHpUN0vpPQUBy91b+jfiQ9k4x/f8xLx7g3tmHXfQ4dG
7Bb7t1njW3IYnK6NeLAgCUpyUaUt0yXMsy0q5lckck+uIkhN5nI9GL9+PwhzJjnc
txZ6cOTvBMA59PftFX55x5TJD2eXhqCyNH6OKKhgGHx2C1nAbpoITICVoC8LDnqJ
GpHrej64DA7w4sQsxOGw+k3LT0sQCjmJ2yhIE6PortXwv7mcanlh3VqNfwKB44vc
5MHHeZfR9V4uY1XfC5ANLl5paikgUt94c/a3E/fvDdn/PPin8Yg2pU+JIDOsdLYh
VdVXtYVc6Pmj2pTnpz9ANa5dkchuN1Cc1IYU0wjXvoXesRwbZJBEpf+u2GCAUSiX
VsrL/Fquno3rP91Mk/Jk1hvhGPCFGAKdqavH5lmDWVQplWBIiim1LXrsO3MS0etq
4Z2aEzOUSn8vENJzFnsQ3o4ez3aoqVjXJcQW4wkEigYkLo8h8JL5m/h1qajo2+SH
9k0Fitsiauet8XgneFgdTD07WTbCJXsm2p0dDCWufbPOmJ/rt6sTRoMp/F/S0pNo
2BZfkO2ugFDH8Z2TGSLmK6x2WEk5TpnItbn38qEdDOtderPzhnLAUm0jeC5odP8Y
oRc4qenWMDbpkEEfxuB2atLdbTOBhfzILsqPlgJHVN3bRfF99mLFh8TmVPHdNLNN
UoMBrR+ua8N4Z1dRqKyBn3s94L1o2tiHHbKWMCMbdKx61E9G8XHO4jQ5aT+oykMT
JxjQqNqp1yOeddu40IFCi9VYgmVv1rR8DXr6XfnZNAM1XYs9V7eHoF/KPjC2bvAB
FigxzHwwXQVeot6UDO7Gjrr5dU+G/2bejb5B5LaNizEJAZmloRmoydbJQ01hwE5I
ImjEkoJ+lOcgYpzB1IPLGNXUyZF68y03MxHCeaXrScIWEg8sxGTy8pWj43byBdrD
LVsqQIvKihECcPQlUcjgtptJVKOhDiCOMaRgufAg/2gRtXQHuC6ICPhPYsHUE61b
cQZ9/ZNCv9pS4+1GQ9afaevPr7oU2Hi8c6cOYPhVEK9rPDg7tCWIHm1p8lfxVhYp
cUtIsGXuZt0wfSf7+Ep/nQXnOqzL02vzTfJk0FDIL2S68ErA81Oj8tFVZ4xQjhKg
YXekifU7KFRrz01NZ7qIuKyokDODKnxKOZ33fXXefbyE/cCbwKULluH0NLlfhmph
kqWLksoYBTO4NTE9/4E2stIEeffW1wc63EZPEqDYT4T3iPRk+QF8cYuiLqZ7xNwr
GbPeGZAkNp1qEs28UEif0tsYHL6qOpZhKkFXefWuI/7Epqghb4lFbCEo3DkGDLRu
s5JNITrIIfx79EpVhlsb+wUnsWghUTaGzuWXLxBL1MNUw2RGb3RbZP7i7nJLGSxh
VoVa3KCu3AvAKGurojXONgzsZs1mBBtwqX6d/W3vTMcReHu5HW8+DuHy5CosRoEJ
BDprtwvy/B5MHnRZYlRHG26BJfkTX0GkyW9674zgAD2MRDV306avbL2o9gfzI3qT
9mLT3utRwQ3u95DcTzRrNgOo05kPHHyJaDrbmHwZVfmtmV4cWV8NnEXSV/9axc5j
degegJ4hN3yoFDh72F7JcHKtcRArum2SoWLxhcYNu2F0QP1DUo172n7gsJOEsVMd
MLMz0AQjrED52RLZiro1kUdqgSeBRmG7dvbi1T5dgbJvFWQgUV/3CD1+W+ep5XTd
On0B70qF+Rf3kNvVUREsQSuRHgIzQrY/mmdEruew7VdwBPfEiknZrWaRRlmogUaP
dZMvK31gTzODn79S0HcKhSYtsvEF16pB9RhnkjF2cY/JaOTwLjLijTRNtDc5xPL3
HkTbm00cNEgMcnH/0xXq0CnbJ//xmMSbhDYq3q50PgY2ASqMsfIl8tYwUk9UV9Po
P6n8PV8ffQEiNql8B03OUExPLAixnGPQoPeFrXZBtIGY4BSOqn9d9Fq7vavEC7LD
yveGFz1RsqibsQsmqC2CRqqV/vWg6ZTkevzEusMZ/MC0+kdQKm5sw5S20niBpaaK
cc5dGXKb0ItTbPe9uOe3AaFx+Xxvyb1tNBxs03hfnFbFy9HsovwrM0x9Unn/+Nal
cR0oWCpa0VueCPC/ZRk9nrpdxB46krPefH2s/tbn7Kq5z0WXShxLk23MhaM7EimS
EZLPe9TRa9yMDZ9mu0iaLxa131SzdgZNMqBIvkHw53aFw4ODSuvkEeip2kNzu2E6
227iLV9rH8KLvtHfg4n9ckVq1hq+SwxG9j4YUG5FjSlbEACQR8IiW0Dbclb2tCxK
ZrKgbDBGyeVAxOLyaWDhw1+v3ekgaBTiynRmiq5cOCSnIKnat8vER4rBHcoEx41l
J4Ozy/v1pgi5eKq81bkrXvgtDUUotYsZrMgu/Bb9fhJsFzeJosEuhXAcJAdYkv9B
cW3z0BQGOWL/7WSPKElzlAI9aEl/rBnotZ9XoLRVo/vYdI4HNG9aXoKmkj2T6V+E
Y7h1/O5mDlQvecXMLDIXDokyLHYE5gpmXw1irgqGdnWYgWwtBRKhUZPph2zcRsMt
OSY4F0RroMbco4sxpLdAuRAd+LCyki7Tx4jedq9h7KFvLpy3K1I92bTQHCwsj+hR
dRaVbzbfvxQGCWD1tcaVORVhdCUa9f/bBG+1z7+bDcD5fBzxAJsn/mqRemLXpRa7
YNv3Wn6f3fV74yOvc/qQnujP9CCwKKTCd2dY4Ij2jyGALZc5eYoLTJ3kIKBYG3d3
9Z3NDumSx2Cj/7sX0qdNCleSLxWUQ+imiUqb+MJwQyMO4m24MeX2YckGndA9fCJP
2DUx0c3ecENsrxDj7KnjcthwCcUkTmDZQaB3RkZGBekJGHXp8YydkQGaqgpzm2ta
u1OtShEqxti8XYhyE++1XtTzMszEPTyAW58hKkNnfBLIFresgbDVqvh5OpTQA6H7
KfWkfIWh8lQ9ogiu/njb6+JOLiJhsfxnh4lO/ZF5u0jjlMeQL4L5qowb+9uEyIF6
nfRN7sMHXc07KuKJJ6kv0aqGWmOhMeVuypbjtP3dlImGYgPqpG2MjeCyN+p0LzsZ
vF6tbZw9m2qORrS1qLFjvk2fVjtn7EGQaLoFEpyCypkgKgK+KCJuQDReAULtsS9c
6i0BxS47rmM5/Eb2Iqqqj5JCCFFbiTo3Iz42bak26ZqJ5/X1kY7Ta2CJZfXP8Dtv
ByCIuxLoA1I+G/wXX2Dx7/LzEywJIlAWMdWipxJdU8ePISeXBUuClkxehr6LosSf
M5jsjrQk7zV7TU2vm8faR/MMpKdP/3O0Xnk7+NJixrbwZqbciJmfr3xrU6S/6BYi
38jv6hQKfO0U9FyYrFqLuulRJ9f7edKh0bSyp9HiqLRBlyn3mOUTslgsCT72yq4I
fcm+54J0X6kdMTerG7R2+N4yf/G0PdqhgFD+wx8GJzvGgV5E4WWzqZa+IWGiU0+a
FtO8Q4UHEWSOmDrWIxJ+rXjmdTyDoL701L2WCF2yZU3ujwJCK5/Hvi4TvD0NfBPl
1zOTzVDPcCG8OabDl2lWT1UD1QrmDQ3q4dQ6Rb69SI26qNWBpsDx3Pspb4y7aeIB
FGkL5mFgGk/S6nURYgBnC+XFFuVgNHY87FGvQzZPb5itCoRtUUeAeD9KDjuAo7Iq
81hEFTa4UocS+50b+J7Nfuc6IfCVTNhr7qeck5d6hZMMC++Q4UbXYZcUB8YMSTDP
cKMYriajyH7qZ/Hn+XZqOK+UlxDmC4eYm9AUQwRtu2h5ndws1wGPpy7TZIjZDOg3
a8NXcqZhnjqA1r96DeDCEWwwGL9b1JcpKOc5V7dWX/L0eDXvjFePor7AOdIBTtA7
GMObtWCLwCjTio/KzWKM3Nxo3nMZS8GWf72XH1yyiV3rp1KfY1DKSCX1q7Lk3wEd
igF56tUU9E94eMkDTI2R/JX16hW7waSzf7De8zJH5yIH7xrCixbUWx9wCNF4KKrK
so6rDxY6FgHDQfknuQO2cHzyEDi3/tc2HZQbIUi7xi/X+CKrJiyTNzVr7vaYA0ug
bWQm5wQ6yyArzsfWdGP4Vb2FgFHfMAouGeN7sfW0dhnZbdZtDmdfHLZERQnLGB8/
gnVQx+KgvXjFsMolHQsfBLhSJbFtL3PSM6ANl257p2Ek+/KwWa4HTdlPblT8PMNR
Y9peHmjq+62T5pYjVwUqA7sg5OIzWsx77SgzramWBEEZ41+fOjJ0L/sFKKjAbgJZ
8f0P+iNWxFWHa/+THy3L+/6zs1K3/IkwpSSDmvhSxTrbCHqZFBw+Sj9rFFexynJc
QT6sebH3YpWK16snGjPUDl1v2MCvYdIU37Yl9HqeL7bWs8fQZMFSFR0JP14/t3p7
YAwLLGU/9Kq+OhCE8KLcVtqCO/v1lQ+8YYGOX71viJ1F0PWNmFlRVGWVPBkUY8Hl
vA/Ndj7YB22sK87l53ysTF3dgTA+LjNX+wcVoYcAA3qz/9IfbcJuo13fXBn9sgxU
rWTnwDd1FDFqx/GwfNOTjHV1RSCXc+kKABckgDL4qrsNhAk0BGZ4kTxLFajFDnH7
v5U8aVaf6TTY7xW+mW7E4bQNPb7o5eJmoqqx56UUDPslnHucnLztU0YrNU5/Ad1e
mPfFG6pD3r9+9SwnDDXyvbaxqDJmjfb85f8QWkctmsrmUcxFlrsIT99KGodG4Sis
y1cFFQSlnaEzyvARIz0uioG+F2SmS/TESAGmt5/Iq/n8WtLcqp1+4qcS0DB11N2F
b2/oHe3+uzfHWd6GeubpuWD5hXRZezVMyeKXvdVZDQVpQq2IP5asBtl13Ljh/Sf+
sjWygrXD9LeG2P4bdyOKlHc6dgKwTFUYsMDeTfVaHGjWNiB9KgTfXtTq4tVV6F/O
CPPDuG1HfBX/0FVeKDel8yvVy8QZufPyg1FmWnTPO0YivIDDHOtHYMQ59YnDXrvg
fyICm7xvXLQVQJVw/IUNySxCIZdvkCsqx2VROOPcmxaGxapwMMBRsXkUaKASHY/A
ax/9A+yy68azajHAlEJxwEycSgizemgWjjkwiHDKS6WlxWwPwzrrdnWvca5ji/1V
X0NIZydtKKDwBsOdqAWhhHmc2969NaWV/wsGiTR+zjrMee9LSvERpR+7PL5YUWzp
4FdjnoQHpTzhj/Wy712GhJ1fWafq12+P0RQ+x86/Grb2FEiFuFuHhX8KPcVtAEEx
9B7L1wpe2M6uNWZiyu4kqKnMsuKQ5vVPsZi9AFFzNr9MhA+k+Pg2i2celYbBk4+K
ZwLPgQEs+M6/slG8VzH7cbldyyuDa+qg6jDF4cg/YNd2deTGl6ELPFge18m5yxXw
sNtg93J3JUy3u/hgyHRcyny5CRS8HzoI73qkztc9J2S3UJumO06cMisJujMTOEZf
3wSD0v6h8EMxgAghsIVvfhbK53I1akKc1qWr0RoIEYKXNsyvLc5RqBkYEOSIFnbK
Lwitqkl7sozivpaAKriayZXSPGTHhm/CGx73dW9uSIDI5UCzScoKQt+5Tr5oYXgr
t5r2C3leIaXis8OJl9Xo0bB/eNcBqLkUj3Bd/XTVKQoDAiuy8YgjMAFn6ZiIhzxI
`protect END_PROTECTED
