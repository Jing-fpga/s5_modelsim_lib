`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
thCx8/A6oIFBoitw2a5oH8AgHpzHW1ja4guscjDLLRGCZQSdT1nAjzMjfmMNJx7d
k9pm5Wu7PudmETm68n+95KZt1bn8bpQIpBIUpNWGUYDeWVML+lq9FaAgxFe0peJN
7/07uqQPcqkLNU/DhN9slsMiDdxy5XNmzOG1Jpv4qgrRH1oN/SV45FrDxTRwzwcc
6KzemE23U34h2HHxOfd3i7leXgguRO01LnpX5T6uwo9myT0qSrMItlwThsZDI0SP
fcFcx5bARntU2BbGS4cJWOlQq6TkcH/R5gjtWbxEHwzPf8QR22tgIm3Z2nJbJ6Zc
M9fXGlZHAryspb4IBcBhLO8WY9us5CXx66IUWnam2VWS/RUS96YXHdGsPG5NPn9a
brxfHPQcHGET2t0kP5MquTK/VwzaCTmWaTMIlHdLulDtJyGljsXnDVnNyFx5sp6+
VL5s3q94cMhuUrbQRXDMFz9K09kg/KM2a7B5Ky1Nr6dicRumVONibDU/xbRXavGN
DR8S4t1nSLe0loOanjr/i5StuCLSKIrYiSkCQoa9suPSPBb5B8rWoxpbTnVMfr/f
lWphMe3ofptfVKQgESjhBfC5xnYiGjwdwb1ilHVggNV5z2VCCZagZQJ1C6Coz78d
JEohOSWzHO7Efx9iaere6VTxYM6Z0A/DF34C0GFeDcqy//fqQoljKEONtbztvUPa
nAJBNHd75IHri8gGSdiUDEBnFLn3GNrdbtOyRh3hsyP69dCa9cmT5wDESc6egIfH
HY4LwBuS4nwfxWcxOzpdbyCOA1EtIwXzyvOwHMFPSI0pQ8jcCACm2goUv1ab0mhf
e7u+sVindudCwznGTw27HsrudoB+gNLkdMHLlBqizmFSZho3KWYgrPVXXqVimgh7
R31KRb/HamG+7VSMH1j5BrFXhMGiNSd4XllSsXMf4xeiEgiSQs0rVjBbti6z1dXD
ZLCRookgmtIk2FYKLvp2CXpo5hsXb9mztgJXMHHQrW07RgbowIp897swtTy9by/c
`protect END_PROTECTED
