`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YGvCw8HFkJFjlxGbr3ijOTgB+pQsPzULgrktfFbdrslTVRmGk/WzVtrE2eeKCbB0
iqfFxwl6BnZgRdQZ992sXX0iTEzYlUmp74xJoSifuSReSyy7zBxDZEDuSrxsEIe8
tMXVeAsmNVPt4k83SRDY1repLGueLg47Dnv7RTIHcoPH2VpkGQiJBctre5VSDzS9
aUtGeD7T4WLvNww36dT9A4vdWUdin4lSeOrLNJitUF+IweY3xLkFd6nzPVRyoOYK
qYUccLruf8DIvjIPP6fowKycW8i9Kde0rjTdxh18znJI8CjrD/06MUMJdyPX+Ads
1N0kiaITxuOLQenE98iWBuyTpvAXX8zagttsM0DFMsRrWFSTTpY/98JadvBiPDfm
Yb3vzgKjIqfZlP0fJsQpnYNDXrcsf6hnOPUDFCyEi2NdAkm8FWvAbST8Bni6uxTo
FoxPKQWxrshUOziMozZKa/ISF5Zc9dCtVF9ZWNPTAZ/gXzxbT/Mb/vBK063kCV31
3Mfk7VIzxPId9GupjSUBQ4IpnBkih8+rZkw9354RSO0WeP93AwEazDWty74J8ytu
HgRPReRKL5x2GM7TVy0LNIGySej5at3+dIpp3AUrSf6/aL+5dRthsl+U09az/o5d
mlYhDkuLk8IbDqLqY+m3NoySU8nuBTxyTVaHFOFRsHleBvZ9MPaPbCNqFZ8FQa8r
Zi4QhpJYmw596dkoQ5vlqG/asJfYT6ELutc3oZO/N7o27rdb/3gsrda2I0ixLC63
u99iCd0T74jAV17fwX8ozHUc9QmTlhKnZyAt+In+vl+DEyi6uXPEG9US3TUwuK3h
vzZBzPhJsetTVSzV3DZc5yFHXyHMhtNh+L1LbRuNbsmM8ramuHg2vG6Zvbnygn6m
TyajtM9JpYmf1CJ7s7FGAc3sFgIUIEYZxtPffm4rm5/WS7ir5ItnUG77CBhOy2IA
B4AUYgghNzJS3w3aQOpE28ZLPl0bfBNVjZ60HRXTM05mBYWFt/x+yLYcPwWJW/Ok
`protect END_PROTECTED
