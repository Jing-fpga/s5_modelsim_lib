`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9lkstgpNryskktuvANaTI6xvlCe1ubtdAgBCpN2AGuGHkoFkXv1KimawqtJElLwD
Ine2ADuKpaYgqZbQrOvIOHkVxaBPXFLri8xRagZhcUhhsDKnwIIM+DSZuNGlz2rT
QKaICQxx00I1/o1XML7Jg2goECNMJBalyJcZOs0fVY1V2bL3lacvCP63lZ2QIRYR
wiCAzCQkG8MZG7uhAaDbxWNyyGafIzdzY/vrunf6m4wEmLcAUJw3egcfW5BiYe6f
uegFeGeAKE334OhZaYmEq1MpW/cPy2gKvcj22BA74sqoCOJSLa1mATlP0nKMx7np
ohxm9sYGfDuNodDBmMIIv4kQr4JGknwjnaUJGqsrij7CnzscLQRkN3qEgv7YxuS3
3sOoejthHbTPWUFyuqYDXPNltN7dNHhn+Hyr4d/gzd+1VcsiHD5+5E9SBUkJDuTH
EmGWmzSYl6mfgg7lUu4JFb0AygJ7+MHiM0D+PfXkCqZNGL/aa85gyRxUw+BuSLts
VWx1hWRXxQGJ6zEJjXjSqXjRc9/dBJtET691FMRmqHGxQhjd4TGnM1oO/oYeMwkH
hiScrfuHGdRg3d3VnQMk7wLE8zHzQT9NkUgyDRiVbQNQ1qgM4tXe1vSmbmReTFog
JM9+FB+aNB0nQjT4GoU5GK6Hjgq4KKvATeD7e9EiLzrBjCDiielRu65zY91xU2Zc
2K9AGsb2QjwL2VgKk2JBgs4wZRnca/TrUQElI4VIMD1Jb3kMDSEtDRM7SCHwu6BK
vuJLih6uQRqqsjOUzTe1Gg2RW2JbZD3nCvU72cFOfFNYpmgdygeYWxUbn2kydfKB
CL0/dE/WN58WqM9M0hqUq+XwE1L5w+d4SxQWnKRpbsyGUlj2bEYtEBnbwx9xHENj
SGM+1hDZEvPEgFX+NTUyK4LvESaQ6sNL9Sy53HI4svKVSE1u+cyaXVfsgEbjRwP1
Qj4F7qw4sxgQmRi6L0oTTeLQ9VqveCiz4mKZ3giY9ygSwIWUBmgB6aMvgvGFd4X2
Pu0YVvMIJuGnajVqoUHVRFK0zxsulhi5pLPxSWDPk5mIjnDwlZPeyefjkDs6/Iz8
ND9ibHGbL8kjxK+p4Q8HFFL8cMCQhFwYNmmOG3n5X/tXldPs5MyRWJM0wMWloCPf
nAOJQZw9fxOcwb9LQ6luiEu/nJAD+MmcfmF8niuNBfroHuja7vO4yvVjK3O70ffU
UVgUpfeBT5ANRfLN0VTtDenz+CRI+1dzxzPKGxNf3dguFTA3kUGxVECPOzxiDJQK
FnNJKMPirpAukaydy3e1eAvh2N17YFDL/sMQ/i934gShUj743FYrlPO8kpPEV/A4
8pKz/bsQRQ7zmfLdqmh6UegsK5WJzUDWcH8ZX6OnrmkhBTXkxZyr3b6GU/Jo5fDo
2vgMwC4rNmvrbJnViGVplzRhFfZeB7fxdETRFNudW6T6ontAAzVNQSjCuiqRFf4l
Gn3ljnDKg4fUEE0SNjjVa/eMdWDbzqqXKlLG8bB0l9SYhUghqwcpqVdp6Fg90yky
p20N48QJ3EDNNItIuXTKBpL872H2SkvG53UYLszjAZXWkE4nZ0VGTKRWys6y+8xz
jBYJDrCbl2DMI6F1AfxppzyEtnsuW5mzblIYUxuKoujhYBsV67QvLgWn5JvNCjNS
W55XB6arbOqzRNWfjxwEeLUCzUqUy3m54Vtd2Zndnu1Cgq6aFtRBpBONF9oMXPCV
iO9Rlh5Kj97ZFyfsNdfO/YzcZKX2oArU4DO8amMJiFrtsQNUbExi3XdPNkd/L3+3
ydt4Ui/8o8IMroc5cQkmj+X75lM8LgsoMam3FCPb8fSlhBUMU3AQU4vPsVDNmC6T
HlauO9lOJWmNWX8JG22mUzYrXgQZxL4MzyLa8gsxN+7f+kmHsrD9FXddNZdGGHVm
QRJaotPAlm2asuPAlk4IcAD2Z/QJo5lk/9m0CNecE0pRS00AXcJeACAYmWHgZFkA
jQBK5RsrEscq9WuTl0APWw+qCqL6k8eKRxGF6XAas0b7ODIAqOO7M/GrnLC+vrRy
vPehq89kJOqHW19oYaava8ylnXgqYvbMqqlmC01jq/UCNRe6WH4WHHnUHrG0eJAB
vL0XzsVmZw9RcTHzFKer0PPAcPHY3pv1vaHbsgd8MXT+ga7mmyUtAWwpijSQyc9c
qEqDWXzSEijIfoY+9txkqBq2hmRqcdnVXxmJ5oaVxrpqzaa9+5VI3Zgjv2os7hZJ
TxAT/x/h7ieQX8aZBHsDflhRqIoLKJPUiwl7UC8TpCOAAErk0qJbWQxppegJZ9Zc
9s08+YJMK9TQS9kTsoeBz+w9faLN2e4wqpAt0nELSSwST5dzg64fLO6jLmwyQUY6
ujN1AbKcVElrB63QXRbUXtGa+4vMtEln18/XzcQdIVIq4I7N+FWj3jz4mwsmCGRj
JSqRYuSTnioH9y3rhA3xKYaN0llsPlh2cdYoDQnNsr5HoMGxfUAcXwbp1DuwK22o
zSm31DiDy/pVdy79DCT+3GflK0R9VSox0MO2oX/Z3kl+oMx6d899s7XHxkcwoetf
3cf2OAYNhwWafD8oB4hjKFiboisSZx2YyEPRA4iD1VsIyXKjmY5UdRbvuUxSzUbR
q4TpXLfkZlFc4KiD7p7+9zzJrNtSWkZPWL/kcUH9xCNt3JGBe1aFYFo+zWvFCkly
8A0DFErce9Rg0vuL0EkF4m1oGhDMMbOoV+G1eOkidMwiZz+u7tSKCOdA5NnzIOsh
61TbUt8rm0tlvwBU61Y/MxwMny6N1vMVqUioSL68V5vNl28cQSXpkN1qYJvhbyv6
bvOz/33yrleDWuPoIyClyTTArmWQjidNIK/TvCsql7pPin5v/M8uhK3FVKAIbo7h
luEXjQ5oOXEG3P8U7f16PSl9qU/IVOo59+MfMlCF7QzsBRboH8fe42ljqtd1I5yq
i8ST0DqyMqrRAPQ+rC9oNHbe9soHJYaLhgFAKPKFe/pTLlrFKCD4/WPCCTBGnpiF
T/C6Ac9sV0XLoR3KNsXfRauukmXkwIUCPSzHqpHjxr2eF8RPSTOd2Y4TfSaYlNl+
HmKgdno7sw6x/CAROPxeJYiJLvu/jnj7uQk8dYTq+Nz9QzIJ85kUZbcvb/2golgE
AbSb3yso8X26U/2lGxVa74VZLQ5g+qye+38lvBMO+Plry2yFTyXLzHw4zrIZTmv1
9DCZEAGN6dSxdN7gLcNbLKwBDsFfnN9/rwJrNuzICquOEu65uoTZZWA6VE5YNxtL
UmbwUdBexvfkAasPVwYepWXDTSlARjAijdJG1UsqYVyU5fpYMusOCaiQel/rqGxp
YPnLgNo7qvROV7HGdr+N0fvrsvY9b47TmsWI5v5AgrKDtZx0yESmcUbU9N2OqJo3
f1dolZ0Tu0thmImPxPEvCM5jeb3CAlJCEGtviUFjfJrpgULRPmg6dk+kTlLKaubw
dz/bdpaQYgUmssLzaAUn1MFH3KkJ/2DaF2LzmISTK2W/g3/Uh/tJZtIljcq33B3Q
Mlb5eJugr5oSusMU7tLg1nyARzd8mmIFzoetBo6ukFzeM6Y9iHycWk723f/Rj7YB
wQvxFuDemh+RvVx7cyWsG+5I/d9af6fKA4Zc7iO2Sn0J4QmpB08IWSaN0I+T0cZI
kuybVLkZvuT+LOaId4jeruUsv1dZeYa46yNSyR2RVZV/Qy4deBXC3HxZCVSYYVuG
+qLeNxSRQJsuisSh7Z7FIUnJ4ihVgmTFWtURSOm+OH7LHG9EdgIKfAC3xZAGvi8K
j33LfIODCYJDcIl/CjO4H+ahyfjHQW+Gf/qR0CW78Oa6+iIcW/Ws0pFRgkyNX+CE
VJz9ehiRdtQbq6s6MnEYtUVkx+plkUFQ0hVdW7KesliRMRmu9ZAegec+WEXgkT0s
ZL2pCBZMtkTd9plBLX4k0lBFLw9MT1hDke9zVCzeL1jFAqHTe4B323nOR7Cj51s1
V62U+Q9F+VRhhU07imylpHbAnpTu1+DC4MW8Sqbze/EQaGiU2ixED0lNfZ/9Phv3
U92R4U3vG88GdX3QftKmFPhDnmyG/pg/a1pwPTbwk47E0QhtyDtzFWlDNV3j/L3n
JkeDIUP77NajhCHf06mBd2msm5AgGPsBtcb/ctquUSwJe/LYrn/fkbK3D0A4/Tvx
iq2HB6DW5T+ufApJboCcOTvltdkDGZEU49U1V1VSCmO/ZT5xHfy4TzrTz5DwWwZj
eV9HSs7mpgw5S56HSaytX7WEWCkB5pZ9mF8Os6bi66dzmMXei1G+wZp2yq7gAINL
HxnVEIG8QuDpmkz48TS+k1Z3yXylhe367V8qy7tVEsptLa79yV60SSrrhvGhAkn8
UOEMLZKR+5OqLPrSId39FTTkS3hYqVlFcRSmi5fjnqi0Ru3dnE5jHdOEFeUDVSIs
wOzmqhrpnGytn48GTeKRIQ6ZlpjrFNH6FXnPBFFe62syOHIOtfiQo+VgNOMi36rI
0D9XWAa7VGipocJzDpwHLyhyTXJsevI5ZgjyyvbYFQ3n5HNfBjT5fMwJ5breTn7a
4E2THSIV5hes5WvbDwYkLe/WhaV5jMq1l4u65S2eehVToVtegDbfA/hqzfvOnXQG
v5W9D+WmANpxnbVQGsB7Mi5TuQ1DF6AlyTCKbS12dqUDNF3R9xvTZuk0areTXm5T
gup6cQ5ikNX+3RinIrf0lXEkKXqYh3h9gxyXkQwqPQwfiQusncKH1wOLcCxfx2lE
JK7zcTzhVhVENAHwYzgEaVjDD8cpyb9SPL1cIJAKoQ1U2FSN1WmyldPx3Dg53+qL
QcDknjP2wftS6edesb2Te0htUPxEA2xX/ZajMR4T+3cE+wbBoZyR4SsoGr4UTtLt
mXCJSPeYnqYaDPXxlA62fwH/K9Kb6CNkt1PtMFKpq4bFIYN9q7jE7HDhCTkZguSN
k/TPNICmDMFwSsbjmVMQnOg7z7uLFEqwUVuYDCM3hq6FRIphafAr+X6Gt67F3mDc
fuL2k+92eysR1lb+XuAm84IzD6HvZYgpS8wsJ9gdL7zZvjc/3Jd4cvh37+QCKDoD
Q0F7BiMiR+KWJeqLdb80rM3BSLcRKFodeGDvJRE2s1+X0lJIyYd2+QXdZfHDoRRP
pOAxi7MO1Cg985aDYEcQ2nsKwFuZBrB2MCbArY85Nm0WPfOAAXBIQYHkpmcGIsYR
T+Mg0TrItIIUkFBur+L33V9hkEWejhH8OialyLprlS7IOG0Sgz2QLBtjl8QLpXq9
xtAEIiPZtsAZcSxKdchWCucCKKRN9JorpmfAwmGxSFsWf2WBw79zM4xIVp4ZPTAo
UIVNwG3IqH3jWLfYoqRb5rzV3SBfQc5JT12xUz6/hPBUROL87trfwgbCurNP4j8K
hIP9w6EKOThnpULIqN6QuauB4gRcyfDra5R4kWWivAZ0TDkv5xv6tcw6OIKLykes
VbRGuI4PGv6fbZdvHmkF47bw5vYofbAUcO1Dyyl7L07tmFF8vAey6ox5UcQH+k88
ehhM/PZBYfrQwQgsfm6kmspXmSHcIR2bShZlOORL0mTkl7GH0sn3Hta4CK1seEoG
MX4LX60fUM0/TLaCCq8VuvxOl9rQgLXZA2HrLA+95tPgDSUudpVDQyaAcLD1QiAI
cOtRm2gpuVCSdqQ1UHEsjXsUidkdl4235A33/pnTLWUovnn2oCfUpX6Wdf2h64/V
XnEHj7Pmhpo+yJu9ifK8GbvaVAwU0vTJu+skDpSwloaUkDuEo2iGGfny4aG1QxBu
PPGw1rbOKRBaGFjatrmR62CL+gdg5/ZNi1qIHW5zvfk7jTNFmdKsBPSUER6Ubsf3
FXJapGQEzPM9BiOCYK4Y8mDGPi6V2cs9EWYolUruHXZzk6fhCzjlL2V4+Fp5onXc
GG7y7icb9UBoOFk5686VRbsKlf974ZPwwWekMJv+fmpHVNV+9Q/V1izBBuhlR9wm
8ev8J43Y5TZ7p2omAEJi3rDpiCISGl8eGlJzocox3LrQuEJRJonYf3HAXBBI9RCs
oIC5bKbHY17ZgWbLQUwSBxW0o9WMRQAn/kx6JKiE0PPr1jxlz3uhL8TmKK32XFNf
xrhy0y/EDjh5mRw2uw4SXc2U0YA5dymdSxGTN7FxJmAPw/zLqJxAUGMff//hpsrv
jhqnpVLw8dU/eH6JpwxuQmVfyRX0hBmN5dviXEeOHEqwIbYPpTNrzy3c7GfyZgq8
AqzRjLj1HlG9Wbs2iBByVRwBiXNvbljDwF8MCtE0PItVKDJp5ZzgbUHPHBD90F1X
6slmAQrxv3ZdJgJIeFFa6vPu97tsCeCUmTKiDsyvy3/SBfKNkPvoW2TkffaPrTTJ
sakqctqhff500q/Nc1Ku41w+5Joxm7zXUlOQH931FechJaVLCCV1JIhJyYvNafdr
GHlY5obt0t04Y4MDXKM4AYIpYOmpCOS7bm6bI5fNDm/AQrEhufdeNF6UCBUhtJiV
FSr4YRn9AFFjh237xJm8UvPzlKuQQl/IXZkcL5zwINVrnIcbcoNN4XE1j1gkkHt2
vr/D4BVeSdXjRKYNHpmr9Q6BnKc0ybo+5ERJBsdt+Ot0lqbooQWQr+AqmhUH4ib5
s33JuZTrisfbk62EUROuCAb1nGdagLg2SAlvKZHVt/YDh7hVfCZaXkr429CWmwBf
+MJK0N9P9jG5aBNXMP1TlGpD3y6XSJ/TlSXjgqemYZR7Y7Pzl2jsVBYKcPZ9KmPd
ljdG2XWB2WuIwyJ4IgCbj8vdbc2zp+nPVhDxoNzaIDNmkJJlIpSFeYIxdE2Z+2fF
iWEqmLuWtUNgnwNqrb+6tqC+rVlFbSEty92JXxAgD/DeHSk5r51nUyHiIiIbdxGD
y71/6rgJsLAm//eFVpQMdHb59YXr3IRDezjYZsUZYtaI0E+7yQVB7Z4n+Tn4/7jM
5Le2XuSorJKS1sqNrwS8gUoXHr7vv41UV/nhboPu+fMNAsZNbjp/1OYnMMSNhPvq
YZU+/9kFMjuNeuZRsEvqnL0n73JceuEyk6S7HRiwTJqt833t744eacxdxd8W8NTz
ll72dRu/gGT+AiDl9pEGa00G5VvasOSAKpjhcXqzIXKyZyXpb8LL3fvVYhhqJMlc
FPpclQdSwHnKzY6I+8AoI5gQ2vLM7GS5OG6ODJ/Yb1ZVq/c/CEqJW1G9EJMWI18P
`protect END_PROTECTED
