`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/fYlCl73DSpmpgAGYT7sJCXRYC+lF8z818lK06LAy7sIthnimhrQLEUeXZZ6wVfw
4XjgpGgV4fW9wnNUJqsvZf/V5pqQ+a+r36ONNw4kesdnAmRsnki9G8c3QG3WF8Zo
NKDQnVztC1J4l+xHx7c47fQGjIBGJR+wlCXK64nBqqExodYdDRVqHZ25v/dOexe9
/GbkNyfv6jobnHBcgZZT4snnYRKlLA6G/miT9pKYKO2q1VL1f1FZ89Mf2iH2w0qb
7L1PiTTFFSYSiG7RctvQvA7TtjBG6EFOhOTu2+SAC8j9mGIdfqWpwDTjJ/5NCZDi
q1gwZVhrHfbS53G1FV35ut/QL+IMaFC5jjyjuSwmkSN3zncHzNau0kLhRqsaoyz1
tAoBwO1PIswVwbFXuzMsl49IRukjBAbFaBayS93+a8iLzfXT3ekP69K7egJDXZIm
MMQB9XumXqq9+pNBnnaH89Q4glc0XehEG3mL3HhhVoxaM9xdyL2GEKsN0mQvJOM3
KNrHU5XQwIKBbj3+ovOtb+sWjCD4Gz57KB9EhPs2qObgukpY5V0wI0SHhzXDo7MI
J7pEAeg+O9+A6/PbHqU8/i3SEgkxphbuH3WEK9UGE1R418U9l5Mn+pqGFctVbMQ/
wjou2rrgAgizV6v51VgtJmYcgDPSN8DSnlrHGhjzKuFadeKigE1dPQi5Fp/0Je9j
IKoo2Cj4csBFPClAKL6fTte434FEhaDGqo1eMIbDOTwe3Ny2+eSOw2SDpmBP+Ips
nBMqsThGMMtyzDtAQDlnrFXDayixjYedR8qf3f/ormEdRxESNI7vw0KZN+a9VUu5
IstLMF5Np1rxgXNdykIE2LqNxpfLEvYvo9At5bo56nVebzMv8oV9SYctJAVMf/vf
YVyYJ64HIo0LgMql6YVShqb5R+YeJfzhHvkt4hRQEOlNspzA4OMHE+YowZJvO584
Rl/2DKdxKuROudJAEN2WI3DtlcUUEo1xQ2diwt6+AswUBN/PfrHqjxy6GrN7lBFx
TiHwaeHqx8EQmGedkum5zLYCpbVLG6VeA4V7Wrr02szEOebVp2Ib6hWX7+LERKFj
N1HyndJ8H151qC49YqVXrQKIl89qPTCZ58sAl1hNURRhd1nk5B+yFOjANo/FCr3Y
LPJd/doWMijah5sSmf7ZefwlzamXc3HPNzMqx0QLHp5MTgE8DRnXkT06oUG8TEih
LAvpK2dUGYP8MNAHVXmSN2T1ms3k2m0cm4S4/yUyrG7Hie0a8vfaXjdTdqma50fT
u63/Xf3p/KU0sPNgefOlVjTY0E7OBiOl9Rkpqu3VykcJtrVA0g4dYKQEF72qM+mp
boa7VtedEz7cxTD9xuMM1KPzcNJpMVCaBnsi+gaqKfUZ58wuQ1t0AO+iqXXa336y
DJGjaK2aguTd09/4OQnHeHopC3oObMX8hPiINIRLMgFkclCw8xu0iDhGWU/owQAy
mw1kLKWTOI3PXO+IRs8QUJ16osA+QrJd1NXvDYtoQHg3VFjPVkMz/JJJ8Af39eLa
bsKCY4nl443FdC/R2IVWyDSq4axadOR/7sVzO7HSD3YX7wxe7B1JbUNPeanaL3wl
pS1CfBbibdt+ZfmCFwRLQSKbCznjsDISsCpTSSYU2JGuJwFlxacKawEymt7jsJzq
gkQ5DlkZgnL4Pd2b6J/9wQ1YVOPzwJ4kDtYK8MRlUplNcisp/YD0aUHdkKlSzIwF
qKUaBK0stNMKa9CLM3QC1S3NAL+9xSh/w53aheeJl1g9q+AZlWP9rQf0QdNSdf6h
`protect END_PROTECTED
