`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tqMSVC1GNrhGwA+/1Du7EWqfzKji+F3bSrRHRRGmQLmCfAbOaT832UtSR6hZP3+D
TOZ/rwu2kwtDAgePeyRc2By0SuSDw244qGR/XKq7gcOlb1RlV0abgwpke0bh5LEs
u31Il+c9840GWgupIUdKnjXP1EJaylfgVdA1mNHKkAKKsm6eodQxpSN7wRz/Kf0H
hvDFwKWiL2ILVRcEG6CI3pNYJVmTfGirlOllF6FBGM8UhyYOpOLo4KAFKojVUB/g
fXWHor7Mq6YEn22B8Ex1fFiMqYuqHCs5GGKfFLOPMAg3XB0LZzbpzAwiLRsINtMq
RgNpecYyLUZBh32euVlY6uuWjvuljTL1/US8oXk1gczQPqfk1F8c4Yx5NDNZmQYZ
kOZAaP1YO52WhAB8NDOP8k5P/sXustR3BuMiDrOC+zAIaFghQ05Mv7UqhOvpXLdw
7POxxHap5kZ4q/Ms9is66QLmS43SffHEJs/Txlbcltzb8sGV0JuwQPPbyBoLDV2a
0o+CpFkqS2S8zMbfe7bM/ry1/1bzU5MOMpfrGnQx7mvGAkKCZ7X+wsC5lOygtavp
kwkyobUujLEbPOB2w8ssFg4ukWr6BbvndI9/z1mgwHhZcWArYaJ24C4MZuTxA7il
p7lkctxx4ZQFS87eQ6tKbO7k8+Xck2LFHs9O7mrYj8tU+//gFDT6pHdcQxvO1+x8
10ixzL09q+DY28PM6X76suZpU3+ywU3vHRKsIBlKjdgWp5c7aO604/M5RY0PbbHT
afNmkZpdS3uxRhXmgvNi7SpAHu2RhQ4ncURwDYFjU7tJ4fulbrtKexWg98dfXHAc
h9FkK9+qmivG0bfPmu/zg+SywgKl8GnwdC29xCNdVYCSRpEuY6jpCQrhoviluf3e
0l/ZA6JSsE9vXe25y6yne21VtpPFJcV2CPK1pb4FlGcvMp+YYT5USn6oJsGz5MPJ
pNpQL6t+dhnjw72lkp32SKpoPwcrM9F7eVxNm34maTDYudJD/ZuySO3NCiuj0q3j
M5QawXMr3xxoZeK5Es8ccmq0fAC+kLJxxFffQXpynjajorZWfDRC0lEFE7zYrcI7
1BWPskUIZHywY0h2gq3Bp9gQ4j4d2gmHt6GeMPU/FBGxltO49yY7PLToecgaoIG7
EIn9Uhqd8tnebIXMGbAQzqZGSJ3ZTjW7AT9u6HMLyDoLO7mi/OwIT8FpTeBLxDBl
MC6M688Ntj+pOHNjkyIDbzRE+Wu6W9iGjIr//M+HFibovycxDZPT8wPgr5dCvxBk
abXehV1JNws9CswE7ejtAeJAswOYvI38XyuWYn+jcrvmoF9uhb6VFVTVOGOJK+dW
iJk1f+f1briUD/fplePnWBd2AT5m+8tieBUvQ3XK75E=
`protect END_PROTECTED
