`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u0li0RP5j4FTE+s04VKXKALQxICthcFLhHOJlo82shIXiL97u+RllEk3DSWs+AEv
EQ1LCtjL+4zgrqhxm3+wMmsCWM+8VTqO+lFis2uO1zDCPKPPbS6H8jdHAvJEuaK0
S7F00EOGev4c2eGxt4zXMXjF9rvdWifOk+IdqtKR5mdvp+mEG1uAA8tNyZChNRJh
ApvGTXDCL8j63mjXxg6hR2xTw/XBE4r9kA6YOjUzYmPhMgF5AORLj3JxCdVYoMd1
tlpXsn+tjTAI61o+A0C0ZU5vFJUesNdI8wm5V3DU2n4uwddFeFMhTL/JjZtJ9rcf
4k6Z9Gjxlj2PS4YyOHrtn6Gpmf5kRzSG/7I4ZaetDR4LHOeY59kwFqjxS2hQcl2S
u9tOd3JEUD3e+TkIorb6jdF4TB3OXvVG5zd7/XBUQgjBK9MaOTQBa5ckRhKR9Ebx
Wsxtf4SZa3srOuApBhpJBe3LfERcJqZ9hvBbh7upsdTE/O5cPDpntN+cduTYutri
uIlQjQbobeQmkN1bCukYUfpcH7BNHWbPCnUHup3iEBmz504kMeTaVDs5MNTfs2Vu
6nCiROfQiaP+YY/IOwqN/0tN3tVwMmYcrqVfoKE57dFstlHRmJB2G9Ylrr2jBo8T
uhkqUNxpxhZVCd1gA/bxuCy2/9SNplTbfOlrU3YjcCCS1LPoivO3JsXJgve/3zJh
8rN/9vAkonDVb2TgwFj4CRdFcJbSBPelrYH7DobvLddJTm3hoG9/9a7B6HYC3Oy7
Ace9T5/T+Z76T77sCl9FAnMWDBGDLw2kxYI2aYE2DbDZYi1XRsUQs60fAPtKbCer
kJLu5DHWWMUd0uZSWtTCeJCc3KxuBDhlGP3kkpJtSqEOAc7EDkeV+oXuMdLlMXbj
cpNYLQZM4N/vrhD6oirBijZXzhKMAYsgOksfZFoW4vwVuhwhnRmdEhHra38SYJv0
ufLYYKb1cztI0qFxZBaWdixLixStj80Rcr9w8zV6JaKR0r4ZS9lEaCtHwRKI/NT2
1QH0ZXI7Z21ybrdvNT/IxIiZ2UiWzjTgQVjncQiqR5PjIzKW1MEHQRN6TUwy2Q6w
JRFNqlcfO+y+4UDQH+HztYuORmYagOuVheYXLxrV64DPT0RY1NlOMkD1j+B9DNoZ
K2VmTjaV/45k1xPutFnP9EOnkfQeA+4k54cW58Ggo9iw0FepHzXobidv8zb7ClDJ
tE2fcyXLXBTzbdr0yphp+qETzPC+PreMyp1+caI6t0mwVIvo3kgZ3e51MfGHj+Jw
4y69gfnt08Cul5rowdBrMD5qY06u2UgFKtzfH5VYtpqq3ac6Z6V3v7rzFYc09cQn
aiv3Ncmk1YuqhOZEJw3Oll3yHxQFWUSvl8MqH8rRiB+ofq/4sqLBePzXe8kiDnfa
BoVUTRiEXsgnS04cPVDil5gdLN2t5XNL/8FSPit5y0DXVs8amjEJEA3q77DwFJkE
vVV0NbAJmVUcaGUjH6+9LW0ZIdxHROy0DO/8pyqoy1BhlxphBJLRhkYIqUrklA6V
u1Kvnsmy1IGqDi0JMUBNppMmuP57jZniBu/2xLQiSFVVJrG1EwSNYd8QYGRQN9oM
3VpKeBVu/S3vHCQSj22Aua6+jlspJdt/bJDkmh4qCXZwsv+9SndYyNt8w1RNMS7W
TLsdblG12s4K5wQLUiwHCVHY0HuMq4GfDhuKs1NeFPx10VwYOx1Khpr+xfBw3SHv
4T84qKlE9e9WMQAhtYgpeV6sDbdaEweJX7TDOdbup/f9DyUliz0BynDrXGn9jYoB
+oxSnuGI06JUaOQMzZXryX4Rxd+1Jq0B58T/HHMZ/mf/K8z+xRDpJD/PgAXFJGR/
HBhmTf9OIpEp921IX5MZzLABaUsAljFuILHyuC6nk6pVIREtheRRELmtdaT9Pa56
jTiC+cATTHi8xnESPLso4c2TcyZ2LuJ4tSPOTfgcGIA/Vx5WBtYrycMek629wpd6
7zOI0GcJ1eQh1zz75OgxqgzXXxrZspSiWNoAJkbptb8r6KZwGZYk6c6x2bMgX/lm
j7R28eGRdT8cDIZvovmcCoviaHiKoBsixPEwjoa9H1TzeV2s6qfhNcNBTYHT7alx
916pBaJA/hWdEYR1zE37MnGJi7USY023inh8qitQdmE+s8ybSvyj7YNaicbi9ag7
Djefa9YWh8zi8XfhvqDJ3KXr2r+6U2h+Zh3N10+9dAORGA5O5QxoxVVmbf4nCEOn
UzRF3II09ptVGSlpHHNIhAsRwerQ6hF32oQiqKAOxF1GaCvv/+uL/p3xKB+vba1Z
xt+5qZvRbNQeyR9p4Ws9/ytFyQsNm/kDvJqYPc68BOg4fK2TnWtmEzrhrhMTeO23
KGs3apgs0cm+ZRGajkPtdgXjS3SpVZx2R7BtVFGcdvFJUjg/PAcWATDrQ309EvOF
BlrnNY8oC6LIJzWB/prrn9sFjQzciefPHED6ChI0dxIJRGkaFXTTgSctfaUQcrjH
JCxCbxrbUbXkU33WU2vnm7KUDjugR3dVU9OS/x0/T7GzBeDOfFPLFF18bDKV6OA6
dakaBnByIvpZu+2Tn2nBdYgch/z0ubR6yRfqJp8g5BPz53kgVU4IiDdPKSf0OAuT
bnVzlKJ8M7H0p75aFADeA7W5XaLGgrLcOSCYfWd4MGmKA65aZf0HVYvMLpQFZf6w
uKEggK4rQjcnmAckagvebJUuh0s5HVxj4/arpOOO5PCdg0gV0iwuvtHRDCDyEXps
gsqThai544pyo1mwbHPd6yDwncShnSl7gNe/V7ONGQkuJSlxl93QAxS3zoErDF78
SRjibOfV8Y4jB5+j4cjsb4cBtmPtJQ/mKEZjM0LNSa1N0lsk3VZYp0jCcH2S+Xmk
bA3U6qylF8XfNtzc7vTXNY69wdSWaeX9a6E5FmznqIvxL4BaTlG0+j8OhxEZpePS
Q3xNSqJc0ufANwUx1n/gogA68L1aJW6dN6USCEUkPz8z/lAvpetRXgkYUF1U1BuE
S3iDeI+8miRw87GIgK3SAndaShRYiD0uhtH9A+1ucGt/oQ4Q6dwIKd1i/DpVXJQx
FnfAqetLacSx6utbQBEa4HOkwGAbdCBWbrxWR0MjgVGxFxKl7pBJuQSlN1LUfHAK
Mk2Gj3FLfInC5J69Vw9uoAxYaVZzYSANhiWx062S+h9GOwvbRVJ9Ls2ReRcfNZ8d
MUb7+BtUSSJjaHLNUx8ALFZt+w3rwQPQGPATBW5pSRQ/1KG02Nql7ANZZtPZqAaD
6h2jUesaUROWIEfBJac55ie4JiXoadOlybtwOrZdl6X/iqY6htUYI61SddNYSfRh
I3prCQ7QrbymKxEVy/Kjt4DUbmcw/iScQb/qmJOnhLhyZNWcNk7KpnaN6dhUmYrE
g848b80toHBQjmLxcc3mjixi1iI66hUtp3DpT95KOWWeIiGBG9BsgFQzb68xwO4F
/LPrQFUuOvuQOuwl7kOQ4UNAQNHw/ck2gfEiEJQvrMgQdXBsRU7urWzsgFvzlrze
PTgmxYEca75LYOCa5sHr40D2PO07PIPQnekXgqtnao4lN3m8Y+F+2DsC4f+EqvTr
inS4F6P9IU+/B/0362aotD00kAEA6X7rpKUBkrcYafEN+gfs4J/vkCIZgw4g9IFG
ub1+SR1Du0AgMC6JYnmgjZ75ue9k/MvlHsMSI5fCIw1W5MO+MdowfP0j1vil+nXM
7qMswW8+LghLEU4RjYiZEhnmJzL2EEZdGsiQT4JEg/TRcQOSwvnAa7f/Z3pGwLAP
O9IA5MmUQQXkOB/4xDfwcmORTFQXr3GgjkNIRuW4eoVeqFjyawVMb8G5vi2gcHke
lXLdjYm4gTK7SKnnXEO6fjE9m4mjxMQRbt11dkJifJz1Ms2h9BlLQSk7ODnKbqBy
zQZiU3rxpZjHw/ctaMjLOa3hUM8Lm4XGfOsx8jFlRTGeW/PwyknH2Q96CfLVwoPA
cAjyO+lyvpYpdQG+9gAvISHrCEpa7TL1DRkMRrArYiUSz29+C7wuzSQrML8DxWry
Jcw0V8qfZ9/hzDhFMgSKY0v3iKkih5jw+vapFI704x71kQVeB2zY7indeuM5TNMb
V7cYe1GcqYNnGX2u3lFk8hoL8rrQ5AiZfiMkJu919Z6ar8Kl/p8VKtXYUc+sqNvR
xKKTUYtz2cIMEEtkVA09qOblG+zo6LGZDnVsSHhtouC0027ZP7WL/FOT8ZfLqEpo
zq6hH5Y86DF5+e6YPJkUzpD+6BSD82I0bkbq8bbPW47voEeoBuQtlgIoYo3xcPSM
mOTG+NAgZMv7CRL9CAxIRfcJovwXYofXPeIhACKmKDhUoLFEr6NYSHDtgOFOe+tg
MfiRltepAAIUo3LVu+wLuQZSooEWpNFvjswv2vU3sJlzco5J+VcUOmjQeOcwWvFS
yvKJ9I+9X/HmAB0DulMXd/aMyhEmCCOnGtLYXwilggPMJUulDkX8+/DfXD98ZqEN
XXLYYNDH15bfFPyTyM+sem3ddya/0VwtNYWnJs+c61dXSYArvRaDtiKa2Ro3b6e/
WIISBYL2g4DeQRZRx80hZ3EsG6Wwv6GHXGr9vWJZccHZMzpnsJTS3DUJI9NyM3VY
zLRPHxQXcS2Dy3dbLrtFiCP9HKfKqmHf7nREVHGC+XQZDuDk7/GNwPSrX0fp90Da
lqLqC8Ny0XbfswTeqk/CHkAI5ASnw9f1LiZxVL2308STIsGxJ4e5jnN7pDJab33S
`protect END_PROTECTED
