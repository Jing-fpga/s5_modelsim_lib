`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6haenX7JK+Huk3FmUgk2KyLIRmR+ITqxl5QKdImTrFDUVFQkiTY+dZOg3hVjtA61
7FjfwMZCuDJJIwahFo5W1Lm0VCVp2hO1uEfaSsX6VSy1ntW7kgMIQ2G50TTs6jI8
PY2R4y4MQTjm6KLvE/6f3aFfQDS+dYXYyvZfV/S9xsfsHg19BLnQPBNHcX1WbC2n
/ChwRkB0Vt/Ky00Elwkfgkwb8laoWtGYpwPhHZo8MThMmEaSTCCrlTX+e2vmhgT0
ed7mdvb4bB/TxCW0KxPPOYh6Pf/xIhwQgmcdVN1n02gelQSWRFnlX54Sj+EN4tfn
FmB8tVWzYxqKEb+glZQxRjAuh4dH6yxHNVfFvcM7J0zrFYRkN86pTv3HknXREfrs
w99FUbQJLCLZ4DZX7ir/YhVEfL6gTwUxaNF1KPSeMK6ibmsruS32LKH6fV4krZz9
OVn1m83qeRzYekyi610b5ezlePw4GRaF9Y6pSx39NIiDDWJw+g0t0FWFLwv7BAqL
nBTRGvzB5UzdanpAHtFrCf+qHASGfqgxGSbK1ONMXBm8aCdP5IjkkVPCeSHec3Up
RI9eBi1ME99S2SdtZuNhFTYs4kBRt10LpupqTXxulO9bSiPCgyuVt6vUjIh+affV
A9ac/8V7IYBgd6XVhCpyKnARMael2CwfRm73chWgmh+T19aD7NVyVuTiQt5DOiad
B3WC2nAVuWoUmAF5u5LuPHfcNcifQrM1MN7ADmisAkcznbgwOmT4p4wO3EIAeW8J
FWcYYSCmDDzKqnu2KDFHcFJ5Pap8EgNHB+T5I+dUKPrsPbzAhTAfDJ2brEXQ7Kbs
IwvM7B/EEQt+Xg07N9E9essfcdboC+SZ8/ehZbOBe81QX4cnntMMBoBjoXXY2hJM
CuBOmU+2X2WmHC4QSMj63UHeatONS5irju5UzljdW3GeZ8L3TOPFWZs7h4pxWKCY
MOWnCk65BLNUli0Ime0IqnSidlE7c1k+71qkG1DKdO0hL9Fkdgam6uWnfrM8WtAe
pu4X2OqhWaStfTEnHmus56vMzRUgb1TzByqi5lTrqhiyTQ/Z8Zstr//lSaxmpnY1
ALR6jXl+mU0XdQdoSMaeNVt6KzXt2LkhSlAOnJeA3fQyzy4KcBujVSPXcasC8A7g
zw02Ga0aza9GCN1dGoCpqcWgZZiTkij3wQHuEO5GfOOoU5/1TMnvm02IUxkMw0mA
ogCWldAa5fGxJ32yQockVbef/t+qgwV2U7ORpI+y5J8jXZ22jXDLxbn+HnCSsjvQ
IkDlFjJZjzn/1241lffwX7oFqjDR9+VIsD0/NvrKXr6xsp4c9onpaoEHl6cYVNSh
0VgL7X5M6f+OKM0QV/Z4wNu6D8ndGqDluKO0m/4v1m7JCjgP+oIuRIzhW8o1CW6x
Z7gJqVDcP2QyliGI4MLgcUJ0VczB9zO0XrKiqxExc/45SFKC3ip+oXbYebcWhQ2B
+6+aEbniN823SfH8RRNOVU+yYXMBfn/iNC9KVgvyDwCJyHQVqy4lrytnvewbWqg3
yBnWBWMzzcwuL/xGMn+jsV0DW5rGSbsvWyVGdagiZRCglK+9wWfVG8x7pYxWDgWx
aKWxtvdxsiqui847rA2AOu/61Zs7BmtbXGcrBMc46W3kX5H195LNhujbDvo9++pd
TcPBNQZ/uG95jC3BZpiiUzy7edKORw2az4OcjTwiqdcDOKFjonm1in74afqR1RG6
nERTBa/GZ8PKuosI9AZDCk9gvL5YzJZyZRoYKIQ1tObV9bpQ2Jwlf3qM0jFU/8Xz
AUo9VhgWtfIrrNHIx6cFroesrVBLAGnJTJuLdfDkzr820R5oCbskYwbNKLctbDCf
XkrnRxRsAuLynDOcW9/3jg1YkChcrg7d+iMyS9xS06r192jnCW27JULqfxgWWhSv
z3odIM8FwcwGfHxGvDaKG0PZQbjxMKhjg+91A3w0vPmGvUC03gX8qf+8lq1PzHBq
kDs79kz+QlXUdqmA1Nslub3igF55zb9I3Vq/wc+ig1Zajf9jIJF8EfugAT4yxLQP
0FDqQiwxfHVwmjL1dW9obLCIYFzhevi6a/01EVxxq2LjIKaerZ0ESgwjtU0vwNtL
9/th/zGWvg4OY4yoO1CeZATEdzwG2EVihUEiwWBEI1MwY1nJq/ISFuliKHP7jY2a
r/emciOp9R7HJslpJBICYg4AfdD7DoS0M1Q1jNFpsnXWAQm3p7qZ5SvBNhl8XSxT
wFq+vYXUsLTGQrisMxR61wlTJ9MdkasO6uzPy+FUQio++eZzgv0sAP/L/2q7NUa7
AN4w5Yjv0gYyf7gUAFqV2A==
`protect END_PROTECTED
