`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3sBXiDpV/Mbb67nSOkkWbsLGxaJ75pheTgngpHg0dzrmDol62xWesuq21uUX37ih
fY8b0t0CXlIgB3vtZJscfZ6cJusi3N1/oSgzpoZvSSxidQ31QmlKiOjTPmbNzuBk
mhYdfzsfZR3xLZjOGOLo+6zWGSZCREtM5UWqzb/F8zixTj8YVUwJ3zZE14onXeyu
1szvnFWsG+hyug30e6V9OXPc4tMMlj1OfZhw0HWPOaCFvnrkOLyhuopM3eUY3vzr
RU3zjaxCy+sjta4T7n7U/gUS0xLq65iP2VbZWIlN1vjul93JiGUR1kWhArPtNbP5
dCmw5Buq7hX/BzU/LE5/d4NL1UGn5YJcrnM/xsLqJy3/VUBMiQSUQWsfaQPOFiAH
mikcUSXbO6EhJXWCT3NW7+uN5+FpUJA70N6N7y2IfX4+7li1aR2RXs5ef2JCRnom
zwi/WrY1fsV5PrrhU5oVsBv3x1JeWQQe6GSPQ0t3vGaQYXE/dddrym60J0zWRWuS
zbyRkelw/kFvBTIrALvBSe41onACHE5t8c7AZPBNaTSb1T01R3QNHX1KeKDcM9H5
U7r4RTYI33y0txucgv9eSZmouHm8Y1PWCJH0MmfmPZHPd7c3+7VvbzQ+AviYuj8m
elIoPacZCarEPGpkZ5MTeGEPPTEuFTcbIDZoAg0wrK47pl4bP32znz/TOPgv+bfp
FvBnzsybbBS30RTm0Z/NfbLW+cNBHy+JE8YmRfcRKRdAeFFA3NHMIYDliAPa2Qvu
GNhb7VQIewffvaWm455IC7OS5qUXI8LzZ3wGWqp8Bh4CQE12nyALGrUDtecTieBp
rM4sIN6yl4kZiLVbqXSaiwQ5W5mSrvOn4/v47PBSTamr3BSwVC0/kkcWaybULClK
M/BhzcTu/7QXPTehj8wLNsTxbjA17OGjkWxQe1x5+54eHRvR3ggfVAWLnHrY1Jr+
KWsRnB/Oq1/opL+C0nViMxxLL/idDprT4JaRENt/U6HuiodayGlL+5t748NvI85r
2VQszZ6Xug/GZek0SbIcOmuxqrsIyf7kGdmDcOjdvKYPwzWV3wuadn/+yR9Yt5bf
d2bRNahhoPfUqGu5UD2OogoyR4aKEdptlpvHKqsloVMtDptTp/g4UTMjYEuZf347
rwTlcHzsfVP060lfuKvMLCdZV5oImYDoTvM57GiC1MPcTyiZTafqCbBGv78h313p
4bGfBQWtMUX8y+L9ncONcPWlLA2z3sULbjO5ZrOLpWdj+zrItP/WKkgB1kZkJm/O
Emw8iMrOeXL5Pnc3zuLlU+wC2GJl1yysRHAhg2xQn2i3N6i8Rbblm10rGUykPYRE
R7IeKtKD6bhunkds6ODTMgsadn1YE82eseqzFKY/VS1myyQL3cZbadvJLpQzYG2L
bjJUHU1cFxp23ryR0Zzjov8LW2iJ7TU5u/rsdW7F4THNOhVd/aC8rGW6RPXMwyCz
RnpxYFCUB709QIe+/sWHGOT1KHBo579I3jiVoifj2cIfr350nmG0y5wnEJtmTJ+/
mHbThzPRGTe5ce9RXciV6wFEnfGQexuLLQ6fGPKlx1vOa9EhAYtMR6fVXYhk6KMT
TC2FAp8NkQz5jxXtPRLZazS1K0LLMAk6BOxBm6w3KCwFKUq6Q7Iyta/dLjuRaKX/
9pAUYKAtalQdCmUuTwnQ5I2iRFAR4wrgInUIGOAV8jTTu5QR+m+KS7xNEttOiRB+
ROJUTo9BWcimYr+y8Ex3ksFDccyiSLUxq4dh+Pc0e3gvmES0GP5FU4dVqxKdMMcr
2JwqN3yRyYG8ivhGFbFpeefK4d6SgBz6Zchw94kB2h4R3xfIs4aqoIZOks0Z8T6s
ncgvL4AcVVrUhtLYmfvOZYxqrf7jgWe/ObMzpwSeQXk/9OQSu3xXaK/wxMRmq1Ki
mJuqAbqxJtqQC7XMH66ZgxlCoTRCJlSHLr6+cy6nleErp4F1YaH3UZ0KCjmuzIUK
kiYk9Kqf7S+h2rv4ydIQP6izGnqggVyXtG0m/7BaOG0Ufvh7gS4zj9ewKPU4SeXX
LV7EZhVKROiDiyE6+x0miSab0QmIAD8yqTa4IiiI1i8HDZpdsKgERk1QCztC/Kpy
j4Xxe70jwuZFWkGCHgKxMVzbd+RgUj1M2BnX8UE40qKW01DY4qYDqEE0RTTy88AF
kpR3RpY3oPwqlbmgktnOUYm6px7t9cMtEDLxsSAUDsRtggNoxzHsxZkj8Wf7fNIM
XduRe9O3X/6yuexgS1G+X3C8pAXkk9qO0sVuCrNU+MkGzdg5FajpLGIMKt4DPhjA
4aYvKkN7MKuG817T7TCrJkyG2Y8R9GMpRxyqpS2KA5MbozUCXSGrylPugBdbtLg9
HodVRhB2LxuNBYHwPJCB3KMBR+s+3ZAAG4mn708DZbNPkqFnJhkem8ct+StnhpBX
5Np73RuizXfgJhd3PqtS//oZUJiP4HrtENordPMr3p+NISBLngr5ojYqh4Ky63rq
xIQftD6Ll5pG9q6P9vVwRBWo+4XOKFVWWTPjrCXOav94JzduwyEkg09EeltyiWgC
gBayg1xJkQb6VPWQu9dUmvxOuZSzrSxgyk6djnEHpjp3EyaV25Ms8tZ4c1qUADsj
MqMysZ2cHuf54lCscAG0uRqWAb7CQWUxOxee2HGRrWdHfkXNFo1KeTUT9FukyENC
uceAjVi3dOk2zmbdteW2d5PBmDQUxWV4XPJM97e9RqKfOvKWqHFS8usGiBtHTAr9
lS8Ll4hCApE5gzdXS1kX0vcuQjzINjcoSWavhc4V+vyn5j6S2xwKPr6LLSW2+yd3
0npSjiCY6n20ohVfJ7Jk4fNokz9W9DU2+2dWJDHcHWGdgNnmclxL6Gx1RjPgkBrC
AKUev5gu77ax2e4JsAUCVf9qbSidnlpjd3npvocTd0Kainj6mASc3ZO+tehtp4Ki
MU+1nBp+3QOdcV4PR3xx04+HCaNoBv/IJ9Z4YjSrOhxH80rrpn4zLsXiNxtNC4JN
4GaNwGq/5PLR/D5Q4YgoGBvyOYbLoRu6EDfGws7DM1mAHU+1iy94SHCxuL7hG+kW
QAWLIR69uVOOwN5YdBz9sxQwGq5LmomvrshKER5GAoAumfVaaswVY2oKhshvKtAj
jr4jMKRuK32rnjlZpumHaRUliGaqZ+tXtG/uuQoWdXi1y5snm1Hv8XsVhL/ohoxo
M6JDwsBVLqmMq1ixZ/cW77ysvWp70WFhEHvb7IJ08njJIyNpdm61/hXit16G8W/s
Kw1uCyQdksGq9lCCbE1stPcW9gPwlsJ/6agpN2mshDk7sxHx30iJuendzg4n7VIm
cVOonXjourNxrKwrv1sKvipLe3m9AtHwgEN2ls7ugaw3P1IBxGocUCoBBKEdYtpK
vQH7a45l1YmWVni4YHXfoHSkI12E7OKSZhq5l7fSdTHGx7O8jCS7sQds47P60aZB
TkanXntmG3hd8KM2A/t6goWzNGd8Z+g67MmiOJgj5fQ26RbpKpkoKCuyf3CrytjE
N073+iilu3zgmeXGd6N6PMiY9dXSzrJpVGDruW57QuSMupdWYIfaeTAjjEMl8Az5
`protect END_PROTECTED
