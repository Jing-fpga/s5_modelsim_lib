`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/DjIzsg7NXhSRCXrDq4rQxPfOBX9pxhdM1psGyE8X93kpKTKzZpOXLwYSByPbUZ7
zMXLmM6nualfDU71u6yGix/YHea0V55XLoMkCCrFOfyOAAaNzvPicDoBtnR826fS
nZt9J3ElX0R9mdfRcxHEVHNU2WA3lZVjfPifOmvXOu2Y6qYmeHa+kQAprW6w/wlm
LMZobtv3k+sD7EiclcUFMuhhYtkY3AWOPyPpaqysuYgHMW35ooaczNf/dCLS5X36
F3y2YAxXeESYh7ScaYfDds9Oljz1ioof1eRTK6Bh72sJilfL1o91w97FMhCbuQmI
bUGMtkuFrhAo4bqISPEx9Ykdn4K0incaULE+phb7F6i3xRJ1oLNruJF+jYzgD0D5
U5C8r4OdjwHv0NDNxe4VNCJwIGtFNUCFZLJU/8fa59l3grxuUoz1uWXgf0lC6sFn
pKd+XUyIObcI9WrNJG8qr9sSya+81wx4KoHfxnBcNw+1a6kDsyXV73QhrkRsoNLo
rsrPp9GLkmKm1nE/TWtdlTeugNiKmLxQjFtqToqmcGl0HfUbIZunJU7y9U4AXXld
m2CNxqxaL4Wdmf05PS8J1zfcn85A/PuDimMc1V7KtjA4o+0j4yfqnoO2h0FbHAV0
CFtg8ui9aCyGV15uyI/HMkVEjpOORYXww/Xu4lJd6Fqg2kXZA6MKev0wBmLfiY01
ms1OqGWTM1YrMuRc+Ld1UkhrvoC4qUNxwa2AL176qW+H9qP2Q2MpFEjvKiM1/v8k
ALsopO6hkbAf2zyXKnlFiDFJ88BmnIKFWwS7qm7DZepowFUtOIUBabTb9mUILKTq
CKOQea6fK0CC0fgsQKN9Rym6Cs6GQ0buLFlkPUxgQgGEEdkTou2qGkPqFAflhqP0
CCmHsrJ/hRgyDfCEqlUz3pCslirl2VfE2lXqq8xgVOTIwHLCyuVhXQS+W4bHJgTq
v6kDMIBsdQ1qftyMNcHTbdkMkUF4WwwGANQiGAv6dkG3bDDxo2G8xSVwQQpbTsR+
rGXnkEhr1xWHOiGWH+S8TGf/oFeuxMu6KX1li97JCRflPcfk4cS6/6cVolIRqaXI
ECMmBH5RxsqZJs510AKp+ZQ63C587s3/L3ghXhNcn6o+f9snOPPP3AsHQQX3tXmE
xhc6lP36FZ5xa4ywln4h4wbN9mVy035c8tAUGGIsz/oj1l0W36Qwl4+U+i2VscDi
vX+q8ujcL3Qke1mW0ufkBi8C+tFIxDPdkbnhYPkzOhstzuGjL+c0KMMPpiLHo989
+/s7G1IU9CukZVpLwMi5Pe1uA9ihj2ZACD31Y1r0i+Y1iGJ/DmhyvY/c2yRfiN0K
LVGKe3hbWlZUvjX2X8P7m/8wO1tGVyafptbStJPBjE9H/8N1a6693SMPYnaYnMxd
n8FtQ4qCxngbbgB2L8RU+kIkVt3ZqI7DLDrtmOR+Lf85ikvTR6ARGwpTY3C3Qlzo
IWF87IL3gJ4dxGIc2AZG8O+t+2fPmN96DQI2Bj42bse0+cNtQXCVFBWNbXNphBxL
cC2kLgDCkLRd6VWuSuIrRAJP5B+cUuEkzEvq1mRzFwYIxTymU79h6DGClkjMVF7Y
fEv0qgg/vQTtKK5Gu5VW02pfip9d3qj8LPJzHyfSZ45y5pE9cMuZ2/HyV3ykFcz2
4jvWJ7Oj3I+Tp4G8sBvSsb+BFrG9uyrwkIpniWEOQScgBPi+XzaWIHwkxnZvLPMV
WPwIhXdHB74husO7vhkMnikI7kCxKm4Eerpx/tgT3WvNTmhLIJbyu3+PwVBrdovL
xGylcSi6w5j4VWLp+VUBKXMb0vh8vhoGNyWQ+fGH5q0tQLzOw1Wun3GRF5pGJOdl
wvB+Gw9BmB9AYbmhwiW4+9mFwQZ3zJknvqSlsI7iwxmFpcQ16yTGsUNng8LLhL8/
CIET+3AWszP21Uqwjm9njZFklsr06eI4NCk1q88t6m6H3f1ja9RJKecg6YARZL3v
123Y0wzSiuTPCLwwY8Qevm1FZBg7iIoh+UvMB735paaYxUAzr+Ec1kJswTXu1Rmd
MBJGaDkdaBc1MqsDCYxEyhgIxD0HlFOs3dGJ/GttPfxiQ2xADrCyivZtLbsDzMy3
VY5eNLCCc0GCzhuFfvUMxAR9GkrPyhWKa1P+L0c10CxhYGymf/oanQ7mLFsQKATF
rWrUS9NH5wPhiSfirDbthH+U3ZnIm6fh6Qwja1q10CMJ5MaC7dl+I8n17/5lD04l
9g2kaax78WCZ5mSTXJrZlRvrSbfGDaaFYpeyOrbnIvKJnkvq+Klq/YuoBIT6wo1i
xgDW5/71u+DKaBhTlMiVe0laZY5UYbEjN036Md/XoYaUEB0J8bi2BJ6VNJx+s8Ct
fgFb1xe4lMzBQ+t4WcE244TjJqpheTJW0EtL9nd2aWhp26AFqbQOuRlUcWKI6V6f
Z+i4ZLHwccOfhLSBRxbcULVpxwe8TEAf820i5+hfKDUuvAP02OdC4kLlxkdDesWa
kjPvj1Df6mAsR3Ml3rTZrY6DvanPwvGEKJ5aZFdI3JJnQW+Eo8FJVjDmWRXo1ip5
I2Cn9NHEnka6ZITRrAAEROcDL+YFFBlaRQC5IqPtfL5OkYmtJ+TF9xfWglb8xXqr
F+h3W1GfrV1eyYAdMtqfaMixolBtpNvXC8SmyRjzG5NYkCJWq9ZoZphZKuHV5kWn
HGu82I0dFWVvSv6Un9sa91O+nzSKBsxvPzctiZ1Ok+L1Eudq3zUzXaWZrBS9m23x
s08slaYj0ajmv3RQh/JU6/cLfp9OWdWAEe+FMZTBY66Xyh58WX7Qh2Tvv1cUeTFQ
gox75+FIboxU5mgkWV+AArPN0p6I9Nbv64PStj110pWMSW8Olqyd2RksRWxm3r7v
NY9Mdemgvwe8vPq2LghBWg==
`protect END_PROTECTED
