`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8mYTAsJYJfR0gtPcJ3DwGdgt2rP6wk9Pe1X//wD88S1bsV4ITdbO4Oe090L4eTUW
etQ4OG/XkJYPxMYLn2uxRcE9LQQceofWjvgFnwNx/Gk61zyinokVXipP6natORl7
zRespKRJacmzKluB7y98RzlpeRAltncTI8SkMW/vSNLhlm9COI2Q7BfW/Ol5KOMl
E4C81vm6IYcW2ZtXF/dTjjw6zf9zd1XvjqJ81YSWr4OUwPN4R8iYZ+QmE9rL23K2
eaJ5GYgRTroimYsnfRdjERauwN0bumn112V2Pt2aSg9u0B0HxYpyt1jlGbf/sCvZ
Y4WBZFGecz7opQAopUgEfF772TI5C7rhXZXpC4sKrPyBVOTgQkxbwyU8Y9oPn2/Y
W1Z9nKAa6dN3x3VlkMZQ0Y8ZyaFeA6xXe9QhGeElpVbuJMzTqxw6nd3SMZXqMLCK
d4GXypplIMFfCAIazG6sldM7IUhgvCsoahBcxSvn05Q9kuZbRE4E5PaB2+RTqBEY
fvEYiZU02YYLDwtP9oOl9HxDc1RFIgnlZ8PmvwOcExXejRjpN7XkjKQOIXNCMeL+
Y/X1lbGoWI9d1OhsILY2RTa2ZFg3zePEbSqJlFvhnsS44M+tztv1l5L+Iz1MIZ4s
mQoVXPVwHI28fwbGcMqFMD2sm6p5gUq3agWmsdQa2jnxOH0IbQctQPGxfXVv2ylT
1iFNfqw3r5MXlfPc8gHGyf2iGPCuhbxVWnRVB+FWeUb++rX+Y8774r3Nes6446Xv
cpmFsjrg8xABJ0yTLi0ks1lRLlUzC4fB6FlfJIw512kcYskZNPaIA//yhRNq/U4D
Ml6H9fMTqmgUWV1Y+ktE6dQr+aIjoIs5v+6gBcu6C/pT2G9YwEGVHcgmORdk6YkN
P552RhlU1GL8iPKVOEdUJazC3Bn451/r6akSkX8waUk0ZvErdSA+tsmzGIz6E1qV
lq66YNWsMtrV+g9r46nqDl3Pxy58NXgIIP+HdhUd5aZU8zR+YkguQJlFV/M6w9tm
96+oBYiWz/+VJSSGxlmWKCW6Y/AkHlULVKcIFs5faK+s0wcAoaLlNNZ5eZKUtfkv
5gNjCtmzqfcxSNeD2KTeReZTs3EibK3B+Sg7mU49tc0WmzLyWoFFXNvNeuLD6z7J
3NTEvkrO2GX1NVYk4wLt5/gdLdWC4XcM1AW0ZaEKooeGc4pyBiaxSqzs4rpSOsNw
TP2JNvX1cIelgGBaLKkL/0ZwIABWLE0gDjsvbzkQHqdQnRsmrtEIDeTPfzn5MrxT
ZMXkITyhcWr+r1JsRfL2Kmo0+DW4MyZzo5+Y/PvQb6kdvQNDmO6szy8eBhtengYR
ihjUzMfAej7eCEp4cytm/drMp0vHLfTVPdo/GFUH206PSOWVihHjPXHl0OQDw/9C
qjIGDRCW4UfVAHV3ZDSeQPY8pz3M3f7xHlPGrkKRvP3V3XSbZyeelFSeBegH80Lw
yn/rnShvamnxY883w9utEQ==
`protect END_PROTECTED
