`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jdl06VKQ46XpnLtrvYbofDBeWXGrAZWTVIhC/FiBvbpFZexGvTFxfQHMduhsaRj2
PWaqvUQW6w6W+m5+O9yA7xuq13DwOvYNwSxBFQP4kwxt3VAIs36jeUnJC07wrVgS
CGRsSysWYOoWo3FYSr14DBkfydZDLW6qXKEJut5VKhW0Siq02wdL5fo/54gmrdVy
xlH8+pxckl4LdFeGzagExxI/3XY6lPZ4Fj3jVWVTvol41WGubxU9kg8QKvTsd7mv
vymsnjRpmotZNRkN0A52PH7ktW5JwVp8Humt7fjF8wS1PLg11n2bCi+5TzMBVSiG
+aBxK8O1Yj7oCdQOTyam2YM1ycwFwIBNLRv3l/L+e4X6j9gr7Cg0cjtlIGFs8zCC
IQrMQYB6L72beejx78g3LUcasOWuN85mX4uo4exk1uRRlOm5w1ZT39lnJWklDe1w
z7iev+2srxUO3EDSpXPlrxnhwd+vgrGSGnwfFV3IizTnCfimRdQo/EWkOUJpZUp6
`protect END_PROTECTED
