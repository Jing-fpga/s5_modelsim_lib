`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
83EU8oXFJIevjAm7O9Ez1DbjEsWn8/R8unBweOfe+o+8wIM3iGg0FHgD8IN2wfrW
cWW1Kr20z3NvMh6A7Chlu0Y+GlcOcEY0C2Pn23VUfdkGArnt5r2YfzF4bSPJFiXq
tOrLQO9/ARvfgYKBrpBFnb+jWzNiu5efeDZsv5YzdIBTPRf96p+sM9Ul/7d+pKbF
B0YAvo1TprIYlz6JY8aalGTsbXOCfRuQRFmvrFVJ55xsgLdIUkDp99b+y5u4K8kM
qq5Sp3zuupmSkJ9/R5bv+fXz+cpeehGlPORw0zoemxJ/i7yu+COv/q3LRpChMlIH
yM9wky09AkBLC3QSqg528O2p6WRXILr3NBCi2iJleNRj03Wtk7OZ6WMLBCpOW0Kx
f4Yj3txNA03KAShxcZJIAr1+XQWEH4XZMoEuBQkn3RzMV+UExYCsKTy8MDfOrC9T
ncVHBxkthLFIL8VE3wpFqZEnJxc9nHv+3SnQclNTY5o7RPwPhYZ6nmPay3BXO5kF
hlpQBiH16zyh0k5co3l3pbJsQy7Ri6guxcyJEViTgChFRRgt+WgIDRQfdsLCT5sx
yTUoOHhUxjZtB7DzfZGmW1/4hzaXOzRaZlhL18ohLU/5TuOxyAgI5e5SrS72TySk
p/0HiVcbt9XjVeu2TIukaAvATkGP06psJoP5trkyhKklFJ4f6p7N0EC6wAVlWjih
11SadrpRcpuRV55cqE5MV9OboPOThVXfumk2VWNP1ya7temsM8dgWE/lI3fcYl4H
mFapKE5j8jZSqnpSGEuZerOyxzuiLE9KFjcuxQBvrCGoXajix1H7Ztyo2AU6VmcS
WYMfeITYB0V5jL5OkB0M1ixdhVfnWeHfLYMQ6W/OlQB7qFnPYlZV3/HbHV65ZURC
E71n1z33Bu6onW5WMQhTN8YVmOdso1nzswTYiVlqkEfYszeU7DDo7pzAptfcgTa2
Ek5cW2ZcEYon2csP90u0k37MWcgvPUW9O9Iu25GRo5dH6l/FspF7/JxPJxDtjmrV
OMqXiSuG/WgR4YhgwDbZEUeoYoVWMscR0+C7fLjqQgsr/VGjMyplsrDQhMtuuaDu
UcpDyJCf23fGyGWmwkszwcv0wyxFxdhncZzW0z2bOf2tDdoELwHIEpSaw7gXYOy9
oop8jfJtT926HO17W38d8Kq3RhWmm5hWHMbtfMvBNduuv4KaH6W4a7ie5lHgm45F
SZanlg4I8S5gbbLzcy3kLmVMLmFp/FfTDkd7wqW+Yeq/qm2kB8Y86cynzvvH5ggG
9GRtnXC98wiQup7U/W29P7L08B3tdCVes22o+wh++GEo/RZ7If6setYnNwHsXgKQ
O9iqNGtwROgMHPpIQiFwWHz40akmBroHTxCXpYDLVv8LEzZb82PItltlv/0/+NNd
3KtoJKD594Pxv9Tfh94GDTnqWsOo0JVAoHOPSiC3X7QvFdM9mOWBmKZs0AW3y07d
6j5iT9Xgzt+fg9PISmldMCgGK6zojh+28TSVdXvNtXcW6kzgQg8L3KZq0zONhhKm
`protect END_PROTECTED
