`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JCvulIy+6gi7kIkg/KYm8ouji0Gy3Gp6oHZaj1ykFvota+FCqSUz89cM8bKws96V
DZKW0yVYdKAIZ7nAh/5vQrGsOs9jpihSJrafnWlJL+q8DIQPo+tgzcjnlHS8Nhcj
FSjpl0aHtfj9+MW4tiRpEVsqLWLn3Ct6N9WCeW6JSMm1fdhjI09UHpUCXJHjgn5f
jo9Tbx3S373GU/z7L3/EbldcVO83dMDJ+tG0MwJ5or4VL/pKf/udnvtsqD7U4kqE
qmgjcN0aCAs+FIyZn5+/yCKTqyE/Zi0tM5+JfXd4uyuNv+6l/7uXKcA0xp/LOGOB
hm+dZzs8R1j9X48CPXjpX2NJsRt2rhS7+OvqZyhNlsNnN2hlmzgFOCabHxeHPlB2
ZmrUOdWt2CA4ZSHicrGHjolN4Jje3i9I/qK4tvC69v/nohG6YXWclapvBRC7FNDP
IOxRoS9l3BucrVcc0PqzyU3HYJPG+kapQfO3tmvh3+0f+CKZ2Z+ogWliH1HXYSqO
hZz9eFZa8LPG6FFCfS7Fp6NLLGalUL8pW1I43Sa7Jzzj+GF2m8afDkcYvJbdxxMj
sGCrPDb69uf9Z7aq2YCz8v35RUCWPazX9sPWFeUAtVapLoN455QciUQrc2bADEly
PUisR30631MmcfrBrdCqazsSoK/b+Mu4J/qBsebhX9MX5JUYY1Mm52reuccpJdVx
dUN1g50mH6f78gNWYd8CDhiFIwqhTW30LEhQvSzYKA+uU2dkrdeHn+NJ3lc9QnxI
Zc4rrCdP3Q4tpq2X2fqRnCK3DLUbs4hToUqaXzRamSquS769b65Gwg+4ap10R+EU
ZaL6iCckt+BqxmSDWmdnTtXQv/sVnW46EhkaJaGJE1DMFx1N5QX+9Gt0KQGfRMbP
zqcj1FRN7tRxb80Ot+t9uqv7PVvD+hj/dhr6c+HI+a4=
`protect END_PROTECTED
