`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4af2TRZ1YojTti1kxEScyfmDPfJK1kJC/geGnvQLxRZK71ovZO3UZNwhQpv+p3DL
qwbAsBKxOkNm9n0lKbY7z+nELzIDRbiE4UzNciItwEpgw0RhRmWHMQjS23+lALsG
lf3qhrY2SPBDXNWICtvlkyqzQOg4mx7FH7b4LOpJMSDmQcRhTC1Rgfu+Kp/pxBwd
rGpeqg9zrkGStiJ27kKyh44cux8Ib16hCWZ+XHyds1jBF25zHbHyv2zZVKmxYBHF
LfN1bZEZ7+G0Mb0ssLn6yjI2GzppVzkmMb41W2XRNw3Ngs6WI0YbzMj0znixRtdR
LAgeec5+4LlrnsDBh2w8WKufccPD4VwRbsY0hAbB2MGx8cqEg5OIlO3kxMHla44g
dSzsyeyE7YFXrpBUcn/XxQeVQtcW3e5BdxJFz9dh4MdokaEHVyw9V9EaLNjjtyss
Dy3IeY421+8aUaF15+YgP+WJoaqQ00kIAhBYZe5MTVu7TVmi9SQ6TOhcRYMlAAOx
m9Rekmv2m9vdc0SLDnD0AEX8gHmf44BBl4xkY7FmaTMeRwp594WQ9NKVZMKGw084
ck4SiAQl/7JslnY1j4uxZgE4mVt8xCwNp7bkLoxrsYWDAA3kZ7q27SCTWLBn85P7
iEuHAoy7qmM0N3QgoZTiegFG6qk2Tz3HFIJNOrTwOguZe1c8wuF1VHrO8P+vVEEi
y86g8TcUgeg0zoR0i/rVLPV2omeLCwXT40DP643vDlFJtSG83oCdzLqJo1bbJY9B
9xqT6pIG81cfTQ6Bc6VHeEEXYGw8ULbrhDE8DP67a/xZw83EBPjfW99eBVcHVKC0
`protect END_PROTECTED
