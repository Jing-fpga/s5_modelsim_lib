`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t/udK0/QKI/2dsMppvPZQ/Kas02Dj5ETpOftEs3nDy2x5zjmDAD6TtI0AU1z59KP
lAlxgrbGmcjTN7Vi80RdtULh6EfGHqhsP0byrwws4GqCJbWWODeZXbQspV88S/M4
jFfZ+R+XB9ed6+M6luXUpORFs2gR1attyaFXDJ4+H8zx4ZGYN/0+fZAFYlRWNsoL
oUTt6Pz4Em34l474HQyK/kA3cMR6VylOETyNt3KXkm7mXJ2urnegscQk6Vniah/H
NOOxMBQBt0jXN9Aq1qM7LHpN9HLYRQLXkdUOanNqQ5qYtcIMKLzw2LlqPxEsbKg2
mBQRdReZ5taleeGuMw7Zxit85HMeBjQ6Q93RoEmbhJD35PMIpgCpggoopnyrsSIb
kzkr0uDcwt45NwKxzjcShkB6TfQjoc5ernUQdwH1w9BxLo03mHT2Su0PJLEeNM5O
uZ/YNFA2Ug/NWi7VKaSI+juCBLRXCFQHkHD52uUnNJU560jx9nrVqLb5FXw0qk6t
87/k+bE6BR59bXhLcp2jH+SK27b0mHU6oCsu4/168RtCYvzJa5RQAjCEzOJfL0UF
v9af8c1tXtZ2T2dzERtBqkGHPQP2eWtn4ofsfJz3pnnN9U8VJ0vgH3bBn/QVdmDn
raWy+JxsavQ59jiw+IWKqPfWORC3ZnUxggdya/MPLNjH3fQF9XPaA4j3CMcgf42z
YbYteuAR64HQF3eoEVrJLO3zExAb0d8kUrSlKq/Gs38CsaRAbLFQJzxTkso+Eg1G
qxAR4R5924kXDV3eyjfGLU5ohx/eQCSuLyQStBIyiTTp2HWuV2sHk3c1fvOmuEgm
fN247GLAzXH/LAHnA9bqncAtqUp0g2hX8fCadXTPr1lyu4+wvxvWI3unUylyOL24
lEx7QHdPt4lWFEZlHrcRIRGcVIIVfgoSbJDELTk612GM5e/KjDT/XYWSqNarhHUG
dntmfMMC3y5Y/exwepBV7ZboKyu2bj/3L9x98OUMRkuCG7FQ20oO0uLwlxvwaKm3
aQOK7wJbZwiQMpZltCgZ7GyKAE/lZHjyJI+2xtRZt0pCfS8i6jFb4ScBVbqym5qF
Ux/LEJ1B+ywFlAD7GYWC0Yem2pyxscJxRAMjVvQpZqa0qXq0uyCOAFt3Q3J/v8LO
u2my9+50+4G6RaUzFeOYjiV+uTqFaZLqe5FbH6UM370PHaHhpigT5ZQnbkFmW09u
csxYua6lQDHdBh6LkHpBK/nGsHmuGpEhBtTyHT/hGMeCWpGV0L1uYNTexp2CnyY1
Aa+iNjskNJY112wPqhTq7S2qiNO3SyLge/a16vKMWurRfcnUN5XEO66TcKqOuZD7
hO0u2RvhAfecTVBruu2AeEsdtLUeSnT9mPsSJ4coOI90NkhuAEq1OpndX1iY2baz
edeQG2SHBtpFCMDvn3IeCUS2IoSlsSGx/F3BcKv60f0erFxD+efoUCIUTALyaW9T
ZyQgDJHNIiNWMVk+esN9xm1Ah8sy3qPKl74OyI0Bb1q0tUvtGR3SWOpNnHekC+jO
ihb1pN9bGjbFFHsq7NxfqK6vHUITOGkwFdFePAfGMyTvQel5wT0s8xmO6uqGGucm
lE0x/gkS5CE+2ZTGG+BY+qd06YKz0zq/firVWyliJIkOdZwgW+3E7OJ8i9fXBl2E
ZeaswjGzWiBWufi82qQWKfwY+Z16nJc4sScrINc8CETUZGoce0wX1pD6e0Xkscx8
OYM/Gehq5wGNbKDhPc1rgKiEicWpjjIZZAFod1IDmmXY5s+0IQyjCXa90wJQr0Fn
4RLp3Eds5DFmX2y0aRX/G8q30pcOLlqplby0l5Rmlpe2moALf50C6+mtgjYhf1up
NZl0KU5eKFl353W2ZgdOriFL3tXdbgyQG+20QFaMRQasC7E9TL11pk//7CPoAp5C
9pR8CVK3VQ2FRsTBOvxVQXfYTl1hLCt40PJYagQip4LfzSTqhJn8wFQjTYALYSVh
mLJjLCEyYSorqm4VR8IRtA6LG0dLYqLrcNPQRyIHrYy7sTCKJozbRh8QEyP6AaUc
8bKxgPpgtSE14D1P3aPqerzkBia5ekj/sM8uWXyvED40k6WqNTLK/PlKRPAcC1qx
HCxas3ITdhZsDoJ4ALhLpRlK9OMUJU+Ow6sjdJXZ7wpZY3SIwz/K06x2A2s7LMPV
o8y21HJ8gMRcC4FCfwsY8tncXGiYrwXrqwQeVfXFF31pzChwOMkw+wTNNKc6cNHh
CAHcpON2ICP9y0hHleCg//mriYhSx7hDzZ2VQKdBXL8Rn9FzG8bwcdj4iSJlWSto
`protect END_PROTECTED
