`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EWY6sGMZ3iABeOhgHdlH77vflawyibXfrF+rTnPWvZn2RtE0fZ3tLQ+D7qelEFps
lppnodu/kZK1QtqDrNtAb91n6pUeNGnSjA0e4C8ifCXlnFl+W6Z7/JE5Zwtuexat
pmw04JbDWL0q8lRb2jKH2dF6O7cFt/kjxeR6aA5bEHOCWuGVIdUNqvcIzqg8eusH
uexICpi+XZoa1Yn+3DEdEGLqIeRB9wk0WPn3BMJuIpcdd0bMLB2CzNFB9qL6ug8O
TJt2i1O3Mj+UoIepRpvCGlovtxtcxz1of4+Bw1CdHYRjGRdlfnv1iwhef+XqkupY
Swt54KvwrTg0xcRuz81Z2cmIBjMvn+3cCqxd92RZirfHjF2/XhvCZB55YC8rRVjc
`protect END_PROTECTED
