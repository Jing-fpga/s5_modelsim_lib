`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KXHKnaxPI3+ficHnw8nYMS0FzPckyeyjGK/8uj4voJQr/gRXHw2m/XS1t89morwT
9X1OQqCMm52Gpkw5E3R52KV8/iaEzrGvVZgJ8f1bV1yxm6ivAgsmxRSpJXitveZ8
HYXgOoliLIZjBnQTxei/wLEmi9ZeSwkmbKdmfqbsDjMBK9eBKKoZxE5mmDBbHw1b
VXirVsPx6qK87QOCqaQAGusaSn64Pr5ZjhuQW3dwGVJ6lUFEAkxBnSMYG+8iuIt6
YmGpXzqPwBM6aeAxxPXC0rxjvS72dVFzjuaHbhQKzeC1GeRZZV+Z1cIWpENbweiy
Q8KEtDLxaRnJImQqcNg/kfbR0fpkMp2m4XhsN3x2BoExzFaN+/+oxhwa65A4q0YG
hwioHzODSFz74X/tHAIkC01Y3mq8GqbXH2lxl8+WQVUwFwRzBKbUpR4kPO+RcL2O
mtKzXTXhJlmVF9bpLT7uClQUC1goH5FKEwVMHF6jGNg0X5Ts85FyXepGnHv8kgfP
F8Qgc1JgUEBsitJZwzTHb3QrqUiW7Q+vbmXd5mKxEamZxtBzvM6/VmHUALgEoiqO
OF9pZmrGm8lZzvwPg4qYJS+Z2atethczVQ0H8lgNgTjW8oGxihOJ65PJTIbAAzFs
2rUbUw0XpzHqLOvL8bGXxM0n05UUl++5T+NgtYqnKh9A4sArX0NxZNFk4C+o66h0
m8IfJnME7w6X+fka8+vTCaDEzAc+bidsiZD9UD6+dsBG74Aw6PKAtSLij7acGfAT
0V69h3ywB9ES1s4evliQ6E+sdzI+joeDOJwKdECgdjUkIlwey83SuWLiKzNReWLh
DWjT2/vN2a5DZNwiIg/ztZPVyYLw3C71aLm4wIKb+U+ELmu4d8yoIQUMBocyoqSZ
f4rLbM1WN5XTveAospU9hEte6ckSBmYoKuSR2wkQ90GNJAJmUX0MpsG1cBsFmNCs
vIur+7DayW3zDyQhAeTnkcRj8TDtvIy9SILohR1QgNg0n3vEyI5My39PHAx9wwkp
3eyr7/5Yz3JqeJl4zcmHUxzVyv6AWysiTjzdn5YzSz7ubBTYPiP/g9mwFfwCkrBM
V0ppOiO0I2BqRhz817Lg4ZKtZkC37YmTu3vUMM9n5CuDtqaDNV5efuYOBbjZvTFu
bDeqbSc1vzMqKO0E0CuzzLgcz8GIaiDPyzYxoUxsYmFblTZ7y4nkIkenL+iDJ39I
GKGBkF47Kq8i5VYyluZSeO+HtC4UMjBZogZWmZco+cYUV4dWt/r2JktV+W/KOmQz
xWZxtQm+adH6TBlnP0CfTYGUFismoLp2MX+6RYaLBYX+daVRRzBFyBh/eADaNPrB
SlqqgQeSmPr6fZsJTe7C4czKuM7FgcAZhK4FqmALkCjwzLn3f/gZ0w/VJ0OLrv1a
oMXr3XhU365YrtKJRkU1XjMI6tN+TFR7jEBxfGLGOpjs7qppH4KacB1ydz84gPck
kSp/1qOairHL1oFKTiIqvnbezCBd8qZiPLw1VGynpSIDRvq7o/9feSK8hrUJENyZ
NN/GlOFQCj0WVmx/fW7PakJ53fHe56HUvkIyS6gvy9+LWFK4pjtuVdudjgzq4r3U
Q5NSRrT604CRXjl3ca+zMXsuc/DPq4jGTrVDU23H6z68pbypagjVImjSE8+EbHnf
I4h4TVSLEAxpgXO3ymQpDHo3LSJtnVQmEpNabXuu+6TivU4+kH8z+UmKmXZWeOGH
FMs238pEPlbDZ0fB15YXHAFMyXq5EiVc0b4qiO4nCA4qMSeTj3Dr1WtALuuergym
v3UWy9bIn905Bq5p+nklPzJRst+8YmOSrw/ErRWo5dpPO6XlAf29xYQX2nGYOjqZ
YQWLuu2g+lKW4ct1alOg/BEAUVDQF2dEY7oeQbppMuba/BXerEhW97ES8lfXlVvL
yyFmCVUGmDY8xx/ti1mA+WNn/M4TLYblYR7UTanm1CNPjPMjtWcGQKjL4WIxk/pl
/O/gM2p74lyvXcBJD0oAJkDer+6lM7A3bbhjHj0ZUdFK4DcgniQ4VUYjxxNwdoM3
xpVXkEiKPA5qkspQWzDBmDwRSANEik90b6Vims1Nhxs5yHo39wOWMTtHxDkPqQmS
HQAkJZ8m9uKXrucqw+ycJ1QpTriTTqPHMWVbDdD3pV7+YYRH3t3AG1Q/imfCMBje
i9Fe/YZDRxDHl43B7mwgzl4EUifcqSEQY0/Lp1SjgDdTyYvms0p6tFimoA4jEwxE
sHDeYRpC98m4FEL3B5RHMYD7Py104bCH98a9JHUWNxZuz21bd6wiRtvTNXJWguGb
8pMqT4SBR2tM34E0Iy7j3Li1DxKcbBNbFsnm3oEUlffSeDT3K1K3T4rU+WuvPibT
I70i5GADiWfkTRTW47k+uZl4Nown1Dzyow/rfuMDLgN2Zfk+fWYZWBVkcOzPH0Tc
1UwMLRDffRxOieeF78fZ6LviATeVWgRs1/+nDEH7U05u+2ZYnzJaoQrp+MaLv1Zy
roAEXT9HOuyUm7SWfEM27A0M/lrhHhrLcIEj/8q3huM=
`protect END_PROTECTED
