`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mgtVo6Dubc9KW8Gnij/csfxQjoWYZn90hmSBJ7l04y7OYmQq1BZnRZx/6JOwljfA
1aEdxW8jveJXUJAsNpe/WnRyUkc7HUNGkWdRNGTV/zA/oeMb2nrV7vaguFfQIrHI
dg5q2xjQed86r3RdqgHfuyw6HlZOa2mD9z3eaTWzEw9BidyKHcHKn5ZkhTXVlnCh
l/kXHdWfVWw+2dvmFSLWFAlqpwwMqFQtdROc2GxAfLyOTR15tRetaD2mP50fylL0
vf+LL13cnsmw8gdAsfmSsg==
`protect END_PROTECTED
