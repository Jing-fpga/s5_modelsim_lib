`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8rGA7HnZ5tpfq8/zgBmA0Vso6dH2BM6Rb5eTtJiBrcKmItURlcihZvCCd7p3D+/Q
O/Anr5rhUm/TuwXMeZYfSpf7vXaEsEcoWW9w+jnzOZ+UsR+wLjzi2ZU2SmaqMyGr
YW1uQdDrK9X1BfikeiOvs8Z6JgOzQIu/k3/Jj4MCvU6HjNdpbRhVwhE495SJY2PS
QwZ3TyTbLyYzP0Aq2e7RRXJ5vykJGxxFeA7gkUsn0JB5uUy9TQgDh7MN8XHo55sJ
WmuBPm5BN0FL2mLa/Fg0tKDAYf5k/8r31NpB3MZMIBfJkv+5p2d8stYmyNm8B0/P
OFeY6WKomT6W2fWxbylNfsYFrIAIGjus2SkIAEPfcXjga4DNHRtjlc9IWqIt5eDC
U7QrbqSQTtAY+03R2ocMh9Zogl3vvXC3/ZRb/q7oTFWXFjd8TO9HG2GmJPfvHlY1
gkOvVBJNybbVeja7/n+apdDzIlCdsMibtsfzSsA4PkKFewcNmTpHnzH+UBtRbFNy
qH3rLpYCt6adIxiiO29Z5Z7vonYzGVE//FIWu3z/XMxTVln2MA6VzbjvwofacdjV
HhIXwv6G3FAPC4cUTpVHVGBzIYDatOSTtbNgbmOVThbqqrFzjMt6JMXRqH5Ev3Yz
u/3vTNxISEnJPpx8q6vrwXp9TOK9Nr3qL3owZp+TIlxQyaAgBmx3t6ps+4crBvCc
/d1V7gWcMXsR9+N6XRESjn7TffBu0Y4/iRgAwIkqKb9A66k7xpSVnQ97UMRo49cW
U+1Go1inUpJQqfqWNaSTE+M4Xn+h+lUFGAPAWYMstP3xwSTeVdz9lMTzbwfcJk/s
91qPatWfauPvajJuDD9BRlST7hiuMSCviWGjWWPraKbPC4JeZ+6A7uI4B8j0SSly
POid6SSqZ4mKk0mCdbJsOoF1k5epIWIj8pxlPnomWZ2DGzRnFagrGtOVQohOK1uv
NYsvJoZdClmkoQiyYL1oADMuBzuM5ulmlacn00lVpxDcSqf81PZsjvYZllMmcNZD
Mi2OyNhmJqnBrHyx2i/CfrAYsIbbp54c+Uzvqg422zY/0uafKmNTwC0eSBYPDc5h
pwNElmT8fLC9tGjX1eid6m4s/YWegDAuenRHkndEivcbelY+f4TLaoUs3fq7QbhS
Ga5HyZ/xjm/0Ue6ssGZFDWDrtfCAlMv5Rq9uvupWpdOa0a+/XZYKT/ZRAdSASiJj
nsHwYnxnm0cvgkfE5cBj8hKcx2sZOS8H3BVk/JpLo0DBAncsJuhwf19+uH2o2uVA
SKiO8YH5RF8bmnf1mDDuc9YPYubCFuXjDS4y1Gg/KfkbWpFbPwkjuneTqmyQk/OP
ApmC+xFUmDT6rafOEdN7W+8vx+D7gZbSilxUf6Py8o7DIvgmrGDxC2STcCt//O1E
a+pXkEqehCFeSSkmabCey7E7r1fgs+aiHoCDT2RjAnUai8GmhEoYCkNhTYpn4y1I
n6fhyJ2UHBiNBwgBtzsBfuVTQaawjYhPHBnrV2fAlpeOEzQRfMy81asOb3bNI25q
QXVmeszn+3BGeN61Qp3sLAVIJ+jGVvu3Iw2I5S7fR8K4PHLnJnQVCDvBcVpGOyzE
jiN2ZF/2rNUPThQzjAff6Kgwyo601K3oItaTMfQWmMlVga3m8ACv+hVyh1k86tAD
6DGj0lozO20KE5MtlZG4rYW8G0v0krXLwRBrSo6GfMeIpPfsW4ZBNkDZoum3Qx/R
2nQSEOt4mnguf/leXhtXYErz/2hZxWhTxFLqMmQkKxwVULF3X+BSfKmkNr2GBuL4
IQToJmzcwOF+mNL6rHjUChZokW965y5HKoQA6YZhYEg4vQl+yuobU8FIYNq0YhnH
yqxua2VFkIv0yFlFFQOEGNV9AxNfPzrHoOMFDrjzxMHL3z/ar+V9hhFfGjS3RXV3
euoFdbf24+uE8EljPcM3GHZ6cr9JgP7Ht2Eg6rVQuhd8aUF1CLkksajpEpPVd91g
K/PaeBRRJZbTydH6degKm279sDBiiJw7G1Cc6msMCDeKS2JrSu2iLIEs//s1RIUi
bueEHeWOHUk0IqNh3NgqTuij8SmP3EIF7cslZcA4l2YEeSDbWBK0lLDY2Ad9UJJQ
ZLEMQxrEepeZuDRqPsZuWnjokFQq7JDsABfd/W4yqO4l3P4JBTiwrm5UqM8IgkCD
D+JanJNFyHyIhwtROXweGUWU3aaoeWDj2OTN7yVw6dfm4nzZq6lGOG2JKNJTjmIP
ToHrqMVS8uKhkOtJOqvRq8BATxThkxqeTVx6k/caGezJpe6xqHHZpukJMobUBtIA
nGeftcpZDj2o5zazEzc18ZF1fHf1hBxeg9CkBdAIqgcbJIBmkZIh6XTeA3sKI40j
beq1r41EA310CkDqnbgDYAFuT9fscJdNrF8Ygs32HkXhXxK3EBg0GtaklmFWU4j7
jsOYPRkv/RcCgNJBGHQ46+PYCAbJejvf2dFMQVTa3uucbTXF4/LN62I/BYDEKFGm
dqLNELXfxGrAhhLN+vPp3IWVsxkZxv9DUDQxK8NLkEnS1ENZICprkWeAvfzDw+uJ
XgswKuJ5rCn6aoRRzcAF8+5qIVYRGb+EW/Ol++6owOTooJ6uq6nvBo3MfoulaYQv
FEzMG+9XqynMGX/3m3bKQcAuW0NGJ8ngKoO5C65hOO7D0/EKgkhn+vN2U9m9OiRu
DxfiT2gYXW8rHOVNl0vxkzzYWlapsYP97wEigSuKS6Xfb+lnx7GJePrYOPZA7fq9
fTM8Qv87x5su9wEM1LJnL1YsJofsVkR1jfSNcNozEnolm5lN/PSU0eHvNYeD337r
B8pmCHuXK9DfNBpn8n4iRAJIY1TYkl2Cll1X3AV2uuLAIp9LAx//9MOnH5kkWCFL
c0vEID953lxo+VFN2M2rowfnP5IKOXzQJ8Fbf9OZ0/YwuNuocpnEi1SuKDDcP4d3
cbZ8ohhVp3ydGCWwUe7vbUI2JLV8NyptWabo7bdDn+akm+Ffnl7ZEVdmrR8eAELn
LAhi8gcNoSNb28Rkr0Gokm1P9OxVGafXWw8aun+CuvmkbuSWCajvV0ct9zuRbKIw
QEDizmNhvYR0T04GMboO8BiNrblYal3QqgmsVhr3KilQ4yeMu9DCMEFrUReEoGsh
1Ms/+0OvFN33p/lDWF+g/CE8twDMx1Q93Mx+T8rdxCaE7kyGbDLWF0BU2KXqA89Z
vGgBw0gScV9F7DVzOCTg5TlblE+GPE9tmH1qXyDhFKuDcsZa3za3ax5ZuRG3R3B6
cJEwR/vDHFvDeCr6qQoCRjxidqCRcPNybWlRWS8Yay0pB/iFP21JI+Dx3wR0fiVf
Cipn1SSJmkFYCOebuSHHkl1IoB2knguz+k0ys+M6p2kLbfGHiGuKZQ23spTVQVdg
EbUPrfZ7UFIvErfjrGcqcBoWZ0bDQwVDvkF43VJLyvCug5+QdMRyeVeE2nvHlCWV
zx4xhgmu0UEAHBmpUf+RXegy07Pzp4BD4nvvlWpu1tt+/R1supw5kum+8mMMolpW
6wtY/DrLVb58DVMBozQrISz7bf3OdY+/K2exLHeADaCUE6xg9QWMM/xZj9kODH0P
QAblCrGmuiQsShL9thAYHxFwYb0rvZQHt0Z5UW+dg9XPRlkd9FEwyTKJd3x8C18S
58X7+KajndFnCs1SP3lF+nSbZuijfHjzcjdt9vtbnCZRGX1Fos3brP0bX/rJDlWb
W9v7MTAAUtuQMUFsgn876jK7M60puYjWD2ey6ip7W3aou1LqLtP0UQ5pNSVaAhxd
lqewQp05xVIvqnFo3PC9VnuMv+RsuQq8FUKNB6RCL9GYoD+r+zqPUJ7OkPh6WOyR
+WAlWsv6bq9CyQfBnBgoyvhzAu8uF6IxYPzQzsgFkKLX5HkE+yQ3JN8s+D6GmrVK
uv3nbqCCGf9NuRV9RAejGhdlbKKyutiiQ3T/SnVKJZCzLhhxQqd2p1x8OnZ/lF0Q
+lHaf3h1UUQ0+FuAIfh+Kt/koLsZpScxkr5PbwsRcaajTmrTC+xOh6BGsHdzoFRx
CkFGnoIqXF32v2JuhnsvpaiuB5U/95XXhc01YtVoK+GQWTNz308YYdHV9Jwd9CZB
JYMhAJsxIYCuQjGM74MiuGSZA08ARLPbP6ZzOtUMZEjAJn2P1exxcqW/nog8pA5i
+5YdxObfjzXSGM7V1SgUoi0AcmA6nG/rwTB+6NCDdcq5ViCIHADSNg5do77UQSmq
NDsr/awlEV9TJOB8XKQ9NLsITyblxATqBZj1psIhmPPS+88tavm9+rgiSj/SF74X
c2m7rD0MuLCSFvhXnc/h+vGXPtone+u1w0vAqHMP3zA1FtSgP+Irj8HXfNvljJls
MgsIRtDPsGQ9imQ/SJE3RvVpiOstFSGBtqE7KzRIdq8IaDhsYfGqwG3vf6oRTddj
SWl8sdB45VikewoN2HA6aoxl652kt5xJzNiG86QE3+nL8TACRJyxANUf8YU10Nly
INANgvNO37SKTwRM2s8ufccZn2HaqsTZ3/BgJ4Q9ekt2TdRxYfJvVLNkZcNp6wIv
KTrPLGmp1a/vGQ0x984dnDKi/bgU7wulC9XC5b7EgwtwbUYcR/qNUs20Mvusr8ad
OaCJq4hmWbkgu5y1fKDV1YD+zIn0suw3ZIXZbVGBN1nVFGpEKLUcXnSb5tFoy8U1
vaTFs6mAjsU/GCUc8C69ilmIKq5MTvg5orMnRpkwWYccS3ygW8Fy4NMBRRCqiSyA
y7mnrLhUesY+nPUKNCMSOa5etjaq1iw+ZtplwRdBZKIxcyYyJVdJBYVXAnyJCYwA
NcPI6jQne9XUa3e12acHXAsdE1eh+wvWZyTMrAvLB+tYQ4vJju8eVD1ZzTqzjAwl
YmO59ndTecelLRHIc8IphUtba388l4+z3KhyFshKpc958SGUbvm4TT5baOlymV5f
MN3ItuuWC2ggX0Y6GoiKHlHnLcoeGD/9Nn8gmKaT7tP3M9jIndUztnKXVRJIyueL
PBdR96SlAKGVPijId433U3raxXRi+E8iRj+ezCJduaTLgD7DkzU2Uwdm5qRPSF5o
9xbMzKy4n8uQ75piAukvMONtEs9dJ09l6WByHPHo8L9fSIXrvc186C3caBEB71C0
ZP1dJ9UmFsXLltzXkKX6SSn6CZ4wJGe1MY6z0c28YV68Ouyh42ZBcAp9xxsKyVi/
S8CxnHpUVTuZyOqZ8ptAbnMSMrovbgVcXnODUNLgNDYA2HWlQZq025UscWMZlBYU
MNiAn736xVRyMPH32DgBGo9IesY6K/spxB5EvghzyWJSUGk+NOrU5L6SYjtRtovE
lj+nAINuUVsCZEYYEcmNY4ro4buJRVIaQBj+vV0BH4lAc8aN4jjPwpINXeJsOAbA
b0Okguzfd64ZWlAlgYDUwvLWhm6T2RX3TAUgWT5rNcbVeI9O8/RUvSbk9Mr8F5sT
9T5XT+p+2cUOUd2GGeYH9dG5ZXuBhnP002FqthjGDzE7h2KLXb4bibCbXiFk/yW+
gUat3vMLI3K2DlP2jmBYil6U64wwGApcLu9+ZuArXGWc0pT9+zsGJdphQTX7zZV1
EUQ0f6VRDddikfDDXE7i3Z1QgAmgUzI67ooatsUlcM6A/YehbxF+0u3zapWq66ZU
/j+JBZust/r7ufjBo/c8bJRS51Bts3+Mfrf6crcUz6a0gmpGnA56k+Pzn7A46jZB
8ZgDtbDKCEojIaAroQSVvllohhsCBI8YVaSbBo0vLlOAKKlGBwKvbrcXhiv1vbfG
AAceOCgP93Mwc1A8JwYi6AzRyz4J05vKWBNB3GH3FPEVQXefUxPk+vtyKwWruWjG
YX52vDuUTUtN8E/UPbIlAtLwLisc6IWTLYO+XlqQofcd24fbOZU/F3hkCYOQO7pI
RKLyeKSKMNDKwlO8cwfQvKP4uKOQirQYASgrJYPPoArSVpHNtS5rksCaG7RWQfqd
6Uf+o0n/NLzc+CEtUmvc6V7rOHF5DPP/YUn5DI4+zW8VlxGd87zM0sfSIf19MOon
c1pnKaC59w18svshF3bPOpuw0RnDNBShD1dG+G6+Rz+amVkQ/ASBA3sjmSchzuSV
AoGRk1ckyVfPWMuTTj9oAxWS7clkjVsxyBaw8CzVW/IOZdpwEa5xIFainhe2g0vU
2/4WSw9THaK4CXQMRSEA3JzD8ZZbczukPduau79OfWkKJotaK5u2S8iuER0e/XYi
Xi1KS7tCQIergBmQmSp1o8x/ccoUEdsNtPdImgawIGvVA/KTfljKzk0fZ2MiCzmU
mOPUyT9K4+Z+fnTyfCyWEwjJxbzkFmXPW+6NauYwOSo0q69DqlX+2d7Wdc4hyiGx
QHAo7ad9py4pLS0KU5iNWxazXw7KE0/xUcTsopKMISCvmDvHYUMyYvwne90HW7CM
rvZwp9yt+TDEigIwbE6Bh1+MQ07NEXDWrjva2AuL1U6ON9MfZYPbE5s609KaCCBw
r1hW+DuNd+QWtnKPSMx5wQ6G1x+oCgNI4HzR+462B4WRS1VzIOKjVFYMDXaZAXyr
BMcshHx9glHYkrNd4L4QIgP8S4L3UxRFakXd9OzB9sYA8nfcTf3SU/47OVyOyr+K
yZdYwMbU7boCFD2m9P/OIMeVaV+P/DdQV8zW8oT1PPP19r/JxRdBolfsXtrbSEO4
9vGARAvLkVBDHLZb4E1CXSWI0mpngqMS6ip5uTG69l0STUgoLiqaiaOuHZn/xLfy
/bRMWC37VDVG8esm0N2JhfiWj4U1fJyUgZOEnBzYuaM/HIuyPg9Dnk0Fx9ns4Kvb
2R2eot0wfZWJksRq3//SQuiqlKCdwXf3W3R1a8z69+RZ+Ho5KNY6l6ZDZJazvkCG
wQ1TyM0fUhDrLiQqf2RGDlCF3qXWmPyIM4b4VK0zucr6vf2xaymskv+5dlwqgvKs
oJ8LUZFNJ78q0s8YYXJOSTQoB5vIc5V/aRbNmsHrzf5JgBvVJqaH4gB95u+9A4qN
0/A8opQ0VvQ/sj5molwvZZUw882Czo/9XieLkI261ciJxj/ncrhY2n4fY7zfSBvK
FgxPX9Pd2U0dJsLFRaabygwsuN2PyaTG8tE03gVpHDpO8PgdVffbzbBQEWHR6cO6
MfOCK/xzMEO3R6s1mIn0v/U4jrGEK5GlFwDBLTrAoDo=
`protect END_PROTECTED
