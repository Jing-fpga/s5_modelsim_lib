`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zgZSVYUI0JG8AjVC21+uKIooXcwxv8FbETXw6fuHov9Z0CsVIEf7QIuh6h24JN1v
bqbUG5s6fO/tXDW49q7+JorSvc+mHSXaiyjPDgu6VRfGiuWOFuYcNLv/1RyViD+l
HeRX0x82EZMrCK8S3y7+fdvcw/+pqEArk1WAUMYVQvwtR/Zcmz0W6LdZg59c1rXz
WUm007qYd2ZI+x30MeEWr3OupnoE0+3KQzdbqKD0D7QKj7nXe+BfsEeJc43ahi48
Sz/mR35DeisJf/rQYKO22rnA3pRvUIujl5gY4OKL9+DqgcKqrBHUulRynIringa6
AAmdPmEvNiHf4rgtJnP1hoWuL/02ppQBPwg5HUUHtYYn9YYDBL4Wctp2Zhn1ES3y
4Qnqr8UBoryo+4Wxcw/qx+GFmgpQcfC+1Z98WDZkTNsapuBTqrycCdHeQcAWYSOm
lOUDMFg3B6/93QYnkdjKfKY3XeOC2zZRGPlztJH2xo4LTaJ/S8MOqs5MOtm26Rrj
bzhDOGEwTd6S4FV6W8f0j9kFztpHofiuLWoeKDyU4bU9fM7wifwV/fD0BU+cyCxZ
TkvvCmB1g/LpCuWhsbgQHA==
`protect END_PROTECTED
