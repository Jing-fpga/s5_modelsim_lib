`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bxbujrVpW/xLZqFJ6xxAerqMHUiyrU72Gg0vqUwTvYiO7gVBPpOQ0zDnQBFRybtq
r+sSLHKCzXLwIC/9VGNjaBTkZLphxb3kLiA9kOuez+kQYsjEtepp3ENNRaq8SycF
2ka7o3lCXluM8Q4YmQx8gSWES6aCQGQq0q3EYOKPDpEZdf7jikfM2SZc05OHfn02
hrMYJFXS1DXmwPdIOsBf3vAPwGK/CGFnBCBuaW2C04nlwqXGZHzfxPvcA36EWTap
iLYUbZPgx5zfCBvENdBEGrCQbsZRMYf8mVqrUSOdz+7MvCdMS7vXLhmog6e/VERb
G8aIJnOnMsuRBhAqAGqvqAJmA+GgM7IPDdHQxX495qeQKIoOSn9x5iKSTThPqqJd
DEpLDZEhjTlBqS4Dc7gYCiQLvDtrmlNkRELSh8QpyT22RDCOGo+BbmNw78xoa218
5cMBZQMwC2gkFI3ePfKmLFMhRXxacQmi3c5LvzNN9eOiB2kKzQLbYQaMG8FW283R
Oky/4+mvYloXtmkY+TQzYSqAsrFkzkdHqdOXN/FswdT98m5EX0UY/ahp5FKnKW11
yZAy2mP8hCqP7Q0GjzczQGg72zE1VilYLAHoGnwUiRC5nYsHtVBcrPSCqr22lf6M
xtuul5bdkE64CeduWyR11qZCW82LV7o0KqRS25P0gzEBZWkG2H1yz4vFBtjZIDbL
xhVMIamsZoRX9iivQQTu6KJ3HHgV1tINlIhbfDjMrDwsbsK/qJo/jNTw+VLie5AS
50qywZs31dnmncZP8dqR/IYNPleiZr8hOiqvZNQ+jbge9dRPyfdIreIjWjcLbLjc
VgbaqnBDe+9znoaUeGC6IMeClOXb07Djj9AX19LEqa8LocnLW4ey2/v9Tdabl3FE
/cWKnjOChJB2bSb2isi2Q+nG0YOyCvF+EkzV477+rWhsJ/uwf93NwFEnOyu0Xdtl
ZIIaWycNWARJdOQVCNY8o8qYFqGs0uV7EvJFirosZeNOnnTUG0xTHLkEJy5IW2zi
tlVpPrxrdnEeCXDiU3Sl6EUKFWdUKlySPeeRTjUVBjr1H7rIJQMq++uKBn6AY8+6
S5kW78BxdGXhtdmamchroLUQbQxEpfzm1te/8XyHf6BVQhXpdpBLmqCrXpl3AVBV
S5dXy7N/GlK1ZZ7wN+gFpNcCfPECKxiofzwCWZaHxNJslIXq+mj8k1TKgIaiixYl
zUUC4XHrYPiKlkjLzqtHXKmA2NTVJhf92A0SsLip0vu1VDbypg2FRq8kJn2VoThF
uRBuQNKBEUNIa62d0CDmrY4qgrw2jJbxVV29KVM/Hw5mxLGzaNlsY2wWnMt1v38R
`protect END_PROTECTED
