`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aeBxFREHB200r2MchYazQNhtGZAbCBZPoOuVcoWSYI84He+UnJ4jenuUQX5FuTrd
92jQHqAX52yNnNMEmAvXMN/ytWXtiiPSJ2p4/Fd+0BMLHNa2x8qqOOQEmJ/HN5qC
CurET+IAeKt04s3G03Ok6d6NglYb3o3jVbtdbjldxElT7yAZyt9Ktef5pOUgYlUt
jjtWc09G614xKuXImTjgabTQ4d66tyNtfhhibjP6hQfmOSocsVpH0oMclF4WU+bU
JNWi0pUoBw7lvpnSKALArZw/Ti772/CVdSoOvE2ZiZo0m8ZWG0bSI9Qa0iSD3HVG
rJv95eQPhxmD8fdK9EuxQd4xqJe/srmX+cFDisJXWIwQW6VFxEaVn62Duu3GZzFG
Xv4/uctqVl6Ns/TojA9GtCFHaY6t9KPERfM5OdUG4dyWIRn0oswlsw7CMcOnHqnj
4/kqMamNOLzGORv9sPn7aLNF4GhyFtFcXD5wSJiapO1qtDNmZyc8kQ3F6YXHDPMf
PAMAfVSowU1y9xz03Jcnp5xAeju2fnsE/6AYw4XRrgcTv2pdQ4P8xZnKco20+KZc
2ebTUgWcbjdD4v/Jvvu6r8THhyz7DcRFXPYVndC02QtpWsZcndzlNHMjSfIWBWeJ
JgXC9pkhtzJJp3Pzk1eFyXjLR4KcZR/BLyUtjGYaDWVCuoXjrg+Qa6iTc6mDwJfS
XMGkiAAlr8FmMHCZW+FAc/PWNu2DmYXpsQxKn1JrDV+aG8nQXpKmtyqP7+EWzN3Y
jM+/WQnAfEcWfkcksR2a+v2SKjzzGt2VRN9E8z7GD6nqQ6xMFrV3u1+tea5MePb9
Bjyk31MOkyl2OCWEiw1PBEUfuAgzebuKwP/5LnoCRfl9Ckc1pEJTbFlu6UBbkwK+
EP8rcOA23bAiasfbuhHWZ7PPILk2nMaNtUEqixIDaCuxc6l48fACjBZr7H+nTx/V
DN1JAXTZkcqmGUpBsLcY8jPuLe6Sy5IX35XePVce9pu7GJ2AcIddekSZYlrKS+aI
//kZY/vTZ6nHWtjcmroxa4VKSq0p+g5iT2pIYv/epSM+ffKHcnBehe2sdywEVlkC
xInLLAd0lCnWSvcfFJHAc3+0HQc2EUu4lfnr9AGahYd9iV3wg91lR8DFtCTWWlb5
BhvlMuffkznVRUPXjP8+aRqM5+aqMyyfUwWoSGuVbjab3JHuhgY7OVbzyKRTdYa7
MKAmCKaM6TGoxhm/ywWbRuM17ALRM3rGt3NoQHXGhQH32Ejjsfc9YDFGGTD44Iw5
kHODmabH20ZvwKbft7r3hoMrCuUpGbwUixVcQwk7cykNfpPkAYOKRVWyEcqrXMBZ
mrjsYSehWfedAoeXbIdXX0wfbZW0bSNEkLTNA0ywsqOxrPPiY/P2P6k3Z4NGe7f1
zkZtXYKC5vDCCMhDUbkl+GkquAAZ1YyipFmc+VZBJZip/7uKwi09sVx/6BY4Zh5t
jT1Non27Z+d36uKTHutXkFheVRDFfXvvbJ0AW0JXu1sSGNv1eA+geToecOTew5Ee
O9zb97E4R3jniQKCfcsIn7/YiUYK6ghiEsJcD6mTNSMLGHX4qQ8eM2bO2f8eUjmh
esE6i0cxhjrAPUZQ/8ro9fnzGunPeTIAqJGa/VlfJcp1jf8rz65Va/nJ8o7wo1B6
9mTwv4a6Jd2k2+jJU6aMeNcVzps02tWKuQX0b+GIkEN5yU2Kadyt6ILWv9BAr9S+
SDIp2OOpmcLA9YqaM7w9HryLcttPD+KEKxzd8J3r/P3yP5e5HCMmFlpA49d2QTz4
tnxVhmOaBE9nrQAKyp79sUkutwG8Adr0V45n4Vif7D/WZo0dRo46KR31ed31oEWC
`protect END_PROTECTED
