`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VbFd/wvoFG8D2pUtEXpJ6qRx+ZJ1CnMNP6YqkYiDGYt6OpqMYk526EOOam40pmzu
SuWNC88gmx0RuRaYztTyKPPwwTY1bTKIufwGk7KgsPyxUvpahXAiSov1q++nwVDh
OxmiRjxJ7OaPuPVCUXnr5JoCdQWn4kXsbQZDL7WmJqkK2r/PhIougsnKT4AOAjNs
oMmwliktVvGqBI9qZDUpD1j3+necZJDJtUAWEgKoUAhiEJk7VJdfxhRsMh3XNwgP
EQWWEZk6k5EjdvSlyJEqWeUXcqrhD++Fv4zdoxmnuPMA6wz3AGlzBWFEixt3K2pF
AH6gqTtGRKTUCJrNdfQLi8hlzn6XDxereMBclRaTRFFViqDSEY8cDkE+CgDcYQ43
vIPBSI0nvs0R1NPXoQsGJJD46MluW/KndeXHrXjifplGN9I3603EKqA0yeCn0thX
xu+p0cEhlzRpydMUuS+SzucL+BKXYheVEPGZ6fBhrWhs06t5/gYhHh3VkGsbu6Uc
7zITFOAJysQ4V1Q2x/xWCC33f2JLXWijqTxV7+MAQnGrAnLXObEKtkuZ/J99OJ7W
zqISiW7R0K6i5G6TY5sstMfBAOSR8EMDeaTl6B9gjlbMK4QSzvUVjREwgEX8q2Go
55VRF4WzBLDjaWMCZjQAvyxuNinDcNiuCuIfQ1MCf/fZqJ+O5U0Vj83lWIG6bAWV
EP00X/ObinNYj2UN33G9lXJ2oohOyaxbqgHGbRAdWgEFB5PF1QfiPneewZNTZgL1
NvSTKJli63emwSfMKOdmN5g8II4YCFlyihLKng37F782EtV7/V2W6jPbC2ZihRdH
9eSVU99wdyxjG3V/0Ll4awb6YZxMyXz7lqCiSwU0u0RW+ESq3s7S6AIyp+IoDskT
M3G+KdBsvz9hwomi08LPzY9XjLmmeJ85xytCV0uaj6qbualgOot/3jAommNdQPcQ
yet79s6yDeI47rr0kjkK45X0PkLBEmMbLbcgx5fxGPnVKMYhvbQoQ2OkT/D5tA3Z
ohq88F/ZDhzGPvcTwGeqYlF/UFo0Q+mrM7uHzrzcNgfSdLvMNFkgcqYJOHd6Wotf
XwHJHGWZEjPIQGraAKN4Q8cnDvhHsabJwEAyZl5FlKMnmr6qgOQPcmQ28L7do11v
Qpu0J8uvVtt0KUBjfSiTpaqj+ROYDUs3SteqttKVPcUQjlAxMObRKSBRZGMV1U/U
3ExpTChcYIHzM8S4pthRafh+PJhCB960i/buhJ+w7Zrfffd9HY62h7HDGYiz5kxn
0/g9g3+F+lzYJdR33bryw+1y2rceOhgKwD2v0WhWqnQBwo8of3aCvmK/jJaWlyMA
+35fp6NvRl+1lmyv+0dqB77L5Q6ssfm5AhMokR7cy5/JRO9USobZlgzz+a7XJFHA
wzHJpOJLLZ0mdOXMpxc4QziazSUPq2/fApvVGCkmVB73v8L5xKhxRIwbCVziiGet
oFYAYXks4OX7AA6ai6nawDejApO2VwjaevPfTqKzJUnYVwfpXH0HCEg1WiG/ZRWa
`protect END_PROTECTED
