`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ALmdeOsW790OeO5uyMiZufU9GJ+tNistYA5Vlgkmyb0//UnHbFJo7e8Do9zp7+Ss
mNEi4LW9CUCUHB4TfzwI0Ao5ztDNAXytOj1Y0e5WaELgZLLEEl5wx03IEqMqHUrF
zESLmdyl04/mHxd11dh+nuBFz64nPAA5p32qj9jPw2mLXTbpbxaqY/it+K8e6fRO
HEXEQnjcGpWSmYE/SS4UlCloHO6sDUOZ+oidjjc3Rqml/7IwfT4FkX1QgrGv5qxI
LwxYfwCfWlFDZ2g34HtCcMSt9oXO5YOBi1pIcAIppv24d/hifkN2AeoDqNaP9acA
2+BnVS8QHYv4hcK5xVGIQqalK/VmWeOqqfmAGHgDJ2zMXJfxpDfMOee/NFpPye6C
fkYunF+ruMmZPkywusy7mM5+twAJBMtHw4o7BKsLECo5VR+evp9lfm7P+kZluBvv
zXTa8ViIuxwY2A+ASXyczUYCe3CokZ+AsQH0d9sn6bWqPh3y8+rFY4ThhkdhPqMQ
R/O4HPzvjx28eg4pYJkw0tjSKMhAWR7BRT8pYl1+qiw0vam0D3LJ/ivLoKaiZ14K
3GJsEU/XO9mN4NcsqWwdk2B9iW1PANnUubMH3uuoTGafYR0EFLqJ2Q/Z2zgEaWtU
Sq0iWNpbMoifaFYMP2VFz/sp6d+sSLBUeAQKoFraaaPK4gVI5QxJrU88SfXTt93K
npWFW8dg2MMekSBWLKSlIRtV6W7isukpwYcritceGBEas+z0OIH691kkCWJFtRbM
B0dxQEuRY4gbufLRsWH+ix+5XCsMnHBLnHzK2L8517QZkWo7tSqwazThyMPisRIl
6QkSsmdULOpiBcv3vfSrn+s53/+Vzjsn6HMrHIUZUges/e1VKkeK9wfGixo0rXud
h1001YfIUeIMyWApkuS0rOzE5ypkqRLTEfJvbqdCc8kpq2JbnUobMP7eWdYI++Ef
uEqsYB0xYZXLJ+1cbgrZ9pqolZS6G2sEk7u4r+l+SkOcKbT99TVaanojll567GEI
sIdMAS6A0Pjf5emv4oJsyaRnxDwvWfBEwlWbShMiVFon/Zpb9GNVY3Hr/efm0b4i
SIgIYnIBiSLPgSHkP9alByWZzjf4BgpC7820JDuuriENQFWldGJhZjjNoHqjg77V
E0xLXx1coePgKjTJU3JCQZR+5e+FKYCUkLn9FSfPI0xlYAjUtuziN6HtsJl4imz4
UGyz1fDrxgzNmjWFyX3RyaAdZMzIMSok5DqwUEFByv5k2/LP+2rtL6GqatCYU0L4
Nc54JBoUuidY7oB9BwAcgjQlFPBUaCQUCaq4HwYNLSeyK1ecsUXdxEJ6lk5sCVsC
UEKGJvP4tKKrNSo9Zpl5JLk4EGe/KWGHdO3W78V3ImUJMZZUigZfmT61sY1sw9Y5
evYIt89Q/vagdunZFa/XiKpmZDZBgpADvTn/lYSaepWbGOmNUqKqohv7HcmpKd4q
ZfQW1uZQUnMq5pFzuxlBfIEVn1G2tbJ1agYpK1ZJxBo85+EEtn7L/l1iDu2mluGs
r2rT6Ol5rT1QDh9BR2gN1jwr+0X9ZNaan01SKaAwTfW2tSdAM0cp7eJrYcVqDI2k
VvJOtbjN1yseghpDwOmpofa0C7WnKtQ060oPxPotMGawE8L+wlhB9JPTkHkmvuOM
32HcMn/J9fd6VHrZehlqcd4Lhx9TnmFl5swIZt6xNiW3/QEGRVz/rRASMXigwK+R
JX+H8klYTHtwMo5Hbsuip0uCubVL3eeROBk8xoZOYEIoPjYg6/TpmZolmSwaUgL5
zwci2lySSiC/RzGJgQYUXpv/OzyjqXqlNm655/GzRiTAq0AoJo8MKhhaMAVAkESw
gz8qBlBEujfciw8jmVfDwUKi8RZjSYJvMJdISnC8jydl/K6f/twO6HQyVg/SUd3p
C+s7jvwFJ6JG8vmsNuIxX0hF3tqiyZQH6MrPAB0lkUloaXVVVC6MDy7+B3qpnWc5
dxmdJDDXTj4BqOxNLxLaa91OaNUg0M+pEFrfejAupLr3Zl7EH2ySDh0Wbwydy8Oj
PNlQPsjQzP/C7PCBv4e4N4EO9VZZHOlmRqNOawKkOzKBZ9glRcYH/gSu9nTCC58W
o0TzIlstVmF/1FGeT16YCLVUrX8e3bNzfIVObNy7xSHOzHI0Ph6Yt693ifkJe/RG
UKrXzRSlxAROuMV9rkvQvstZgXvXd6ko0hqCG8KRqrIJzzcBLJJWx3VJuEuG9hDC
KAUl14/CN+7CuoWLIaExG39cySP6X48RaQbbvnwK3Cxte7U7S3Nc2obMojgQ12VM
YEew9smy6Kmu3EHSlnAJz4sqKGNNwb0YQu+3cvCb+8pmwZ/vh7GHZw+ZEJdUelGI
ITzB5h2vS4spZlxy1/9jXH+3YiBS5OgKUrMJICcZSWCH0VoqujgTS0n1Pq5vYCOo
z5p8pblx+wJpXFnXhMRjsfiYncjAQSVxBhiPiRIXHm6aaGccFQICiaYIN3YjeXLz
IkcGcqNQ1D2sfJe53bDkC/Mjzt0k8XwiTBBKWCgiBq9B+u70nfvSpiAgJRKXfbTG
57Wgrs9nz5uA2ikb9lUDLCQF2LprY2GGfajP4R8dYFGDdeT06RTNhwloSann/d1w
2D4yfuldV7vnmhyG3ifiBHvZgEp256nCZtYFFjaKXnAQfa3R6gwev1Q1RBAKyJm8
nkZPfjMRM5Dk3q4wy8GR3G8mk0O9ju3Z8iuVzFzyFuVnmcC3hn7l2u7vxp/vrwMw
WB4SpEjflItLdnNK0miFSJUvc1Zhg1Qtsj3/YB/BWFh12F784H2bCAP9wM3vm/u1
6Dsc6HiNZc+l8HKEuzkB/I/qPhRk3sWpmin/6VubDAln6iOk/0Rc3mFEuGSKLECE
JgkaERokJbq+VMcIvp7nzM4+6EuAlv1cy2wTSyod8qxvK9A5zuAtsACvwuhJ7qvw
bGInZefP5T3eqA/eg23bnaGea1GG2hzGhLffzPitcbC2Sg4WIIqcMLm3Ja1ZQrNY
G7KWXOyU++ZAGiq186bXydNY5TARxqPQUhaxUACUefROZDSzKnL0olGv40oElD2y
pIFCalZgs1CJMDeR1k720IpdXMaQk9vFrrXwl4rmmUjscOAxX7z/paLvJVaWWVc0
Fkjruva30IE7H4V+2VtjYYaUuW1C+mPBEki0nhxDozHEjEYrTez4CFkf6++RYBVE
YD6yXBDQb+L8uxE2K+O7Dq7c9ZYPNPxz1FZ0sMuykcE0qr2BGL4c4ypIfqDjGwhF
CNLVldhGHiVF/4xplQCr7t5N6kIlxQ7Ebl2JVinm15+bHdLArtD//uTxl3DQY8XU
vsGRfA62zJDZjxEIndwlYNEervt0TQaNhGLC2wxPKb2OG/CLnkDgZK5cRWJqN/mR
2NiCQlnx50r6PHa5jtLKVYZ8CGYOPVUeadMrb3X8agNbuv3BPzEfF5QmI7ysqi/C
I5CQHxwhsL+SDsn3FeFxllyGfYVglZlHX7ReJodLzqfKKVWwWV1efRDovl9x7x7S
hQ3HyQuKxKhyqWzdvnS09yq0zucJvTQgVKGdlH7THI3MNaIK4V6RdiTfSIyFGnFt
8SM0bLSL2NRC0+S+fqMK+/FmGkCzzJ7n1qknOhbOwnqW6dRGrNsfkPY2ydEQjItR
HAuBETzlic474gA1sUM2wV5z287hiuJ733Qmof/Bq8LJ1Iy2S05ij9Vk2bEjeB8S
36vydWyxM7rfyyhH31S+zcU+8RQVjWvgJ4odmlDJ7875fnT+7I0xfhOG3TU6dZ2L
qnjG47EREwbeFx76xznA2Hkqr7DYP6bfJDeJ97bJFk+zKbIvzlPBRvFOUuvLOnAD
5PaKq4b6CltlKeMk7g9kSWuR3JDZEqrpUQlM8CJzy1ioUBoffRyuNSRErRniFYfL
0grI7tMAgKq8Xx1wTDlNXmeNH2sWXK6HaQc1Owipt9VvEdK6nv3HzC6ZZmnPJJRh
SY6bYKDWg2A0/Xs6aMrVpJkKHSi9fdQXbLc6qd3Gp32gDjFHUhKK/TgJIfKZCQ+F
lsXCFrH4U0PjAIe/Wx8CQJzYjgnm5Q6e7DOm09KKzhqLrbrW8ee6qUQof7dobfJL
/ELwUMQtWjoI849YIUp1LDLkIlcKN2BDH1GasJ54KJiWTdxWOOivjru5NmHGjM8f
xiXbhR3elZsXOgTa9mNxO1xn5vVhyA42e+DkklT1/8961cdFR0MmNwfsR0jYSBKu
cL7BJBM72cCsBQN5RKNnohy75hPz0RxP3FAejZ1LhNXFn31RoPiiyi5ix8kOtlEC
7URYeNJog07j7dIWmO4DbJHMfAvUUUvrqdSB1hQvGwzVJKkfFVO3S9Y+8lxfGDec
xwYfbzS419uzgGLpK69zMBCWHwrtZdwOWl0b2hbWyL+yiYohxARmqMMFX6FX7Djz
84dmbEdsYyUP7qMkwLbgFqxjpTqgKR47M5iEi4/JOWj9pZ2UOT+TuddMzkpiNFKw
Bqj13W27CxBcBvJxOHLBOATJPVSRCx0ls0uWP2aKs/53iR0OQzLEQ/EcUllKNJ96
XNAlPh+E4T1DEAKKm00LC+64swjXq7FfqKCfoTQyjZAyFbmGDXiIGbMsc9NxsM3r
cMXommIrvBIl9NeEY/jICr9xZ6/y8VRmGnFe87H/YnQ2bfH3DJ2l7YKTKOqsbscs
vdjjbw2aH6ea/cf2V6ELvNn7gzwAbyLDLNeKSBE8aa5g+VSDwSfyBKNznXrlVObQ
COfkQO7rw+hOWnsEf+3U7FRfcccHNKiwlAcpjtj3Fw4J6ijVtCOCfvtv2rVFyncY
0cG2gzH18ZYWR9crRZ86H54YNAS2MvvEV3KH3sygYLMzTxdB3kR6eTF+qkxBk5iv
bGFNfsiJ6kf6SXdGc94ZSR/tAmCLPPRdRPIL6/LdtOxiGi9v465Msy/xqCd7JY4X
U5bJh4BRYmU7SL0GVCQWURfH3vAnRBybS1ggKdf8k4stWFn7VrOjgsuscp9Wx4Sq
SSahjYXdj+tdR0eKfaCCrl3slWCGNKpHQOKBUwrZnaORVzAPVr22e51UWwEZwMXj
5q4e4x0WMT61U6qLkbLMyNZjWJw9rArkbDImuaqf8YIdeCa1tjvR3HoXmSAQTQws
HjV/njyD+5jssgYPaNVf8G0XgjtXF98dBHdhWYOBf8pwmnqldrJ5pWRKhwoS/1D6
HdPLXGiKznQkzuofDNSkah5YP/Ha85L0h9rhUWz9JWUhdaf8vKtmrboK3VkzDMrj
sYgQL700LXolBTGJoBUCT2AJ4BIjeuBQ9TLAIRbCkUN08tcfduRmSpWadHdR5lOE
wEcbKTVRxqadX/ruMFoZeLgcsYuIKLu3HFK4+Ig+jneOCqq+vbZtgK8roRdSGY4c
aN8cP/BxQNiR3tmT2D9y/XRRaIhAmTXuvXSsZjt5BASrHLRfAw7GkFiurKZHxTeI
zjG714XofdwpXUGRRGLufQO8sVsk+n8n6TkBOugeb46nhhSysDRhMl7hZBAMoCR5
tOhOr+j3Tvb/abK7MfUHX3OhLR0+BIeVBxXR9ZFQ8p0AKp89I8OY3rCMzJjWef1j
+B/w16rC4WPFcyRu7EGkUOS3WZokMk7K76/+/zYcxhT4l4rueud77Eu6vG4PkdSa
DDDQ2ujPUE9kofjWiYGqZRc4F6kQFWqEYAS3QTESgAlFmk1KmAFhZ+HGLdAlN1FQ
YChpePn+xn5ybSl/X9zdbsf4Wzn3H0z+hMtJY79olJBuuU+sdFApjR2DkOpMVutC
Dsz9MWVtVlj2ZdTnsrN6TD7Z1RRvzh3eek7iHPJDsSihQKFkGpxNQb0ALUJ6pGeN
AgR34nA56njITq/0nLuVPx8O/WgVMo0uULMOa2qV1vf93bF+m11y/ViXsIJPsDbE
aOMnsKh3yqBdK4EWDSHoxA1NxD8QdhUgcHuT8ayjO/c=
`protect END_PROTECTED
