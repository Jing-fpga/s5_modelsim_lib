`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pug9i+wbXP8PaLV3qbgl4zbVnf7p+0638jsUE/0EqvWvc5eazLoXC59d0BQohJAI
FneG9QoplpKghprA/0xQx+Xv/uG1rd9uefWFmKtBMl+bCp7nT/9JRj4sS8lQ5myo
7pCylBZREZyoPHNDtFGsuOPpMsTieqAb/rVkl9h/mNPV0skd8jq5GaZOcOXV8+rv
X9+yQtS9rLjfOm/+gv8CdTCZb3COsx3f4jsL9RZoeRM34CZUpn5WFxn3KiAiwdm7
/fYDu+NKASeLrLCLAhvaRCHtzrZlphtz7Te8Cgwq+CjqtslYcyi/Y5U6LvceBjD7
2k6OsvquyeNS4I76cdNr0JTaFUcnhg0Xzu98djQOlScC+UpdrBL+RSOZqStJDzHo
r2Zm+pcv32cSVvTEQ9oMA2xrrCYHyl1eK65b/ZyARZbWBRhBCkRGyzcC1ysvXL7b
UYKuGlhGHjMlQmrnMNQahR+Zim+wSGa45fda7XoEdgIRiYEI6KfYo/LYGbA3HkHE
R8M84MKMcEfTy5b+4H8dXS2V8ecGT7+xvRJVsK5kqLZ/fiW4DD2c41sGXnrd4mYx
pz9MqsSYZMIHF43SHzJDklSlv2CdxS7OfFGNypOxaMUoNuJGrBqLHgUcHOKJEqfk
J2FcOIdS5P8tUWty7Q3QErPyXpLVY/G665JHMZrG9QMAWKNDGwhiZSxg1gAuLGZB
5PVbeasGP8ZShBlvWHlBxCfhCre5O2EtCgdwmsenWYr777utueghQkW29AwJLyzG
okiCRQTwKRn8KAuyBkL3qngkhBo5bTQRmE5K+mduVn4QFdqfPfz9vUbtd1mE3T7j
xjZly/Y4GSEIq1BNiClUZ/p3EmoiwSSQb90qLNkQPMP/XLsYPvafpAXcku22+fPQ
CXcEDgtlO8s6PSLxpJXGPw==
`protect END_PROTECTED
