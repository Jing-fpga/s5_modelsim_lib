`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EOzQ4FRbJQn5KPUEwQ7sdD6f4ArSgUNj/ElJ+qzqzQk3w7vg1tMO8JvyjrzE9EJX
eF92wWcc6t2LBrDeISIbAnxxIqqr5hphcofAylQIhjwPMK8gSnkrBJN3RakoOIZj
2NUFY0MzGJ4KeV3j/mT3R6dGG/t3xPVVCr0CT28NZwrBkD7QOVCHQJDDf2gcCGEP
o0EHJbGXB/J2uvSqmTjIt5C4OTQ+OFOPan/7QeFKFSAKDrzo73REXb+g33p/V+Yv
CykKBsM5KyVwrFnCbWLVWFaS8RDmyDabf9v/4jyHQLZTkgzUqOTeBB7y25AcMWg9
bE+HmIZbcFUFQ0r0xC3Df9v8ZGpyREvmgko1/UUvtjQfXgbo9LHhHL1anCcj4RU8
oDF8yN8Fh6xSo2g48glmTZxRfDCTCgw0kMU3G4+zpRFU+wPu/7kuE2+hjxXZDjZH
hgtjTwlZ9SihUVIFRcjgq/59kq0WmD+X5hX9Il6FPVnSiJldrIdQj9TpR1+5hDMF
EwLKZ/u9HprXz1+0HnQjuTad2g5bnK7eRKaL3Z8NH2yS4t4wEuPomw2+WM9n+wkp
yA1G7SZPii27wOXDY7Pz3IdD2HVZm61yXGvxOJDjs6rT+VpF5MPh0Qz6QHzJBjRK
otF4K/R3pb65up3YbKG1W7Jj/72qWL71Bnr+Sh3w3/jZyTjmqyWCSE1V9Zr/7vZm
Y5YyJab5x2+4DDgLgOGZ+u3lLRInZoR9KqtbxgZR0yM33jmN2AVKMUC9kTCGYdWb
Ym4UWxB/PRWgAG5NtGQjs+FUIECoK6NsiH1iSMP4r33kGuNcoBkYkhAqOolYH2tS
acdKfN/819HsT+X98nsxnw1pzlQ+TAW64acvXMbZkB5O/VnZM7mWrW3seC1Ojf5v
qRwWeVsTWQL12W9zyEm0Ferfs+K7VwTw3TwAVh9YnNpNnsDG3evaMkq8L5T2gY7z
TDy+2usMeYsE14YXYO1x438q3dYxHvXMN2179GGljlrNnh7dcoE9K2ai72CCZIAF
Q3zkAUfxyOggkPBIPdmckMAUJdLkar3i9DB3Z5FeWkL3rENnDizy68Cft+Tbau77
o0PtmtQrdtrQuyCzJO2ICHbIita1tamwfhfEy4UBueHodRYjSHe9Gkf4Z1UqnRX+
fmP3q9iIL9e5fPO+ITAn2RpcMkWnPn9iyEz0Fti0V1N3xgh8edEAQRu+sRWHdk0g
WoEQpJ6xxFBjbx5RtfBLEBMaFK6aZ9KEFNb0peM2ECJSKTaJddwiiWRSX/AaU3Bh
hXgkl2xaybq1bV9Qt+8sFoQoScIuOW/uw8Lp9ESxLhgk8Oi8LB8nePtXWKICSI8C
UIH86dyCf0L0LJwEfpyGGxx/gOmZECRmr/I38jVHln8mbnpDasLqGlQIxtO2ATU5
NeG09fQv923zP85HoxcG6mzyygzXoz4otc4kcg+T6WbCnVxryIhZ02+0vdz3OiNX
4UnemXf5ZR9l998lrZ3RJeD+dPIenH0ra3BBxYuYSzg7Gg5PJebgaFb3+PJtJd83
u4qqISKTbpCFkWZesOQmR+DRCXBIMzBSN1x9KK7l0+yB8loIqe5eCEXfnWsn1Rpn
KKZMpwnMt7QZPniFHvEa89ELMz9APj0Fojy7hSJ18xnS8e0iAkUeGVdFMoOpJLSn
3xWbe02lX4j3q9Z0RaPTaV08YUJzGW854OB/5QmIjp4ZE4xyqJlkJ/THXOOTgQ5x
moJYdnxEIV68csnot45sciwzZDaJzB5jFsPsQpMAlt1BEOzrKSR+4cYCJqWve5rQ
nA5Mu8iLVcvSmHMgXFupnE1axWajd1N0CcMK0LYlgH4fsS9hFsKIfxXdADaxP8a0
pHoFCpO069vQoq2l5C6jggpSDgLvQ4AjGV23MevJHI2oku6HR88vchjYqHVR7Ymj
IuOlH6Odqpoic3gjXhKQLHunQA1JLdIxX3XVLEdvdQ5D8NSmg/kslYqx9rGA/Lml
jOn4ccjsKY02yZurTRc9Y6PVL1Vm4TgkeHS8qtbDrPlI7hKmmVy/N7T2VdlhW3SB
Gx+McntFC7ltt5b97+Mm2jSCRggImxr02wmQY6lDOpawJmGpnS5sMbiTUJdzQzAf
tUCuBIRu4stZ0G4DuKhE7HIud77o0KC7LPTx+5NZ9slw4b07JAMfkBtfwqHLgcFE
i/DHrCbNiMKXj1dTOcmUfpqpq33MoRJ7tqJuJ1vQKjyzGkxojd8tpYnL8IYR4toU
NFms35F574lUzLuN8ekH5oF3AO4VTLQSbsO37EJDi3TeviXUFfmRT5UwCt1TL7vr
YTRuWOpZJ1MjpyfGLAkReUsRdXA2h+rP97PqEmCiRXBa+3Dqi7IK83OB9jv2qzEo
7mdGeFHzgJdc6QhQkdVBWvcc+9UBpZ5Dn3xEZTivd5Ezl/hzhSkd6iPaO0IPn7GZ
iPVJL6XiBNRzUWCcp7K6+X2XaqZr9ce7iV1OPDiIFrXCI8i0AhQkUU9g3QpF3Oez
zXtFn351kSfpFn1MHhTwvkp/XfdFMYu+jM2o5yJJMk1zdfrW1uTMdlHapLpHQFFp
7pPZXk+OwoR/aykd+JUp6IA90hdecezkbcqjpuTIbE0OqW3oBoEpE+ysl+99Gyw6
5rJU81YnVarkN/nGiKQL5bxvAgq01cjJ1Grb5bfbVafpnoi+a8PLt8DZSCy+Rhkf
NbLZOlgiuuvjF4ysGZOt2L/bgw6zHvdrW+/XUfKiC7CCww1+EOFtLJ5ehAbXy4Cu
7IOIycSazGCE7ZwFKo1rUH3qXb9wIAP5szIyacn/w5hwbuZR05Lp9iYol8X2KoMk
dsZ2yp6MxwaRoLYEEcvn1fNUmqROhkYYEWJs6jAJF9lCL8wxebRG+efYTNLYEwGq
NPS9U0yWRKjaoBdy4VHOW/jTp6mquB+oV1va0SzBeC7meeyk3ac/yaXonGXQYcAQ
mPdC+3UQGbr+FBzMBUeHUZE0ZZIrEXQeAV3VqZTXJi0YGt9g1Ei+VBi/latO0uFQ
w0FEiwGakBv32OJRUHjz6GI91R6a8Ye1E2ZpvWIZp5b9BnxA4pXEDgO0hAOP4L/T
4SOJoOd3j4tEIPRs9f5TyL+rCQOUO0v3cDu931gApM3eIMBYQ0M6zrBgWXwv7OVA
KovFF4nRIoSHWcP4DRxIKYBQnvpRPVeS/mJwC3fCL2l6PMPjwroajS8guzXy44DU
EO3stVXPsEVgdp7a4RARRfzbkWSRu1BydTzL1BhlyWZVsavPQxYugtQAY3mcHNvD
f+Ws4ajCha22cH4BnW50o1EBbZ4uZFHkl6Kpfsjoi3hwjfv7bwG0yt0jTSkl9BS1
/Gy6kdVreJx7yegnjWHU+KtqApTHQjeYTv1B4hO/VenSefg8jDfs7+f+dWbVQ+Oa
sY81Ow5umm8eKn3+c3UfIiuoT9k+csVWmtcyI+rMfAa9nPapKCfWi3cdNJkjU9gT
F06PHY42f+JREC8zFA+r4t59//RyzL19Lsc4nkBlCwxTBnjOlhX6hyZ0JbIYbdZY
Xgjl9t956yGCcFeAg5koDKqPMr2PwvacZH6FqgCNywnkMQDUJapf2wAjRHjw7Ha2
l0monKrsHkBAMzB+BtMeBlIrlJX9EWgmBF2RWQNt4c/kAVAnq70eZKcnMiFpIkk5
751LsjQ5uRalZTb4j4+PSUAHJPULP/eCWUiMY4erHgHCKtDp7JkqRqybknzWW+GG
QNSCeIFUzVFOhyg1HCYgE4EjKbgvGCQ1GXyHSrqPN1KVWVAbgW1vl0BFtEBcPVwE
+LPFjtpzMgPKwj2W3slfrp/dKWzJKm2Stj92JdcnqHwriJz9gIS/1hCeBZLFqSCk
5wSPSoSMW03/X6RYX4nra4Wkm8BaWJcpN8vji95WZcB/gkMI/20nshwQitDHcz9f
p6VXohhzyrZRnVtv/nqVkEaF6Z4dyM/YP9wx5Nj9oIHKcKA3kBi6BYkgVpB4KhGb
bu6J72b0q4618X7KNVE4DD1ElJ7/r0VN8u6uyDvO4ZlcLn1FtEdfa4zu2mM3v2Hv
vVCz0UBT7+toBtDEX+sam/RMhJcpQMOefYTJQTNmX8FGEFjtB9nvsACXJDt3cpBy
ftw3IAfox76sW8F3Fpl1ZlbYco/o+9luNzJJ+23zN3MUIgtAGYjrGzKoTZM0zOU6
+TorxDNbZmivCQOiOtuXNpuVP1wqUCBUZ1CsUqhWaQVqKhCwUngUCZShP9Ma2eZR
ewAJI1oNTK9QF6hD1vxPfXR1fVP4/YCT9vw7wjPBEsfWle4ikDChm+H5wc+QnfFq
SVX8uEdR+wuEA27jeTty2QSWwkwUqxDEC7xwDlnt9FSOJYwsmkfhQf4rv2zjFR5o
nxhWRtOiVMW25ddRlqQh8FZ8Cjh1A3z6KpdT9zcb7Mej9MiDQHIPzo2V9vUF/Ec+
+cBVX7VqZGWs6bcHYm3bpR5t4yYdlKN71UIMVHaf2P3KpO8egUFEDTuTFJq11aVp
WDv/8zdaTKNxMA7slUhvjP83eqk9f7mcAyi+gakqzgIp7nJSw07cGHenxnBOCMfw
9t2+l9bPtG8CdBZ8Npwgxd9WWauo4h/WqbufVF/JixVSFdXyqbJcSAP4z2RDUVQZ
le7G0fQ3G/GE9yRnBI7Zefu/ebsRlyBFxLoOpo9IOUItTfkbeY6edMUGCAu18bnq
PboqWBFmWC2pjE383ySdnK1SeEzJDWJovLYJXocSdfMTUiiS/6xvpOmYKpjxoixu
X5hXSd39jf4k27g+2ff7Hu5Oj7mmTXTmVg+I6SqCmonhbP23n9DeDAhvhYXowQNH
hJ10PrK7xWSFCDrRWHsEnFlUbpnNamQIl8xvp308RerdNwGBPLQUGpTar6R5SerR
2WL1TyphkYnKn12a9lSO4DN0tnKiZl2Qd9clgT/d0Hc0cc+uw5CPDsAD2YBGmvJO
Iw9RKZRxp7FiMlvNe4N82Dfi1vWhnduZKWX3umQ+Zc2pTDh1fSZS3t+Nc6KU8bW3
Y1/qCe9+DYtQTjxIs13QXgrGZD3ilpdZmTrhAd5J8odhEFQIy/RB2LJjb7IEAJYB
1ykdzaQBUdFUzB4T7KapvvE+sy6wKMDToRDoJgxQmbsCaw6g1fBPgB4OvsUWVK+v
L8UN+JTwnSBRs3F14rd9uhi3qIbxnMomL8tqOZGkHc2n5rDUGWt/EC5piL2p4CHb
ofXHRfgj2He9kkq1c0foblezs4amnpAdYqVZcVWXSe2Q9xIYRoikzpqICK9dP0AE
oUd1Cs8qiKEQYMW8MESIi01zVi9viLU8zPBOi2L+97oLoEbjezL2UE1AV1JT1rP0
N1exA9jahIjTpUYeKiNpAiC3wbDB9qC2+PE9hg+kEQ14MCk8C6Yqq8PxK8GKqarY
OlK0mqR9AW9O8RWilGenCdMpsBycu0aUnE0mleuUjufxEQ+E4dip44GZBU/5S1dt
7AeQYnXuqmmtyHqh7UiJbH5JAs+ZMyqB/I0BGsgo4yrEujeCEtmIwWkP0CPHBPNQ
iq3DdbyRdaOM2QAmRCLhiSsCkZYCcxbdQ7jULi/FJx6/G+x/UrvnKshsI54FMvak
XCn2deAkzMNuNHHIaBdueqDAOHN+dmbvDtBZrGy/pg+BSp8kv8/EI+0FbC5DNue9
ko4RAwB1oW48/2kMTxSnY2bfEiBdP725hUC6Ej+dF4aRMK8J27qx/QJJrtSIE8US
jfxR8+G/alZUI9EqolebInU4s8jdIhdFEy6rwyoGkTV8ZLI5HtDd2E6pZWu0Dc9+
N6Z1DqV4PH+27F0sLGm24owzcG45gkD0seW6YGJ0npiBGKIKuQOE6XtIEvECyund
GYCbjhYu7tDZBzZytegTrSEtO0H7I83FgSEgnxV9RJocr02wbmjUW3fOUMsx+fGR
A4ojkIw6Q7g8nDHkLnrfmT8l0aEy7OceWCOp/8OKRS4Zo/XrCC1Zp06f6sjLKO47
VrkCq/7esNc3zvjuk84xaBucU9lfVCRvj9hkzBQDkQEV5GRzsMQDpKA97GZ7Zkyj
AA1YxHALDKjhACeumKNy57nwhs6KwO68jHOJCTwb5His6kIAx0hqDCToctnie6st
5XhgOodtKu5rWneB+E0WhCZpvXQwGdqstSay0PvSo5J+xcXNlgfkHpSYqLh/vspr
qZnv+AC61RReSVctevYjXvLdsnXPro4BPKsVSQlii6xIFiDHa3eLALjbVhSKJbRL
d0gjC5pIVt/QVplVO/dzIGtga5NO0eTJoX+U1TddMUP4457dnCL9huFWvGfjZYYc
PM7WmOsUSNSpvq0K95YIM8tmvsD/TZRWZl/qVictQpbMtawOo7tyKmKGaWhBrJRd
GSlyE+110dyOHANM/r/K+P8OTpSQfsxMd5GerVHQpawimZTWacCzc29GZh7VJa/P
e1ASes1A0D4yyP0lQu0O10yG+wvinXB2dIK73ayYJY04nvqDux95EqXHImapfx86
VyfPmrfxXHSoeAmCIkcG9r/fso64vJ0/gicWF76gnPIyYtCDVKY1r8s+vqEAbkv3
EFpvCUM2BjOBg4sXZzB46sXQjHYrw64zXBJ8sR2BRpmf3T0d+3EnDVcqfE1Sq5rn
q8pdFeisWEhXU8hoDdjpie5P9D1M3tUe+pxGFhgh3SRWPF6VZSkMd7pUR/5+r+Na
E7SXQIYQkLgj+U4tVRUoxirMwyqAhm+53F/vmaNUFLI5cHEq1fXiURt/Pe64Mw5x
9RsLEtqDoEcuig9LsuK4cebxf4dB3nN81bYv+Gw1haST1CyOiJiNvLWcvx3r+C9S
xWZNEIPm6bpO8gEjveHKuY0W1TsDEGl7O4cSNLOi5t5SY8bfla7xmga8RrVf/12r
lcwdNdZ36v2PKZxbScRyG/VQlzOHcmYNiwO83Z5tU8Q/BecuOshOc4wOcQOosRrH
ZYHjIwYxhVEaUpBOowZtufqBRwzcKGSO+HYvIDbwnj9Xd0xAHwpCyVBMHxXg04lu
Yusx1441T+Nq5qzqZCcr/yamrEGVr4qpYINdLeJaq0cYouWRbtT7mJOxk1EIfR6j
DhzDbf2CpwqLWWqSD9KL3lI5TIp6cWb4DkSHdhLock3j1patnpgrXWKS8U9llOyZ
9datnZezz1UXiCVxTeIqQaXDCgy03DaaTNBLLbnAVDn1d0t7guf4mqXLFYoi7m4a
UmR22nRvzMwSFGWj1qYAt6ML+b4W9U3oKU9MPW1ERFk6EeCNHvKqRZYYy3yyahMA
QaCyxjMSF6VrRTtfIii50uNgxjedjpuT0KVySr9Ra94SeXSxP1XGNQd51GMOyVGG
YRPEIqxHwVtmmIKETKLqfsq3JHJHqmrCkoVBbqkaH6yEu80v1JQnB4y19hmVbGMc
NzWkr/HpsaVGoYfsmEWc3j2zZAIMaBaqJPL8RH5bPP8ZHftKvImQ9KOXocUZhy6z
ges8EXv+OBaUwTt6BXfwn7SwSi2TJTlQBOZvnFIYxz4HfcL8vcvnaE9a7stwyEzE
Ly79mqQFuzzMGZciaw99Jchl5DqHNH+PWLvvHqtYzXI3TUtbTzUkDlPB9tFN2sAI
tTX2Wev935jyQferZ2jLjl59JqoMlxWWAr5RHrbBb3Yl9GhCYj9FTgciZQs4NF4n
GCVOmvFEsjH8m+HCs5Z9NtbR6eQXvRPEPoUIpKySw4VMxhdoVVduIF9JEvtKs5So
9LHCMQjLiIHIZUZ/MAZym1/S5oNC0mLWGjBtfBOzJql8vYcxlP71X13Xx3d2zXW3
FaeMObhpiZ5LFLYBHE6vFayVFnRov4RSiLk3yqbEhXh2YYdO8OnqP83Vz2gQ9NE1
dCHxv0E47xy4CjbHnxBJcwkd5NJ6wfbOZ57IhBNEPY1H2ZXJjh/JBaiqt9rVf1cw
86IrwCE6E2GgXSlO89rPpdP+lMBBDN5/tVPOqtyuAg9Exjl7vrvGXswOfqiEsxfl
t5VzUNHKpItVJgon5lWP6k/iOYbko4kc4xyCbwZqX2nNws52aYYWc5iNyM3mGO2J
UlW2H5fuOs91Izf4rr3XOTU6Op8QbDm8v8M3n0iP64ouRWpvYWOHdnAgVKIfv3Lw
B1+2vTZm6QbnjE5eNmsYpYohBC9PkWMLfpsKv/o924X9YZE0tFT6HnkAWLJzIwep
4YZQx393uimHJ01YrruCe2Y4oBzefRyVrOf3Xh0dgwlOMFi82OQ//Zc7IpUKyXNE
QV/nnlr9nXnJ9REuA1uKxag67E5u6QIxjsNlRMPS+3FM/3z7iHrIin3bAwMFHf4v
VCIpSYE/APP599rbPu0J0K1Yb8KxXf3UawHIzn7wWXy0dahROf31guZsaynntBmP
257pi45IIs4xnX2MYbypnvHH0lcW+UNZoNwAOy3CZvOQ+mcACWGxmlfVzJIO4jKj
asTWoAx/Q0VMZL08AW98NNDoTwDtQjPrvTS1bAybfe7HI0yq7ROU1s1dG7N+gwwF
fZGGm0ow3C6pnjrYvxgxZ0oS2pJA+lNDjWLTkWrT/2WFGB+bnBIrZPghAJqmTrPh
rYeYZh7xv3+JcJ6TTscd+2JPr/IuATa9vgdekX/Z/b4akdcuLAx/aug12ngrCSyA
LgWA/HpCbaMPYyMbS/Jd/YT9S4ftTnryuxXvsr/QpKIdqwXdk9jkZC2FeTk8OGF4
T78BREH+btj/A0yct13L4QSqghtqpAsHmuLX+trzgVoBPZ4cimksTnOvWr57PytF
Fd2NnhvZ5+0wRum2p+FL1xL35k3lBuwt8KuXx2z9YDQ8OCFcjsJWfwj+b2CGmAL0
4NP6lrzTwuzWvLcNGqg3+bh0UhaPkU7jGSakyCbGhcwR7H6jgEZAYwQc/7ntil9m
ZkQKLXMqKuHq3YGwUwLKiqUrKH//0Gw81tq+BVkaR2+rYqNOczW9JjHHzyvWEijT
sdMA/BSlR7HVmqq3C66RA2CDpofXh7P8WQaKTWiliqF2pRFRLD4mky7InFAmMvaB
fJvFsV+ab9ENmCgOCojeRSLim2ykOxF+a1FkNVnTKsHTGx1H8cd+4a+EprBLcjEZ
ewsF7kT2iZH/Fke39/ORw3yVDYYPKDh7jEVsJXk92TptVudsvZtDSCAPS/RrfWgb
03LRr9I/Z3fISx+39vqA6W/NTM9YrvkCfjomV0g0I+45yC9T9o8s/dY5pS6h+WSk
QOGa5bhiEvVG3wIv+qvhpULLPktujbF6DG2xnF3FY3guTwCPLNZUqCa4txQlX+5K
wrrSVKhYT5h7a0RJSlVz+mT7gn2ixsCFRzo/9hpVQD3GEe4kX3Z15re9qMGBnsUX
IjOYD0Lr8jyZLkfT8VmjlX1aOZS/5ZiOjUhy/NLKrDddQ6SUskBQxlEMzPa6Bt08
tO9G2H7OAw/mmR4Vq6Dx92kwp5Rcn7pAibInUM106ynFWM8sndwU0afrSXKdl0H2
`protect END_PROTECTED
