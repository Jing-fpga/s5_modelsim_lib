`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PDl7F6cIrrvOErEB/9X9LtqU3RMB2tIHef7VJPAhEvsknRY4FpbZ8FJfabFjYogV
NP32KiO4DMfnadLImFg9sX+n/JPRCoMJjRtKbN6VCK+N9yiWkr6DXxqU+NucHtu1
nEY5pnrvyrXCRqUdYcz2ReZBApfUzRwA4alZMiqdPbXNiiQ3oJHVLAu9o6YPuEdD
go+FiWBkU8Ty38pZGfr8jHTFvKLgKSGtvWh8zX7TWBd/bwk3g4BCbGEvr7QT64JE
kr2MVvRsfKXTsFUZn5jtFNevuuhQ016DMQtZgawdBit0NcQfYukajKsLc7pOSviG
cJLnVC1tfzJpWS28xiv8fJ+CBHJ7XoTTGTTZ/w+5l7pg1qtvCNxK8sImGqVS7LFc
BoYvc2Sv1Sz1ehU+iFgH8WjqY9n8gCEERbZIZ84AxTTJh09kzWSA8tXFBUhGOEsG
21c4bQFhN6e1m7hEJzcdCg01ZVlblT83KF45jvDh2D4UiQSxtPjEMl8JIBtQdQmD
fIRrhV2q8/+zPPfiLVPjD14K6TbFIS8i3AYjfBUO/TPLm3jiafZamLuQMxzxNrva
g0viTpQSn0Xqhe2O8KzkkEWR8F68DXFZbfa/W44V4z/sAas/az9rXFZ1IZNX+kP0
3SKQrjJmCXzC7dEHCi1PCwd4ycJEuQeL9iYuJP30Vw67+YBfOl6pCL5823kZ4RNb
tck+xNTbku0JYwJAGWJxD0La9iVNmPIiIg0QuLDmATJf3rKDzMKwkcPc6FaX0oS1
0CB/nEA3S6aMHc0XjUAz3uiXe4DvYejFG+l0o1hiyDOALt+0K6xICPatZLE+ABFz
ta+6ho+f7DGyLwZnp5SycXVHpNxV7lBrHucK3rASdnwZZc/5gB058n8cN2kuHlGt
wLy640J+Cm0zM3SsaoHLFX+36y9sqRxpO2qrLY13Ygww4HNUY7GJpkzBKV6UWuqB
ndZ6yaSM9tqHVs6lgCevstcGEJ/9Rd6vHEdNq80OVnCdQPxKxrNZFQ3dxJ0+XN3A
HkTB+LU8fDU0+PyGDpKPio1YynGoAPfLqO63qC+PWx+slBykvENKtX/kHVtIJ7ll
NkbRLHEGhMs5X7YyuY5+hRZMVej/1dCr5b45W5KGgKuCVxLYz3uMnwkQrKzIUx0w
vh/Trfrf2donYqmlCjEp/5JA7MVAGmuH3ooJGMWDxrsYmUdOeT1aMJ3l8N3VqQKq
83UeXjnrkEiQVkrvQnUsd2/36I55rVWWjSHfVLdpKEKPEMDL3H9O3uAoL4ryZUn1
yuL1diMQR/Ydl6m9kGu/KGP/UG1UQ18mFwmhd9ZIqkVbKAecHa0I7JL7Pok3oy8D
uITiucBOVzp9oQjdn/y9sLq00+s+iFP5pF78ax+mok7I/qjIGLy7+6NNgZypgzC8
ExtiJL6rY8JTC8nnBSrbVGyPo+OViT+fS270nDWQmh6qpoEXEJxfWt6z5xtDqAYM
s4ZkFskveyFomuZa8jizlN6pclJ8FCIB8AGBDs5IvSKEfsbiAVRYEJtWAQRDT4a9
NgAaqzgQdNJtwIXrx8JIBWsEw+WGzK6MUXfS9HCKO3PJ4/q6uDv7stunakgML53t
pKH4btj7Ygv6kK/GK75rOQxvFCSRupzlJCCxoAzgL/UBnvKnaDa14JyepyZShYS/
NxJFUQi+lTxAjZbXxcM/SYo3xB4oOOrO1240vX7xLXNd9Bsj83A3qpZ4d5iaw0g+
ryDzPBqmsWJAZWS6XS9WqzLyHYHXj9QpFwhM7LGN4lKqDf0zVX6JjGqOWca72m4k
1nwP9ZKTpJNj41GfUdx6VFNss8OyjZZZOYESGxgHHtOGyuYlWoRcZxcQSRFu92/g
2AZj/hQcp/BLdhpd+9dXtcZ2tWelwk4dt0pksAdZxh/xpiNcwwTZ+JF+rzv005RQ
V4K83zO/52m5jo24u4cOxznVuQV6Ru9JCQS9D5WPWpPyvSshk71q8PF13LSvR0Q8
QkD/LfE4zYiEOvRb0vyjp58/mqvXvOFz/SY5usIwMhgcffeuc+gWq5pQH/QqnQja
Vt0Fp7+wg9g8f++Ularj9DG9UI7foHGyC3DIHqYwIh38lfPsHevaMpFzGT93dFvB
36pco/YN3lz+cUFt9fTSPhVHrjqB4RHqmEbdBXP1EI+p8V2RVslXVQo5232TnGLu
/kARiSROuvelkZU1HmY2RUvpJUU0hR++ce3rs288D1WQZK/YX23XdUlxG2j/CiHZ
DZZQL0lF5sy3NVgsuzrEfoSBhJQiu8yV7Y033j9BZm48ZrRCzNrtikNO/4CM1SW/
2HXTHyzv20OOKYWGsPr1VivfkcHZFcv6rNFvb8NQwhyfRpgFTH/KuorVyyh5CyBA
Qs/wXN6DitkacG5c7/b8t90peoI6xNH0CISwEAnwJM8NzEyDq8H0Qos6r3qXHmhL
z129Nmx88nOBDYy2i+qqFbqrkSzkkuFRKKBjSjzhYnnEuOoh2oUSjzuOtVFycHNn
iaPzj8RkZA4VWOLztgGldTps3cR2XaDMvEOJfYO57JF1QkQRugbOXz5cQIsj24fm
2ZA90Maxdzx3sNv+zxOKblf3N3U1bD4AbYXBw0B52PtoZmVZnknESWmk3WQSh+D1
gWSsH6PdtMF0iMznCwaTVMBWvU6LkycLrbmOsz43XlZpA7qRivhF2CtaVXlES2Qt
yDRq7PSgHIN8w+1vCMff4Hhp4Atnq6w8WTV5xzRpS9JQLUhE98Nlfmm3pMHM7XhM
58+s2F2ihUl2itsCareuOOJjYIDWKdEE3aCJRoqcQS7EVyhwvf9WWH6McNSs/5DC
phiCeydx1omRYdkvjjWTK8lz3OekwtfuvOk3Xlyk5bk0CdK0cGNZvsG8D9Qq+cMd
Y3EcIU/0o30XugRrtzc0cYn1VfFavqVO61Ib6nJHuWpyUKBvyIGomguJsQQkamEy
cRrfsHPXpI9IcwHczhpirhos1vIIxWCYrwTR0bZ44K/HC9GR8DwfzSIznVRSu0Xc
b/eHdfihPWrUc8+FmzJKhRSo6BJhigxPa00nZFZMmkHou+4ryDpW1ZzA3VkBraMQ
QESZ1Gg7QP+GY2YVAvJITdZuTUeknRANS9Pz2DChD3qAgAbTly94rV0OZD2eQVHc
cP1PLKnasOz1nWzN0intvh+Py0OnvMTnqb7quZLnhr9IREl3pseEOeEgRQt6uwo0
irQsnsIwEC2FNji6RhKNX4OStcTCFwLQjvCy8Z3axvrYa2Z3kXtBPcWSI8nRsId+
58Zesc60cyGbt/rqd+hH7o4ilR8WYPFtV3xEUQXmDI0kGHiuOPWwMQ2sMseWPBfP
Ie8m4XRX6WgvIpdJZiDFTNBA4hURZg0uJYdiJ5IPZwFxB3Jy7hXvzdmOzOfXpv2J
MTnYd/wPUhYf7BNsQ09puOUxgdjc4vPKd3vRPQpw3qCZ5PkiUm9XcbUEHaAhKfPf
oYSGMWx175YI91F06WQGfMVN1PEK49yFLIhOZI1eLML23FrKQE4yf/KThlk5nvM9
OQSG/ZyIBjQbMZ8FpSy8u8bWxNfhqu2xdDaWytA3001xEWggz9hUGLmux+0lDhCs
wyhPea64vMJcIq6nb2HuhW4kEshBuOythhOMNTrync3ou+Vmgz/7cI2GkTNh+iF0
Y/cGrnXDJcA+0gkH72vwnQU9TQ8zRR22lDyz/kaOH+TuCKo3DWIu9FP46lOX7JTE
HwNC9/Mm3ZNnivOB9EgSoF0r9WjljELRYFOs7dUk5jfTeJicQ2HTa+1q1airENaH
`protect END_PROTECTED
