`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D9k+JKVlCoZyLlQcQFVdkI0CMID2mayO9wgd/GpAzu7YrvBwCzhaQ9QgAmvhlTwQ
oWCgAlFSX5z+5GkcQmPWQp/gMC5zot53008rcXPTq6hqhulL8T106GhC+GRI9MBr
Vm49YPiOt7cfOv0edNcAsiRmw0n7PFJRJQx9w7XNiaadYfkZs7+yYHnBoYjbcR0q
ZFneOaCoGj9flGX/hRj4qz1tIkM7vpQSzMhwir8uC3pF5fLWNY39u65WfYLIV8Mg
38qLisTeZhhAxvdIExYVLcW8c7wr48/DwFR0VoIh63S3Y5ahcJsHeq4dl5dKjexo
VH+9xsecVe1Kd6L9hWRyr6AU3zem0GB9aym5xmH7Cj5u0JoQrROzREOxU8yBji6+
z7csYYeJ04KTkuhldsNn8yiwFv8I2P341pyF5+uuWq/JTy07NyFm+9jSWnoO3Sy0
YZBibkXxTTIhI3uQEsx3jME0THKctO5DXEPsoxRyVauMINfZcl7Q6LtvHztWUpy3
OmTBcipiRwSsQ1A+XHcJ41eFwbbAaLv/v7GBpZnG2pbFPd0Ql5yNaUaXv2IH9P6l
ME6nG+VcvsN2DgkpC9bf0mIvnQoIEoDmLhHt3GwvqAErzehEDk5C03tsLtLzGp94
pVAN14nNPbzZEM1eCg1+2VCYOC1wT4mLzxZwLM0tbdrB+f/TykssR+AfWS3Y7CC3
j8ZLgdHUCkitsPTs11Hzi9Bzt23CBf2BuApsGET8QdHhuP0eu/jT2KclcukRuZKj
XJezhsEPd40VXHprJzzgHQ==
`protect END_PROTECTED
