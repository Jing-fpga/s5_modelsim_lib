`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aAtElW8BxanqJ8KD3hchPrCsMyGmwZ2NbYFkBVGV0EsxAQdJ7Kvb25FtQWIrz4qk
JJcsEgUPXHnZzLjA5F4w3VvLtd3qMagpZYh8KG5bBvtMmKfhjUeV7rv4IYPOzEJJ
zqpzbF7qSubPQb9ZdUZIu5K1tJIR9MC3I+icBs0AkStCL6MEAGerARh+WOt9BsVi
S7xn8mmi7lhK+1iSqml4x3ThyMixYwLOrjdEP/6mE55G6TRDglp1Xb2jpnflZxmf
Lu6qklwSQhtfUD7jDLNlRyqPyzgKMF6B8P3VaBuf7WtIg+Q9fqDq7zOGR+05xH8G
6P2Vk9FoS6O9BojOSVuZW/QhanRVLevaYXXDT3UQfwQs6+p5NKh1fDzhiit9+seO
Bz+WGG8cpFcN2k/hh6TrRFlNqNzNdXVCUK5P3Uf+J6oRI41Vds4FDWu9VTek4eHw
NyUDBL8YB+dtHA3yuoI6zoGc3YV6jnKk2euhfT9YNka1a0ajsf5r1bnh4R+bYZ+n
2jEcrmUDzQYr3u2CVhAXLJg/CmgfneNJtzE718fhxnUxXy2FdrIyP6qP0yf4OC9p
25Ul0wwks2pxiPLjtDwD3EuxWkR9maJclQVQJY47K/qWf9ZEFNuotodZOFsr9fC0
VBOfBjWqNfrmGndah5qrgpySSObmklfwmsf2JtRx7j3UE8U4qMNkL6iBLngdLh2O
yN4yt4dgpE9pGTiSluOk/sXTMgPUtU4u1HOAh/+LONrGZg/fFTPn4kwIYOdPnoH+
K8KRG70iI1i2jdLHwXxBY67F2+5dW9CiBlKNZ2HC2ZBxIFSi1U39jbdIRR9SXrRO
VVf0Q7d7bHrcvHbxTAzoXCAPKjIk/LJshIN9H595CX0I1eEb2cBS/yH82fiKm7Q5
/ewdJUpR5lUZiTJxrPS8ymAAj5qjaTKBqXBQBggLuwFhyzUUNyThoz0g/WSQ+PMP
WNCVs/YfPQPvih5NcfG1MMCPBqCW3li1q7tJ8U4Dyi16nZ1uy1lgKupyPnfxIBUN
ialdTnPwuIiUFTzfLwJCgL+4b2VbsTRoIURS3PSLu0SevAOvSbNRtpVZGpver1ps
5SVe03LdeoDw2oxYe0ROFcggca9TOyPNrMy/fPfssFWrFkDF0hzcrH35tHJauVUA
1fbZMd/Z6j1c6gEaqHPGHT+PD7/2kT7UBSWoCs9S9W9cWSkTwKHqUbL5pPqKuibX
Os8TOGVLcU3AyZftsfvO7veq8TGvGPJaeXRDLOVD5a+AbGSsnJRhPhHYgEYDW2Ux
H9oKgBQiFLFKORGO1tu7FaDQJmxkBYMJ1CFoS9n1IDY1woNQZ/6rXfxoN4PeU+v9
kdhvFG7Sx3qHPUGzj6wWlvVZblmCKgxyk2yt2IJxHJ23viwRv8ahyHiO/tBf6X1V
SfUMnCgwaptOcKFwGT9KSmdcfazBawjFOm9nsu0XiZuakRA0iNGlb24MRo3Ssfo1
fbjeJwc+e3Kx+kbf7Bvn9CtTH/WTdIqmVjQ+nt+cS+6mAhsUvtRzRjNxBngSv3l1
QKM+ASWKuMOZRflbKKY4hFSX3NvX8DaPJ78ziV1Gb8xkmP+v6wU2rbONVbxl5b2X
rnSGLWxC/qpJQzt+vQ6TDKn7NCden4I2ZUdoVejL4ZaP4fZ5bTkDAaXxvInQjQjz
BLfU25Y4Nzk6xg5HNxoPr2mqqZ3D4vRWQHtKxsqO+tVWhEWMJzA2McXoKLKhxrcu
zcE4XSWqve1yPmEYYLKylMlROzHW6fv//E/Oq2V6OKZeNEyzSh1ia1moiRP9j733
TriNb1ZghhWpqZkZNQCXBNhp0wCi/KYhRyK5lpvBoaEs0PBqXut9tHfx7YapqeU1
fsQgmEfSwmyrAwB8O3YD9kl1JFjygWUxgLJ+UqIX+1OHff2A6wzGWY3p0IlBq7tq
FKUZH7RTguZuRcjictV7KqmG98IUpSFCQvPHjK/aPxoyP9kjip9/JMMyqhFVfwXb
DvycXjsKoZPASty6GmbgilfOGa+cwKxz46dj5A1+subw5X73RDi3QLQ0zCOtYrLH
/6vIlDSqdlNqB+pUeXPIs+lEjb0YzzlWKqj472Cjr/nuHyelx0Jhhv1zlhuEpMHr
R5gGpjZRAn0PbnpScQ8j2PCIwmv925Ebcy1vnu47qxZOoOv0uT/5CgXkDT+I+ZgF
ppEXMfToxoaAPJjOYw27tX2jli4p6GnjtS/bIRx1h8MxOI+BauJfBbVSkZgZcKIL
ffB7nb7/elAVX3BpIHX8uCHMFVaXn5hl8+qWMTfnKjyPPfYnsCQC59RTbzmEEQ9c
IWbqOcbBawrKHETTKMhCoEOrct7nVJSh7mC0PIGvINSf78ZIDFzJM2Igy7UmnT8s
sO8HbgWl4cbvXGa1nB0PyRJsu8z13FRBrHTUra3dqhsWocrISVeFCDlUaTtNk6Om
QlC14emIGLjEdvX81Zmcd1iJcPjnnO6vPded9W247DP8haL+tCfHcJ+COqLhWvli
hThqfmGLXqPIEvI7PCuyurtUFgb0NAHwFEHVb+ylHqQ=
`protect END_PROTECTED
