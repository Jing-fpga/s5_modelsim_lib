`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b5MRABefv/CvUi7+M5N4LyKtwptc3B0SJ6hCGW06TGIb4MCuUEIn2q7xf21XCgrM
XnrXiurz5OhQhKPQ6zX/XC3P7mSZOLb++6GMtXvAS1/tWqP6IQ4XIYDf6qK1o3Ac
KWI1WKh03sgsl9GlYdE/vK/qw4E7GxA9tXp2LKTZq3TRFRICK6gHn1PIdqnVvgn+
DJL7icVAzzRTo7hY6Nej3MaKnZEaMQuh3Tso+Gj1LDlviGhT1F9IdA/E/Vw9XM20
SXa8uAh9fXJZ61u064YnaLao1kRhWn1oF8E6G6baOd1kwuebKLwabrQ1alI7/p5T
RPQiLTft8YyzdUitjLinkGNspWRQ0t5/VoegWf6gPYrcnubF1fiB3WUhChGs91DD
mnAan6cdypHb1G05zSU8CA==
`protect END_PROTECTED
