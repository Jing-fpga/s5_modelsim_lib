`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ptNeayslewimx49893iLptMXJNkGzFKVL24iaVQLD1O/tmLFszltKe6ixxu7Fx5Z
UmTWR7eVMiORouyt2m44lPtIEhufH/bBdeZGxtI21zh8PHUGu0DZsx9RXBaRyML4
e9/+FfrAPus1UZalxaCvgA5nt4gO6D/ny+9Qy1dDxSHkWzItu7QFYpE42DyoNCIN
ozbP67Bjofy/rwsLhNYACRtC+G4aQhs9sNHDCUEhQOiasmKL1VV/AO5jE780xyjo
aXaFetfNPgM9xmvVsejeGVvGqROAV6dAVrt0lhNA0EopGPsBozCi3dYN/Ptwr/lb
EoCJjhsxWfwgw/pz/HtQlhLSa7ZYfUhes0azoyDiDSYV8jemU6ZKP26LIbp/wu+F
6Q0on9OZ77Xw/7zncJFTXusP49pLLB6/9iLgLdH4xNAyZdmZV7vWMUlQUfrbnkTx
w0y49N5NQncxYDvm7gp68Mj0IbE9PABWt/7sEENPWiXN2ueMuN//cAXT1JgVYRyR
hkN4nSj2bMvmqpPvHnhfVVFJiaI8OhDFDmgMlqc00RwbaKCqOtL8xg6xu7dZ8c+E
zIJ7xpeH01cXxPfcaJtQ0HCt1AXWq3JzG2EvdeDbnSkC3Ok5bBG6hxtk/GkaDO00
6TQ5ddW1Hu466LCMQf8MMAGe6LQ0e+cf46DKWGBxBGN80Aq6TJUxqKbNIyXkM3WF
o6obwgqO1uOxSHVfYb3PRyzlLYqyd7/OVT9PBBd4sLnxBQT9e8D7IliU4ENzpPdO
PzUpxUBuDTi8Cci3XmQnAKyD5JYlI4V8vrBly6Zh7j/4VmPk3TGPpVaiDfXGYt0S
SYVn0fXXzt9BffXb8AaA0Ws+pCsH/gx/iIK/tEt8bKhGEvLoTTNxCk7H+HLUHH/r
VBm/4v469LTzppJnY7XrVUim7i/QypawDgeye1XGq1j4Y0YyJzVTI1YFnk5SIMBL
6Qg8JTEHoNToEFjv8BWY2pJsUNiAr+cWe83wyUKK8KMwYBnNvK1ncmpxDXcQhddV
P1a9fZk03xYA1ZdoRX6yDrIRaBRm1/ptFSazAHy0MDiFqfuaXN+lpJHQGQGSPx+m
XuZEpfOGwkgB5YYy0j+aeYgD8a6HxEZoTmHHCU3bpS+dk+3tzmSBS9Pe7Kyu0Frl
owuyA/SSvxHlWNCZOlB69OlhIPcLV+eZfGCFGbNBLOwcesp3GZ6pFRvj+1cn+/CX
y7m8ZgSqm18AbOJCzPk+2xVjBRQOO+dalqqtnavxVRHzwLkxP7VwBII4Ck/9YmH8
pQ8oobjlOuGHneT+KApfg97ExDPMjVFig+k0xeXS+s5j0KWKLmu1Gqk+dzuT59ui
/L017B6fo229yJqfpUeYc57fqc9RfBT44eddwz1aJNDMFeCbfl8j8ZE8udbC2N8F
F3Kj0vlEYmYdH6MadFU8uZxT/EuVVePOCXHJIepystjFkBnEq+PcwlOdtvYY406J
5oLk+5VjlDtja+sq8BrxSMgXYhfHTCXQiL9/0KnKQrTdLAppOwZsE8CKG67Mk1g6
QAcpRckknmzBmHPkDwZfh/enuwq8/hbtAghwSLBUluwr1OS1CtgdI75+tNRaob+R
ScJdtfXrE8gu9YiLVYrYNQMLCaCG6zuBwhnV7ysLl3XS51W1y8E9JLWg7sF5uTWD
YMWY9fbMRixG/IUxoqMXRBEeJUDwgAlfvxs4OtPeQUlUhP1Ow7oF56u0bKd6ZYME
VA9RgVAZQSo/uyCZJewZ5dgGnbYHIMnttMAXlYsCxRVnt2ad+MF4qq7ZKnGZaNkx
F+rnq2XHHoxWsbkaa67AsFkcu9+AuRwwwWMZIvL5B+riApHfjL+pwOVN/tD3t0Di
b+A6gHw9L85am4jYx8c3SYF1ywkP6B3wtpCQBoC5VrOX08XqHLCOii7i4SU3uXqC
qvktMFRSmzDky54w0PzuSPy6Lsr2ci7q/dJ9r273zW7LBDny1mNZVz62He9r+1xE
KCbT8WzXjr/+aKpQdQBlI4H+vwc6BbbedP37jt+FFRnFC8gFJ4cAI2lpesbG7NLH
KqNuR/OsgSonmJKwlqEjR6uxm0FXQ4V/NaZKa6SSF2ryoWntNUYR5NJMFITNu3+E
VEJ4fyWwS1/4//ldc9+d7OANrM2/Px5EAohuX1pRPE0=
`protect END_PROTECTED
