`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xsK4mYQqG8gEJO0L5192LF6EbLsTZWmj4mMuWqMl/8H53lgN83QVxToHzLWfO+on
J0Nt9xeqIwPKG61jB4TX1IWxee0LkNqknUbXwRrnZSHmUWfUm9Vhes2c1fudqtyr
EFiSf84lKtcMkGmInSmXkIaGpAHLA1jcBuwEzajbx1CSh/KxNNQrcbD8SMgV5wj6
7QAt1ytV6GDwfCSCDAagcf2fWX6ijG+x37YyOizzzOIwNxzaLNVb2U5vdKx9ySV+
S7tPgVh443rwiLdcZ6AgoXCiv470TcuUH28yXjnqEO4rHDJzVI/bFmEayX2JN/KC
ZPtdsT6RSqV5DA9oPjFgvTBRuZL9wVNnDRrjaGys0+5KoY5ZbOZ8O2pqUVfZVn3y
b0eMCGglrN66FxNMqZP2YbpP5sVSlSO4BhhQ+7vDyzWQJucZsaHpW3JGKgMNd3XD
tViD/qVGU+FwzRLiWGnEwHNYy3ahIOzchYOteg4xPLf5HCDMMhVjvS8qorCEhAKw
hM0rSH8kVOACcju3ISKVypjOWUoGF+jSQi7911GKXkqRmcDXPTPiaVyhQF6YMXLi
dhcb4EJpYUHuqNw7wGYCMscYeAC06RD8a2WgTWSbJLjB2kmxeqmZ8mxDWzURzxph
DNSBxC0qTB97UZWP0ruXfTFc7QLVTe777Kuxb5QlcmnqVJl1nMSd9gexrQTKA37Q
XCn8XEyNrbKKDKW1nGvkHfxtBARlL1pwH9yzA7iY3Ur9roHcM2ZmxrgLo93QSgBS
oN4ZfrElVBRrS6GPmVZoDhS3MjSWKQvsi2Xfb/vQ5hp4WXuAY+0A7sK5GNJKvMKY
N4af8IaNeek936DRFQ2i6dpFQu8S2ox3yAXA3fr2McK6bQYhQKJor90aklr1rHXU
Saw1Z4BIywaZedmu3UJzHaRQFz0Z0CMTglLoYAM4gsTGrDw0oBpP7GbP6pxbYRj0
E6J5513NZAYrzGOKThCVW6R9wFbe8hGaCpwomDRHWozy++kf7TmWjQ8bpZbsTSQ8
6i6rVrWjGDBj13X/y7GaehD5o9uqybcTOegP0cLKI4hTPsbfqArDJw5XWS4/98IK
VjZNgJZYflfP0QacwdxoQ6hE9dab8weRdOzi8GNAegWtZe5rfN/a9FUY4Ti8lZuF
dRYvyvzUDACi/7ljsMSfeySf1XwLq83JWaaEU35Hu/Y78961plRCqQfPC4GHOHAs
dsdqDrNfFYzQRqVEQlTu8NJ8qzxlZgLtYwy1c3JKROLVeDD5px3OXOl9tG2ClS5b
+wgxuMVnNGsHikFNXrwFpx3vWPZH4AXHtBtKHxRREi7S1hi1sFEALSNBEBU1/7Fr
eN/qkC7jO0HWp5zpkl2mi1+STx5dq2c9HyzjTeIc8V2ZQSsGWv3XUw4L8liEMz/I
7qq1IOQpPmam1KfdoTXWLhy85WeQ0q+coN8nUQO+R/ToBdJmaY1rxh0Dfd6QtKm7
l2gLnF9Ll5UhdNu+0iGhE/LULfB0jJqVGXngOcBr0SQ=
`protect END_PROTECTED
