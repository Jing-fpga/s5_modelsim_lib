`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UZQ9bGxTitUphYmoY/7fL84lp8nNyo0WntYlLIO+RwUC/untMYpiT9L0vpTLlLta
GHXRC4QVOMMWjq75vcIJwAqe0niopSPGmMNwS4d1h/TH9A7YfDQVxg0YKBK1GBwP
aun1/iUj00uRUFoS6UG+KWHMlUmdWwINoeMyJ5BpRCAjs/Qcm31fzDZzn0QriVBY
alyXPdY+CyOxog0c/ZUmz+GU1JkRM3Ao1HJXmjyfsTeiLTrtdYzIfRvyYajvfNSf
bHIRcdI4SO1jI+5NY1QXoubFrZySDyw4cP7mgPGYkZr+sCh+ZaNdzFIGlzAAPKvJ
5pEP6qraDCkaBAuFgOft8PNcEXv9lieSJ1uCf/xSJtHfXvJ03/9N/A8JB3VJyxKh
Ptqo1EHwi+M9/CDb7BI7gdMPrzO072Q8fX5KK333xRMhxJ/gjdehwQnGkmNLU5BA
VdyZkRJWbZlM3p66mR1udQsumAcn//m2VR03lsRInYSq8nEykPHItiaJ41zdm6LP
9BvQyDs2viA76SPocvYLrYuDh1TYHnD4GGr6qHKevqJ4Av0J/TeURze5VmCQZgpj
OrBpMxqx34FyUW6qQxtKdLfSJJ3VwaZa7Jq3PnaW3a6jxx9gNXEq/uI+RwIJcQ7L
lkw6mcySIj0p6bkmOg0qcvMzuZ65Eudx62a4cZ2k7WvOjs1HXdKprzoU/FtsqXif
vokiQuEOHvfdzBILgRq0FneosI7vKq4ZtEUju2Sy7c8YdOg/njTLJKoUjo1KQPnw
c3JjKOUXRfhMKmfO9o8EinzqUxJB3EhzL++U7y2RAYDdAo+IXDJPTyf65KM0gPsd
BPZk+PD1fzBnYrHisXIpswHX8CmchhQMpniLymQlMLp4WaSQ4BFXMUT6q+UTAepc
PmyX+/RfkUcylQEIbY20xgtgpvEiybe5GVqg5R9irFiXcO7cCtSyjiCeOUznAqnC
T0hksgXabGV7cqegzbxoWPFXgbJqlVJx04JB7NNQJHjWMv1glpzmuNa8dSigAoZo
iB2SA7DaLvgqr1LGdQc0VBOeno6wE/c27rnvtDiyhy1n4kzSyC2xMvCsOTXjlfcf
uqoxT3Y4nWly7EkrgQXmaAd8b05r9+nyRV53LPkyUx2Nn3Aw8CFESI14IPWX5x7O
PnCpNSJr9TbnaXy1ToT8mQQ5rN0LJ3KQ0EkPkGAHT6nsVEeuQhqtFLIfU/BeqbMm
rILuU4kwoVuSLcB/fBlahoMVbRsk4k3qtfOkfOYfle6Ay/dmY1vuTnz+G42/sYOQ
MiXHFLdSfsWT82VO3Vd+NOYMoi65FGOLbqWa9HsP2/XIO7x16IwD7iCn5rNP+YfY
xKyERHOanRIxXhuMr8vF2uRuzJ2OSJ5OATlhCQnnT5LI+I7/gjJ765Bm4G90AAD+
0XgPqyHyomAQw+tC7UxoiBFaGNdtKiNK/OG+Jxv7gbbvyzYMa2nSEA7QAnzdWQoL
dYMuWPUFfIIRYjLS9ZL62eQ5jCdVfrRp6aSFCyqkXWvse0X7V8YXruD+gHuLKzsx
ogr4Zzz/zhlZg0eb9hjKaCbolsgkMyBkMo9UhjcMhJDNxF2/WxUCY721U+G2utsL
yj+73vN2t3wSRNqGR4HJRUpVcAH7tZyp00tZhfzpgG/4oMPA12ijra53Xl+3ovMW
F0rrHR9WtYbMHTdeQvoC6YmkatK2Qp+BSasmCnI3JzoN53ep8F5MmBDQH+ybexRF
TvZi6kV8C8BLGgSDVd35LMtv9QeWPZUDb3LONDN8w1ysVZIoy6h3BHlYoCiy2Yt1
mjx2fMrzVakrts69fPZIcfJ7zkBjP1Pq+aPy0YWQ54xMo7g26MmEgMYoHtHl7/ec
`protect END_PROTECTED
