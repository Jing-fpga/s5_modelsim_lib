`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v7bGlLzZ4gLcYEL88N1UJvGEvGjnBhQcw10ChczRr2uwsv3avirakz0e53TV/p3c
qlu/d2WTlngBtScPEO0GBeURJNxuGlKywNWMFXTHkpb67A9KFL7Lt0z9C65n2EwU
sxLGuRm1J+6wTJufTwcNC7GNzULJteeeyRJMR1+yssLD2PKdc4GCSgo0aAtjqn8l
83vIi8jAQH2sSNt4DLhCR1PZ5AMZ/8yzSaGMUiULBIEIukhoE+H8uh0SStXokM16
1QMaIkAiRSIrntjPwsWbezLRz82T2iMyiVpYsetkp1muYfJ3sTjSf0syFEO5J8K2
VSqKiwksBPM1RIwkCr8ZM6+CalNgOPNOqus1IKsnP51U1WJU1Z+NAEhASQQyV+8i
V0oNIwYqSzMOw7ZNr9loKpMZOF16tB2sbXiznSKO20fKV53WnTFUXn4dfUAMG6jT
VwURERH3mUWueHLoIWxCfbhfV/LAn6u5qtuCu1P3u9q/ErpuAz8viVu2BuTF8nAm
sRD21Kbsc5LVk3Lr2SIMP6xpKotJUmOmuSb/qO09HMuPZXrN32RcJIc9z1NO7z8y
JjJMyOPtXy0dYqIvltIlQjikz+3YAHVNhe9+zPUx1qhUzfAcyAMnqJcJMuy7UZa0
ZuLLW7qeM57wWUlzvNdXfWknrcxs+Sq6wP5WMQDzDX8Bw5BoeRSiDoerI7J+ueN5
Zyl4/0FkhoYWwVW9nLZQ7w4vMAdP0aMCxgzF5CrxMOmwxY1M6qLcud9lfUTOfCC6
Urih+R+2XVsgufT2+TyzsIdTZazlEeHxMHzdddTiIv18SOr+X8GL+/6P2hvcsswl
TM4+tx/oApEK8d52hACkeD6yq2MPtlUoTWuosOPrtXpi09wwZJZpi+xMEierdpHM
T4dHj/D1aLDM0Y23Af+Zm1/bppHXiVjZhYavfh2zXECFdsby9AtMS/s6uwNANzO/
JmAeFSsWK3sfP5ELypXzRgeI7St/UqzdhaE/Edr24nA7tUDWf7NF0IXHwyqtCKhx
h0okGdK07pW+YNMgtCgLTdWbHePQXQYDUdRxllEREDKwDwb2mGiVeSzpBp8oIubV
`protect END_PROTECTED
