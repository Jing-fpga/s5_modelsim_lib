`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KyZrq+PbI7J0cPRsciiUNt0hPFAVHVzOgtaqOFJHNRsTSKJjxvaLtApODsRNVqI2
sMkasZTn4rclK+R87wwV52QcXocGkg5QUc9Je0BGuABgzsKxHno24C5pVuruoIzd
fVo0OWpO3iuMw8LmGZdVjV4C0hSYxyYRi3ruPiKAZ+1MuvW0ST4PQAeMrOgC4zHk
j6uCZHwuiEQMu4qpRLS7PlPHDY8nVB0JTM2Y6j9hV8IfA5o84kX7S+gKylFqtaEW
nM/BGRmvkPOONYIStyRRqTr8/GQKbd6u9AfLL3DTpAoOGCLgcI48fOeacP94ZbnR
V4nsFMYhAn84gPo869RTazMQLws0wc8xswbtSCjV80fxEndJq4N9sp72S82z98Xi
cQ9HfycVbd3vUSHfs5x/0uMpPNL+1idIx6vnzAHthABAlCAi28QN8lahVmq1IPaA
fhLJys5gJRuq6IRF+X/SKH/F42ghZK9HLEo7h5mV9l9U+kPmakUHakPLAdXaUBaC
RzEwv0S4KHXxYXMl09b1dNH6pdwyWcvd4jdoFJ5otQ9GnFmp0GcIZSz0SD67bL8W
JoE/5SygoZs8SJBQ7Kw/EWERSjGTlKuQ4TTZe+mO18TNbtsppg25jr6aE6Pjzk/S
C3YyXf5DeM9ATyWf69sIk3H4vcIa6naT7EW/ea+SSv/btA3Um9q0Vg12vc3tetsW
xPLIZrotSFrVTwV+Gze1F8ZicYACEGgsrgGjtirBc/S/587FxDbzWxdPWXxzZEp+
Ki9/lFQnuWks4oPAdDT8fJ0cKNeQhi1hWd5yTyuWECTa65SH5hBfoHV9jU6J4O8Y
uLGai/Ttub9SdgOo4nOYZZfBvCpmkj4aw0qPy5P/eEpUS2/K5eQ6ML14UaAHOSUN
pXYKAgg4XMrQqb6Df3Mk8Jhb3TQ1wrLc+/HdHgIHlMs=
`protect END_PROTECTED
