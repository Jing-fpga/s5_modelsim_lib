`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8fMvf956BLBOAoGawTpzpyD+1+2N9i68XGOjrgmrKPSuIBZ2AV1aV078EVtkSQwS
BlzpPrtzfemU9nHuQ+a9KE8RLfpTzOVWXA1D1UQRHN0Cfap3b3q95QmuDhsnp+1y
S3euhQMcfXpusf3saJw7qfWeuGIOEMeO30Sj4Lc+yy5DaLt9jBj5IFn4UZyIjffk
1+lStbwFjgFq8dA4nbPixBnm8i8dkyaSpfdpMIKfuKIsxchBIAv7Z4Z8UHBS/IAw
ybUUx2hsZp7fd9puRBHPEiJfuKbLhtAB6ik3ZxLnGXDWQgIlvaIL60CGsYeWVwMf
sFYkdI6xnlJRilyHx95+A/i/xnJpmrt5Ns5KMgZzsatR3rYLjeymI1GulAUzNQCY
zj1/NYbeE75/TT3WOgwzFqLFkTvPbtUYDmTTWQ6Q+llYOd5HM+TcCqHYcf6TySZY
P3JAOj1CSiBLEiAKfDxhma//1mU9pG4FHJtYZ6cFWQI/PnScZVba3xBIJZaztchO
8a5ruktTBBRUdMGnEDEIZ9WuzjqpYo/KnwlZT/zmk2SWEn1ywepsFN1ZgCECKvbh
Zl4u2eVhD0H76MOG5SD3+v0+sVKdsK+ArZvMxb7OBINOY7SzGjxWHOg2csyjeRZl
4yZGrPR4JnUXbEvkI7uv25+3B+19FaeuYbtnRy23fu5O8YdyRF3jca74cNK131ne
7fwXZ6ka5XbbasCfaOTni53Eylmg6B0hp92IF1if6TLH7wIiZME6eJfLBolKVaPA
gMNJDfh7k6P0fpaKqp1XYkqDbivAyo7c9FSVY8qq1sXgV3QaohBYGQU3zsy/UUiF
fv/udWW+jFlur9AgyQi0ajBk+4OxXvRc9bhKzC6ObGcFcgrs4QebkJmQsFsyl8gt
hbLqxraoXkRwWM5D4Fz9baopWRmRQjc4KlvMLd8WbFGngyGC1pe6LMPz59Cz5Xh2
PwaMDdXmgX9yTLW+UYjqohkF/HPJZgLaBqHq9t+ENm43BA1116MUxBosy8VGajN9
GZ95d5gg0Zj4R8Nt7hXhVnp3HHgdgL3subxhqyK3lyDHIT0Jwe9xJO8wZm7w1DEE
JQwNMOUU8t4AkNxtFXG8Hjxr9vwdLm6eWoesF9TVJ8NiCiEsKHu9Ktb5GZzRRZfl
Mfk4XPutSFMPQpX96P01DjY1FHMvds7By3DRZXvk99T+XjQqVAQ+vgCpFFMYGT9Q
pYRfoTJe7kmr5zHES8znehBEacukjNg/BomVakVH4q5z12V7TdRDplPGb4wPQGxH
ffHkZtImeZZP037Jd04g+/pFZ117Ge27sknpOKoa8OuyGCJZ5gVYMAW5oRzNS3kB
a+XFne9aa7O3StHqdrc/lhm3KLFXDEd6EqH5HSPczTlhdJ/InnjEEDIyf+YfoNPp
XLMKMdAnYaDi2wb+F7vAZZvOrCSFmTljo30PsE0/qiPlPwZtywbnUWZNiFe4nDKS
b6Iap/Bok9cTRWy9uxs8DvmZ2xFU2tSMzxbLf5HdUKu2ayIiiOtIQLdfVbgU0kCM
TQle/9pCF6noX9SCmjhXpG22fUf28Qcrojzp+KObQZ7reBsmKJlz9qifbka7cKA7
0ymWE/dpeZyvRjdytiia2Byi1AkFRxuVG3oqovXTmBrELW8soKzteMc7olt6zkrV
IkKTqD2z8Koc4Z3T/wjjlTx+2YvBAcnyqSkxfUQkhLxYD57ykZywwl8DXsBpxcS4
HNOQZ4GOdHm4BFUKfjb4ObGe9dsLUGLBxld+OSvGCTUZn32ccAkgraEnzL7VivmU
mLcU7mQ6V0Td9HbmDnLEQbCu41896hSbaDQmvyGHOyz0QjYS5BE8GUNKSRrTfpSf
TCB0PU2wooTc0fOVIPYzLJxezu93lBtJbqOSu5vRtgZwEBcx92bKdY+hMGG5LKc+
tB6zNUj45dU8fvXzIV+RH9kF0faBTiYwG7horR+TMBFARygIl8L64I/bKEbsrrSB
ZA/CKSeHakzp1eRV1jxdD6FJu2u837+Lh5qcBMns23ETzSWMR5ZBzLRoDVMCaRWe
GFiBwRd+l6Dsak5vydFO8iLe30rjJZ1dlmYtFG4Cr1zSMTvwvXU575ITOU2w1QDV
oImNfY4v96DytFtkeHkeBY1CZBaHHDVj0Sh3P6rC59EqiNZUXpy/wJT2g9qfre+H
+j9kWm9peYkBYchvavM9FaqKCMkrDQciwiEuanSMEd5KRMvgYxVrbLy7c7/shNBO
/uZEgaDFHKAAQHoKzvj3lM0VVwtNekXPcJ9U97CRh55jj9zLRal5tpAcwzLsE18u
yuu8heQJolaUmGX2dwzMv2W5Mk5x9BerMvibtkfh2NwE/E3YGsQMDhPCGV3RNv3z
piJ50j7SbxQTw1LkOFXAMOzgY5O6ezrzS1BFpe9OYdnMGzUYiYDLLf83wovXGM+J
1sms4IlWApcx3/GSbs5j6wDs8dHlM43ZP71/BJxMYGs65m+EFl080bMFPvuHHUPV
NS3SFdsaGyypybG1phRaNAHHohwOM2EsvnIcZAp7e0tXlZrFvRCpFoE/KRmdL/pd
bmxlsoiyaNLOmvcvwULubQ74PE/xtgqSBfcTyt9jwkeTQmiAKquywblRfOE3Cs6w
UFGs+AzxIjZR9fm7UAmqAohTpstlKuJoJmsCFoSW0S9szgTd5csDZeASXoQ3yFFF
DcoptLL83pMm8ODYgRI5/x7KTXqzz4KZbn2AOfwtfA9daa7gQa7JITSzuDH/bmkE
TMR3BnOq2c60um3y1rZYv/0n2uIBE/oerXn67Lt4vgNLdcz15snMG9PufDpoVfPN
DlaKJwF9nsl+NlxizyA5hcpznf2N55May2JirwsjNknN/srLiui/Rp/7C079E3mT
euJf6RHmkmrVFid0a2Lkus3TKboAn8rCCan8vbOxxHaKg0DD+od004fsa8Ng9ksL
nDt2+psZIY/2r7HXZHUOuoOSLLeoeefJJf/rFcUGissXhDWozRQpAl1p0Oy7Y0sF
r3Nwl0UfQZ08uyh1S57dPYbrM7ofqdSK3CU5EXsjpZa8bdexXblvOcsA0+/3owpF
F9nmpYRrBLTdhTUMQsZgh7vJX43D47QGPOR88W4823RML4ShJ3rBHAwrrmDg6bB6
tyFdsSJ10j/b7kSxJ4lM8w6OHsscxodReZcHqxD99EY3In38I7IefK8ZgWU72/73
ShdzFmwnxeV2zMX/7Vsc5QIPqWEevV1a3Pf1PChD4qS/3D/4H0aP8D+mZb3Vl/QY
yX1VAnZMeldvTcHZZMv9F4k0fk1FuJv74jgpwYlLvlHvmItk36CTY9wKAmYeOWIz
Okn+MlDc4LQpM0rd8qMeJzNjlvM5yo9850LQ9LGqZv8s6ZJFqIPqe0yZsXnDoylu
Umis+1QbCxAM9LyjtLcDkpXY+ILQCUWD7E+0X7HAatsRMQ13u9UpsIqJrReVcYQE
sXQiew+6t1BBSuoAEG+3otzedA99S0jCiuia3VmWOuYI7afoSiPXqSY7XYBKGw+S
V7MbofKyJGtSSC3H0Si8KXl5UmBKQGBXFwht3DfBg7ozN/aNoexH7cVh4s9ovSfJ
`protect END_PROTECTED
