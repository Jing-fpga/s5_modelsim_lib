`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+rSbQqtksjFDFuu+xOYEPKGNP0RcBN2phpGPAAsq+B8vImw7Z3PvMV6ye4Y/RNTK
3enFozma/x8FZkYwhUjkHVTobRTRjgOqGH5GY5aCXLG7QmY51XTBJkvzUklpTj0M
BE4RA84oDH0wXGZoRYO+Eeh2SiI7W+XYl4CJCn8DG3UwND+2bODp//9qVDmVPzCG
nL+bg2iBd9IJ5Y2XRPDnSFm9tHCLJZWRG45XAr+hLCsqydcHcHAV36Iuo0A2U10T
uDRbf3JZQ+ryK//h5ntsHpfjFUSE3BDyafVe/opujzaCQn/iylPU1qGpg1+5LBzA
dRuCTz/8+wP7kWCOSpUpnkmSdN8NQbEt6AD1kky5qXPxDeEkySkBAzdyELz6b+yO
lh1mdDNrXcB2sen63Fw2Ja45G/jvO7Z7tHKPq8wsS4IFcENm49ULmHIdlWn7j8EX
tjk+h1KNh8UZm0tL5bzLc5JT1eu+1rPNvbSeo2n9AzBPnolwAJPoxddaJ8BoPSAF
yQ85+SI8GaD2+vkcvaVMLT3zzVwfI+eTeNrC6PEVOipxRly9HVxSQAYq2Pr9PFtZ
3/S9O2yB7fjDYZwnDASekDryJBiiuuyPZQuMxgvHYrJjCHn6pM6+N1YvXur1cjjD
BQsZIQOcyozlqm4cFha0I0xjcVGM65QPSqzCi5OcwLRMsVeLNAE6zlIUyHrC40Q+
`protect END_PROTECTED
