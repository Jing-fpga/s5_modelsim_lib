`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
20ej71ZWSRte1moNcOBStbTAxpyvjpGS2bGsqbBowm0l8tGHZJKwtwjlSqzEE+ah
jEfclUamWLEGK6wwgAxWo41G5sEgCbhqJ4uS3b2xbP3RZT5/6/TFrIAqza++YOAN
0Plom3Y3Ds/FKL16a0AIrtyxQ5HQzVrkzerVkDDGEW3OC8eQ3DAkNmnOyrsWovZv
+oxBppnxIfGWNBKkDu+zR3fYmDrEYOc6uBdaT++awEMjAuLAiwDX+ClzWAYENhwW
5urNwvLL/mC7Hc+pXzfZrEQ1uk8O4ZiymXDyAZKz3oB0Ebf689verGuAwM7PR48g
jlGsFpRFkNc7zQA47MC4UKr1BNtdwixcuWCYAVvYwUVR/H87KmM8UYBcHV+CLWLH
uuzAet8TJ+BT2gmtB1XzGNdskuvAlcH93byReDqPa7LFBhcYVqla3LUx3Axp8IM7
IPqhdDwwFcb/qu7mkCtUMT/XXSkhXJtg/UBc3XfPRAJwOsXV1tN6emdlgHowp1yG
qO+oDQB6k3gFRIhNCGnIEyApWIa5AKPs/gSslliy4j1vkXHyglbGeKoNLCh3Fqtm
BunsnbV+6pbCRxYOMolYi6OutsW6U13wxYdSyrqxkm2DGpDrTVRJTVKnssjtMkwn
eVgb4svBJLLKgYc9bkRYQxB2aBVLBY05ZYlJh85nYWO9aWw8BaI8ZWREK0fNVPGk
h2+4Jn7V3KUQpmE7JK4DojdtqlAUYbzX1d5d7RzOUVugNjk0uvZsSITMVh/oS6Ke
vgBdzijxZYQjsvbY0W0/ouzW+5E52Dv0ok+6Jcc/5mhdLjVEHvDnPvDjDQhoNsDt
6l+L690XjrQYIzO3+NavFFe91jbkjOq2skfLankpzvWxTj6K0pK6niZ2ntPsYZ8H
oJN1Es/vRFflOMd8aorgXT8j6HdSmqKYxkVU8mT0XNMCfwQ51vamxMxV5MwkY4Yp
oDGw9/5hl3m3qpP7WcpKqKNZLVvBzhcjhzh2RONL4coNZG3SjVy7EyIciOua8PAZ
VLQSEMazmowH5hJ2GIxKvCUQSHSzCzxJhiE/yI5sZMVsn1t5jiew5k58SFQTG6KB
8ygWSLzwdW8XJ1VgbRBn/NS0Hcmwp26WFe471AqsVn4JmEfrPe8Fl3XA8zXVbLKG
7vZ4mVaqp6CTHKbQWoTN1L+y0XM0s500rSInF2/hUoYT5y02JY99zYSVw9olCVrh
xuBR/5HeHXz09D/yH+1WG1XrnmzrCwQGYz43fPZZ/12jlo9OocuavBLKiuc20bwM
a920BcLIT7A0W/AozzqT/kfjjXWTbSmtnh5sog+ox9r+fCOYmGZBqdbR7uq/0vwc
dMGPNXUHzf4QQeYjOvKqfmjclKZrKTjXR1GY9VozKmsnJTcKQ4wQP/fqy0KjXONI
S8yOvUMnzw029r4+eNiH8ym5ESEv0+9azOGXdRZgO8VwSHv7Hq4/qxYCB1fgfZkS
9J2/iW2w/l7Je++Yi2tDt8MR7StvPqAFJT61qUkKXDN84vLZpV7N13V7E5pf0rwV
YcuMjZ2HssQnKfa/U0DUq4QBPgWyay7+uSq7DFIFKxD4yx/usyXct5aW58Iye6Hz
oT9H+fVWYkjUWbkX3NPvknZegqXaURBjWjY7Q2m8vl99S/Yy3ibvy7mp5d11qlTT
8ggwVLS7S82VPq9ZJ518ncvPezVeC98jm/+T48YL6lvFPKTWwGscaIy8qgnjZ3nn
iwJESYIY3kbildX+vZRND70DcY4mE1xXXQ12hJOG6I8npjCWMZCj7msI4au2Pu4Y
Cwmlrt3zd0tjMRrZTRb936kqXheO/3v/oGogT95pVoCZtNO6tJQn6CTyze4+OQUW
Wz3Y6UXlqaLz/UBPhyJNAvUQo/OdE+h5xFt6FQrMOCKKJxkqZQlNtRMdAlQrMvpm
6cQ62NYrmpP9+cfyruIaYV6coM4WYFwh3f5umtMO/Fu68Ixv+B9xwK4/1IHMEQNp
n1u1fZwMeff3YkSKkvioMOFKk6ajLaIUDponR59RNvIZU3I4kIXsT8T+I1MfJf6j
rY9cld64eNuWFQniPdJh0kDDf/DJJ3CGAq3OZ4uQ8gtWXRL8IiOZzIP3MmYauAdw
xYuhDq0cqSzxZL4mfpp7eQC4xViBNbjvdTf80seLSUx2UCztVODd0pq+F1e2Eykh
hfpGS8NW4nVH/rdTFlDDKpIoxhhLlyJ/LgLKwtq+baHpCipi3/m+cHH49Qa84iX5
fWrLMJzoKCP501k3DQEmbRJXo05/Qgks9qS0zowj+gsAbJzqKANdZlY6YWrj+3PL
Dm9GeBDJFIoaSHip78diIGF53PEJ+Eq9jh1a3mkTXhUTgwQ3iB9jsMfdY70wrX+9
nIOlSFGG944uZqYXPRiOL2/7hScIg9earj87AHfuudZv9jTKUR+rauMIAXwuK1dv
yBuqp8IiPJ32ym4fSvD6HsJLldFnEySnSOxSIc7/6gNplRzRbp+wR+k+JTxl3ttn
2Ywta1SAHDbS8l32uWtqMe8WKplFMM6t9IFJjnjAKR75RHArlOgYSiF0UzQh9UMa
0u1i1HInLVX1FESfM/0RzpYD75b3WF7pXZ7toPem56dfGZV22pSXfvMETv3AjrEi
QaSP4br29jyC6DhuIdbRoH1hr/3Tqp3ZBx8YBx2ICetNwMJ+aApZFvkOlqVe0HNc
2mQobbPdI/0ylVAnf5oaTHGyNUSUKzlUf/Vw/3Ya/PwwiaHHRkaH4DtMzp4P0g+U
trEHujFozrPqsdel72AeUb++rvDlcRA4zsoZ3id1Ie+ck7nRff/bXnhlxc+ZFOwZ
wsg5Rqj2JXjGpPf63UFfCo90g30I56ha5Ip8HgLVzunYODFlEZc3dNDbn6V5qAd6
3Jh0ulb1pLAhujUM9VrqeqCPHo/c/4xw8z64POKLDpkrDnalEFgfoSZPDwniFFhM
fsGBbkPSPO+2nkIari01lH7yvBHlenlVWpWiWbCApwrOQ4Q60qjWeAV0dA0dop3H
/Vqft8PHML/ORLMkrbmSf1PlmMPutsUwodhiPZ3eRGJDOpcSN9BWFic/xI2yvKh+
uLYG5XmxYUx98zTvJMQEtjOey10J4DN71N8B3wVIghI5fE3wRCjpS5vjjK5RcmCm
2efBMdPUPSLjdbYHVTea3FRhTO43Gzn6tCFnnC0wIr2DOvy5hkiawX6RSBaCugMZ
Q+jjIC5hPGqBUFAL6+ScJUsLj8Vjhg5V6YnSSiERNdkFrRAd3przRW2ZR77qdhfk
ddY9NIvLGpk8XAjln9/CnCiEBS8vyvrb9rNi/1uwj5IYh/qeHJzxeJj2NDjxpvYo
7VGwZO1pB4decSuInhZibVh4/IN4svQZcLtVgAVxLxANeUNE88HqBgFRNI0IHZve
DUbwdjRpmJGCKbnDzU5Jgrtq1S+XXK0tzD8VYCcAZA+oMWGGB6ghZX9pJ/CFCEcP
Xd4IlgFXJF/lcHjw6qf4AKnWYk0/Tpl0VtThA25o1N8U/Cm6yO0Bfup7Ib7NyPXm
6VEl9jbC082h7onI7EerMgXLegw8ZwG8oB+ysvLovuaSJI16gHCVsqUWpxYiHshT
2Up1s5nJhU3GHVcmZv9hYohQ0me2rXE/c5PjOF8cqiRQF+xvnK+iQQa9/F6VRUZ8
hTF4gfo1rrfL2pVdcXcC64MySHRY7fSoOupcy/1B8wDsNaC6oSHf9MnFWACuRtBE
sbBxwr55v4BClpFdZbi51Q6A7J5wN8krlvEUtEM2lmVekcnIl6UN3U+ufQ5vDN6w
JtbYdp306SJwnIWkvwxZ+CauDtui05Fkv4L6RGyXZbnvSw0YPZlbSA1Pbgq/44w3
dOTFpwT/0tfT7iwjPh79rnilj5+6Gh5d99IfzQNjG+LbJXoyuc92XXFQkJVHxXjF
z5R0uZ7/A6K4l8SMpG3qVmWXj4n3FxaCrmUGiBDC/BXrlmeSqH8Dhd1VhtFlEloG
ytX/bmG2plIEbJpY6ojpkpdKMxX0YeS3pNWwu1goocFpDwFA1Hx1yKm/T+QSVJuU
hqIbA5bdFLZRJMy2iCNsDaYcUT+P4v5Yjds7Y+3lgbpq6TIMXnq5wB7beBlLdabY
JgVY3T7xMJ6XsrnQ30GP0xJE7Rgv9Rk1peOLd4mrmAUWiCg6qjhJErcHaTk0pF2d
T+HW0Jorpb8tTQNHVurh19INI99BtwKkotEI1uisXBxh3K1LaafettoR6I+0Vgv9
Yvav5Z8tMruca0u6mvQBW/tflzv/K4mMNpyWXksEW77lKvvAEMwJum+i2OEs0tq8
BAtwHSlS7jFdba6+D/l+4Ah2IL8sziT1/wDPuQmfRDh6xyJQYIrjKLOOM/NiMjqW
gHYPSXYmcD0LW2f0AEkpcJPqASsvS+TFeOAvMfdPkV/BqTLLfg6y6VFlSa/m5ICJ
R3jnFlwGWPrMaBiaqcmxKJPp1z67ZiVJXQtbmTbU63gyyhkToAx73jwMmeVPOpZs
cVeaKgcLoF/qGG80iAbz+5QKKzv1TrDnF/xNk3+rnO3jCuBdwK5qRGL5bxduSZU1
QU0ZRJxOsd5/m4kivOdCUWeGOHWFTMEFW+t0wdIiv8OXXcI39GOUApMsoOCVGZQp
HRyS6BDy7kE9szCLIaPO/onEjceQdA4nA6eBpuQPrQAyk/0ecLg16v4J6urYqnq8
bJPvVAOTPzqs8soKDcNXtsxYEOeSuB96pKp6wYutnm2OJ35DkTksuf06kgcLtAZ1
m7z5cAbvwVisWpKl9XiOR/PM1H2+nKPa8ou+PO8hVeMD66f9HlkjdPqqkOjOopV4
mZrKgcgerjrRGmehbqWcNRPe4XSulxdXP0Kaksck7wjtkhE0qLn3avjIn70F7qlr
JCNzIKo73Vtb63DDW6GQGXG7GqeDwbsLdSbgsTNzDaPj8QTiTsYeoXWo+X9Yvmv0
imiczLnVnwMDG6bBs2HEu0tymavDNdxgZa99UlqB+QHAJUFPOi+myRFIpHKkxNe5
rZEGlgT55iTEnTBfGR1bpow92OelmoqFfm9Oi/q3n2H81tAXIeO3mpJOPRY9zpbA
Ee/yy55GWkRNhGYxfa0uzzofrOYo2qwjgBtqjqNaD2OxCHGfpWwuuw4KuVh73iZb
wQlcS3Yhac0zfHjTTZxWYQlLg+yhJ/fnMA1/9F/DofRo1819O2026Rx1er47kUWD
JHp89Qg4UCvOhBRAjplztNRO4fbzJmc3iFEjQNvexvmWcRCA1ubmG8394B4uKmJR
QTziK7vOpfw/3obE9N3raNoSKFlOoVrJAV+2E3smYBdZZpmiUPugtffQhvOz/tbE
+Wh2v1uvsCBQIbk20k6rQVN4zhMAVl7Z6VtPSSfOBO2eFvTEHoLUXCNk0sX70YcO
Kio/TOUK+bxssSd+4khaD/wcgqdJMF07R7KU6zu19CgxAtG+m8gvVlhx3z5KPLk/
abGAp1ijfuRzyl1an9NDjkZs0mI4hwKD3JuZQNooOzjm6vfDu+dWoFaM8vKZZv/h
eIwn6QCvpo2NUATKLdHiZoJB0zneMmtiF+Qn4vvhWUxWqpZFoMJGh+XR1bmW6gzx
b3oLp8tapJZ/GL6sO+xH9/yzlsR78EoHhpV9I8G/JrNRyBZAUL2VDU2qBpjGabbV
4sB/hvrg0kdeO8IjTz8CWFA0Cm/n6IHkQOZ8ikR14u1QtV8/pUV0q+ZsYcjO54WI
wvMzdSLBkPtNfepX8Ys9XxpHhNrNVBbL3XtDAszYjCD69tKJ3YxTNYUzsbP4aUjb
DWmcxmh/EdgtdA9S1jjakRVipJmyhaDpXICKF/7+nTivePnqHblCDncWHmRZsakZ
uU9FrTPvlX9/4O1onFcwCXuBOyg9FlEZKwYRV7GnHcsw0vflvtTdLBta4553jG2L
AQza0IaUufJb+O9k6lEigZ70NyERzyGN8wL7GLjb8PSQEMwOM10vsCDGPW6iV7CT
v40+k4bRevd/w1/4B0jqcVB78YqN0gwiC5knjIrqkqSLgHiqvq5GcNmLIihpxaWw
SIHKiGVUcw1du+DuoxMzyt4md3Aebn6p7TdrQN58UW55kEAzDFOqRQ3dulaSlOua
8YPG+VEgzuogI1iKh3q71i5J5FPdQNs+ZKCulBtXDVe4OhsorS5lbu44p5EnE8YQ
/U9TvLOdn9x6DRb9sMQtPoRzvMolRe+5z/Fi+wt6r3WOEdabo40DZGAM4bPm4roB
muHL6m+jQOeJvoH/AXQCBmkkYDAyr2RR+/i/TFO2WS3jgVE8X4CANDVRyJUasIkH
mi9nZeTmJb6twMn+wIynRkrJC51SXcfrow6pS8j3YVBA1uE1Fki5bnS6pgGU2JjE
R3ML+WIjtl6qMWJqhadg5iVjOmp7Mkkz50rTVqdVbRcyl9IDyOf1EyJtYPeJj5YS
c3B4AxTtOG4Yk+CrQeJ/DkTFqyOcWdkyK91rqmA65BQVqJjlAFuCNvo0hDFUcvg+
c/88M98pBbd0n1pHXDZdQz23ycWvF0YKtNjFwAG8F+RwUz/lWtXFFVdsTonz14Ua
USpoh9Yd0wX4+t/c7hTxKa6rxEX7yjJz1Y+hZA0VSLqpULGWeWfNjHMBY6BvK5EC
BsTZ0cNNnyy34PrlC3Y0mYAvyuQ8XcBAueknDLYC9C44lhE7Hf8ilh66SaMSm5k6
lQsBjD5k37r5B3+4Tgkzx4hOPj9c2W6H3hz5UEsQnfxZ/q4vvtxi57X9AtzLOBEz
GFicBPps2yA4EJyhHiYJY2wcUFtz7T9OZy02J504uplX/mszndawdDJX664tWuPe
Kbyh1CqwkSDhHY3WVTo6ubMFc4qNZmKDRrsW4c+8GSvGREc6zMv1FLbdhLzCOOzZ
JafAyZ6fxW2J4Ph+LSnYibRqlpuLOrPYRFYkypjVxw52aYZchffmJqkZdbSwUjva
lVgyDFU2LwS9dS9B5r+LjYqbrKrK04J0CMPhpriRL1lArzNH+PES7a9llrMB0hkk
6hRNgQS7ebvR/XHlQCW9t75RgdaaGGMKtasa6NGAagaZlLbpnuzLITu/h+DOymE2
IJLGS8GM88DCblqid2vqwYE3WbOF17rvk7s3s9ieVQlEkAU2+jkS5svEC7hokKhJ
tt9J3zolwpQQ2hiUXzki2C4SQMGNi2O6ZSQ64j6pFPlbI2AfSkJLhxYQXbC1gObR
0OmD+ZL3VLXbvb2poHBmfM4JnoEXPRswh1p4dT3Pk93LMX7WaXRHljv10OMy6i6t
9rM5SdCQWfrstaRZIhq7NlVTvBKSCvHTtz37S+Q8SZRQEHOUU++3wfyeFH/AHmRa
HnRD4ht730RC76XGTkzzrIC3j+LEHVlRmNAfOPSA1QF/YNBFa5bfNFZ4v50ytzfA
X1otqbB7LWG+Ou8DjHcjecXvSfnisjJTeN90rXag/OgB9zzYSIxTt3ElFrkSo5yi
wmBwSlfnapkOM1I7AClNSfIS0eFmQoBWiGuahZQ3OvJ7rniUvDOub8s8ylW7wI1n
35ulO5oAxFNxiRPxjVhDi8NJP1iVP+u1GeIge/IxTF5rjngeWOxdp0dqY5QLZMeA
fVr7jQtogD94sikFygh3HjU5D7fddkhJ/zBqz7pcP01rzaD5oevbAQxfwMOcZrlf
gZNC5jMibBSEga+UUb6DqDRMWi3ubVHpqZmiQxxgwiyFkn3OB62kmQT13LnUy/En
zL2g3yBKqcv6A7M7YeDNotoDrvB1PjTLSXtRiBRTqDd7GC3uGtHBMvLoEysM0iU2
DDJrAK4ikTcRhBKNnpOiC0TOnazyUndTYFzKGsmck2GESTXNCQVBAwvvh1K9v5T/
opNJfdK3L1ez4kap1hLy0vB/Xfr0lrIwX3HiRhtey9KNRLIUqyT7VE7gGWE5X9uO
PMyBcI/HGoVMo3UxhBPceTbcA4cHvpzn1+jTaUVvHCkgcjXe0Wg5aI6jYGhNkRRR
LC+ouFiHpzq9QxYq3LJaXX3D8Vajbz2pAdmJAevCl0x/BQxnxqziMN46EzzlqD9Z
hkituk75KyWZrrVtej+6SvKiPhxs6NxS26IPaMe8HpNK4vCNRVZSTFmQahYnMnib
Kbzbg4ABAQgfVc0NMAgtiI/UekhsxarJA5yrT+UldY9w+1EZpXayAZfeyT1b0rI1
QeQshlynV0aFEiHCErEs3hUFHjol7/o7wZzh4IvEOGaJknpVOUFFUvnmGYz8//n+
z02ws7gDiISj7x528oPAbQHsTqpqS9ZufErvzRTNsEkxAjTAhnC7T8KpUpST7jD1
mAu1jIIba7/i+LPT9orXkEnuQ7Vb6TfQniktV9uB4tOL6b9L+vQhmwqC6XVpHHSu
KFV1zZe5GjUoSUMMisUfWnTfjqa0b5cC/ZdciAG7kjWX3itU27Ry5U/Tx/xS0pyj
7VqVib1dT7F9n1lLiRSvDDCg+07mXeD51tw+ubFdNOYsCYiflIKkiUn3ysSqDNuZ
UKqnvCopDscsCzqmdH7KXBQ60mUUvUySwN0xJE/r5xhhb4XznHBhdaS2sv4OHaE6
gkCaskn/DKPTvWdVFBxlpVYf1/MKu6WLjv+Pf0XEq7b5p4KqpJAFFRjLuk18OEXv
Js3/HKkmr+GPw0IMJjtIgHuv2IMdvELwAag6irZzUdKDoYHJu7pYxig+qkyQGZbi
sZpvKtFFOCHKWv2ncM3BdUpt6yTtOVVR21bAYZ/u3aC7ERJIPxfi+6s05LARhxlk
EMX8X39IVNn4RCha9aEdl92lADh+fxPY8icSYxKmPz8V0J1OGpdKN9ve7w+GvwSd
eof6ePcc60bIGCDaIPw2zMusoxZJrOzX9IBRXq9NWIW/hgL7fliJE1xGoliBeVwS
h8EOSogZOAOERz5M2IRdP6WuMfu0HGmdkjIQ+jQmWYW23O530Ia4OoG8o2kBciip
k8XIUQ/vziojV0aWYHTRZd8cKmanhE4eIPYEsXrbPYgO0gy4SemKML26zjC7G6iB
Mn4O0Mnk2i3gZ75AN/J4VoszszcvrDwHOgsqU6qCbD0Ub1o7ZiDSdLxXwwa5EjCl
eHW3A8k9dASOSa9UxrDwAIRYOPwAgn2x+96kME0fa2yOfzUx02FclNI4+SUlyKqk
Hq0og+JtZe2ACxCPljv06qwsJO/cDEAgQeE8P9uR0ZATe5MViIjH48Qy4Hrai6v4
Jq4SrMl5Zv9vSV1/61xR2GJcgVQC7SikVBd8rV9K6ZMAxrmG4hYFKtzJX9CBVU1e
wH60kdsMEfDykD4eeKaEzlOmweNRXANQBGhfAzKceXssOFCixsOXGojHUTllN1wA
NHOoARkf2Kansk2do/T7Gl5hHLVp0oGfvL8MWUz249ckhqZ2pP7pm79HOWW5CrFk
PHKI9Kb7Vp2GLUYsknyosf7dlDKPzGUovAp+9sdP7gm2VXNJdv/X0ZQ8jX+uF37P
okreuto9MJjQG5Kb6KoXmKnuYgfvtbBamgI7e05O7iE2VIDWshIfXwT0ccE4rrsE
hW3F0H2ot4AdPgbwJUYDfOPoatJPh8f3c3D6AsssfD6vfwZZ+8oNBtqZ/MSD9LwF
YT7KVSlhLLzCkv1P9qsTZyIDCTP+M7xLgubWe7nmBrHiNGYnL8A9jEqmypnbC1vK
/qvT75fECUPqO5PkT4IvBei5y8Z2CDZuGj1AAMWMGqpBCM36hMxaaa9Kmyx4u/yj
ytGsOCRvSUmI5pYULyO5cdo+8nhfXSrxB4KFdN4/CpCFq2wLiCzxjAqppAYp4Z69
l7v4BZMTu2wA0zj+gPqxDIje+SOXYu4Or44dUWJ9ZziIvqcmdThBIkvJLaYr6HAa
xxc7lePvww7n5/xXIsu+M/WAVgJda/y1UL3b6QYoapHG26UCqV+BR20fxbwRE3/V
JqQITulksSWmnuBso6hbpyDsSNc9Y9cbz3TmDGBjYbzLOW9+EfcNcXw5RdBp4pWZ
l0a6A7zJ1/hKGJAImSfIURR4+POv+HfwnoXPxbikuyzUZkHM0rmZkeBB+4Z2Za22
mOTtUhLXWKZmYHi4cPcoEvDjUfxPh1cOdCaP1pT825GDEdlEbObqJAMrUGuErGSK
UVi6zyyeJkY5FoPlyI8xmjSw5rhVRX5GdlHWW7EjxmBujY5Q4DglMm+xUEt9ILki
dabz6zkHpL+H0H+0K15GnIwjH1QNwru6x0pi2K98/iFm0PpiE3Kl3+LpEExruXD9
W3GOTOZEykbBK4W+iwpR45R5cLqP+7TPpvze/ROxAVeJ+2GiD+dhJ6TovVOTWrSO
WnHZpmYhVnmNMAIGNwv+j1JUqBIDVEvXsv+3oubY7DZ9uxiTZ2t0J+fTKXeSueCh
qUTfcZhxs3HywvPgskjSToiEfe4TnZWA2ikYxNZq3to4oMcLpHk7g+Ym1sjGVL//
k607AUn1NNMk7pDQ4iTp6QgkbyDdlXOw0nE6+tW/dlJeRb9xR+ygCAHEqfTJ5WMS
2xwWfRpJzeNHjel60vNTI1zNKCC2Z4xg3xbpPEWOvrAnQk46+YE05ZAIWVBdeScy
/CCgoWp3I/ijKjdBcsJgO5AjWeKPsOYj/b4nguu180yRl2Q996Pj/Scvc/1Rb7TV
NB1y5FXuGGl7VsZQQKzL4tcjNMmEJ1H89C8tn9yQ1FYFoVMr66+DIMkDEdfzRf3J
hhyqIdNPJbAELm1zJiMA8tRQv1Ttt436eWdIaf9gtT3dv0W92WZEHm4GzyUOl6XD
5SBVWeX6ssPqDpGJe6kOvdeWdaAhV63EnppdiG4AbGlMoXAvRtgvNkqJZg7RnXgM
f3n7aw6wo1QvNIsX/B0IlBvLEcArE1LFOW4qEpvQMGG//OjQlS6CgVKp07clpdFS
uCcEDmh8QHF849b9CVU5AfGPVfNmoUmPapdxnkz8haHivoheKDmIOlW3tnsIHvVo
yeQ69wylBUoywLi6olxH8JZhnqYPfcM2HolllrN1CBTTS0uif14jPRENnJgb8fIb
ifjhWWSMOGJM4f76PKf12/I0ub4S//Ywhxm7a9IkWo0ujaBIyzW/IEaQ5jX2moT7
Abftt7TT9D2s4kvmACz/s+6Zy6rqe2yZ18IJ8WdDd8QwI4sZH+OgKkXRTRlk/Ebd
xXhIgFvPNVK1D2L3VEOhpcZTUiFb1LlnZkLmXIL8urxiFUHuDYrLvoVA1K2M9BY7
wjpUVAhef8F3s3hz0CVCmDmjbdiRav/sopl/ieFfqN7eg/MmME+6bwAW/Wlz0fKI
zHhoE/ojf69Y7nj8/7sKFved4tFGhLjig+sIdf6ZgmLAtfPEASVIUroGTBYd/DK0
sdZQWeC9nPBM8Jkjx94pAJPIff+U7m/3NXNRLdgrl7idyijZuBnie0dgt3GPXBgf
bjK/1F1iU69cmviFOBmKMx/ivWsRO8z7ZIVGIJRv+NRSqxI7h+OCJSQ2Q12mw6fr
nYsPjTEtZbxADuJHYxcGMvxtabg9E9ZBsi9vcs2LLUozCAKenNN1z/HvDhsMndRN
FvlpQcGpdKYYhzYCbq7sp7TOeN4jSNAHZPWvIhR9n40u+m6l22j9YJlIMONqlcKS
Cot+FK29LD1mMyByi5JH8P0VDRJpDC9+bHnkf/0lEMcddkv+Ks6bBn2mrgtOsmk+
daXl7/Md22BQugKusC5YPVkzemlQSv8nFJgLr6ETslKBZw4hsGe5J5NIXUdunD34
uRpEVk794659ZBkRkVF72CfNwYyjDUds/ZIScnzmo9KJWoCj+9LDhp+XXqjg0Gs0
SmTIAqnSy5MgcqqHXH70pJN63pavhqy4I20yj9j/yssP1CSoQe4pA3ARPa+Fh4mm
SZ/ddRSa6MpZp4+g0hJ8/j3I9+QjNH6vnegfuxfiHeN430DBPHeus5mWx/EE5w42
5KVfpfYQ1mg6X/p2+gyqoltxpTzDfB5a95cHlN/v5Ab53dU4+DBmeeF+otK6alzp
kp2i7Rk6W9KCAw6otXMDF/RA+oLzmElcp+2tIysM8CNa0WWB1MWPittZRwMsnDb4
OPrIRi/r4IDgO9e9J7s6GrzkeZcLYIakKw2TV9Q2yKpIkLJF7aE9lfSgv9DqI1Ht
2WEftK3IqvYtnee/kT7vhH1tlLovcqfKFujg4kwFVAILZzVuJ1MGW3mDFDh/Y3Sf
hd4LtFPijcadsuDH9Pzud9mQfQuppDHwWseC0dRSZ+PXxSRpVEK0Vn49qy/wiwb6
sEmXCS+O+slyQEdflYmjIjCsVdoS7mHAbiV6y3Y4Luvyq/6KSO/J9Mg3Ndy/UP8l
5umX3kuUw/MgtEab7ws1nkzggC1kCYbInKmAF8dqzDCCQNcIjw8/HhZIdebbX4vz
CN1QenbNexRFUyK6FtjlIGxS4pPm/RYfNGuzjmtOueVy6tW7l7uWBNbNafn/J7xQ
imS6o8cX9a9FLGjhMgt37HdM09F3v8+1Kdjc6aJegg++SZmkinbngBZssaJaTI22
TtRPtTpSXc6QvGFcJSqi90wJi2J0rkfHFnwVRZoeHhEuZ6q3GHo1yk9OmOOeGVLO
COecZeOUZWbN8NWQKMuk36FYwuOc3XbtGO1F04p2yBlX/h/+gC3kqfNxNaYWoDSo
N/UcmTZHyKmVsc5nVmSUUfkAXRFD6OWwJ75v6Ofyf2JeWUiiSGkSoCbg3VhSpvqM
JH5HYTQ3jnujVXfng86Yc7PB+JiYJPGO4YRNpVVYdLS47zo7uFgiFZHTDSHXX9h7
siupYyCPFrt2L2JS5/b8Al8xYFECvz9D08zPZCDU05pxWt4oIZ7vXDMwfQNLKhTF
+JD8rbhJhrA/8y0mYfUVS+9Q1wSL3dLkRoxLTUHcuCR5TKdz2H8nYyeBWaTZTCtW
oVATPn3oWSeKfhi9GKFldOaQ4vMKmvBSJXDTEgs2V+6G+LV0hmLO9LCyMDaQimx8
azTdzJ5lLBbA/MSHdRVolP52ax2GrR1OpwKl7TGgw5lA8CkP4ZwuroagG7PiFaee
wr3FnrildbDik2/w08PZMD2Elg0o80478725Y7vSJ5Vj96HaS+Nt4Ftxn1vb49Mr
ZHobCRKOAE4jvJk3MQ5QWTMUutr1pjTNe++TPFQzABg3GKNLzRPCiZEhL0sYTFLp
fhUTH1kJv+YhDR30Znd2DtJTcIZyUtj+ohCJgCDahLvY/CcQ03sc+KmolpRKZ/Sf
5704a2AkiVqfSjgHSMX/wABovtBVLXjFss20nHaLE34oyWaafMT9DNgR4us/wlQ4
8104pYPoRZqclWy7YYKgA7wwzvt6+90KNy03OSq97+VRdieNOI188T/4/YzThA8h
0pkiVIgfsKefnUHbcXqnQw4ZX9DS9p4orUnMb49J0MXqufhZqyGnZkSyPC+PUK2y
GtyqQJQynOvZ5zeLmDdBrVMXxLE/VPJjg/q9MaOYF+E6iZImsk7nW8rzeW0WGGD5
IxR/qcXWJipqohxXFn9nemnCLkcqEcNwB5KPNuDnA5qrpTZSV+VZnQzIqg4P5iAc
ajoSzBk5CIQfcIMUq9Qmk7ho84yBbQzLu4SNg0GGBf7UDhwIlI8bgzQeW/Z8UTwt
XB6bOzzVHQl7F4Kfq8OUpKY7idtQwq1OAPFKMBT+fBkpSjibqbAynNo+B2raqVgu
zXdIcJ+gSUq85jmzdFDPckxj6fopssmCJbXynHjkkEOtVZAvgjKT+MnNbdIx61UK
IJqMksY6RDR6Y1m4p2I8mvN4d8MiLnfROY7NX5PVB8ObG3epN0awaFi6noqDQpXj
FD7ea5Lfv/GAxJB+5BB8g7X1LkFpTgkad+3lVuOXu/I+qMlX4SOZkQNwULkjAfBf
KdHcKir+tEcNaMx97s2UNz4CYf+VTjPovm/bqc/h5R5wspBQCxEMBiJ9hnuFZYrd
bhroQHa4emKS6rOI8BZAnveRApSQKBsRRv+8IK77tnkLOT8bhCy2W/iduP/T4uaA
sYq4hTi1iIDWxWLkGrePiioemnWo5MTGD9o5ybZZRyoENSDfYr+KuiLENhJlsWEb
dQsEy9rPrK2mLhjM9pkPQO2Q3zCkpeyI/W2EQddW5IinVkNQf1/gHvNmeE12nZqs
doX6dBrpGDkzH9UNPFeNsmBONcJnMDwbAypV9m+1k6XbvkH7VKyAMbyMwsP9W53Z
7PfA+5Siu+kWlukj9RCbVKmYmExhYh9+WZnVbmU0VUV0up1xPYzadf57cY0KhF7j
HWDBLLESLMQDWbJsJ/Yv3QQ6rkJrX7H8X+PBSwP4sq4Awtj0Ur7XMiqfRO4orMMB
iJtvX4mL1rfqycyDRk+iUlzFOh5KSZ/FCwR7ojcPcUM2lI7nhEjck0rVY7NO5wJU
D9g69V8bCzLGIV3izBEF6pobEqdwIqIuJayuozFo+tsWsK1ogL3dAebkNOH2yGyG
ACUhg65PwWCMntrhO9sWUDRXfrBXPhlLIODfiTi1v4mQFJNaeXpObsY5bBOymGBC
esFPNfSet8JYe4q5rRr6ms5vU+WXHkrm1LndgDY/y4lvF15VteHECO79C1chHRar
lZpJgKe1FXs+mlfZ58uTw/BZTQrM+C3ZNJ+dXJgsL4r6zQ8ZUYMWV5l4t69c/g+l
k9C/wMg0oULh4lF31Sa5F7OJzFPlrsRzu8pUUXv7LIfJrxvfRrHZqOc5lWRIMQqV
N5ifrreAnZuFeWS51wqMlUmJ/3EgeOblcsDMlQRPBjGwBdOYELM41HgFpfYjjGUt
JlEIzmhftMNdAdl0Gjc088JZDxqHU/IjBbKuzAaSZa1wGsnWHkH2psbjj9ADgyiV
Zq1XL+WYw9soj6uSBrba8cWLkcB+o0tWaQliCPS7tW7gnd6BB7HWJURfOMesL4CY
+IY1j6/fFYka2Hr/PqhDtwDU7eeE+TejDGei8UuhKJ89JtMtmSVw5TNg38WmFcXD
vm06jzcvstisHDQepVYSBxHaFWJPuoh199txgr7KnGr1lAEn85v6ZfB7/WHVv9DH
hC++VbPhuesBgPJyuff7xlLMjtvYxqBkKejYcJ3m6FV4IYGpWNac06kRQ0L7Gk2C
XaVoGlA+5kJXsEM/jQd+kgN/MgJFRLz+SdEsYqGH6F5kb9N9ikIcbKvN8FgZm9tu
K6cKgTYQ5+8+M2DdvMaYImUeQIe+gUZCNWxhu+dtcbp4xaPBPgIo27mSxNVvznQ1
V5Be4dyhnS2fy4Im6U2k8NSVzkcJEczQV+iIqciiQwDy8zG74QQOd70vSRkL6ZUo
5gjIKlTYEJvlC34qWLszaOEetzN6D7BVruNDt2RbV9hx0r8L9UypJ+wOoKY2LqE2
8qI1xgKFFoizseEzHdp1Tp0UxCir8SyPphHdNM6JQEwiGagBcJSOYQQzQVmftmGy
hK2VL4/nXUJJ3x77rZLkJPLDhJ50g6z6nvpXuTB89pC9gZUDb1mI8OY7uDORYJwl
127syyTTiPGsOvzcgf1TyNwlbBbEilX1S9MvNeBD2xw7qVhz7jFoXO+MQEoSICdl
H52/gkkVjoifSu2ehLRgaKIrZnUxZ5twre4CchG6ybZEN/4bO4ejVS2dJbeoQK9a
Lwn5zqKrvLSJxvBrD8lcT6rojtFHs6wCdzoBvSS9pHRCsxMWaoclMEDIXn+oEIx7
8Qb606i9Dnm4h2ic4cNYEc6ttt7g/hYkgiJ+iE3hOVEUEE9EGh/a8hd/fA/Up5Lc
MzZpZMhPr38MIXVFhsgBuAC3KWqGz4X9H2qjFWSXvEK59vKyr6jf020rtgO3kN23
fzaoFQ1/bVGrwsA6D3mpClTWGZ1l/1et2atLQQR9MVjO6GGHUpVh9mK0xyEz5f+U
RRdB/a9e6Ije0+przxjiJZfPjhDj3kxy9YJT/emBIT2Ul91bkGikAy21uLRiZgcW
vhDK1z6tEUwwnAAoa/qy/6SkBl9bSUx5j0o7QI7b19pfJprdHPlkys9snBZOWVQ7
b6TyZ2wykZBjlDuK0fJxn3HoptCqUP8nF9v/3yRS/eutW6pdoLp62pxsyGt+egf5
9HUmfzryPar5XIl+ZUQ86J2D4Wept1nVJS6w3nrOSF0P78CdMtzrvCu6Mllz+j4e
DHhV6VFcPtrFBamT5CL/wfO5+Ig4bBStmsax2ArtcE8yI62DfQizRoqXhjCQTHb1
ypvDcYuoKyORmfTm3rflTqVavDvhugKXAiTCM42Q3ZFcqBgEvuJQCDq9+bqN827n
2syTZrvQBtkEADaCxITAHJzfcW7r1s8lxN39e7WjJxwJnxb1p25+tEEghUlvL1bS
9DA81Qgsh2U8TiREDYUTHb8xaTC1p9eoFH1HQ2cqyiZtGOXVjsK0zUdKyHKQyuCC
ACtkM2II0w+G+YbQnN4/r0FVX5fb3y8YZf63q+mWm5mxNUrzeDlDmRxm8oH3WTWg
0QgBQlflPtllRgpG0NppD7SKqEGE7dw8aqs5QHd/xDPsAVWHRFhGe8eptlpUAx32
O5SqDEn/6WsgoCzoiIZM3+IRtW+OUTgBCg40IXmJAa6Jaz4VHhYBKXwiixG6fATF
X+RszFa5hxC6gacoA0QKZ8AN7d0Ftt1eirFDMwJ9C5cVfd2vwD5i37W5GYEPHMve
iL1fVA9jBaNgLTmXx+xlGlW/FDM1+7PcEzcC9r1HYab5HPOgwTkFHBw21ygris2x
A8eD8kImua6TSBNW29uVTinAiVA0/pzuBaN38Y0RtmlM1/+WgqtbBx3/52/59MFc
0EkBbK/WBqp7dZ43Pq+23VbzQaeUnioCThLW0VK1L2pBc3+z8NtxGT7IIJPdj3am
ZcpfPtYzQVJGak4PBHiyesvuVvNtLB+Z7y7chpeEfVMdcu9J4VZ9cgR10Dbkl3dM
IY2LXhXVyFKxsS22BiQDjWALc2LXve0FTJk7qDBi92ZZWzDF89jcATSB0N+y0n0X
mYsrqh1bphY9NnrIetKcHpXrrlGMBbgscwEKTIiQgH9ZRLGlMLbeVe7cTiB0ub35
zAa1pbg3AUcfBOcmTOl1epuT2pNi6dOz8yRsji/z2UknBdywW0oIgXtFpNAFUw2j
IxIIYfAnhOqgKE5i+7noRIrVsbBJJxwc1djjVR2pWKWG+iL2DXNeWFg56IBX7ugn
2uq3BA/mVaBufqpNGIfgcWkD1AkRZcrT/By5w8kotPusxVyzP8KA0UMg3oLeth60
pg0poC00MJkRPSbUr3LHx5vUG25ZHYrYtyQSvLp+aWVV96mGKe8ailQmnTsGb6Rj
IBYTVTsl/U/owz5YuGe7cEEbi+E29KE4+5eukG0O5Qbv0s7nhD0D/rqVLhiCbseV
ARDPeqrUq2F3k2LQlfU0yykbd/0GWf6+wFnyMlApoPybRueTCW5Nh/vcB0Ojh+sx
KDTGV1reRbNkhJwI4M996dsKe4vBv7dxKyLT1AVtXYpd3CqL+sLB4sZBP3T7eVPg
O4QqEhbFPfZvcvRQCcXzVzN/9ZW5g6pgz+llsrYdPKK2VRYWt+9x3tBKA0PYLmMY
8zgWAmPD9tzNoyb9tYNqDiceyJfFuvLwwiN+ISkVviLmkCEVRKovBVNR0cFnCIjV
Ok9ECMCZRj+FyxBvH7QB1BRyQDOAMg97frXDWBqDqgwgxSSWdC177tDoJLbNo72T
xrZqeN2LEPKqCZMtH+thMIw1qtjqwvtJfMPOzItia4cxfc7LISOWGoR9KZKg24xi
ou9sGDc5GawT/M3yw8rmkSD3o5Z0Cj6iQu1Hs0Td1ntQHS2WRZtn3+vxxjZpvXgj
uuJBbQhUsvK13CjIt6wjdl4OQHM5S+MSUFk89O8Ff4LEjTGlt/ldeZIYq4GwMgSW
L9s+ko3vdudoUeXFiPTNvljAaud1IoUZJV/QmR5WdSQTd3Rb39aNkBYgE19+dKvw
YwmBqvty2x033ExYLA7TWyVXyH9xp4ew/nwzRd2IQBGLBUrDUOjubUUUSH5bylj6
63tNKSr7a88U7/EAinh6NTXZpf1yUzaR9afr0l7AKPpMyaCuD7pXcrQZYs1R46ez
pIiV65jT1ilz0z6z2QLh1NOgE/M7ZXLrBx++gBixqvVhXgnmhiVHja3ZmgrnZRFn
jb6CyRhFiDdaIMkM6BCjALo6BervTl52tSUljdQ009K7+AFJZKhCeCA9uEonrWHU
vwU+iwke5GLFX9JukCtgCcJ3Rjq8YJEyg6uDrjDmU3Vg5EwDr/OKHWr05Bulbbn/
scfupI3+7EkWcrjqg1yWu8+CK8Yhs2nLBn52HtintjnofIcBr/M0yQADkCnKmhlp
ZQhbpgHyPmRRIqeOuh3gpE9tGbt7sBDwGlCuu4LyrUojo9GnWdTbjN1UqJiuuVbb
RdLgHxaBIiX4ayX+aBg03uTwYotOWjYD7hIpJ+GsmuhhCLSejd2VVOfbCCBabvv3
nrGFbOn/DHws5Zz/HySMPcahkG0qs1kY2KGlQSAoj+zUnQXUCshq0J6F/2AMBF27
yU3aDaI+6neH3T521DBMFf0rVWav34p7BLKEzGV7C6KWDHeDeLH3foKOHH1xNa9C
zhT2cOY6yfQ+sPsz1Hd1gIXfBVU3axHYWn1ZNYzrb52jeVuZSR+ISPg3aUceLiLV
+zVvNBL8ICE/n+m1mrVDk/WnB275A0hVFmOY5IUlwryTKZ1/fbq61kiMiS5i59RC
Auv3ulM9WqSCmrGP9zVss5Gu63VD8dbs8oqk95LITjTWpHanHD343+y/l2wrL56A
s4ljT+DVOqroMbAb8lw7yveTM4cH+VSM/SPazaZbGo20dzLqRjltBzOF5qz130El
84hc3XFsS8livyfEPnY8BS14yPUrY4mLLPYpEtUFebkqkGPUkh8WNAXjB8Q2jYUc
GaRby+1gN9c8pGvSekjuuEVj1pyZf3iwuJy8OSIKlHQ=
`protect END_PROTECTED
