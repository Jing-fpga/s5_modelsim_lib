`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sNUwf3TMRzLnKPsl4n4Tsv/wpQLL4RZm4hjyzzuKySCZGd0FwyyJZFRilzF8Egkl
7ZBDoysnef27GaewOF5L/stPZxMirZ10TmqMuE4Us2gM7Y1Kx2opkvZwJLJSxKhH
H48guIhoD8FjRcUNdowJQkTnUU27bIfGE+EhC4LFUNcHD97SzhN1I60LGD1EuKBL
cIXYk1aTR9NZ/AylRRYhH23IvYOH/25uoP39e13UyblAdRUADC4KWVv91M1gnX/x
u5G/iqzvTf7nk/UskSSGyd6ejV2AkX/UdDgBrbHbgabnvb6Nu7dAgZYqAyDjG2cK
NcABUnfHCHEe8e3Aj89ivZMjPelvvR3vgqWUCHmaTQyCqvA5Lbp4db+RfFfSsLp0
lG9sUfx9BJvsl400F49CcuVZ/M5izTb1KMYGAAH7zLqKoUQaG1PC7j0B/F20imiL
LRrqEMsth7e5LraxlryT/OsOMO9swhtHa7oc1Ns07qfHTbYdQyyYNy5E0oDgvTZZ
uI3S6XnSxEYLcCS9ApO+aJMLxra6VYWj42/ouhFNHZiVgYWz8K5n4gIEfgLuEJ6f
t4VRaxuoVVBuPp8VZVyoPG21q2rLMADYbXFfSXX/VS7ulJhM416xHyPIMwktU/5N
Ep+MbA6OhKcfMl7YOQebpoqGmlOcckx62l3IVIPVCTgBVKHMt0quL4G2VU+VwzkE
xUoFwWo72BAsdbHZdB5ltEJiOtqku5OAF7OYRpH+yeghEeHcBd5mcW1lqLt8Sofl
b04iC4Tk6G5HYZBzW680EucJH9/UgVMsZBu0FY89whSUed4hR8NPb8RM28xy6NNx
h46CmGxeT2NsH18zYrxYhEbIV7zXu7wPKy+rwQBtYn59RjUP6Sa7yS4YPTV2IYyQ
7jB73Ih0mkOt5lg8hC0KPca2JBViVpLr6bWZJXY0gtyLDqMg1CApsnt6f9YBl5pK
0XUqdQR4TpGzvZIjlynXYy/iKYdBRlZgFgJuOVSKpcEoYXF5aL6B9cjLBnLTieTn
thOn2dqMQw1iA5jJ8ODnSW1kvzssIRSMgRd0q0V+/jVE0bQ6+9FABRX4v8OjUbnV
uNWuG0hHut1PQVjEM35fne6T7fv82zv4us34JQWn9yXdppL9j0SN+o/plpG6B2mZ
wHrv/iTiwUB4ez7VWP5tSQ==
`protect END_PROTECTED
