`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fW00BZ1VWVbpozOs83JULHPM3VHZGPaHAAsWCb45vnZjxA/Ephsk7+/keEgXU398
FdEwnUY0EGZFibg/1zNYV7bqmIacBooT9iQ9NBg2UttoxZZUcYLKvlNTIp4fXI0e
P4G70dO/5kkovaFkllkJxiPy+AOJlEiGEvYVcDc/JWy3wkXP3RxYOz5NcsX4epcJ
2HEYCe4FBbEyHAJqb2S9JZYnHwk1pFa04iuKHKN8f5m/5yO36hDxEoxK8b2kzvGE
+D6wK4fMdfTsqzHn9s8kI7lGRxqlXIu0NF7zJ9/H53t8+Q9sb/Kq8t+YU2VjUIHy
EXoDSiUCrFxdr1JIy1MHy9Oq5AiNIjvpsARacmCCHeKhsHhz7QVd30guAEWaqrnh
tZshMnSyJs9MK6DbGCoLhNxvlik6BkoshTxCCBZiqMSdkAgxji94FOTlNiv42Y76
hFm2F1gyFaNSSt8WLDFHoOdcEgmGWw6SgWn3GQMYOOttqfMNjHpq6X1t18pCwXEH
uL5h+focTLbEw4vjN1K0j7r6gPxd/ni3cUfhEhGHUHuVx2zdwC7k0Nplv95xP0SV
1fLQMI14uU9YsbkOsfWF3zaoz+1cuRe6icoGDUZ2WW1SjFZUMFxWhwdpZMvcmwsw
RWqi1kUWHPMU78vJ7ljwRUtX8TFXOPANoYsJ1cMTz0owqeQ4ArnGigZgNP46dKfJ
S28saOVrFmYGt/uM/mM1x34VWzuNZyU1zg+AssWibZeAEoRg+bgodc0ohKAJ9wBH
2RSQopXK7G2BVH/HrPYB5XdyCruU8jT6NEVhy1tqeE/1aeV/jSI18YKiGRJ9Wafk
ZOrKyNBy0qaEDHnbFP8bVJ2Z2ctn8d4PzWuEBrvMg5SYtFOSltJ5R6giBMk1rap8
GEiXrbL8v1lINNXW6U9etFvZ5z+wjbej7GOXsHbvTFI=
`protect END_PROTECTED
