`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h7qU6p1EznfIGNTG2qEXjDRFrduvBkm3vMr67FGAqxEBO8SIuHrbf55R+5wawzHg
KtwdIsscr82xKiKETsa4OsOkC+mozzzfYyWFot+Acrv1Ldwth1GwpFFuBKXg0yIZ
6a05z0DthMs1cS3B0FXRNJ3EKlBE2mR9/6tjnf6i8+KMeg78UFllufpEU0I+ttdh
JdUET9/O4eYFX/2sOB0KnnGwDWuAHD5T3Dd1rh51vY+zARISEU6dF2ibE/5lkpyi
U2vRdT9WOsx/3V7VBC+xpMp+gZB0ISAoA1ATIPY11ko14/xJPlwdOmQw+x/RTbtn
1dPHRtOzIrG1CB7qIH5Bcfxz+HygLHCAsxgcPIM7qFrR4PN2oGgjt4VtrhmgovH1
viMdBlQcSeNgHP5oQZKlvveAHCqO0iBsCjU5Qv5s+SK/D+sur8z4Nk2FHbS+md8/
+/BcmR1p21ZGRiynwpLCVbvbm98Q45MZCu/ZndDDKjmYToch2YRHeMzxL7NlrsRb
4fDolrGfc4Oe7V1ONFxQcbcs+/q+q9wRgLVZplq4t/i7/bix3M9A76CbvztPGNBR
H4FDV0htDgNobSMGU2K/VkcN2BYWN0roLAkd5M5D4q+5AdnAP8DDy5l+itoi8Zva
gknCIYHW4LNjm9PLbNze9dYw4Kb+DJkyVWZ+NNs2UZdVRPwerLnZc/DI1ooVBaUq
s5glPvTPNVWEMvaD4NTEte6MYkX5n5D4DjAOVytYWHd+ncUYhAe3vYpdGaltqqlo
0gngJhwxQvq2J0JwwWU5DWGJ0y+M6OTqjHsSQIBDV5otEHUV/tW7wzWJpUwVijfp
73JLJtZnW4Sq9LE73enprs8CsW71LZxthy+e8y8sXYNaqzZ9RZ53TNka39Rn4Stz
U59DmaAqW/L2pdkNmO3lEWTBwK99vnm5r0B1/H5Demn+vShockB0Q8jmONjqYRER
qwHAdVwobGLiUE/65Z0dHfT8nKHZ9fPh5oBCXKxQ1EnND50VHF8Y9gYYRIEzxnnr
rUoDLYrIVhElbWbRABrbTdkZLYUbABQ81fe9NI5RZQIdUFiaAydJ+OVmC4J671KD
EUz6ZA/OywImGvmmO4KV2Ec1+2RhoHXF3cwbDVPhhI8cuLIqhi81LdC0uULVy4s0
dRBfWHV2phgPlQVnCiNp6Lk37aLjcSkCl3SzPWGMo3gu8SkUcjChJ5mtQ6AozYJ/
NGo7Y7dMyDZu3ACCMXCOru2JGNCRaZlSRuY0GYJD5h2VY3P8NKJhjH0FSh0y68pM
kOhWIxM9XJtfXfU+7VBR9iqlzFsxh8Dnqosh6ov7kK8lhu5aCKJL4/uPKeff6+9q
9M+T1Tmp6S6rpm3J/LHnFqmxF7y6rXeeJEJFuKpwObd3Z0j9pGHaEV6dXm38VpFo
AWptNfXuRP9+2FMC1ZKR/Db0kBhurxe9BH5BN0JkmigsjJVgXYCzd+VcC0WJbP1o
9W0N2PqLG5KYOCMdh3pxpW/uoFuyKUkl5sUzFP3iXfZn7UfWyl3YLlG3k0kPD+3Z
Md1tQgJvFxgsHTnNyQGC3LN8lTDEMZi4Ul48mfGBXaN3b7/Fxz3rjoponsmawSRb
yPSMnLEWQCKEyr6lCBRv/nptl54W4LXlraxAYE8P971D6T9K0kOHODBZqBzUKAXt
RAmHf5LQu1io6oyk2OAh4hnJiQZbEFjb4w+PxCfwKHHrzzc3P4eNc7tq9VDFtI4/
IICPu/qrTS1teAJUkIbeYubm3k2nzIPS69RXq2EsdhRMG/R0xVdIPpiz5X8grnwn
lY8d6l9+Dw81p1mZFC+B1sWW25K+4xuKvkapTBQJFTGw1LDf6iUxw+dKauTjt9ZE
IxNJer1YuY2jlgSVr5b43B75iVy/z9abruGdq+ZgL2/eTBjQPQjn9YDhGvFn2vPK
BI/paxU+uU8D3NmVz7zB2qeV+odtSqGzVRQ1PWB38pNi/MYQYLFIvNuDid2wE+AG
BcsffSGejCKhdrfyZRS4A3YrpB7t4My5wd/1/h1nXwGVH6fKWN0WBoY2V+z/vTcV
rp9A1V95pr+Hv07jUQKiJsAy0LPHEDnQ1RR217SlWyOvB1A+6ycLOsrLl12kaRRp
8A/zDuFPs3o6syYeEUI+ISrCgiQVVu2jFc8WVILmgiIGBd5XqwHpvw5HTkvSjMuw
u+S5mC1nfLkniUuIKvXgHoMTTowbL0Mvep5RPJ0DMGe/XVdj3BR9YgbLGf69FELf
S+XiLBm4sgUG08l+EpUtADp5AUMG+qqyN+0CfGEtZlvZueMCU7oCrPSyOcAuHNwt
bpM2qauW6RCrnPb6OueenalZc52r6hx5lEfpvrnNZ9Kn2Bu6DZ5VJgzptRZXYV+A
GHUdjzvK8uMp/pBdsZEI/1CqsEjcq5er22/79IP/WfjnbNT01MtG6/q4HcD6odSm
UluZoZVY/jUjVVGJ75tEDubJlontU2a35k+BEzSudX94eoKtZDbRwW+HyFRa797t
uUJOarVkf//Hou32cSUr7ECTjneDIMT2SMuhEBazojyVWii7+CJNeqOkg6EzeLuJ
efQ/SmqXxI+3bsiz9RJKsfQ09QNvYrfDdht167x4FyvbCPlYN0hay232Iv+rdEpH
eWNsQAGeJ8J+cMb2eq6C91FAZEx/2aCmvNB6kjQAgh0zm4hj8a4ysDK5w5wRn2A0
/sFltuHgHt6WjC57vdAzygr3Q9LcOH05k8Jy1p05bcPL+3j8CUGpQ46qVT8o5knh
nRbfX20GfB+SwrSrG9dzts/c15W8yScCyf2rNERNuSBDP32jAMB2/uN2ZHL8R/5/
g5a1j5AbTZfW0q8u8J1iVA+USm3f5xpF+VRjp9gNLwjKzOdbWqeMddu5BGlShbcI
3DG3hyUUqXvh3N+N84/H7kzTdadPrryy09myFQCbjipAYgcZX2h9l12pP13qN3lR
SL08wlXfevdGEQyNpd7/jlBN4SwudHFjLYt0wkLOO7UW9kScUFILY3e1IEwkSLq7
vJivWPp4T643g0/8hdtMucndnhW2uk52qUoR+T23tsPOpD2Io5VFarWGg7zn377g
KFWxN3rIn7qKig39KOd4cJ0XF8YcIClYLXyxhlMeDV7qEAtqrIs4sMW5agR2pCY0
YW6taLgWJmVkMf3F1yJBBi1Rld9LJ6gGcgyazxo+dAGxX1aBtllwLnTegCYd7P+5
kKfietJrRnDGFbqkaBsJubmswp8AlsycgLVzTvloiAOBcl3YFr0elauEq+1zFD6G
u0USgRfshuoS/Z0LdiL1kHvUlxMvSybg9NqhZPj5hMhZQCWQocxgVO1EgyfVfucl
RpYKnSBABfrbNuSh7AeJIaUs6DYAww08IxozO1AlsbLsfAZN+0769e3vS1PjiC47
xn52hYV6/htb+PSaXxX1D/ezwPkoaLEX2mVhVquaEke11qgVVVdBTiyrmxhzUP1T
nhnbA5q2CmLv5bBLPX6a6IbofCfGdov3pH5gGV6Z2oolpv6WPmASGv+xXFD0I/XS
L5TVuAJCU/WMK0COqNhIgavaB16gjCkLNvqg6jsWIyE=
`protect END_PROTECTED
