`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ql5woGC8b1TL/VsqjHNIq2fFi7I/kHTC7x+K4D9oT2F4YRs9xFrEkSYN3R5dr77G
IeyGrKYCvauuLuNUI0WY58b2etMcJq2eMUQLLnylcDw/TescTzE3EC7ikzeQytGL
yqLRdBQy0eG0qiXP8f6rPp5f2XrAaQZ7OeADHFPOUVX0algpkgjLLDmDUVvmlX2V
mze4s9jnlekBOQhZ5YvZMUaYB0FyPvUkpXv9j43NHCIQlo4mm62d9+3mOi7U0rMR
yfD+CRIaBS/fShb9yiS+GcrzB8UJgNny7ZHeU5YxXuXNooPxhRrJo63ExwwbzUX7
BL/C48afynFcP65H2yP8H871ocsjF/yrhnIbrQ/nppMqhoeOySIzcLGIzRmtxePn
`protect END_PROTECTED
