`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
68ugywiY/zJv61mJY4FDSa/fG8KE4KQC+VK7w1e2Q27goB5epYw9h3NUbiaOUbtd
onhKFCAHLwiIwaPeIWWAd9BVO2wtDMofXrmww6KhJr75xdw7TdWLYrHh94T08srR
Tx4vLReomknskX0MkUY6DfzzMyxYy8LohhBqKaXxlgT97mv+GhRaPYxbxqTlTKSS
fIpGwTRMqy+y3RDwvC/+rBK5wXx678KAkE1MaH/kmtREv+T767oU70Kt0Nid6ou4
KGvBsekXZ+7lvZ3O5DzZeDQ1W0VDTKQ0RE1QBIMmzz10f0zRS34K0QTgodxiGPfQ
hzGaan9Ffj5YYkNAVHbYDyXxh58q4oYI2R36m/PEU6wsnZ0bQuwQYb3nRCHtAKVm
BojXVrZDksXCPWNjeBds1t+ZJ4tYpLOsgtSlEZl6r0t7x9zE8xREfZcwTkzyUsXN
guCUS5uthV7CBAefYum+Fotloakx8d7qwFeEfDRf2rGeuU7qEE0iUI5TkjpJy80k
XBSxaRmm3aR0dpAI6VxAVy/nRR8SQ4JuV2I1/rUQ22t/jKHukDwCyz6n54iktCRr
xZbmuJSbMeu/FUcqrINwtDNiQuu6tgya6OimaH79CWVXBbHTO3Vyt4DUmaV1Xuu0
Ds1JzbVsi8E3sSdGBQmc1tLU0xrPW/VqgYuuDTExEI303iDVuyd9ElOIrawWfu9m
M9OisvjvwUcVFUmIeE1WqTBgPUBAOv+zVmm26QdxMbenzq8p9aHAkD2eoHBXvxj6
shwpkJJRzcux2LffezTecgvNFFPgL5VmE5yUMIYufnAkPdDnj340gRPXhB9uU/+m
uG/W9uW5Dlv/Bmpj99MyO9j5bDHWoUqJXoeVQzjIFc+E5Nx8EpqkL3wBCFDaR1qh
nYXNmQj3d5YyOFSycePKb/uEm3RxyWw+2NHLhSl/aTgb9BvHvcm3fMRsKgJnHhnI
GzB9WWP33QnXvtm+JfbAvCQX5H3jw34FC+JKdFjFNncO2DOXYAKJ4m/MnMwPD7+v
2CJ70dkjQH8NTxxI7rLlPd7j5xrYMVclIJL5pjuqhIDKz8FBl+FngvPogUceiQV+
D1ITR1nWMG1WDENLIHp8nnaozX7UnAKtGEygD2R1b7ipbGhRTH2j0qLELJ3swx9/
LXFFCbKj49EDhz6RExoXznimu9YZH9sjpRUw+GAGq5MNeCBMGPOK6xPfcMSxnoG2
5LT3UrxFyGVE8498aQsUa8bgfP0fE+XYiklHSVzcseLfa0uyyCpkyeCCbtPptBlT
vOsBQakrAc0WUWqfl9B4G8CvM4JzEpaECL5CwAZPgy6IxuDr2LXOyQ9T9OJn7Cl3
mRWakgJc7301oZb2wm02RUFYAVlr4GwKAXwW2XJdBd0/prvqF8CAUlG1QXDKN+Iw
1RwV+4K/JhwtRpu4rJgRSmKiPBCq9RxFkkFBONtmrXn91+SqRM236DxScrnG6Jgd
GNXMzeJxUA1RQMZO2AA8GgDl8sS3HMAXZ1ycpEtSr3IpOOTSZMrEPnlf/WHIs65C
QBWqgCbg8Au5H13p6b8mlbnmVz9OMHJVaDQnTumVnbCuagipzBxoyRPBKipvYTz8
nM2N7/hQA+BV8rURyPGPbmJnrgpEoRClk2NcSob4bxbDiwslgavLB84EQ/uoM0Sj
mDRb+leG1guMRSZaR/5w8A87W6UzVabHpn3BpmUYx7Qdv/yPJ6w86jgDqlVPnkp/
9MZvA5OXrq++F8KG7TyV7sSZT4ek2cdk7EgYwp1ioYT0QzGJxWCirV3SLD0DG0Q7
250AUU4KFz3cG6nIsB4qzHZ3kolYvsoDtch2zDsvjnqw/RkO6Z5BbE2XwZUzTjZO
LIUrs+2oh581q6K9Z2MyL3kw8RnVAs8oPL0YuU+qbpi52XTxr2ao0fu2WEQEmAkg
wkG+xLNIbLwC43mnh0DiUj2HqsLh8qBhvIPDFg6Z4ylyGNF2w0smD7RGfj5S2cD2
GMM5mEC0jLD7wWpm2zY8L71tnfwmukISeGMzyzXh+vR0GIARw5VeG1vW/NA64tuI
L0ac8GDmMJOULK01eno14Kwti2yTACeoQOXZyJ5hAUhJisFVB1O70Nv9RbtfmKVH
6+toKkNicJJfHhM5bNaSlTYZ/DmeQ707seYdbekS6siEfV/vCvNiMS1yJ6V+drnF
`protect END_PROTECTED
