`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rV32KbaQeoVI2Koa7TJ5GsaUUZk/lfbExqK84bEPb0GOIXHmTQwhkH4Hn6d7VWYT
KU89ysenBrzN4DmQxpxIFtDUlcVDQFlo9OBML0odsr9SuVIhMsvMDpp8FgB/3TJl
RMwriy3LiInJRq4z2JjN87Sd7i5Sj0sR4Ik1a8G3gQ9qtmYQISVjtT4LgjSyl8nj
BmuBYCbC/Ot0HlDUAFwxJQkHQ56JTtPuwMIr4HuJSr5Xvt01CtL5mU4H5EE/so2d
4ZHlgEeiPpePks15Ztajs6lJSov5HbWLdZiD6CKVFasHgMHDAdBDH0eTYUpLJ+QA
9/s2ZenaNec7VNRjcTYlBBwcUCUal1cX0wsbTruK8z9cu+FMhRQCvfckYpIZN/Zq
ACUYu4nhgdcUQfXnlnTsxeHxzgkhYBqptJ7ZTRzGLXsjPpuARvppSKNr5st/81No
4tiUrmFbha5uz5EuiWXQfgyjeHDg7colN2RFB3qXsoBetglD7fm7ZH5CHNsvBv5D
uK4TmIWv/Tl1FuCjewd7+OQx7YO2P+6fOMjB1B6YgrFTPzg6BHLBLLrfNeqKKQr8
CpQhzqblcqG0nDUCMBWZYi+0XCUidlfN5kVVKTvFzVCfmQeMM3MJcuABbRZ1brC1
x1xoc13LIgNIXBpXz24uOkaph5Awnqz7pC4tslKtp8evy/cdonBSUaEf2LGybROn
xa4f/u31Qn9daC1GgiLRLoYQMYxOvOgiJWtJ1RhOV29TZGhEpZZ6nScsMb3YuNiD
TfVOsOxu2fzepXoYZvC7pHrg+7GaZGTN51exIekrdTHjs9O+JgAOlMrhK2a/4w5T
cJLjEwj6sj3t1sofAhuMd4dB/6+j/pUuFcBA8l1csF0sKKisnpAEfeUctMErHMth
IE5ogdgdxRoSaf79PFnWs8m98SowGMCL+QlODR4EgboR+4FLWRnU41wQFWB0Wi4g
7w2l7wfbx1tYieP2fKbdjfo3P66IOen+tWj0sdiKmsDEAYVjRC9rpJsVHpE+uZes
R2lHuXTj2KHcIuN8ctoCzA==
`protect END_PROTECTED
