`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TV+mARKr3fIBFqoSFkYupugfn7Rp3aovOUI82HI/JsnKDx7HGA9zZDpQzGwysakD
mSTMFrjrUbjD9H9ROEgWe7e/H/D9QQ27lQPGXaisBTIvxxzgDD+0W3vroDWIVJKZ
T1vgBjKP2tS1iFTyAN+CbQelvZAi9UX0gVrQAfLfm5m60US7tDdrwHhckpsUdA5l
QqMDNjCXmi5ZFwkfAnMc2iwpP3+rMHyJ7l92lPANPbY2S8BTOeQhjhvnt7mDpoFJ
Lr2u366D5Um4RmYSs5EmURqiQW5dL5s9hlTouBVMLf6N0Tbtr3trFSQwrCRMkFkA
Qed5fwLF8L2BUWJTcaWBuTG8m3B0iZM7ZZB3NvVi5eJtZTWi3KT35khBjwG3oBEJ
ZeIx0e9XvyQ1U9ZLmYShc1AEjzZCeBGTcBb8yv1oobd9WcO6+vyxwOf0NYK0QwYs
zL6MTay/Nf8d2xzGzcZO0Iu0hzLkZkh40spTEpMNcXwKEPInuN/CRnB+4+Z9rt6g
S17tNaHLOaTSbA9LC37gLIrmeVLAVdadDkwsiI9CVtBgPRSgrmq3aUw3mfZDRH+b
+cNvbLIyLp5KQWbNLA6YcF5IZNkPJ/zSBYKLCBzaOoplo0hwXNSMS/T767dkiAwU
I25JADW9hu6JZ6UCH20nERvR5kYKiV8cZBdBkssUh85gPLgllpbTVcBPSgXqC6kH
Iao6TrT0T97eLrsvOYgFaI4UMOl1p3fTvtuXNRfnluIAmIH14KIl/zTJtaid+4/R
tLvKFWJRSc4RxpGSNaUDEqvWjFxZGn9jRoXL8FZfe4pkjk8ymhEUY0q13qpvfgj+
1acq48wfilsfvoQO9ckYyywlLqSoI0IOrShrRJAGvboT/qCEIqVHr+4IyOoWW4f+
7IeZgD2B06ZEIR42UvrTHaY3wO8Nlr2AavBDTkoNRySmD2c4nIyDcqJ6KrLISSF7
chDxe4cniVWYYW0cjpwOEpaOJR82U98pXwerivxTcPxBofbVqNWpw1kWBaNJjRJj
XxWgcWyH+4RCptIx8mo8EqjaYOoAYr4B9A89mDCITPB6pcoLBB6N/kQqXL37Pp5A
vQRY3kzqS/Ut9o98pzDxgXwfQ75J7JYsMirD93O1fe1EzuKPW/rg5V0dpsLMkIKT
RZjyDrtbBcqMBez+WVkMaoYYSrmW4XlCj3TZD4A/F7BE9GEulJHClm0/VexXhvac
T5qZRN/AP5r+sdVdSSvaWbJ2X2+MIdjRH0I4FwXfmYBtVMkkyEQ17yMU8qVgs5DJ
2QJK86vYgZlJ9Si8C7LnhvDp2SUPVs8e2UAaZ8WW8WEM83EBrnqv2jpupxFgOlAB
zrEvnzTT4WeqDxN8FPCnmQL9ve+PILteXr1JGRYeVqU=
`protect END_PROTECTED
