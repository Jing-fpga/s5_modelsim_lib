`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+bgHev/uO4ENEx5WkKf/PD97G7OR84McNSgQmuomaxXNGBxsj70nto1ayu+a0tLm
3Anu3ipVr6j5dyIHRhn0r2unlz7gEK7rVbHLk4bKENAHbytVj9wf964MpKHSfZnK
hbfWlHTbwZhmvOtqkV78JgsVTbbHwdso6q8/GEw9aZsrBaQlyGZnVAEcBPSSuoVS
mXtKPvQ1LUHSWs1yZJIcW36F6plJ2cW26SjZRNWsznanjHWYhxHxgPwh+e7wXTFX
OmZfKxr44Zyg+Uebgh+QF2HWCOZpd70XgYqxRemBvyyGQ9pic0rztwv12vVs44Ds
uLBySJDrSEN112ZqILOlDFjJNbtWakhzCPHDGMPjelLGVlIo90kDy1VSGBtp2UCS
bZlw06UAkaEjR7xjJfEX8nf+vUXQVMpPr1/T+nKHbaf2h6VNeN1l8gg2HyIMxa0k
yb5kWMNPPJLI/swBjPTtr5jXRGbEb78uiIiZ2FqjDb8yMEL1ftvJSNbSHYLb2X9a
Yf5EU4tkAhQz8oaPMuAcMsdH3/YcMyzATucYWxce4lnRzfAQN/b6MVJdNgUdDAGu
IDjBAvr8il4ij+16r++/37zPfUAtpfy80RAw3J5sUFmjD1GWbpKQGGetlPrMZA/6
L8rEMe8hlqQ++69xizA/snoG0UlgKlZQuB00qSF1zwsg+jf/EFqz3DnhzmnIUdAl
qNDdssPMrPlkZ4MbeyO2YHTYhuirhYws5Kdsp2VpPX826jmOI2Pfyx81VuV4XGIL
qUoEgafCNnxp6YPh1qUzpLSpAtvKjJ7k34AylX88gszGx/rN133pvXUvRottyf2+
0baaRBQTB09b0RljcCHUlpNVeLiyS+pnzyY+tB+gs6+C4mVl5y1p9NSM3drrYk8W
XvYIbNCO4DB2tTYF4suYIkYdl3eMfR5Vx+uUq1U+ypObErFllC0B4T4hHpHJeN3p
aHN6DaWIXsbNqwN0WtPhoeDuqG1Wfs7TJQ514DnjwExxLvQZ1E2F1rdSJlpkqCcH
y+oYXZYBeqN2d2BWEcYoAQTjvl/w9FBaQmwO6Nnq8pAl68Vl435ETbVhjmmNoiBj
cbOuJoNOVVa4IGjpk6uXOcLgQKkKcFfC+G1klD1zYrAtXPd5DAhXXzuXZSm1RX8A
iqtNEGRBDqYwdSzQcGKQapkVfOJt+XOqYcQYHR7nAI8=
`protect END_PROTECTED
