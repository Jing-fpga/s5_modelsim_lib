`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yBDY65w6BQ+uT6Pyu7bIH4QPrZih3AXoa7wjxb5mkV4XzPvUs+pQBugx8D3YgIEJ
MLB7w40eHahhrAUAjjcQfacEMtEMGSs+cWmhGy7BUUoG0LUYfUA5bV9vlKm2mBJB
MDFsT0eewJPEmLYMRAkwzM5nUlyc81THFqRKmemIORCnc/nqv0K2zrIoFvl1xoxC
jdmxZWWOroo3c0W0aikz3VbBZ6qQfAIP2mxC7zjlk6OaMDBjOgCpQ30hYBjD+dpV
Mm+ZEc5SKlbuG6O38NqdWdSj1NJIPgkmewl6/0MpgsMV9Jln90SK33xL3p9oqYyB
QzDZN+UlQ5ijljAqGoVhxsDH4rpDhbqNEoA8EZMAlPKmRErf4L8JZNElD18gArtp
+cqrZBLOKmrFR90SJKrRB248mPL9XsGrqCT6HHZqvKjSWPD3XOTHQBnx9ACFtfbx
z805pRxltNBDjQomubh42Mn7EUbGpzXtAed70cZnJn8IYZ8QIWDQHDOPLPtrQwE5
jER06ou4ftsoyTYyuw8UCFBYwpIxNLPJA7RjcamIy8sph1gNFsF4OVjzCH9NUHi/
fpT5vLivaSuTPyraEVxtlHrfK0/rNht77foZv6AAszpSIbMT9WUZNEt7BJH8rdlG
7D2N0khDx1m+J8AQBUyzbLEhB1aRL4wCILlcxNPKGj/HidwD7aTWaUOXmwIfSV1V
hQ0raOWheDAsw7bUsICXSqP2VGECDroEu8AuTRrRf2AVmyTcEmgGDIfocl3Lop4k
BDMKL47pihdaFS3yZJBsMzbJXV+VJkwcgco+yarue6tTGFHxgDQHFtMBT2R5jNC4
ExL2CtlgqBHybxjTQHvcncxfeuyosgss4+5C6T+LTnTZr0xxFaoK2AW16oK4CGRe
Mv9WYH5qFMHC5/PE0PiprsWduxWLnbQ/iNp5qZ0R0Ww=
`protect END_PROTECTED
