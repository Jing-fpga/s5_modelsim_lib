`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZSVKUR/LiPQfU7eTfuhrp+NiP6G2bijkEptxfyX5kqIiOI9rmZnHw1wMpEKjLv0+
BY6qj7AUjOC2bacZBIY9+syLkf9S0Wg6cKp4ciqGdLBvn5kyeAWsNGAxM5pjxn2R
bPH1+/UwthXDIBbHP6YzCfI0kzJGe/etEyh5xXd4Qzyx/pveaTHpgfUa5WinWHXG
xXH0HRZPL/TVAAHk2UaMUll2EvCDiAltHDQNyU7e8Rt/ymnVsCTL+oDP9/QHEYDi
d3u7gSrLvHG96+A4QAIvuCcVdelx0xx/vDXC7iWVHUamGhGgQosV6XiQ6mknZ+d4
q3Z1ymQq8opoXis1BE0OubsHZzJ82X5BTPGuw+5h4ysqNbEyLi6N2GTcd1PT95tX
/+7YuSaYdM9cQPVRzAm30ep00wT4iBOSRAVXbgRAfIC3gJaMgqxESNvFlJy9Tb3s
zrF/InghycKKk/N0yufFIFUrCWIzWwHAY8pey9gHfJ8DY/Fb+QpiVzysdvJ97o1h
X+060pPVcTi6902Op9d0YawevBDrMIG36r+dsH1zrktk6uJ67t3e7weBS3IKXRSj
KKK4qqZXvxumT8VFldl7OZBYFlyb1GQM3i75IEMC9/tN1Xz4tWyNDiSuBVgIdL4p
EHWey6nluGRGIA1sNC79bCyqndKGZXSh4ZMgV50vaD6tEBFgz8QgxwAxrBLCpmsn
lVgszEJQxZFO5+ZFaQBLrlpMPtbiAxcGpaFZ381qv5VbA0efhcmjfhwirHK4QI0a
p75xb6HZs1waEg1c/X56YYcbbIeJwQ8nR7Y2Vly3aARjbaifnH4RwkhPOpcRB7Nj
vNoSfSdyjLWyJiNYezSCzn2z7EstusnJCD/VEf80F2sTd30nkGZJd4URnuJHjIQG
s+PftVzsWeKzFX5qD+fPzyqTz/rq7TGbiWwSoVe/OAf2FXrW+5xBEUaw7eJXnIqH
ZDq/ft4na5mobF/aQIlbcNkCr0xfd3N3VJy7QYuxPWsDQA03/uAkzy3pswsfJEza
joIlvnKYf+0B6IRZRzQQnHa3CadYtFNNzzYUk9kM0uOZjjPDo+sMXFxSTZqXvU6K
9WjGe1bQLK+LJetOgYBqpTfKMfXWL++FEO7ee0Te60MOLtbjHSIR10KXSHDX8RAV
MKt+/xgGrRWHOG3HB/Buqg==
`protect END_PROTECTED
