`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1JOs59jVfNVyQmsK0h2dmT2+0pVc9aEbaV2+fBsI1KVWvZ6TN6ih4+C46tVNVGPC
abaxH+pgoqiV84xF2XazbQV66M3fZvPuoRmi5lEowpRIwpBswqsnzNiOR3rw1p5m
HLLsjdm00gwkRa0oilDnC1q2BiIGfovannmRp3KKIG51bEqneDyJYP3Gb++pPlLp
ZN5emTydRVcY1deZijnMOQ4AgKm2U9omnrfJoNxdVHkEfZ/8ObLPqBSifM4FXJgV
4acSUhNjtQFiL1nPH6y51BCBIu4Jb5J8bPppnLgmZY0UcFIGrvGS6fT+Lco6VJyd
+E1w4ijN584eGsFla66WlFYG0zBEbAbuxwTrUk/0U/XuiF2t2L5x8iJE1sIHGWms
5SUfMmkhnZCFKRwwlUenPI7CPe9j3WIgPAx9kHAATwDuZiiX6uZ/sIv4/TIP13rm
ZmR13HQ6ly539lCMQ6W7Nul4aNlFmZ8edfl1YQpKTWuZNeA2ArA7+/EWDbF6iDlV
QlSdla4q0kWpDCYx6BX8cSRnevMT52C70SlX1LH2emJtg5KTs6TfCY5bFj4yLxHo
uqGYofMwrFq/1phPzOeNOq7kA3SIU24F0YXM0j1pe2C5aWiOobajv7WYqiITDwI/
fpRPpD/vC2P52Ra9gVykBz9SYn1FcUWGJDuGLJiekIgH2Hs7v2aUvQiW6cHKIIqV
FwKoq5Q2OtN6ynIg/P9/bKXGkw2DQsnlP1VzwyhYLfrlO7SdIss5Kgt4A9YmU415
pvfpBpRtI2IO+e/ge7Z7MzQWElZEQcp80OpQe6pt/0icLT5u4hQ8NfBhuBxy6qXV
akKSLXa9RkSDWVJcCgsGYH0/5NBCcG0pLR5GC1sc2Mc=
`protect END_PROTECTED
