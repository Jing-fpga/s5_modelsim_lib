`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O8jfZPf8hDnj16Gl+4XdImICKTJTqiGzeZB8wzgA5GkOrKILgkz/wNah/uhPv2MS
zoZVEU5XC9eXcJM8IN6vw8r/7VJ5eF28xjDiEpcWg2MER6zHAyNQCzp1rsK8GEvh
4urGXZpIUKn2pLhqBdySLzU4Ezl3bYRReZdSJ42TDkopEaF17kryRXiROLjL1qI4
MTd0IyxGwjBwrwfJ1+PV7Obw4T+RJIPf+6jyrESE7Y69QosXeCkoUMvkkzCpPQod
PUaJ5vhzF3wepycaJ0cuPaQd7yM8jjP7cbI/Dc1P92AqXHNyS55XKZUetS5FlksZ
VMpaEZJXqxI1IRH2IQ4MQPUXesPVfHPuqdWOd789ErOol5ISZgXU3S9Cokyp9XWX
GgtOqMkJQG+I/xKFf+BrgBiFoe2BxwnkcEOe9DayOfOTuNOFdzSIraEOd/psA4ql
o6w1beEnaWH5LbCc0b4pzSOtsts2QJe6rB5EU3gKhXSqE+DtddiOS4gB1Q+Wbdfb
TMj0z2yGMrxmVWMlBzITD8xaXGVibO0e5Snq9SoAQhxUkHzkBtTHABrZ19dOcSgh
ohI7sKVOVB9Rw19cDTRA2DpyQcUsGE+nFVa4rFMQyvCtLPR+4Nx/sfJ6F+MbmcaF
lU7IlEuQp0ZX1STH5vkUG5/IzZ+l5lcpkvcY+3eCTS/spkEXgtdnT016JI9LCql4
DUMraAK0f29TD7ycEAdDffJVZmZ56K8F0zlqNdJQ0W7hGs2HGpvlT+kRBuF0bbvi
PZHFI42OM0MIdaO5MkaJw3TyIGw2AbbYQeCAQx+JVFoYkd1SamtZtr7A/iVU9exm
nkGkl7kY9grJftrLllczOvk6RWdMHCkTBEfr4NN7G/i1T97+zljdtZWWw5YB3RDc
nPOfNLEe0moxfdmkurYUfhGzT6RtxF7O4+onQrZmzibNcOduuLsshExwBr1LKEGe
sstgzY6iWTi4CzCpunMzXuu9GyEaYJucNkHva1HeSDp22wjkqTpfZhJ0XlG6Vu1/
JFKZHwUZ/2EnWJdp2ogIh47FpffwVA/n7NfJ2aKi8zDA95NZYLlmx/gM7tF0Trqn
eotFViRwekd9EXb32TF0jZybfT6DJiS7vBSf+9XGsIOxpRmoWyFruQkKS9xIkb21
riA3MHNYweTELlBPxOPKVngyHrasCeRFe8oSR/dDA/OqfbY5rcJnSjteU/lvWbgJ
iObcuIpv21AQEJjDgkFe4Dmn5sO/9swtzldkjz65VEp8gNuKt2hAnb3IM0vxydT0
s0uUlHGUw5lz4SOhSqLK3RfQM5toiK8IqJbqbhsbpwVR1MHJXqkMITbGxZn+GwX4
pnhFz0GuOcVzBImh1XvB8okOBvnhvIcvhTbHSa+bTznT1BMZP0XOdkowrkUiG+2I
YgXIDB9eB2RaGXNgxSGzWg8f6QmwoeQ/bWT9gL+kwOekIs1oKoekjkKiddszIMeR
jh8ajdMw/mEe9mHeDZaVCLjaZiefz4GLzPtYM8tJfF4FlucOeaL6q+fuXAWNsCQR
76j1M8ZxHUgR0vVAfhlnfqpAdlcSYtpg/LeY2NUnQWkYnw8Cj3onLNq/OhgzHRQM
b4yHJYizkDI5fLk61W9lljQ5rufCO8rF4LzF94o4TkaF772MSwZV58qJlGM7Gagc
pS3aOoNGGaS4AN/DimOlEGpqwEtTIuYWrCS14+Ub9AJf2r4FDj0TbIEYwLstZVAx
n06AeossmiC6lwzBCxnp1E/sSZniqrTC4PjPhaOzTf8dpQZCYmWaZzOKSElSc5La
yy2oa8W/fBn8IoMSeEq/lNBICfY7YS+qjs461jEIOiVVhBC2ozszPaaZqZGt73bn
V3PFy1Uh4e2tfNd0wpKDWiwxD1L4XQ4SuO6flbeYhu5aD+H5pJwR+cuEsQyQbNvF
bibV1C+LexEgZ/QwOyArk6V28Ymhx9Hvk9qY3wTMi4AgbfsaVkpyA8ZnVgVF0Rv5
iBPr2tqi9QoWY4wuViG9TqyxAj6skg8LTzXYQMMh9DFKs3Qt3y1t3/L6s4FpYyqC
3NRv6jrqnAsVW24nP37b/V8vAC8e5H0+1K/sSlulLHPl7g2hA7PJWggNRg+4BLo6
pEC+iW2KWnig/nj8DDOWFPnyHMT4+o8wGn6Q6LsN454Yw2vbcc8LVoDBneFY3B9N
8JIobFBKBuMUpcMnpJhQ8INSyA79j98pwfqE+lsVPyP3ekdy9oA1HlkDJAYpx54Q
uRgw0etGyb/fiG5xkqdfIUA37270+8yDB8PEfHhmKajAdLJljX38m3+m7rFmbWJL
F/Y69r5usPyO1wLwkKg2lDAhZ1pLftmAZhOxtIrP+No27TSdVDaxnscl81F9ClNn
1zF4qI4mJolYV2cBRha7fmpm2VRAGM+h0OlrlZceAJYtoYzst9YoJZpoxC52pAta
ciwQGzNQeZCiNm3qkP01Ifo0rjpqCJKYrU8NJ44U5zhDtB5axFfO3VFxbRWVk+Z0
Efc891NGDzVXX9V7n0FcO/SOp6CNeA9kDF3jGCVEEPi/rr7u+cU9AV5vfhhkcRT3
6fbVpEEPQdShRCPO9axkBC3sN42iTRXZDLnvRgZcSV2UJRi/+riGTDh3njRWG1XC
n1x9Mzdzu8K8HBcFI0HtWdJzxXNSCBuXmIw54IHrfGM=
`protect END_PROTECTED
