`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S5HPEXPWQ6W+Kr4oGDK5jdM83g4tBROXIAUT9ipLcZv4ab0Bg5U84ZBny0vW9nTz
/DZS9B+QzMASkj7KJ5Rq4usUPHQeRj1WOb1g211YOhTwTu0SMMgzKxe5t9gf09TQ
EKsxfPiGTxwRM4GtYVhVPTj70VyZ1YZsA+ZIh9td9i0wCa2JinJIVgQy7oMJk4g7
Ga921stv+YZSof3FxUCexBca8n/FBoyuB/NxRXpz1gTZIOWJDvCv0izNX9sudAX4
jAZX3SYiX1j+q5y2tg1W0IauygfUn/OtZcoWJDTqXITqFTw1rX7Hnvky+L0Y6Dqe
Wm3w/RhKHuRPC0SjCfqtm7eh3A6Aa/c9ZeSNI1hZP/hLkuhhBpS3Uak9BD3L4kwg
Ty3ZFB/L1FncqqPpI1WZXZze0Ix8QAlOB4qRh9QJvuLllYHsG+5Ni5dA5Eu7LubD
AF6+1QOMRw/s6ruxwgSt5fhp0z4gyeL1Cv1vH2+X5y6KWo68D7C9u9s+752tnrZz
sqVAmH3PKps+wPMpt8DAswks69cJUQ4GD4qObbdV+9uVPzm70q215OanDnbE9JSm
g6YIkfLUdLOGXtoCMJiqFLSzONAcad/OfZhV76IygRgSV0tzJfkoLgMAIhxqbrCq
58UrbJIj2OChYBbMfRF4XICoSZAMrDaSmjtSMIZPKcjiOQQ/cVTJKRDkAWad+hUT
4wx6lHV3IOJlRivbqzoHq1Vj9KZItqp+Myym+YyR1l1z0+Btk0Mu3Zens3Fewuv2
vn7VXa17cs4CGCNUkm4u7nNxqJSElwiQKDgFjlPOXzfBqS+fLc5L1olbWQhYb/Qo
U31oXb+5dQi+1zpjMa/FZ/4rHY/F14jIj4YTcdGhwgSGBS4qgalcVh8qNhuQsxpR
bAKquXpUvO/vnjanbrrsXoaPzSMlhHhbgSn0jjwrtwI2FHyQir532XNsDbf0PmVJ
vX9sMHRNjQEDK6OmtJt7S/ZpYjnJHfTOyLEI0w37+eTztcdvwOtPCsLfJnLUPwe1
2clrV2j0S5x6VkHafcYxSoAyNs4otVljBLleOWrKk6YL9jaXGgtcNLR1yWKYL1Zg
COe73hQodO0USr3Tb+c8xKKYXx2AthUS8xV68FurJAG3MU0MZyuvk0Qh5X2I0ZuC
jw6OoDNPEZPcRIlh/q5A+GGQS1B2bRRMDTG1YWoU/xoFLy2Wj/uY6239vAit/ASC
biFksxHozxq8mK47IAYFa0i+gzju7mH86bvFlMEGeml5YqvDr/355nXvaLhNVfQF
ikWHT7dLGbpbv/AEFK0GItnIrvvabtL7AtatGkZ3a7owMsyEUqgAc521tFvkU/ye
r3YU45i9CZKByAHA1IYzwQb5tcdFmvp+AoGquicKmAjLzR3ZXDsL9Wno+Bp92Vci
x2lHB6b4/0Wv3DkVp236YVnuHvI21dNkHFH19KojacByswu3hfmcMTTwNWsmhlZB
DwsJwfZNKATlgUdnfBc0GSH6pXhD23d2DOtYa4rn5o5X5ash0cp/Th90XTlQ3wBO
OxZ1x/STEb7aXefjrfZeVmy0zlo9fHUL+ewf3aAWDsMTXz0drjF6fsf00TFPE05t
pTOy749zFHJNyRdPNluHSVA6/ZlBBInfuo4QvcLUIh3FkHv61aoSjfAicjjF8p9x
/W6grwjc8n7ntEOjN8xHqschFNilcBcCS1PuRwO5W7evGqgyAVhSaeiAnUgJLyJ1
X/on2o+PssR2vL1Vt5uxLLtOeeOGZVV86CiNWxmSgJiJz5OFufS7oXvORy38n1Um
G5egIy6O7OHTo1g8OL6p+N2zIWE2j1ORNM8cY1pLBpjjWT7s8sixpXzp0x0ki7TC
QlADPF7nS8M4BTlgdCV0uJF8ZZe82LTRGR5q6AwLgXE0NQ8yKOmkYtfkhmHXgUfs
6gisWryjr5pT3gU8e1KFiJUsccu7IKf48K1sSybUH6PU9mwxoC/1UYvPrEoolR39
LWyGCEotcvHx9vsPpGMtTo+J53ukBq0D4IctjX8NCvpexav1dlrKzHzGbDXwIcY9
WXVwLnOWScjcj4y9Wg8dkyg0grVtCnK6g+ar9yfsInpjFrpmnBHZHcAsqIblz1QY
v4732fosfzYFFT9h07Sy1AQr75TBQSJRS5m6rBEY5J9eGxpJJqr1G3Ot9BYhTuDR
NZkP7onTJ26YF89ft5vPf8c/LJ/1H9TcFngbQuK0LiSAYpK9YtTppviecNpvQ7wH
pH4zdDjdmD3WpWybIl+wEoudI/quzXg6PXq9cISB3vMGKnB/Y0N1uCGB1NVDNYl1
uryx318KQ27iTZLhOYyD2GYSTD4f/cTOC5noEK7WU+G08ciBLZ8s05gUr9ZEvaPI
wCHm+u1J0HUzbyhjqHHtiKc00ctb8xYJLf1p0tGJbt4CzxmiD/ILh7cBOZwwYEC/
XHOJI2jV1E0yMaTuBOJ0isdNJSBHgYV/SaNuFIgVGVqtb7q9ZR9jsLqBjrbDM69S
qwnA5WANHFdyL/7ElYpSwucAEmC7Mr6NRBRwS/YJ2BYWspbmcTioHQFio3PmCKsW
h8LKlt+sq0KsZW68MG5gPMCNOsBuzdXWENOwwj89oyVJE1RfFhgApJxGluT3qvMF
zXkSmvslCvGFCCp/BlfUNoPBYWspyz1xjmSTY3OJTrMW+HVdvZk1uKc849lQ9sQg
yeR+3+rzAw2RS7+fYK+gsYKjsL5o4N4Y+fuJzYOoHSvj2tSE7ICfyLg72MQUi0+r
HD/b5BNptOWL/H2dD57OsPMCmMvC8p+kQ0JiZGOtjcJcUlfz3TR9g8VEkPe8JiZu
7FSBdWVMBuug0iF4dq6YD5uM8IWTv9mW+wzV1e9VzmS1WcdkAkX3D5yQjEvPj4Y0
fbgxaKz1LlaoOA53kiuuE/l5fYaVk3nWGZPhaV5nGv8NLO3oUV1RVQjgwas2a9J3
46dLklSFVUD4w1r3cdxH3O1WQEd1nijfHUFp0egpYy9iyekx9+IYUL6OLGJYAisa
+OH2Iak9OucDXhedNaCi+Le+qANuCBClqSIUsJfv17WKecNv2ckE2O0Xu3tp7YZD
Os0K38BLSwMl8SUVhjexwEBGYd7VpV64NrvOc0mYtZlQ9ZP+0Y9iQ8Kw0WQ51nts
RESmQSOnrNkJt+X2gOxqCKVPeSPOmUgCIKfkZjPIuZI3frkbbjvIcR9cQHCul5NS
19GQFRPvOQpdeqSiG1GaGM1RVOp5t4GxxT90HkaFzxg7Bn4DNMsk4XZfr0YvkysB
QV+PIlb65EfuCu8FxHxLZ+GJLUnEsXiY9E70ByVRZ48jhfI6rJmQH3JsUDMQ4NPd
MrOa+qCWHLmi66GMuWXdqhQnaB05hlkaNLt2Eb8Fvqx1FliLLvMs+038KYcVlokV
hJl5clYdV9Py/Cc8z75pMuozCYLyjBxpIuLRb1DlMcbrrEcN0FIPlXMInmhzvLlI
/yCqE929K/pXxbmHYQYtbpixY2wLuqQj0anb2+ADeuKzBvkBVTfdbZkAVE/FGXCT
kiAluM38sUWvCvMhzpzGpXiJTj5dEWEfYRe0dqLArpuDBP1NmEDuBlw/z3pnCS47
SkHPBKAzho5yTuyJGX2VPSiJWXUgEahft+zaXT9Rtj1CEP2HaniYrtsJuTGsJ+FA
NuIFZcesJPzzSCCeAgq5AI1BDBHWBwJNGUHJvD7wYYlTsWaxDDb54oj43guRy1Fh
33jBFA8cqiNh3jdMr2kyYRypeOGjsHdCBuGyES5V9ACrk6PpKewiQBTfbHRlHpy/
xN+Zqlu7u1hhP4HRAGcxQ3Mg9z8iufiHW/jJC2hgZDUjZCMIZzQqeyDd3W+BInwn
vGU+olNoL9Pfinxa69U4VyE3s5hNWgF48TjMDd0+r1cdBYRCWurkv/6GHqkU2RjZ
2veZK0nY9q+9F7DnUI1091H21naCg6l3CWEMFsEBg7Kf3n0NA/HMPkiwHWaUfC/T
fxjP6bfIrVNgrWoOQLkA+SmAgO9EEhkaGwqUKTjeSKOds9RAofwVMIKq+eLwlGKr
tWTpzyPiexVonwLwe0gwaKfwROKC9GP2TxFY0dSnqKlwFIinN00AIydNA/gEcIpy
HYiv8vpsMyUxNOozkSdue62ROP5wO9R4XzahKskhEIddDrgVsNw/MFhmq2+Lsyg1
gs+0gxsos07AZHtwlHRNtYuTqCaDX1ewTTXdxI1ZPfE2xfLOP0dC+NAa8eHTkntI
LYUXX/g2at8KPrrkLiGMIEiPBBbbMIP6p9PFdlIWFAF9Eg9ymjGPwbbxsC4eRlCw
3816JKSWZFWMrB97OOCil2M5XpBRRKyyzuD3adFp99E1obweX0nmDbi4/D5x0Hth
Z4nm403O+4RPKZiLDddt7zz0R0PBeH7JP93eQKe027SwEpiZlWE8G8qhhqwY0lsN
0CCr/AMPbFgP5kOMzu9TtcqVzFD+ocYVB+52pnacx2w=
`protect END_PROTECTED
