`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SiAF7zlPBhNKuKVcZahoieSj6pZZetvmSYZxXR436F+lJRrXWSH0TzGWwCZCsxeu
1VlWuWYX9wBHBXek5O4wQ7JOvIRg5pOCwR3h0GF/aXoXfV3ewf5TYGIIWX6VX6gf
URX9W2yrp5TyoBoDEFdGfEiewKpXCGQXvfkxQSnd9dY8taOxqj0DUi72kpIq8xx5
GK0zSlC2gLaRc45wp6RqxNwmzAXYyy32nHC4Ifc6qDmUsXSnnoqAXT7My04ojkAU
xHU6f2S8MffMfFfu3qqtDkcWqPrFC7sfxQ2TfbUUI6EhDKGzh5Kl6bOdYVpf/+Yv
QdbR8hDzYNwQ/p5lINVYhS6kyuOwkkM8qdKT68XviScoxrrF5MNPGSBge0w+sl+6
gpAvsZp+SQO8J6tdC0w9WGqCkkziXbytOUFdnxYgriMw/Zp+ZqM4BIC4kywkmMkw
E69qvRADy7q+niCNI52vb31j6E3GlMFViYyoM6kpwKVghpKGCGQPK3Ii1ZJvhBjZ
QsLvYj6Yr1bODQExEdebnLBijWBrCBYFOUrvoyQYtWvXuLOUgc+wfBfMo9obKGIH
yjZADozKtXlh1z9MAdWPHwqBK1t+MjmfG9ph97c+DvI8mHWs9lMRgkDQyX+4GzLP
c81Pv9PrxGbvsydkWERaDQsF3COWAXBwB3B6Hm+LWmvfZi4Z86wNwXE11qOfT+Mm
jglV4l7y/54r+LcuyHa+hVc0noN3k696kZ5k12MDGLHoEp7+bfZ7mMzzt7koSjKx
iQzpK/92QomNCnqWQOJGBHUs0B6GwuoQa8cZ9OmFAfOJlioHJkNMDUwAehV8qPr/
RmFT6a0fT4yXBXJ4P/T3ogL8F8uZtWn/IWR2fxr/udgyVnxhCQOQMYB67WOuv+zL
rXulYzC/XZOnQ3U3Nc5+nLkkskCEzI/ZGNLac+ArZDs5n1+5g+Poyi+ExteluDsk
SLvsdLH2PpJ60j2QjhGkr2X7IHbkn5E9+7uQNKVvoplUiuw1ULxhOkv4rbbd9H7C
PGmRIYGId+2ddzrvvTeZn02MolEjVJZT9zFLfd6/IO+5tRSq4NhopbUXN5brRLGV
82FPO7vnedlwR43szElLJC5/7rgN1Kl2jyvJEBKVaG8SDPpOkESfB2QqcmnoA6Tf
nIYAKyYMPB9rnS4my7pr6iMgl7e4GKFyHcOefxXBkPpKmDot8gPG4MqZc5D3ayrt
gVh8kfSlM4jy8LkYbICVefqo1WeVYBVlBcoISno7WCJ49Xg/q/OAn+rtdwK2Kmw6
POK+UTI8lMKE7HaDShi540inZwApPzl5yfAEItYMnp/mA6QfHDVIuf/TZfePS6va
7MXuK82QleF6HTHz87oIXnWub7NkztapxC+fCSHS7Ihxq5h80aFWm8zQCJaq9VUk
I/Gs9zfGRR50DolC62OMpGXCdAZvzn09DcCeQuwy4uP3oZR8zM3EHV3tsCk4KdSk
3hq94NqXbdi8HFsD4mCQ2BguqJJNU8T6X9XABuYLYdAPNkkazpwPw9fGkYlZyX87
2zcuIUGy++wfPRXF3uP+ydZ+qZhPt/37WE9FYTyVMuWeTEDetk2lm/IARQ1p4y/H
lA0227qfN50ag3catlvtnyaVgkenTKS7+M7ZoQEEEpJCfuF45S56bM8CEWIleKBQ
sxDOGMMAlZlpiBLicXM9Rh2celXNfq+Tm0oEFCqImr0Z1YNwz1T8eBO1rH1wt3PR
pz3PzIERPwZ3oEeHeaGx7dgH8G7LOI/Z00RUq1jy1oyexZJo+oAU8H1Y9Qi9gXcU
WLzKx93sKrQc5h/yIWA31m+Api0Fiy8g76mL+p2HEm0E1DMSpoiZ30AJ8/1zXz3x
X82K3yaGas3wrAfLmzg7f5kNlt9ThJmbYebPNdK8iLCQCPimOQ1wV2Asem2E7Puy
TmB8K6oEkCDXAN+r3eDd8fa7AB8lTDq8z/ubSmi/0EvI3vsPN+UHAEIIOhzLT2O5
cWTpF7Q72t+Njtiyg9lSsKgUhzMhwLgkyElNBNDVAQ1Q5a2psqQQfUSW3eezrqTR
uskrPvUJLYgZ3P62WXTb8Xlh98HRMOC6cj4BU2PIxZHrR7E0LHW06oOS/REFxk7A
2heNQQe6cnsF7MgQZeN8k41u36gSNTSiNGvO99B5dE6Re1suKayNWU7TuyK78IWL
D89HI8+KSje+/6Yuhf6/6t+n4dQEUGrkSxfV3smG9FhAKb7rZbv46Ioz7oZQFhZ6
OzoZtAdV/x8T/u/XQivOUfbaVKSqocm4GsT2KSpGWOTMG1wCI3V3gzZg+jilObCQ
Le+CXL7VlCyj+paYPcFylKzQf57ryAAJwtm4eW7hsW1bq/q0feYUeeNHhpiKA3D1
jZWbC6Fb14RHS/2BOLVIIo5k6lmrxQcGj1Ru5ikCqwNZSHpxUvT+n0lJJ5ukV/gD
y3z5rA1F+D9afyiwuLF/Rt9Usq/Gic9JJIg6WXCSoIMWzvV5inkzdUEDqEO+I2sO
NDsTUCl3ZiNmj3hLBl1KWQJipiLwhaFWM/POvqGYl58mpDM22C4dKs8u2V21M9cE
sTFK9LHjGl4mJ1xtf0jGd2PJRjBjBy/IlANJXq3vFhu7JRp8swXmesduf9V/di+O
1pmrYFXSX1fCVWriMQ5VHN544ZI2jy0oMf4Iz5CB996R6cUODNbejmN9pOUM9GRY
7uEc7E2ama/R6jc1hNJVTEjivo6VYBevTkww1AGYu9pUOW8GMAW1G4uWnMrHzWgS
vHZ8l4af+DpVZ2fHOZ/5veXJLMI3rrffH4SsiXrpIJ6+DNLbHUhGdu6hun8lxC20
iTF2BOxSHqy8HMrerQltDfBiB4dSzNFPB691dkLCOKKUb5lbvgkqIeqzcPfrenZd
obbcuWfSU5wHX1YzQfwSE5QH8lzKdmhISXNDjC0bFLn5XwFkid8ndHZzMS7rXOnR
lT36mtdjPdXggiccq44suGzUMmT1YrvYai80GXmwYhoTANwdsTTRMu3ORh1byW88
wAZx+DuYw4myzp2v7aDjMDfl2WVYtgcEt2fYcPRFOx57fF35XvJ6YGBbCMpY0Dcr
1eLLI79HVdA8e4CRbLnGHS3RgW/ingU1Yk3DikfmnAaPBhs4vfMXK/QOoIsi2wgh
tFb4IK54f3ZOKMhU0WmKXplyKbeFJ4geTgNLTCMgfKQ0uiNXScPDXhuk8/W4GoW8
TnAXGMG3ZR/Tdud4WVkaUKWiILZP6blPlz9ZEtQ8xOtai1F9xEU1x1/wRLwS2diH
poe1KU9lK8947hIeki68cQjz8EFVzAThNmCZ2PPf/ojO9CF0Pw2svRUGyWKvjAqY
MgCu8OUxd3jeJWKQqr3Hg+D5w6DYvyh0xP51DmYQni4uedT40fKWxW9KWHL9UdiE
QkiGW6Oq9KPxx3YAfMpb3Bij8eQMERvJ+NVx42TBMdzgm2LQTyxIiz7QVzJeM0+z
`protect END_PROTECTED
