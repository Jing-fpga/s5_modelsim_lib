`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tv1mzgCv9u1Qv/D2dTzuixm5ehrRvv21zcHmCd6tFEBFu74mHadPlXZs67qoN1W8
Mlla1E/aHwvmGmskqVMLPT+QEtlaoCBA41Y0cTmUYcMhHXz+x5hYBJ/e1vKiKYpy
QXrfdCWIRFvlbUHeKmkdKs9nVOHNVrNdqqDof5wgrRlDjNd/dXnQlH5JjJTKWjDz
LFZXxSoJlewJuRlj9dZj8qcdqN8ie6O25LEK5P4eMATMPl39TVGtuV4avrGcZk+t
Yl6y4xiXKI3c+owFOk+59J43Am65GyBeXHOG3y3wYY8+iqIubF6wV5oJ2YZSuG+h
1XdHBB9BcOmnTZjb3q3wSCoqnUiq5ev+C7BrTAf1axy650oji379xAcJHtInbUrb
UGav9SqDa53aN/R/j19uvyUPJJOjOG3Vz+Uq9CLX4lyRTIeKCjfmYZYsn8TJnEc+
blH6PEd4qKKdKo3Xi3TPbvuFF+Kms8v1U7rl3eP06YLipQs8a91d18N8yOpkRi0W
vxFfeNH+YwlTeBc3n5zkEajs152BvNvhr6BEGvnyQZd74B0Gy1uNw4o0xBYroAkg
Gu++fzXYcon776cizs/Mr7dhMaoLE7hgkWi890cgn+KzuGrQta8PVuldHH+/eN8A
SxlQRyhHh5U5144L/smjmSecMDoP2hPMTHy2Xz8987akLkKnbidWhaoMvZvgOh1F
GhR5Lev6XEmyc1JTXoTSzdB8eA+jVgps06sTeBibLKmuqHGmRM7A3+8XF3cG+ZXk
9M8Ex6Dhil+67cSFuEloBp07IwrZSxzJPma8A8R4M+PTHSS28ofFFCpjVD4tjCrF
oVB98ikS7Zmac5MpruWlxUpjRpOChKRFQsKiTMIeK0jAX3rRm7M/ZG6LRBBARHvQ
6MbpdlB9N0y/rkQlI2HhEqOQlh8tOSEz4dyFdhl/qDKMcJxYMYDoSy02fC9DrUhP
WuLSa4mUlUjnlsOSmaa2XX0DcH9jkFdUNqRr6mC2BAFn5IspeOpH5ntaj/b6mgFh
qjssf4tAEqzI5jUQ28bt32xDbXznBg3Ol7Q8SBrSjC8MpO0LIokN5htgThCpkcqv
EEDjEejSD7HiQNSAiVpaSmc/o0LUbzm1Tp3CyJNVPIqDO+zJ3DtgfRyGIpdwHmdz
fNx1Kynd8TYeIsc5MHjgT7c4bqNUg0keTeod5A+M570GWJWtpvAGjDakbJso0VBS
b9ec0un3RxEqaNf3xUQWCbs393u8a1Nl1mmLrfS1yHPWDw/PCtN9Xawbf3Qig3aF
9LDjEh1ssQkCDpmjo9NsKxm97J0+igJ9ldB6iX/8c+A=
`protect END_PROTECTED
