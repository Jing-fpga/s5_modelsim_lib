library verilog;
use verilog.vl_types.all;
entity step_analysis is
    generic(
        UA3202          : vl_logic_vector(0 to 47) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        UA3107          : vl_logic_vector(0 to 47) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1);
        UA3113          : vl_logic_vector(0 to 47) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1);
        UA3115          : vl_logic_vector(0 to 47) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1);
        UA3201          : vl_logic_vector(0 to 47) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1);
        FLAG95          : integer := 20526397;
        FLAG96          : integer := 20526653;
        ST0_IDLE        : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        ST1_GET95       : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        ST2_GET96       : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        ST3_END         : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        ST4_HOST        : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        H0_IDLE         : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        H1_WRITE        : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        H2_DROP         : vl_logic_vector(0 to 1) := (Hi1, Hi0);
        R0_IDLE         : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        R1_TYPE1        : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        R2_TYPE2        : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        R3_DROP         : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        R4_HOST         : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0)
    );
    port(
        clk             : in     vl_logic;
        rstn            : in     vl_logic;
        csr_cnt_clr     : in     vl_logic;
        csr_fsm_restart : in     vl_logic;
        step_rx_sop     : in     vl_logic;
        step_rx_eop     : in     vl_logic;
        step_rx_vld     : in     vl_logic;
        step_rx_vld_bytes: in     vl_logic_vector(2 downto 0);
        step_rx_data    : in     vl_logic_vector(63 downto 0);
        step_rx_ultra   : in     vl_logic;
        fast_rx_rdy     : in     vl_logic;
        host_rx_rdy     : in     vl_logic;
        step_rx_rdy     : out    vl_logic;
        fast_rx_type    : out    vl_logic_vector(2 downto 0);
        fast_rx_sop     : out    vl_logic;
        fast_rx_eop     : out    vl_logic;
        fast_rx_vld     : out    vl_logic;
        fast_rx_vld_bytes: out    vl_logic_vector(2 downto 0);
        fast_rx_data    : out    vl_logic_vector(63 downto 0);
        host_rx_type    : out    vl_logic_vector(2 downto 0);
        host_rx_sop     : out    vl_logic;
        host_rx_eop     : out    vl_logic;
        host_rx_vld     : out    vl_logic;
        host_rx_vld_bytes: out    vl_logic_vector(2 downto 0);
        host_rx_data    : out    vl_logic_vector(63 downto 0);
        fast_3202_cnt   : out    vl_logic_vector(31 downto 0);
        fast_3107_cnt   : out    vl_logic_vector(31 downto 0);
        fast_3113_cnt   : out    vl_logic_vector(31 downto 0);
        fast_3115_cnt   : out    vl_logic_vector(31 downto 0);
        fast_3201_cnt   : out    vl_logic_vector(31 downto 0);
        host_pkt_cnt    : out    vl_logic_vector(31 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of UA3202 : constant is 1;
    attribute mti_svvh_generic_type of UA3107 : constant is 1;
    attribute mti_svvh_generic_type of UA3113 : constant is 1;
    attribute mti_svvh_generic_type of UA3115 : constant is 1;
    attribute mti_svvh_generic_type of UA3201 : constant is 1;
    attribute mti_svvh_generic_type of FLAG95 : constant is 1;
    attribute mti_svvh_generic_type of FLAG96 : constant is 1;
    attribute mti_svvh_generic_type of ST0_IDLE : constant is 1;
    attribute mti_svvh_generic_type of ST1_GET95 : constant is 1;
    attribute mti_svvh_generic_type of ST2_GET96 : constant is 1;
    attribute mti_svvh_generic_type of ST3_END : constant is 1;
    attribute mti_svvh_generic_type of ST4_HOST : constant is 1;
    attribute mti_svvh_generic_type of H0_IDLE : constant is 1;
    attribute mti_svvh_generic_type of H1_WRITE : constant is 1;
    attribute mti_svvh_generic_type of H2_DROP : constant is 1;
    attribute mti_svvh_generic_type of R0_IDLE : constant is 1;
    attribute mti_svvh_generic_type of R1_TYPE1 : constant is 1;
    attribute mti_svvh_generic_type of R2_TYPE2 : constant is 1;
    attribute mti_svvh_generic_type of R3_DROP : constant is 1;
    attribute mti_svvh_generic_type of R4_HOST : constant is 1;
end step_analysis;
