`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EzTvUN199kJTq1qoMmzQnZLevJ49eVrmZ2DZ+lxe1ccIeDS0cRorVkVJBPNJ4RvN
1EqP9BZiL6hjAK+8zHe62096ZPIdMNO93RHLupwviQipa05NC3deDy4F05JrrlOL
LnHzOsxdDXRGn0cWzsaCIIP3tVpsO0Ywb02kaveCCn2nYzoOvmtjaV178YE+ykd6
gAZocJrmwA/Uvk/f/L/2WM6xvJqGc8xLHEK8suwqzG9dUyqTWtbSeib1X5RNoYfF
DZxY1/21il3oZx3BjJJUpT/x+98KkRE7tQZZAxG3dnRep+O8rydZxKfDgK7yjsoX
Bf7Ov4WIJVUTycisVfjhsMJzz2uye3ndtaNT0BcEcMQ8/URQlTPCBbsEm3fayq1S
S8On78YgN4krhW1u38jN3Q6JnNeiEaanCpQA5hqrW/CBO2H6VHCbwjBHiP5L65ed
E2qeLvprFhSw78EZi5+g4VuduI3Mq/fXUil2YWIbHk/Uz1cFNsNWHBofIoPnDlpw
0kAlBbOUSfYlpyt/ubOjjYirr3vWGUmkpyVXr968R2G0RJluBWuzSK7pokd5+GOk
3ND0n+v91FpgLj6nVjRVrQGgTD7zuZg5CnA0BYd6wySfmlnm0yqHrgFeMOyLarH1
Q3Ujus71kHhW3D0HCG67exxirpfzUlGBWKRc5gqd7BkezKr8Jw5dolUdwOjyG3ov
qJXmjr5KZG9OuqhJLlhn8I/h6CuD5u8rRRjje+EjGKaMoNIO4uOiQ9ZKmblWhTeA
z/hgbd29UPUaoJezdFP2XRZHN0ak1wyudcHdNJqG6t8eJc6fsAHCpAbXCJ8wsWbl
GFGv/Q07zpxi03Yn9a3scqVaRwvX/zeFSSapZG2GiqQGG+kGQY80Z/AYFpSwzKbm
oF2PAFuCpgOrJh5QYZwxFDEaCYucsu45P5lG8aAuQTJkSCzzQccWZnhhI1CVy3G5
thVeDh93lXTByV1VjZZMFYPIS48zvhlzNngnC5bQ1j6ql3dbz64+OdtZ/yatmi2c
cBheTuaE4NacNragoMjGkY7ucnyUHZjrtmReVsSVwVkdyIxw9hU1aWO3Tln0ztAZ
KCA30QOsiinrj5kdnu8nZCYREs0PTWIQTOIGIwQ/CUeR0r7K6+Eq5usBx2+8ROan
+LWrhKnknW1nKgyWov3x/z4rYeMC36xM7hWC4jmFofjyHHzPN8XUA0krv0ZkIfrp
vpKPxox5PM0lMdz+8A7lYK8h2vkypCdLDJCxqolg9s84tfzAwylMbMi3psdN0eBX
VEStGzkqVWYEm6byEcirrwtYZsnES+xwl+ln2XOaZ+Igu8dt7altZVeAiHfU0LuG
Y/xoP20NTcEm8iYt8dkJf+7UnWTz7Zfnd+Y6Jt7HuiLzY+bb9KKzuaOT3pjPmpjE
JBt8sZQ9esa7yiSULe9MW6gXNO4NoqmQ2Bi1uVimsz+tJxX/1cwMnM0zDDCvjX6s
EA2RqJIggdIzY3l3V05UoGsEUN6ZbwhTM0anPPK26Lfl69ECzhKO2wyLFq/kg/lv
GYw3ljEZxTxM3Vqar8onkxxE9DJaeRZ0cOzHFHfjO3VpAZwlp/5bskBF4tSm3wlw
TWQL0gKgJB102qemZ5tx5fHrqglTE98Fu/mVtcanIDbFUfDW/nT/CMXoWI5JAf5W
FHcKMP/kdzmYCu/gnNiXPIS9/c3sFpedPhzJNlV2c/vH0uWvwoasUqmTtzVgqwou
RaMQB3KHToKJMzPc1m1OcgaFf8ShWoS15MSJuCaMjs16qP2GLx8aGy1sPhuMfN98
E3hT+zMn495zOV0+aTY/kSl8R/ncFIz6eoVLGD26BkCKEsqev3NfOTEAVGeKGQBq
NiMbcZ9u4uM2wi9pjtJOnOM7cq9FGvG+gSxY7MpK7eiB4oizwpALufZsFeVxqN9M
HMDYBR4JvTqVCsERG2XMDT+e6AbQb8J8WoeI2TV1MXF8v4Kc9nHPOUb9FnLE+Kdb
3xMVdC8GqozXEa9w6RCcSjOa+3NpMv9SK9zX9x4V0SugFomt3PFWHL0UkEJGbZEN
Zox5PR7YI1yd9zttRQ2VFQT20pPXo6L+Gtfqd23Y0xUTPNghk2iSVKpIML+Cu26V
36H2T6CM6niVxBXl23TvZ6rXY0hx87Rs0nXlAEMDa4CrOhOlHQScf2TgOxRC0GgF
9PzGX8xoLWMvZktPPEaHfTEeq42Qbfgp8irarBiw8/JQ6QEfla1cVjQRJO19bLWD
6I/ZU5+vw5npjYeXZ4C//8QxU4rbTFM2EEGS7LY9SbO/CK5AuaNiRVKEIVVjU8N3
YcYlBDPNS39me0K1GNtAz4Mii3gQMtirTNREKmsjUvYXsrMtHkwnTx5luIPm3OB7
VOdhpOYtgFiOJdhjUYmyFbRgOXUeD7Y/dSMuj7oMb1oO2ry7m59/3DNDRtd5IM7I
rDSzwey1jLpLyT6FVLuQeNBSnq2bcSd2W8dIhopqca464kWl98qpJuWsRwq2dW5D
szVjwSL9CzIYdZTXWZ7tEmDJ1UHcR8ywQd2xp7x0KJaEFQW6om7gWQyR5FlMp3Dv
k3W4jditGM/xZ2hgIJpz92j8kaagjpqgNl7ZBYh2lAFTFQ3FEFJvv5xomqmwkXno
OIeishp5rwVkIFUtE/obZRqrwX3RrsTsyZN7YCJ06FI=
`protect END_PROTECTED
