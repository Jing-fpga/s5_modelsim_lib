`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BgxuivJ01Xui3XFB9ISBpeRfbYPKmns0NrrCXRwu42fDrh6aNehxJDU00qtbxoXm
HMW59aqplXv1lAvnW3rdXlnwTb/3gDQ9WEdj2ohbT/F4m/xG5jbMadCBbivHDb3j
sUdCalyhjSrI+oC6jbmIy+xHyP9mm3Zv9wT+XUfHgW7/WkTM6YXIIRlRFvwyMDF9
UAN+0YxN7sKEPtguIsRtwXViwdHqR2SUejQdEmJetmG1UUA7b0ef+Mf6iILyAGwc
/YeM8slranj2pkwXW+3gWP65R14kSogmi52mg6gRTWZPw/QpFe6G1ZWICJ2pWrAd
twyPRrRKAoIb+yuqfwIGMzmpa2ZQqpi/bun2dgrIMkOwosCYTnxs86VqwX7jIQF/
IhMulPYavk/i9M8ocp939nJfKmkIeCkB1MdobMlaWVh7onTCsurIhvlvXK3H+iEe
BAKxLGL+1JKTQ2+XRv40bSM/O6ZqnSzVvXGEBTQROyPqIWs6b9ldK1DR3GscVLQ1
UJphi10O9dNuwvChGsVzXFMWcdxrXIm192RdFBrRbFAtzHb8VbdkHan3ImPJAGco
7cc7Hf9IdnADkjAJv6qXLYoyWlBBYJSS2dA3SATxmthe5xEJNAMPqrAQkwBT7I+q
`protect END_PROTECTED
