`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fF4Xd+yvs5Et/GlW2XEzAgsawuyBxVu5MIdfpjp+vFblafV/63hP+gdi8wzLB/UI
nIH1pryKM680+TDpGLgLDiay2u+IJnTlLrFSC2pGaZQFL6anI2dJZoJlLj74aE7I
jxPdl2bV6DekFtNfjsdO1q9lVaE8UTE+TDFUprDuiC2fuTFsHGM7D2vl4x5fSCfH
jZO0/dYIch12hG2WSGKaGtuSO2Eijr7v72qTPuTiAJOlRm6xpPrNiOlXprOGCwyy
o7jWx3dMS7b7KnLwmfMT3WRZhUt0P5nr59PQSCPewl0cnjxw7kZgAODm9+/2S9Io
41/QDeQZLOVT0MikYWDudSO+9b6g4e6kEtgm6Hw27rWJfN4coq5+fZ6SX7SjBg7S
znYokdVwuwhTGDLmNLA58LCpqpYeIAua5gZ+kgTrH0NHwLxwGfCp7LcF/XnmMPE7
/leLilfjle30IDQb0JwBBgaRxGthkgDVPulZ1+T5txXzupMuoMIm7tG6vlg3Kcdr
fqDizMPvjd7eRqM1wzC0rU0ityRnnDVQiGhtCqpG86dQdVPOp6ypCcYuZQkTa47D
GH9z7e/nycpZ1EXhErc2mRa/jEkf810ZXgNoQ6PORKChqm6C6EbLHIPf4+Zk+8Z4
hcBOhUx7NyTYtXwlpVntYabSp3vIlI/azwdbAzfGGhCAeXtEmTcvhyulL3maWk9S
JRr+em0cGTe9D0Zz5A7EN1+Ikbbjnww7qIx3j1T6Sl5WfN4y2EB9y+RizeuN/RFO
KTUgb8fPhMCqXXxSHD7oOcFxuppddpZov59eWJzFBIg=
`protect END_PROTECTED
