`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W+69bJasiC5/fPqTkORoLNlHMFvrPsh65JdHVKr8Ahf97IH7YYvoCHkp4tgVVr7X
smgmOCfHG4BKyEtfVIlaLL0SUPmFuMKEGCuSfiJTsNh8RF33oAQQX8vyO+R+6yaA
R5K3MX4r2XrOxmN+BldZTdWDMa5hNZm3f5Tf232/ksjUlcw6iG1NjHXdEbsZMIOI
Ou2dAvx8BExHGdiA2eAE02fb6M2iscsr5TUAr7PpX3aC1QYJXFHKFXGdKeTODqFu
KmVDhxJpvJ0TCizz9lt09Rnj2PMjuTvtAGXb2sW3CONS9ZJzssEcYjI4fDBDP2lW
wpFANaslrABE6prs0jMuYJC0LO2HBEWKbkPGlX210ER+3Rv7gqW0amqYvVgF/+RG
559xVozqasYx1DeEn+0iUdXSzp3AxfTbrr5TYkAsuUPzGPcE+w6WuiZFQiSAaA/U
59nIED35tOvt09MJ4eczOVOM09wJWO8mRauhHRnqmb9ksDUJukwAKfmkOkYmnIUq
NZunS+2s6XCOm0J734UsxFdHzL2CUGQDX2ICEptZZimC1gAnYkcXK2eWIyHEzoFU
yQX+mKC2Vj6/9xEl1EEE2AHA+GC/iupR/2OIz1g9FTcgvljtpSQJ+dpN7nAWl9T8
vK+jV5XC/ZUoXZYBUEXyMb9+b5VN6L+6RTSCVtmVIuFijWpQAKX24df32l/iAld5
mLV2WWv/Du0RLdh0Em2nQxuhhkyfhCuh1mAgL9h1BpBBnsdxHJdzoA+QBwNHUSOa
21Os+gklA2+hV5rTRKSBVFRT7XH6OCFNWu5FisOLUxRTVhiw7Jm3aRNfN5qa6qxQ
lXqeL5gtH7H6Yy3RE+JEtqhoP9+RQFYZnqlR8+L0BrCviWaJNIpGy+3CSiRzjzMs
`protect END_PROTECTED
