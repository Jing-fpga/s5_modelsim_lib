`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JUiCbigD2u7nUczPPIjeniSUU83llgx149gR1Zce8WXkseC+EUpJxRRLhQ7pnzS3
0RNEatYu9rX+caNvd+RzXOElJiTTinc7Irfd+c+PlsAEepDDdQSSX3jbhccsARa9
mG2oSfFTd5w8WLi+LjwcoQngXwFge1GdlO7icE7+pzWMOnyFvwBXBrPwosnMwMU6
8bh0y0bcA8vZqmpNvUdLTO8pYKUjl24/KtbUgq/AeqD3wcdkZWNygoljt/KH6PUX
ghyKY4i+t/xmLGB0YFZ77OdYmPbYca4OZKj03KOM1m1MHe3byXTTOhWXebVV3fA+
ckRuiJWTOqy9uBhWu9UWutrQP5LAc1Z02xs+6aU+i54ZaFDIzyRdr49jNg5GcB0o
t1tPbd9aH1h9NaAnV2lhFOmZK7xxWelVjqVNsYmXyWQKf0ZOtYfr1iZiLPiHgjym
kPmMLIdGBC0jk/y0CFmOuN37UbDKL9J0K8Bn8foNFINd5cDBCtC+q8Y/FJ29IMgh
JBAYSmPGV6blkI0ONbUgenhYSNHhq+S5H52pElCOBe1fABl7V7NJs9OiWk6FLavt
5AtaExt7E/Uxz693k7T1r2VJTBKIOcClwkSL1K45PuSemk2qdDfaYToT+xoWH66k
LazZTi+vRqwH6IF47TZ798lBI9EROJ72r3jf4PpOb6pSu0DA/0JHIAtuV5m9J5/+
EMAQaRy9pOYlEVwurKCfg58Rs5E5SfS+ntWt+wCMW716gdR2YXuAl4E1uKfjd33X
7Av1wOEAGjHr4ddpJw7Ifc6f7aOlk617+7f8HCNVGMuIeerJu4EGLt93jnkyJw3v
T06yVAJfV/UWuDKcR4XnsxTfNXa+G2snH8iOaJJyQlfR2dNq3qBkSdyFLZHS5IsH
iXlksxhCT+CB2BmxXjy7SUdJQgaLm3pW8tnq8z1pK47HKbuxsv0/R8sfLCgu/XuC
bzZjYLyoXkKKY9pK6yk8W0hOpjZfriK062LrlzCNGB7hMaSgqkxjMvc8CmtLKioC
Exaq+RyYnA2Ql5phwjoEiua7eS+alHQTAhzdqVXR8Dlw0XOimltUzV8aJVclIi6i
xhoEYQbmzeddiDOMHBUVs4DPPpHvVKBTCE8kSJO2Mbfj6HBQtBio7ojNfGd4195h
65Ap39lheni4DAv2B7ivgwjXEMtJcWLGCC+EiQAAEbLWicIA5f+vuf4AGaPjcIOv
0j4bIn1ogY/PW7o+8hptrRx5CB//EeH9YRLc14l7ukwC+S39igsPykXxmwMuWABU
C17SrixuYrnFVUqxHTFSPzaPdB2Xw3pgqUPL1PV9gCdQdjiNzKH8T6cF4lE471Q4
7Qx63Un7iW5bmTjppueqc2phx6LISFxRVdh2aGE9dHWn0piqkeGvHAKD6xSBiL5q
YI7CrkAOeMKxK8nQYjjTUnfxA9brEHdYwmr9mFe1XDa8/Ww7BSRkjHDXBgxZ1vO7
6CWZKEAJAAILjzsDwcpR/mnxQtZ7wms1QwyFR3P/d4GD3Pn9/DRD6VVVPtSQpWkF
pMGqqdDEFwd2fQQq6Ocp7RECQeSqQXP2nnhyceP4dXPdycJPD3Nkpvtxa2BgEGBr
4jhZDb2QzKz8m8cmjiTzHg3TFVsYOa8Lo3wgrakhxqK+44hisU/IFHq2cEClrJ6o
b5OZSxVmq/KqGBgaqJHW39qvR5+4Lk7GMPDvOrKyJJjEL5SEGxeSBKY27u0wNlQA
SQT8THyueMYDxJavQ0ZaYLRJQ4aucukWYIm8f2ibXF64tm1Qne03aAEn2pJPL0h/
AjE+wGedUjAiEQXSDwO+p/7JKm6PkkTWXlirqJyWlHGeSrb6r60L9U2TFk6kgyXy
9+whsBUXsnUoUyOT4MeCUwb1YM5ylFH2iJ+mPb1rDCeLiCstc5xy6Hr8kcUz2HcZ
PgJUtZxC6wImj8CkuIjQOpAUYkY4ac4NKbdgC4aQnelHsNQahYXvVRI5yRSh9XXw
ranU3CcgAxsihhca7AsAvWalSv3xo8ET1OmW2t0szmK1IFQMvAO+NX7LeerHwccz
Q1AI1Ew5fOEec/7/radDVbHrRrOxqIIQjPJhOBtNDrAdo1NVHCO+djiWDI8Q4tSj
7ahVop5uOWfakOgH8xnx5JvvQeGyQU0ouYra7WzP2T2/EJEEWw+1PLQE6ya7Gt3Y
sepbsZDi14vYlLaUvROpdezd/aEixDc/nCXd7g4wVEqfkctrISZtw6wzFmgNx85l
2VPkCs/5t4BknkYWX0fMqb6ugd4uhm9lz1XiXdND4N9Mojig6uUAjpyqQc8fHpIn
QCan1Dv0qAqTRnFQb1+H2RLT6ilWEHiVyTovxmTRvd8qghRaZiBwoVQBFu4ng4nN
/mBNFNAEztAeRAVKo9jPLAHxKhdp2ORZiR7to/SLqZWc6pmQYOKm7AI6uNQjhOMS
mxxOJRPyE80X4JLjKAsChcR4+Y5xzvm0WPDmcOVYV2QgF91OsiERTWJlc/DKar79
fSxEp18EyYQ/VE7JIdMhF4AXSiXYvkETEgCizCb0r/K+Gvck+/UzvgUauUpEPIxd
24zRhWVbCBYmdTC4o9so356aFWrUclcav25qESmKRviEhswos2KbiTtRiigYBkqx
x3gelD9X7gYylS/hOOx08H9kwjEsoI6pgNRkoh54DbQP/2bfQ+U9sJQGI+iRoaEZ
D93Ranrjf9VSS0+UD2H1dbYOYj7NMIg1iEE5e0bP41HBSGRib5a0KoTYvyq1ebmC
IvzvGXgc0e0ox+9yVoefw4tffuqWIkQ73lsFJd6qu2VPqgtuoYUluf+ruXkyNZyo
70MrErMTTz0AgF6bVpSL6A91AvQn99NEKsuVLnKKZfA2mM6eVS9ZIpLQJ+Nz0tSV
IdNdbFJ8OwcgCd0aiMTf9SHTEJQdE2GE08nJGPjEcTfoRWKxnEvh2fw9hij4YigA
dIuDlXRKinYkX/qoONdmbVbj/x8Wu5ZuW1LVkPaO1d9Mu6LYjMIpF8yNfkMO1hax
4E4mkgarDWjFcmcTnxAqzu7rliYcuJyVbTTuaedCojtGT0BTuVCAR4+wZXDbLA5A
qYFZqd0EAVwDlHyAhbSDTLp0X7nbPa33EumafO4cuLky2N5ZAudHq/l3cBf+58Ll
bBLX0L18tbDWJGjsfAzvJbc8xDDt7o5G3GeTK1Vx/zeln9cBVBR5eQaWtR9JMWMy
5FWxh/iZJgUaKduIwxahAMjeSC/QhCcXnItLLeAZ+mS4jZucQIUFrKNv1z/L2nzw
hTpWHO2x1bH1UQJCb6m4MSb9yWuq3OqYr3lGgtFT7aNB60di3DV0CCXnOHBGjdlj
DMFBW0HFDdK4528sYdvxAFzFRC3bIb9pACHqVyW24kDygf0RiLhlTZe1nepk7Qj4
Nt9jrWZTOWVhHvvL274BdrJ9K6hV2D6KMtpXtlyC11NFCliWf8X3uhbnC2IpvYSH
/8nJOJqIJ8eZpmsPcTqr/3lk9qAhZ8+EaeEoHGZy8hKu0iSOLKhXyizEI4qUmyah
/n1k+9cowJTtfoXJXuXMYxxxug38iL+Fs61ZLmc92hQjZ3iT/Ct6FVgCUWbFC2LN
Qiw5jbczM/btdP+E8Berd1rxHzXJWVUKXTBbNfIf639n2AVp9YFpg3kaDaIvpnJ3
Uc9yzWUOCLY34oLeoNP+GBQodRCGLi0r225jR0YUaF+7ITwL9SQf0ieg1I57LrBh
mvKOquVrZEE6ru/18BklKQdJgCltGedC2ce6s+900FxY0n/S9OqziIZDoEa56rJn
YgbEgSptnxv46Dn4+3PVljTyn+TYbQZi1FCCsp4Dk5HgP5MBly2UM0yHLr9/0QCb
g5ytAbAfuMGE1lLfnmcC5B8mfYZcfdr1U/YJOpoD5eCLh+Xm8B3U7jViKDZUL2s5
S3BOkNXrtQeLPsm5l7g1hpzsLwoNJtSUYqzrjtDPBSdcfPEQzkIEiUD4EyaNPuXM
TPAloTjdETfSw3KxZsaaaCqWIT6kW18em6urfVkg0PSz4yU3Y4K5xXdj4sqHD9Gw
Ha/6E6jP50jbF5UPODV4ICrcWNRo6lk/3Q9JTVqBQ2pAyPmVqVmR8aTJFHNnLyoF
D5ojnAlARSXzRn1UhxH8vtsuGzhfzi58GjwkybSQrO7o+/zfpagLessXjviegQ9u
jYs5f8ImHxEvfdrP1HjrqNcLbMssDnVf1NVR2BfRKpKLIT3pVHEk3smXrVk3CHSw
ZqULYeycpWhqdg3dInZFF3VlhshpFd+eG1RMPOsafqXjT0z8MBpG3eqBm2Jj2FFU
M+aakgnT+HYcuDy9KKxvtMiXRiRaSJLeoXLeFu8OKM4Vg0fjTKySgLsa7Iadoh/S
PJ/6Z8al5JtYIA37vmul696IXCmW+Fb3eCVmBFOfExL0LOLTvjfVhoZXcZ6qeEvA
eJssqbrHcLnSW5uDQf66a14XXmBIyesYBaEilrkR3RkcfCnqxRsfL9jrUEghIXwE
V/0noOaHiE8OSB+TZfZVogaUJBmG7PU6uT7GKHL3qgz3sXlQZeeUqDB1mheRm/HK
3EcXIN9mLhVNUpUrckP0r2w2BtcuLTeFVJNnGWXw0zpJSHesms4hLJYpbMa3CBni
2vFo4Wxk5O1jIMG8prwuMIOHAnIestAieLm8fFVkUGUGLcsiZK7voL34ZzEDQFCE
kHIWIxoUJiPWrLRZgg8U9rdIBJWA9cYkZ1rz7EeSVvRCR01tH5E64PsFwIDc4x2p
IpQXazT+in9BRr6DliFBFF+9Udg9mw+UCxB3211ln0a9ro2sZQw4toeFvwg8kwYe
LVTXSQXp/+iR5s8bkdaHI9zfd5whzy9mJnfkHyPaHx60EEA7tz5ZdUcV1nDSmV7S
1YfV6DZUfipFLtl/DCmPqY5xctno1KR0Es99GJGNNNgbO25EShglWrZc0fkQbEt4
ZyNNEtWQ507s+yyH9sIV6x8Zh1yAo8kZGb5WGUN4pP+zXwhNfJ348UOBiywRgwZZ
0q61Z/DZFx+a6QBSAaeftO1yi3sT8gzmKxioNTPiEO7doLrpaNjJUIjiCi++J6Kg
7shhHhq5lXlSUpTD6N6jkeSM1nZXcLkw50L+vR0FE6UhLBZpBa2I3kc8cEyWUzZi
08b1baf5AnuzVSdcv+kjBY7Chmh+kvtWAyUQ4slK+hLamAbXEw3paDkZFprU4otE
viWeN32Rx++wNpUBDhyOyzaw7tKpAP0Z5HhphA2m7VkmW1XhGYDseW5sv39NZObt
9zCPd+0y0IdQ4ggWe4SA27niik+qZCZZgxgUWJhCDqy8622BZKx+jG8s0Cozc0o2
JqwEE328HOlLsYJIm5FP3ArJ91ZyYh1nKhsLG5vsTc3qs8VtP0BY92t6S4ruV18X
DzM3yU8h6kNfHB2m6fA8r0DSNMWxxs4LF8OqJGmTFOCB9AbXWWvs8gyeZDkDA4G4
+HB0bqLCrdLeRXVa6n/syk1/L1sdGI4KbsW5SbnjvyFehZv7TxcDZpO/dvJaiBf1
+kBUSBIeb603A3r4yCXrpexPBT0hbaiYHTBHj04eFHKUaj39NaFprnVKVo8EU7XK
9hXiM0GMXsqthQ1JCDBSwqWzVW9LK1HSKNbJPm6+k+lJXLLGBPsG6SMi+pXYc5hS
zlG37L/RNGq+MShsRn9vrhW3B38dB84RtKV2yNuJ9loOzhhtI/D06I/4mHig0za+
n3BSXhcOfoIFDCXU5zXuUWwP5LE0mmNUyMEYA04C92MCYpZwkFYPbePoIaxOCfCf
3uHVGKDxkffCCtlCH5mvYfLiO8glfvvD0VcAZ+3eNzF2RiS9gRYswjfBu4XcGiit
781TbTc9Jv/M4JEuSTLdnRI4gk1BVRS9WtaQ9wBd13sjY8cUVwqfrNi0/5LnUY1K
b96FYgNgY0CTKi1DFAcQNu+Ra5JKROF8HXBDvbOnSxYDGi0mChjoUgYWihHDuP5s
+jjHV+beSJVpUEA+2ryraJIsUIEs1Hk7XsA6zy9fUg5wXTSUr1cahg9dTslFudpR
Dq4oD3u96Xf8FY12aylOtJn6DmwZ0sM6JmeP23QOMsHnPUul04AiINPIuxL4fKP9
fpgt5oCQBskRjZ8CNDAM6MOHCV40E3xPcTEpgf0QXCasNakbMr09qohYMShn4NH7
Ihaj2kcsatiYqQtJKKQdlTTn/qt7IkzEcmICfl4n0UgxwytrKudFUdEMVk8zBVFs
5dgdiDRBYA5XqDcfIYLt/31HYIvReCSZddeuc/8oXeFAOi2wUFCyNbs1PGu5mOtt
Df+/vQS8RX8VlFJSiRp+q1Uj2ZcD/d2E8PRcSExZop8BQhQOpx7LkJwOzxPJIZ4H
DnUs8xPy56ZAWOVELcvGdEgzAMhCGZ6/C/NseyGj4rPE1NJUNDmYh5k2sx1ZBvCx
LqvasU0C6v85pqoFR5wUiZCtTZ7jb8MICZM5XEMeiT3iaQnoYu/aJIfP91OnlEqf
qxd7V6+XjhdeI9ySmBfyIfS2ozhNHRq6X/nn6nKNCRALGTdDxNbW6bC4cWpuKEqs
zjNrGM5XvGpLD1nFUjBE/1m6pyAcJMwTbkLoxA9LblN2gWAUMfJJC0rNAIY65t8C
ZDW4/WsDpBiweJ8MPANW5rBs4C/p8Ai3xv7wy9RdKNGQUxtSUPjQTpqoHgI60qwa
d1HNFSsQk1DnRUTYt8lA4mnRB0Wnjx+p9NHLDDEdBPtXLMyAd1hazWrHYI7bnrlI
gmif0bsyhH28CbPgT46aNX6Ya7rO7/vXlnAgLIAFPLbY87LvFOKyqbFkXTv++o5g
4N0J5Aw05vC4tEzi/aqJAFXVJQ8XPl0HYiDxfJxaYb/9nDnL0xddczfdncRKA6Rf
2K8g1s4tjJTscmCjWf4SlFdniGZ2TtbJh/IvxGOOTBDEJDKZ/2iLZ2mj68ymsDTP
35dmj7wXXo7gkgeOeXuMjNORq5PXlovY8xXEQQ2f8stbb0B5yXUzkSqWMZc4jFDk
MRkw0vUE2i6HIGUc1v/Hy2pSIYtvjPfVSNz33x0QICrbi0wQspuxwRHFu5OylaPA
HFCjgQW8Rp6xNhHuQVE3LTTi//Ox9p8f+VQ8mvR+ZZmWqRCWFY1lgbX9mvtDA987
41QIrg/dorceU3U6pb55eU3uGyotY9CvvW20qupVcIGYmb5iOgcBmpHWmEpcKsB3
cI5SquF2sN6G0Sabq/I8fkxMtM9FgEMtV7ABqQtnw+g1EBGAgT9/n/10qrprbQde
0xLk4neVZC59n4TMZl901FpkT83u8mHyfFHgeiTKU3eaqGMABGt7RYClKHhA/5hY
GYb9pWTxUqX6YZEfMUYE9iTLmghwe9GWjHXv6H8PSaPH2vBx2Vl7ZJC90di+dYqm
bM+3sNO5DAD9y+AabgOdnSJkyEORpnDLbsDG3/DgsoatX3Dp8Hzv15c0cZC3NyLn
HJR77ZoY3EHJsy2FX26S8JPJZemFBqui34ZKUjJpdJbqlp1UV2asrj9zZ0dBrXa4
dyR1pYPiOKc3Z5OTKb1dmpPc8ZRhP7ne2sjKvi4PdydLN5UOlfzVKMJ8F4nnzO5Q
ND8tRMxlJAZq0mq0uOZt+/bHG80cpMOD8BSQZ4TntPe9Go6Mafj5slrebPbkrWVf
RvOkRalFhEoK7FM9V11fAXIHDjfRKEJlAyl3KZn7uGtMIxTmBvnNTUUPyeMxeOFe
lkRwcYSjyeXq2AoayV8YazyATgpoNCSkmQVEDBWIn/iPzWyGIMszED6P1Z95DzcK
rLseK6IKkGkaJEvy2/4kiBa7p/1vzJfmSxFy799U+0xFio9WefFt84AmCI0y4rAV
3k83YY/SafX8nU4AYHFDZWp7MeuyBpPhIfceZClbXFgipVAKCicZ+6IFLqDmzrjX
aJKkd8tStRMW6B/QTwKwh7B7TCVo7zsZHTMnkZeiGMCvPnglJ3+BhSmyoF+NDIJ0
jJPn3wwxENNl+6z1Uvoll8zrG5Q5cfs317lQhHfpKGZuPStm9k9H9znaJqj2/Wdg
NttTktrQZ6TEw/qk5dK767C+xAtGa6b2WzjrI8yhTNkSnQAdnNol4ba+90PTG9/1
QB1IjnIax9mEgzMczMsSPTBlOZBo91AiNO5ULuINKCgvrlOoVMyzUMV7lNojKov7
FmmN1NO4up8CBSdkE4mgeZn1UTwuARI5XQK7Up1t2Cf+ZgJ3bC6XrbYgsvPOp9Pv
mjVydS8/3zi8G7cc9yHLKRJS9MrPGZfcdLKBC5ijrH81Y3Qv+QY1Jd/5XQSGJZSk
LvifB+1Wv34oWipJ+swn0tm2gKU8O+yyt5bKQs8Q0aeyUYLcRWXgsvOn2VN9x5fo
VnwdMin0pJs2EttFPsLrA5huJywgTKXNwNdMwna6a90zTlRccDuehpx3Xb0pY0wl
B2LkuyFzA+k2RR4i3SaDl9BW8+yMrgvBL6MlDypr9NEgcB0EcbBiFySY5NiainRW
NQHSvwiHkaCvth5UXg4PJMzB/Qfb9rhxfrq0//cb/WWIs8glvfgCpUtoc1CRT0GG
e8ul6vBZW3rWJ+AWShFt/1KBSVNvhS4/GChxywNR+mDBPEtvj6bwil1aa8KxXktV
i8MoqsA4Ch9XyGoSItgI4iGst1N4sGcxPn4eaNcVWUHlXwemOdOuHx94oK0gNyhP
DeQuurWsOPZL8AlOU8B/xqq09s+dkZkOoQY8EFhcxMPjgU9I96RAE9dNLQDXGIJD
9he95ooZ2Q26IJfASuIAdYuNbQAW/5Nm6Qcuz9FzBZiHDgcRt8j0Zhgt2mvNUagf
Fco5+Yyi2ABjszBBKmxYtMI59nvTbNQd9pg82oVo7XoHsEATyIgyLXl/nqmkUC/P
lcHYTOnS8V8u1/EpPQF4QVutdVgsP7ZYdo6HkC3BM4XfOOhEPFpL91Wvn6L/GD3v
boqz39m/DWWq/kVLnSuunYMcHHOLVq7Y9XtXz0ykY0nz9Vb9ebp0D/e684IPk5Ii
shR5J/xT0NhmyEi9S4SvfYH7Zw5ETHB6AHIQlz4uHlPFDbwS75Z4XqWRWI7phPCl
2uPDyRJuQRROZktcylTzW5+xBC0fw6XZErCJS5pjOs5fVRibwrpxk3haNoEfpmem
XiN2b051HuMkSlK4TNknAWLJPJa7VnNvc5THtfM5hMwCY1+eV5kYeyvsOapifLTN
Z8kRwuodxQSoEW+NfJV4IJsZ31FfVMADh+a5BjC9Y0N4gIiLOCWI+DzwdJEwJqXN
KjNLUgbKz5m8/C7sUVFKl2WA9mc6G6M7/jnrQq4cUBW3n+f4LVKFMBHaPxK0tEyj
UpdBO4xkqBe43eVTnsREwoN4tKaQzgtK7I3jNFwOb14GjRPfgqKf3DCrXB2T2LQT
EdGFoDVzGyLoFalAVmYDUOffgf5iKawsIDtQNAm8llIZ87a9kmDDXi5gmycs1/uR
7J0nXP9FUTVGKMbdYyPJCXP17IFhKVj4PgED7WeAS6//GMCjEvfE0dOa6AHOCud/
oVlOFEoPjZkrRMu+uYbPQ1qog9H/MN2fk9xRR0vyrufCX53m+Pe6K6RP2hhifg8q
HvWH8faF5GSvdzIEh+t7waFjJYFIMt8+eI7WL4TdkgP0xgU6Vs5qbxfimEUTc+8h
kd2s4hC4/88n+H9XwjI1L3rAY9IhFD+ToAxap0LKibFbv3xVhHXS16U4ki+0wQAR
y1KxUaExLSmXEVPtHwqpUNwWcUuhWtv+m9K0mK8VOq/OkUL/h83AKTLhvu6ZVtp2
ZPH10wRS7g3jg50NTsCtJUVhLKL4fxjy6LW825Ou8zOJZQTeo8yHnjiUN+j6AtO/
tqHOlQZb0Cvk5e+H2mEqJevU5Y7hHU+kow5LSuxlByV0mojhamqRISS3Pa3fy8r5
J2cj19rB4uUrXVkW6iPVHNdehKj2haCjh33aCekTfNKAmsjRUIsOH/U+AcnNRFu9
fBkw9YjrJD9MPnoXgmqYmQZl24gSH6sbIjlbceCWXBc6vBibjYEiheKOYbrzmnOQ
Z8Jrz3b7Uwup1+RJkHM/L8Nt9if4n4NdZvRAQpclrdQiGNUvPt3KggIxrNzH5D0Q
m4Y27WCiqekyUqnVxm+V7eYfb9+HzhpourB0FK0eU2PKBqluLQg0r2TqNUcJ2b+C
Ik2qUYffwGfhRz5mnWjRPaLPOtTxWvu9Wcau3zdzYbm1tM2fABf4BWo5MwRb3oGJ
8eVAOQnX8XuBEjx5a/puuPyrxfKytg7u3yNoLAUba5nEoP/VVYnGSIwMtHfSga0L
QUiWtIhyhcCPs+5UB/3AbRELtFUPfhsOqxpwhLmJqfBoVue/ZaqHtLiwXebwuGdd
GddTyqPLVaMCKJBmhCXnuLuDKLy6WnvVvddhEzJMPtq2KX2iPhlBxv3zIDIhQeDN
X6ZbKgNM5tIZPPlS71pHl4A1VEdndnahDSQjo4rJ7XEt6nRiq6ydU2kYClMelygA
kRLjTwsGQpcToz9u4XHHDSWz5Ob+p9xFS7vYEP2bpQFyRbqT7qfCRNqufO2OWOFd
c5hE7HUwEhdUZdGVKR4gZX6/JrayFC1tjmmUmtQka7LpN2jespb+q3Xr0niB4/PQ
mEYzEBrbWD+V9sbC0PQ6zwP0SlhwfopVFVSS0CqH2/LI5Rz6v+Wt8dNShdZFZgxf
wRzz47wJvfkRAdq9ilX3Eg7xI53CRz9vGXDD4T2dKg2kIoyZn0MIMDVIzjvHUAEy
IOomSt+/RbXZA7XdyvCyEATe9YYOpb5S55h5p/9qbaW2/HdXLKX4FZf65181ZA+E
r3jaeK29fKO+ZtMiA/oacUGg2CMg76GOmUlsUl+3+m5STyT+OQTXFJYhsnfQ6Xtv
4LYhL85LIpAzrQ1N8bklC2MpCWf1bzMy1NYuUBfMVf9lcPzphhKJe2345GQpJL7Z
y/MGE5BK/rc1HKMbHNagB585h91jHmTPQb82yBt9+9auTfZtp7iPltNb+iNcesem
hOs8WWFX4H85TqDd/Sc0V+3+OQosLr4szhXmUiVCsClPNGW9It+9GHdnk13foUUE
LnznWmfXk5ZVY9OP8ZfYn6RjCxLGf/xgAibLPZfURKHhSHFj3IPbcYF2hGnFdlZg
e5UG49m66NdLRnbwHnf14AtXCpSfxNqWafUY+u8vq2ZcMnvPK7vZEYamSjGrRB2w
TnifoYroED05eBPoiJOEYmPhODmR2lK9gDHTZt7705Km8/0jXGiZRikF4Mrdof44
d5YA0dqQlKrQCq28bfpTUIi93oPExFIUzVVHISl9yTPq4cGKWViBfx+ohpcjU9ve
U89fAl9UarBuf4LxZ1KcIlgAcqWU7nmTq/KlTYm0hT2wtHD396IeglSewBrXasgy
GNoPu/LCSRnpiuqihdYlKxjGDGqOTUfxPMM2P+qz3XPBYNUNDK4CSM8Ay0iH2bGU
Vb6SBqtP+RDkwWRdo3fUYDVpKOpHO+fAR8n3X5KiDt31nL0/qwbKUbSZNv5eHbPQ
ZiS7DtXd9mj+97YP3d3qfJ1w5P1d5mB5/cJpPJ918aF6oYRHc03mRMLGnFFs/VLs
KQWUgLx0w0e7RKh+vqRE2hucwBTcLMzeRt46JwXYYQPG4/iLpDbn+0Jla89opAcW
+lS5HSfH8HbcrfGJQQ7+DDUW0+3PaiiD541GXR7XUXK7iffwu9rgujWJ0NDk2GV8
YA1ldfWR+1UPugOvOnn4vZHCcvA97Q/n17+Ijy3twN2B7OrTWJfJMeOVRRXBUBBs
wZmUScUxiA0jdjMV7aUdXKTfrgUZ8ONYrFtFuSL1KD0FqWPwZUBxDF6i/luFLncN
EfHUJ2N0Nou4qsgtTYR5WKpMZP15fTJcnaz5Mi3WH7TuhZcStMp3zVLY3/cLa9hk
kVKojCQd2IdECZJPFdDSfgQ2JW8VWDFIuyoJgu22Ka2FIqU6EcABdhu1KfDVEYMe
vuWC/xzvAjXc5sOXgQdW+HvVmoQYiMpCmnGuZ/C5178+5Y1l9na5JhySd/D0dtqJ
m5/9KnQk7jFKcsHxL9igKDuW3Nt41L8KGrsGaxCCv/A5KRVlYejdIOo6i0z9WIyx
7k5q8obrK5yxSiuIYYbJcDtNtr+XMSKhbaM51PQExUzx+dx4nSrnt6a3DxZtAjWU
t2vdsf5EPH8yBVNwSCAmfRENqFUUeiYs1nFZVLhuaYRvTaAF8BTsohRadKcAD8d1
TKRGtig04U8mkekEias0UWKF6GKWy97rV9T+c9gM5Qy9NHn3p+ZwzvdkA60zBM7a
DvD3FSl7PRBZ7g4ne6hWdpyRFOnqrmXVe5YfmtpH48LChvV+1VXJyBkkrsF3smAb
n/36j1FQBo9K8gQ1g50Bl5TywqAbyWU7Vd38FaRjEdCme+e989F5i3uNsV3cDFFH
Y64+9P8rYMQ6PfMYPO0i3cefz/05gaZcVTMEUvDWOkJ/J8e9OQmNyv8XJSaDXP+k
58yWSaQk3GTXR9IHYHpsOU30mOWzUbaJ+xBwruuIGUWHjnCGLZcaR7F8QZB62QJO
69/OypM265ltwE1bttA8rYrN8OmEoY2Cls8kJYw6GereMqL9tO2xJJAmVuGe96Xx
u8Cd6JzoANzakUuzRVOyHFoBbtENx48TQP2gSkLRnLDnhhpkKZpu6KbedAxhtw4e
M5rkElqC1mWc7SeHzwHkHvSnCFC9x/s33fABGcLRMGGZvtTPEZimqox1qClqavJO
EMNEo5KMm9zbMsLlZjiDQsd7S6LKK86d9IqKfI+mDCyJ3+nJxD1hgv3IPGYBafQ8
2dePOQwmSS8k1Sty4at5sIjMc1q/Dqq97H8lLnHQmVwU7stsWI3p04WOr2YnHNP/
je8zjRbVdyAoL87K8zYKv7QF01FFs8AytQpvNaFTvFroYn1uALvKSwPJvlMlY1zI
I6iLxhivqn3Kf8F+NaiISA5/luDFFaGLFAr5NzvK2UfUvlG21qWRRShQSVnfj2XO
JB66kDdthhc6FK9R81pvPmktNJsDVMdBnnJUdUqHz3gzO5BF8qRS6IbLIS0QgJAg
zR9pcNzs0Uc7V76tweqE/eu4205xMN+i2BBARrlvNYh3CKvCYxSID4jx88miw3bb
9F2CN00/3CAoh9YO8QL5s5gAXecjRjED0OGaxUYei2OExCD73D2f3VseHY9vEKun
gFvEBEjjO0hZLXKad9gZrVq5dfVnDDAVDY3GL71OrRCGRRlv/udSCLUoQxE0qh2i
IbAGKP52IlE4uLI2RiNcyyoBQYYvO90ghPfJH/zWFvk8H8UWOgr2x15k1KHWopaw
AeDs6MoZxjKewriB+GbsHCBhMC3udosv1JYRIQcplpOcvTq/MWk4vQmr/IUxi14l
8oPC/FXCWYmAxmSqsRFHL6norXM8aef8934LkJsyPatXJ/7BDqs90AvUCJ9Lkord
cf4d55Aeady87sjkrQ1ThUapKgsuhSgB/MtYjs8+OMUe6wKXp0a+k23bEgGfnIVH
TmXcPu6DRHB0+mBkkpdlrrqXeMNlgGQ+j/D3Hs6PZo8LplE7q1nAP1+O1nxECDbH
ubp6rfiNpbzB+n5Fn7gXe6OVbKzZABawtJRN3RZ7gWPc88FGUMwXDyYae3DL+jDl
BCRZRnLbtCJBw8j5W9Pf+Gf32NmNZkSUEhyIizhGbW2oR9NkxpWqXVzziM6s2+7N
q/ldFMnC/2iycjbG/pRcKyRqaJbpfpZGIeGsADMmiOLFADKv3w/lmMNu+XT2RV0w
7dIk5LgMsWpdJ35oQkFLWUSoLFvLnt/UrLEplDvi33gySYG79cq653jRCqASq1fe
De4iqoo//ggn9IgN5HtdMGlpdR8C3l7zvcLDVqzxTWbK7m0HSlHGcwWpNjbNw2r4
q80sU3VSPtyuVkM/O+ct6/RpM5G28rj4zeP9EP09+VqlKaNf/n9Yshl7wNrobLvG
tr7U81f31GuGrCzhHstaswueobRFNRpjfGqJhS3uTXo0gNjlr/Wh5FV0BPfWdpE+
0X+uEInLWMFdiy3uHI7gEaRmGNHfRPQb+m35O8S0NhXfUHy+8Ctn8oCt+w4FZude
POfqEuLqE5sSWKfzEYLUzd6NLEUOXQfhaVy1T9T8O8/z4ZN7qHgOwAkUg0LrrMpl
HuMEEFfVfTuEf5hKNRYVofjHq4B2CgMqiTWPVZMQ4oSLCXfMJ4h+V58rQu5JYZIT
a2oXR8Bzv9natanawynT/1B6PLDbkerz+i/GhJrpiNcLwS5w6TY0bdJKuFdGaWWu
1Ew7cjk/UKzT5dxAp/pGXs8gGuUPfHg7sZP5fJA3HiWkIRWlG7pIMvi03gb0A+2Z
sMBS2YYvUOtzMu5xB4OFYypT2BFQWWYZo9D2wXnEWvthweI0JQ80YOuC3DBgjVRA
5jLAUs59S6fmRZmTnMaYKqmcxRKJYU6GfGJ9kO5sKla6vMWZrnL5uEM2jrOuDeu9
gzzrqHOD0+RyFR70ufx4wLpdXxEvWNm3X+SRh3njZY6lQff2arKwcF3Qn40zPqi6
WlpG/k7p5Z9gi3cTaoGpm6d97XzWO1IozkWzUp/f1rdERbgei+lMoDQmLfCvpEaT
/zGS/0AJWcTAwyD5RTLD3QLud3jDO16RNfD8F6D4Umo9xR7OcAm2YANlPaouyxtN
wVNQpEEeKqr9JWGNC2X8SZYBtppS5b43ZZ1yfi4cYFezKuf6vNeT1EUfYyeaz87x
XNC7Hbllcef92sMKm9tIrDnLIGhKgRiwBUVMT1kcQ2AUraU+/AH54x5/0Nd5CvmJ
xuIzSse6T5XniT81ssnTjiRvIuzDfu93BfaaKYXat4p615gD56KbSmRBfLPH1RR8
Qk/Z6vHFyQneBBTuDpFFoa/QkySkh9K8TqtWZfm0RPKcbk9ZqTQi9a/6JFtlP0ue
FgDnl0+1NgNYNxrmgEs+RwHAKQVpBN04gQnFbjr+aXvI1iLVUHwDU2ucCY4o+quK
R7llVkJ4O9/+8J2eVbThSTamfh7cSnTm8SXLaPwSqC6V8fJmidg35NPFDENU5WmI
0PsdErPgkgrXtJ1QHeLlC3LzD1+NTFNgIHxSlhN8AW/ZQrg5h4jFVHjwEc68Pa7K
ca0Q6w9F3VhK6lXOkL8gjZdXuhYCHSoH9NR1eUSOsnF0QnXrHEUvlEplUDnmq/4S
kU7oAVrKlkz5NHSNxVIK1kZDVhwA8+et1HgTQweHA2/IR9fNro+MwetMvv4/rv2D
J2izXN3ykI4mkJPtjUYGYaAK9MwC5Q0FXdxHHgm+YcNefnd3JW/Ps26JqTlYqg50
EzttdeMncYVS8C9cV28TghezPT/3EjS+x07gnrgTB4GJVJ5905BjeYhmmPwml4CD
kxJqjw7f8wyXzMBjak+h7Xj/eNETALo/JXJ0JDsueNdXth+GM0r5wvZj+eiC0+PW
s1m77f1+XK8HA0cgrUPIf5MuGq3hCpzYR8cmYTWF7+mD5Mih+Y5BArfWM3hVQTim
VNxJAQoyG8i96kXu0QOJfv9eakrtymCL1OOnjzR30OKM+zrErY+a/xqoduyYtAFF
2qoWOlY6h7yJXVx3iICz/iZhZM8bu3kMkyfsIGXO+ewA4ZXJR/nObB+5f0ywZYX5
HGW/N7JLh6VL7VziteQIvKsDGlKcPfocWtTHPttdhQvtKHGMOcejHj7Zc69NdDNp
ZucarjDn5AtZh+Li0t2aRt9u4a+xfGlpqUvdjzrZuSH8lYEJ32eXARs//10n9ac+
Gl1YS3JtvEfjLTVG42/kqeIhNNf4NhrjIVdwVy3Qli5lgpcWJx/Y5KFUU7jGHi12
dg9Hn9h2NJumj+rumC2+dvZh+RYLd4JLgJQDJSIIZYOBJxnHbTsinJTniXcYhV05
3bh7zeikgeBUvStxMhEyxmTQv/HfpLngJuTwgWE9lDwDRf4aPrkWCQbqfFt3Ce1k
koPyF7pf69P5whkemZEA2t/9eCwclbHp98xuX9NVj7Gr02r2rSs55gE6HXV4ZRn/
wAc0JhLmpzBmE5xcun4n1ty2ozCCA0pffVxYCkS1G/EHpjs92uhU8OQ4X60Wkxwc
o6wMph1PIQhLI8I1qJaiRw7WenunghgV1nC/LxkEVopgWI/NXT5t/308bo3eN+K2
PNpri1LaeLEnvQeW+s9Ih9682mPHr/QNv87m98S4OoUU2zORK+C53kJDYYCBURFh
0NQZ9C+H79TN05pCl7/coccHwqqBAIzAj+1xgjp8/93BE0Kez5r+tliynSQxvr6L
1C9dxUpwIzg2iPMzG2ii/cwc1wFGfoFSB4WRD+R1+Uz687YOIZYm/DIO5lZ8Ytag
9pDClyRj54aSEx2pgrCDb9eejcYEaFGiyRu+NhJrd6PMS1QirKcnsqi9d9VxOpqj
Aat3l98rQd9hAz+MXRVrAezepC6PMISV+n6GqZx6GvaGxsmBs+oRYlIIGEi0JqzF
tG4k1SR168q6SNjvbS51e3JxPP8ai3echs3lzXi78k2bhwfV4/t+whXi5VDE6pWO
cc0A0NjppL63/O6qlm7/iNXWrG/RyYGGKwBftKHR0ZturAFmoIixjRQJ1jI2WNqi
Oo6+vCx0TeUWIXj1OXiws8tjrsVxxKgVv/4qU4T1Af+NhnChuyzWeI3z2vZAUhwE
mH8sbxnAIDO+P/nZpMGg/N2hAwq2ho3Wil11OvraqNBcHd2svn34Xf9iHES4KZz/
mg6ZTVlap80flwcC60vbg5sIk3km/87lC8oM1YsGdAxkKJwTixqMkv1NNFBvgOnQ
jU8GDModZJPyy5aBGNkN9vB8OpbBpn2iKbpXXy4cHJozrzuzMJXvk3ffHfVFE228
PNCfmSWF+2P1V8voxJaw6zCL92j2qrPIkkAdIUr5N6Jo8u+rzJKF+4Y51IjV3N4l
0C3c/5qCdwkvzDKYUfTR9WPLDtePFuBeEd8TrLuE6NzqHPznbGLKWVx39DgkcHPu
2UGbHbHd2Q6aW4IcRfEUwERPF7XO5VBvS1ykMY7vyvsgiP3ps1NrW+v4Ve2hf4US
2qVSsGA2hOk0uklx180LYenp+Cf2kJCGiBgiLrOCQOJMtb7oFW/p9rsa/een3qDd
7AgN7CTOV7qMaiigjfMMx6Ki0RxEDl6aVcqlvuAXtnIjBnfTpgQGazZ5pMttLM1U
Gm0JJ+3dBBGlVhanhEL/DVo+Dh8xg2LT2naASuJfm6C+cwp+oF1PnUnm6KQkGOtN
9QxUGTBQI9ZKPl/g7ret5m2lkjPfhFN/7eYOXM4Vn7GBpkCPPGK/wuPB+yX/Ypfh
iU6aMQSnukj8JfuY/eL9K55i6GX5CThDOMarKMa1gqjBKpnrUekfBBrYjeoPXfwG
8slYI3biZQGUx6xQRrp0hFWFB3LdhLqOFgH3PkSbuVBupBisNKBMnSA40IkrgaN9
q9rmw/Zqng4v3b6oiT1HTrBefDjq/dZk9t6OIYHKtnKTnOLZJFp86pS0/DOyc6nB
nfzUdI/hlBWEJGjcrP+eCwyTnZiQaGSge1WlePmWdEracc63movqwG5d9ivmShSj
QdbseAege3E7INKVSv8hp6cG90ey774p3wdupxIT7fydL7+dHwCzzpNyGOV3D+pp
xbUTa/e4zsb6dvX9cFc137CnZdTDWKloyIppZIvBtT37Wb7zEXHclV2vjfuAonYP
w3nR13E8CGJ+kshE2jo976sCTp7dHlVbx/lk7lVn4m/XqDXiymDn6RYVIP90VfPq
ohE/tDt8l7L5ZPbDfeRn3bls6zUInEdd8Swtwbp7H/8QuoJfgp8ndihFbAsPIVHT
o4lMdLaqNkNvxYrBQf/zd4jtxwCB/WiO3T8RlqfXxL/ypZeg9kKMbBz3lnMxwus9
VN8zfy7+i/MTQsZBrgeAjCBmNgdpaKKzeUy8ihVj8lqlzgVva81TYps+TOHCCkEr
vRwtRSCylqiSLuFUHYe9MbvYzrEWn2pbYnn7/gSYKSjKio/eHm5oT3vellgoXDdO
NbuADDVdbyClbH7nDerou2ogIY5QIzIt/+6//DKewiO+dIfBQSHYe2ti+lAXdkWp
nOu0Lt8EHjDsaJNzxc/jJ7l/MVG1j5G5fH2VT5phYZ/6bdcmtT32sb6/TS3aUc1h
3ow/XVZgZ4n9S1OWiWtajheHoc2MQQzqGPGljNq73Ex+tKo/o5hSF1tjpzcojxtT
3RyiHrweuriCkUDrpZ2TXztQClX2eqc1tLZRB0nCWsKuxxHz79gRsmShEskshMPV
yiYXMGofZ+lXo98j2TRLyPLXA6diBpl/9Sn/3zshwzJNb3xmPZYdeYecjH9wA0tA
E6xT/VmJmMmyJ+s0khfEQ6f3vTAb8ADtNdnj5kvgoTxvwvfulpsOpM9hcbh4ljbC
EuC1xuCrKCBAxzq0j0wz5HYlGfT0fQiOx1TdVBKoHhhkcjYCsJqNTh4i9QIX5T0X
16RbmEcv+H2c45LPeQOXkZQeKHM86mJPztRma/xVHDyP254QOyiKfBTYsO6J1l1t
zVcaNpx+SlX7BrcS3B9aZrXiA2c7v4yYyNbp9XYpABY7aBYDsYc4+FU/kFY06K4O
bAsl9urIZWg+4AsDTO4/tCJvB96/P211Gsrw3J/qCCACoqvDrFValI4AtIpDnLSr
4/vpwX81VIoBqbbJAOjwmMK4giIIaUPz7CP8Q1g7IV+GJW5ghKnsimMkjBHAPfI9
he97A3tu01XbTtzAaSFWmDK+Ist1VbSRn9XbrqwLx/Dkoo7Hho2nuNdy1y4YaKDB
Xjp395MK493O8xPyQ6wH2HWJn6oD+b4Uq/PvVqw+DDm790z4TW7G2yoegU/PZYOQ
iGmRwIpYCKrB0BaS9MZFx+FJ1pkVk7OF+iReEnIgsUZ5O8veTsfh0o8VISXPajYh
BDjrWPfsOwR+AXpi4uGMD0ZZLTAtic25K6b2//nwFBM43/pzXMvcCgNzoQRusz5/
SDGOYGrksbtXMl08hFmWoF9V5aw936WPEDzoFDaA/2oBCYA20sdLgyI7NKPH74oZ
Q0VqG3pNM3CBkanOb4YkKIUECBAlyHkFx9YHNKubvlSkqEiBRt6zrX2xp7iHlksn
/ZxESYdxUDcMHAbCXRtDO2I5cAUWvedLaTcJFHvnbJMWsMUq1jfMcrStjeIkt+V4
N/YWIjGnDev8XEnUhQf/Cq0r7zGuq3pIvskyBEXu0fW/FF6dukqC8hPwtLzFVhXz
Mui4on7+2evcdp+S6Y66HXz2WQNqXaOei4QwZudXjhTtoO+lKj7onTRjuIO+YjQL
eX0xQA3+XtbnCma97qJ13uK7M6z5Loop1tLIqq1ehDvqwNcJQBJD+Ftwj9pFtTX1
/BTLMqTbVUUCc/AzKbYEXOEMmzQreU3Tbk/KJCsqilVsZKFZqQYyGQBhfs7iQfFH
PeT1NivJ27HJZ6d55q/Z9zNDnXSfWD9bekbBjHCnTwlUf1pt5KjmW/yhFNCd1Tiw
QYoXRT4pGNmm7xcl74EE9bfvQSjy4OFtRyYRW+eEBaym+zNsq4us8ZHyS5Q0a87/
uOzdjTApO/bd7alNnuikbmvRJ26NycldLNOUvrohkU+VxD0Q3Cny7JJWlmoItVoq
TGXonUIxGUyUVPsepowpV2SkZRgS96Yn3egGzYKa1RMadG4ADQmKcrzgqUsginTi
afOZzxszzhNfES1vOleED5EVBCFt8SclRXLErMM3VmLJP2BN3y03VVSRrIH/hH1J
c3916/ElFbHhaKQyQkMt6HllVescWH9rP3PH9U9aHxT19e+5vWCvyIVKRjhKOWZD
a6Ar213Uy4HBDracd98Xwzcqh8E7APldeDj3XmQckgCIQrjTWO3ta8/YNYMOvuy6
1xmTCmnOKYFRQ1BVNW/KWByQDbbzPTPjFi2W916RhSSIpBW7Q1La6O77I0YSVA5F
8BNDIhQL1+qvGEkLDNictawMkP8OW0/sOmkTjYLqgiQQ13rPH9dxHh7V6axskLn2
idc0Evqr22E0JfJ+PWM6zVnnVh20MrVZHtwHCvy6VuTAD0rsHRA3NycZT6vMA/hS
MDQtdbJlsnL4RghD9tmPpEeIA683C0eKytNfAgHBhCN8A+YkjY45JBEfD06fTkBQ
S6JwuaD8ZTz5dP4Jd/W5XuaFqxcWwcwkJI84rJHJGXTkDlwED69fv2mYnY+tMiK9
jEytWx6qHQASpx4hMBVt6LuZDDiwaVwk//NzYIZe5CdVHG0KFqTzwDKWjMEDPTQt
vBwvKbbzyCIo/719qxz6qnu57JKAYuGIdV3hT0weXqE6ky+23Jr7uq38rv+essn8
0GKeNMHyBVfY3y/USkBy8ViZp31ChBen9rPzyLwnAOyqevJtJ2TBkj0P1p1hQzFS
9YcZePvxzPE6VULdZIT2KQBRumQxEJ1Lpmlv8zns/APTFYUMg0IhAq8WrQwAJP+S
pBtk+CixheON2QTGSbygtLFGSTFc+qfKp6/8pQK5yiJeEBd47d3QCssHjcWbvSgV
3wB5OBW8kPqrFKeQJVkukritkZ44RFHeIcIqN0GG+habuzyNmYlREGFq4FpX9Ui1
olZ4bK46XyxMzDCVG8BN+EiMBnR8CnlwdZClrvHoeiOoVgWX4zedXNZCQCO5VGDW
zKal2gtTkv0QuudMtK5I3L5GmNjl1BP41sn9WX2U3QzBP0q3gm2ElVtSL1sF6qC4
tLLrbCJI7L+DSsQ7dIJhTmrRFI4xh4aPZotyk403kf34CPnGGqTfQRmykH/80XWT
8tcxZjftHzV+nyfUDSDdxLWGWaaxJky7Qbg0BxcPiwGEzOMVzM2O5teihoN+L52j
zeyA5MIB4Ua7+zxHNHNyzqUDLTHNUdTNBuY+RpFQaNasl6ttmqKembgVdVyi6AIk
uVgxe34zdZRRlKhme8++zpIWAZRAeik64Rag69JBkFF/NBhqLUHXD7evD/JDT1Ir
tGqHua79qf9Ro95t+bXUzW6e+cJ/ZJ1rS9Pr+Md2Tr4zssCH5GluBnpSbNcjVFk3
cqlF8DxhK7kOrb9k8+VsDiQ9G8nMRw2cm2vx0vZkxEIS3idM201fS3pPYse+sto8
nvyMkNbRPjcykcW6gwM2bMKFRWacDpykZ5kWN6WS0f7ZUdNJeXu/hPL32Jl4o5Wc
FGw8pDDZiIUTFuWBY+L36aM2OmDqvNrjb4rN8idu5ymibu0uk3/IskjJsK2zwe54
26CoUOiVfdrrXlZJudn7zdpjeEhuN6/FpFud2y24oetsfx3792Y6NqeNlUy5wzlh
BQx9bZIGRh4sTBpnmkqMFaAj7+F35vMCB712qHLlc9sals4JPWolgornWJ0J8LH+
4q8FLYkGZN6L4jb9XyqULNZcqy30E0s3qa+xuZT7eMdZ1Ot05UYJg944AzoankSe
QIR9xne0fohMqvq25tpf1tUfJOmIE4lRcSmN69nKFEPNI/RrLBlNC5r70T7DBc1y
0KZIA0TrGGFSZIZBMhWSDo4ow7i42PN/mQ8WMM+LJTvJtO78jcw8QSdznEEAdvhU
/iMSig/n8W/rij4WvRGNAzNfDUhKzd+tGTUWatRgBhGd6Y9/ZCsKJ2QOB90/HCY2
NI7KU/+ZOMY/VmZjh4z+cdU8JX1XGngFbgoi7C7WqavJ6KB4KP2/71/+YEP1D/qR
2f0CXVz78s0k3VCk8ZZKRf9Hz/8T9OlZwXn1s5GaLnhA3UiwJ+Am+05+jHu4cbRP
XW7pPB6qixChci9mzZ1gso+YN6cRG9aZ3B85jnw8tFz5CUKQ53mqAkZjpZwVZNn+
6qSWQNtnCCPHvc/Z3d6IRETQHOcqqnfaCNzOGJdr06I9nOLqjxfn5aVX5RwuCVw1
KYvOcrIzZUdILHUhF4e4j/I6kVqVJLs3nHt+NRk0VbCJXsuTqqfD/fISViEcc2fx
8uRPPOGqg0Z5r64l92JTcYb/cheyi8ECZezGbJ3na1caMxE6Kl/IHYd83AB1HdN3
cJFnxK5YB/ga5V0tkGlGtKDbq4YG8yZ9fZq3xmYYkSkRdsBK/+lJYkJGhgt8wdql
H/4r/+Obqiuw5326gnGqGKO6o6ELi+vxqy6UM3MBAMq/3hq9YPjO89vmbVCGmDEI
0Nc7qmagG6n/9VfFc9wXNybWTBspnlJ5S70RcRLtH9JNQ343ZELTBrN3PVTdDbOe
DUZfL6l01jrOs1Dx1BupRsa2tMUt5OI8BKXGTZnJeWtqR9GH7YOKDqDOuFtB3qb9
Bb1Ooym+QNYvA/OfAAVQ0aJq0UdYbo1MiZCRYXDN7Lakk8h9OSy3tHo1VHOF0dnH
rgehv0yLa7PjjO8/vsxVfnMwivfRF2ATBMBpW0tOMdsOt8CY5lXsNyM/r/q+TGw/
Mx6/X306ueji40//SOprg5cdZhpTLF9s90t/O6WmMMDGGF+wvjP2dqTe2M0UiEdx
gvw/ML9FgneOLvoVBX5F1qbxxOZGUva8vMj9up9GVEtrW4/I2qAERctm5klXoOsq
6npDP+mj2YIH51DWeUPvDiQRVVZxICDoGCizMhLzb/90WM9OB80B9Thp0gnXOmcY
d1AmxwdfexweKB7WGbmw/ylLWJaytuauw04Zz/13kSTEiCLtqolicck37xNrAeAs
BHsYroZ9Acokh45s9Q/06g2tejvZhKeiJuhtZyv6uuzil14qErSH9n6BScslyZ8n
clYCDbNJ2r+XJwXNlEVg8ZivmBARGqI2J/os5pww3whmOhghxQ9wgujm/XTZ5C9h
br+C+VKbfcr0RDJ1ooXUpnjMWCKUhY1AqspnDWjn+eqbbJpPang89irWpD83HVxb
RcxIzr2ZpLnprigdYH2I88DAUOAaXDco15zbRi1RmJ1HtThsn6OZHWFd7BDaQrtN
P/UqBzDqTf+tSTTRGku6SKcQo3FEAxhH0Y91glD5a8FEp0+rDOHnRSyXUoKkZgYV
v9znmqqxH/yAn2lWU7c3wolQkOKAb72gNyHgsSyMG3j2rYEganV1TGW2PvtenTTP
XeaWVrcU1kxs5utNs6E5TlZa24+9pYeZ+1rHp10nihIPmwgw4D7ND0yKaI+uh+l/
EpYRVdztJlQuMXRcU3niz6f+3eEeqzswORB8RYOEG4MSsd4PpCLcV/sHLrVDK0kV
3aHNb67c0xyLmqXnEfK1Ivn21k/3+1MZbpRZWXpojSrlcXANI/y3j9/2adUjYScu
ABLvWwyfTE8TmdQfvVgiquLOzYnq/pq0EaIwfwJdfwz2oPFfDYgCiImNu/ZBD9D/
pylthkoF9GnPR+eHbaH1EqICKHZ5oHho5c01kiXCgZbjHDaF8MXqwWjp4VWritXY
Dntcddpg4xyQsEBdJVnn698FZhB3Ks/2IoPKwR5GeBffCGVi5KreI1vqAtbEnuKl
D50026f/HrBy5zVxRCczv6Wi5kucis+3ZfDo8eJi+q0wWObQrVmjaYTqbFOyHezQ
/79MbWtF+JXr8rbMFTznJNCUlOwsGC660J3lnwevTd7C7+zUFV6Yd3gg3+N7ZvL9
zIhydAh0NcgUwWYp7vqDQUUc4KU58q0wnA/9rIgrnKeCg1LmshCTo/D8q839oz8v
VWhQXlrMfDNKhhdiGPT+YRIqy7W9vTJH+6bX1xnBtnBWeaZ8AeQ76wlb/OAnFQCU
9JesfrMDR8fEl7grHQEVmk6LnA+9KzAgsC4NBma9hI+/RLeG28p4rh9y3xFGjVEC
dsttgUbewJ7riAfe23eATU1qpZg9xCQ0ME3X6m3fScLDEkXybUc2xcryjEJdsXPg
QYb93k8YiJC/2ZzXOPD2VZ76eQ1sim/gBMGulIwRUw6sNGtUPpC2lUZInJhLEQjj
wjjlCV9l/DZVpcxrYTKdeVLm5Yw0kZ5JDc8MBRbhzM8rkqvB6h90u5tIKaF3wpfN
VMcrT/L6BTU/lhPgGsU3OO0YSAmTQb5y4nfpZImmyWOU8lFiNJZ13qjMd5TzJTcs
08/yU1zCyNRB855qU8Kx8XhurVnk3/ebPuszpaG7JCV0JyF1yK3q9awle24NzJTa
dxjOqXug2KxkEW8ACLn/7qxHyG9VnSG/L475DkY/Xog3eRz+T/fIOqugU03xEYTp
XkgQy7qoLl2s2AiCoGL1QcAa0Ts0aJTFpIbY7tlo2JHdD5jSenq4ikhR9szBwGGu
OYw5tc8cWZq3+SEAIR3OtpfYRUOkbf+HwZhy0oNWcXQKQCjCYXV5QNAwcrCjS3Yd
ROzw3gXIv20dcpbMQ61Mb11rv2mTPS+Q6LaQMy/DA92DT3IIHbIWXsGAnnuNeWo0
hXjGgtzFF55uuZYd0SRxPIp4bPi7sroeCMgooR7Ht9JwOD6P8LT0wQEcSFPmQfWE
KviQGPY+Dtdee55jStpS6JuBDCQ7ySFdru8G0ZCFn6eiIH+FT0acm0rDhmPl6yY8
QbBtrIAwofWsMQvmbbnpaXMESvnRmG8QbaLiX+O5Gc3H+2aBKBU4YZOTG2mvG/CJ
Ghq+p7/y5B3DjK66eW7NMEzjj2pCiZiSelX/JtO40GoW3SF93shFQhhbglNFJ92P
fTQx8tesIwKpk5FtPCtj2uRH5kgrAF1Rtllll8XE/DaECANDnKHWKNBQop4krd/2
NKybvmQkRBIfdyAvMcLDTVF/ZNaKu3KmmOCS3xFskrcDaB6Gr/Yl4Yj6G78krDES
BE9u/kNRz9Ro20tUIHs+loA/vkhE/MdJn5BW7gW0zWBJcNRTWWAxS9CYoEnzVi5u
+iM97HK87TaZvPL83wt7e6foa5KY5gXgv/rLYibGi1nUuxMfLjaDs/2IOPQXj6xX
l3Nroh3f/qNeshrUhauL7T8DceQ38KFz1+29V8/iEanJrpKp6HWGxhuxpweAcU3p
9iPIl5gbQ7H7WP2d8OSfTiWPGZSYUMcAKTaH2fTsN02paqms30q0kFt2i7s1IjD0
gm9ZAz6xN6TFc8EyJLXI+45EJ4G/YFJWS03H+N7hsgptrxWy12dpvTpucrvlD64x
0CUhZ1ardwNZVZKji8e+/2Ow2Vz6KRWR7zYDWdWBgz7HHnVPPUa3+Cc6wIHNYbPl
dpufzZgaiX8PNEZSl441ymGhhFq5qqmVw2ZtrvYRGTGYrs8vgK8b2c5JE02LdsnJ
IzxDaB2PV3H10uETFgwvpASixy+IoFISlAS8TMrBZEAfET248jR9ZG1gRVoekjlE
GFpZrpGEB+S8ldpaEhp5bqHN1Lb5c+37z2qat06RzAkyr0mAFCU4XN2hfEA0s07B
We9PB1808SihPzmyCEi4FYrELzGtA1+TU3biZfFMFqWOx9lStWs7qUJx/nKfBOr7
Xxqf0Nb5+Wq6ynHwiN+gAnWAYQFsCdeRtkWdek1uz/ntb1791grjauAAJfZBA1RT
6t/OVxW05gXUE/bheckPd1hke/Zd9On5zWds6OsgatHg2p3KhqXpnYpAb2N0Gmvt
yACpaF/INU9bD6ykeTeb8/wn0/BZE9Y6kmlcvWTFVFlxgENZSNpnQOdZ53fh8s+Y
UL+HBQyz5rP0NGnCYsBBkqm87OUtagPiI+T4S8NR8NYQYf+h/pDet2kTgy1FM2Ya
4K9WMLG+KQmr/ATkVdaR8u37WMn7yKGVYct4yZwZhmExlnIkFPSanQFLDg3ln8yW
KVrC2VGU+vOtNbs20gYanYxWvZtQNirX6evS1z3gFsd5dVJRzeoihls7eTfPu6N8
xG9kTBebHKdsSuG/s3/i4+0kTTrSLsjpgzeHZLiaTb0IhsRLOJ2/tyhZXB2zUotZ
g447EKB0U5BhZYd3zmBEFQAXOcjMp+z4eOuZovyi4VzgWz3RCLIEiKY3CrQ9dzsJ
GvztEX4BDZDWcEeWldWfHsmAduBiHplBQBLP7KJvuthMIs/MGjqGYzywYlKnT5qo
yPtgHtNVfjtttXesOiQi/GXstjBQ8Moq5JfIZwZNp6nLvwMVg+tfw9fVCgF8IiK5
CF01es35rn+z9LRRAt+QpECNLnDkTMWu5vOmN2ORfcU3/lfAVkhEaMTRbOnp3nb6
7sp/CJndBd5akmXq9soimC8oMp3D/DZTwsCabyWa5AIpHyP1pJZQDScmqhsJJkM4
e8wFy07UrOACqNB1toyPtkMOHhvfOzUVTgDb4EfH0j79sSoBzs1OF3mvj5ktx4SC
YOWQUqu+drjUp12VodBI+y0/Zf6koGlVLBJLEIAPm6sMg1ACGdpwRp03Kd+O1xVi
BiEqkxSuVmG95HB4qWOktmRwzxBpPrjwI1VEkXIg/sRFupHtO7rTyJymVT27i2BM
KxJFR3bdY5y6dN0r4HuawOZ8Rs51AXG0z667xOoHkqEzY0DzY6l/qaLTbHMi1u+J
Ww3r2BZImPw5fSK3FPeLZ0It0cfuOtBiPeXDtAKtiST92zXfSGVK8ijlvYywCWPb
DPZXge22NMHo/nAcjNS3mNzc8e3LkcnPaSgmGxZcOZ90YgVcS3W0uVdCmztGLYkX
UowDv6v4Ic88f/z4R8JHNT2bm6ka2Wg5getMO1pG02wHLvqv7vGmtUGOYHKlNP6Z
MuwvFPR4ug1ATosUHy96yUvdE/FVW8/8bVOJK6zSzvY1d/9pxKoESmJJlup26TSi
TzsWdg+iJbihjNY0N4Bcjp537kV2VET/zSnPQOTDGOgW2kg3znpZ+ut0PEVw2Rez
PCEs3IabOUiTMhnN8SP4fdVC6yrFo4BM3DuHADonKMAApW25mzSjshGXGAsU/8t8
YCydphtdKWbk/n2tXeuu5QQpn3yX/p/hWUAFsLnQuBpP7xyvZGbDZ62UW3XGLR+b
ImxpD8gb8RgkyM86RJktzRGZgd03mRkfRdxvalQhLH9F8ardN4gsyKShb/3k5SCm
bx1QwSLzoeFMsH77qY9zAUjEecm+0HmfZON2JjersaqChGScFLW84bw561iRQ8Rp
zORSWmSBNEIAykiFyQLmKctTvZIupEWLS6CySnue9NSHJUqfreLVPSa762AwWYg8
2Nkm3ko4PZ+KTxqw6sGPXRbrHErrsFl5BCkqN4fWGTcqS5VsJtnH2OgrxjS/7/Xa
86MxpquvhrvzuakxhOo1jhHMbi0DFdfa/pS56/ItYfSvJ1tIJ465amUvfVsCLX1u
xDCa+WRT83mJZJTPuwBLe20NFidYte/t5fiGA68Ku0Aq9mLYM4QU0Mc4qOmOomc4
PxTk68mjGyLSEMIrCAtEXSDKtY1+Tlh6SqV2Yv2/3SU5ZKrYnrYZkGoAoHAfVAM1
X1N665PdyqcEV9Q8n45NI03xNP60ZAqPVKEU2GC6THAYylo4VxugFhDMXcuNJYki
GQw8E3jbBX28RUEJZ63onsrHYSYekMSwR3uZFpq95G3x3taxmFf4tYna0UDjTVMW
wpwKOdj08UvmJk1YeCz0tKpH4ZvBn36wA5SMvTOcN8YY/3YbA6T7WpDLpIwKRh6f
OXgUgQCIWAl8xP7WmvXYuNSob4LF6X30XrF5UdRrhScJmy95yXyK0Qq35U2RBCTZ
IJ1CVPt1WX4jhMXPjr70w+14LlYaaNQmo4kMidM62MKp54jZjGxco8Jerzdannzl
AT9SQUX32bmsuiXbJjR2jLz1GVxDLz2U10l3TVtWs3huWCVXWuB+dMzQUBpDkjD5
la4eaSwCxs5qLL3c5w2bJxZFxjEsxzPfhwEGm4N9tmt+unkpvAMBOlo889VDUmxm
Now1xjdl64ogZc+HjRj7LpnHVKcJKXI/1MoXNcT7RK6GHjH0pLor2iDCrSE4lcpG
lecbw/J7/iksRvVTeMigtgc8u3srTHl7iXfiH+P2CXmHS4IKxe3jVU/v2Bel2QBc
BiyxaYDRBQ/Ko6ZLvjgimYFjPW5UMvrvVicjY+TUVQSrhXABIu51Ny2J0poavGJ9
wsnJ2LbG2WAsoJdL+GGFL/68svgSHS++JWx5jYjCjCI2adnwfh5rrPT6BXFnUSkS
OYt/prXEBvud/RlDqFcoJDvjbZkpr2CwY8iyrVgAxTk2fUGGXaNrkhyuJo8Fbjz0
P4FStAAIuh10VDRTe8jOoOyzZBjLLoa/D0iBj4bo7PhhcG16i36B6CXH7whNstSj
cd7bWvoK7OIimyoEcfbwvcrBLxzXV1JMjTLZFzBU3+FCvSZEWZ+SzeziPpmBRkaY
HSs4v3HxtyHXDhD/V6mdvEb6ItbxAs7ZzqPNbOiwCls3rtVjh3pXiv0ipL7f+8Pg
n2OxzbH+rLgq0k4/Z6RMDRo/Q8BE3NrmugoCGdZrAhW6qviJE/0/Zb245L9D77jD
tJ0/A2iNlY2BAGVGd16GtXQkQHzq+/OEpePsVoK7SjxUghSKl6e8/GQ3Vt5KiO+b
mhwbXQQnDgfYU+M1tHtYgiInvBLTdOQ4NW5LTZlV9Tu14m/YnT3sRsTeKSwL0t37
OWVHbsgcji+snyTEaUHf0g07CaJJOy4As0bgx+qlCJfm1ZcOZp5GGWWbAQ8UpLji
gXhSVkfQkVn982TWWaZwJ4aJWO2PngBUDEvEfhy0huR8GP8h58Dv3TSoqCNM5DRl
VOypwEfEvTJxQYC6YWENPU62lW5zz9pTjNR+Uqy+9EV6OK1nxGK6Wim9K2IgAVSq
AIlUQRJufXfIVDNyIeYlmEg29PmXg01wRVzg1vp5t7B3CPFUw1M3UIpTkSSqb37f
rDdSZyMAzkKXBl5louuo2LZD7uhXBEqsIClntaidwJF8zN2vv8kEpNQqqZBee9v0
zZVHXsMk8/06KoiD1hgJU5cdhF08BZjA5BHWNWzBgZTswexyzJOAvj3Lr1p7rPCz
t82AdFSIripbJr95tvWkPRHPqoxORrWSKPra/qCN9YSKb8C34s6NW+lVaZr+CQKn
lxqD78xC7z2v3VVdq2wNfj0m1p/0MQodmbHECgHVf9vlstJq3t/+d+ajECN6jT8w
htVrl/2HHTUFGwEJT2Yxr2VXIWu+7wLg+P4f+SPxCgZ1GyBKjC59kt6jtHPEDVbL
by4gb4QsAeCHHZCiry3xmhDOvYs+2qKKy84SQM8JoJRMmwdTHafsSXKTvnml2nAH
TWS/OBU9dn8DN9A690gOX9leBI8puK1s/JpcLWoGFcwZxrj20VIu3JHMhXanVSgi
nYzD28C0htGOzHBCecPcPD/MO/WcIe3MOL7kl1SJSM1zgrACpaLbUUnt14JP84za
qg8u/3yrBAidhLA0ZNunJdLt6foadGZunS8RG83+OGTZu5D3Ug+S07Rrxnt57DaA
q1jAaNL73dIzL8QigednLmoCnoYgOJ6seCTEOpWbAReOcU0MxKLJbSy7U9DJAGY2
MHNNiTl19ddXj3yIR1RBBxolhQ12kasvZc87i7BeIo+5EWsy0uNw38JLSZU9FZuY
ApCtNnoe1Tv115uV6mawQqBW1+9aKchPwXvEnEB8Q7CeWoHvDOg8+JBD3BPZbtWE
+FQxvN4kIDmknEeQ+de55ApoizOBJauTt7FIgnMx8H/bfwzP8u4gUUeb7oV9SP4E
urnyUnsjR9ZiuHsMjE7/X42wuwb60kqZeU46/b1U0Oe3uo1kSlASvHps0Em9ppE2
TTY+4aoy30Pln6F6EaHBNKk5mxJzl9XmbQhjcIzrH4BD1n3jmAQsucHDIZm27wmd
tP/0SXbqlKu53zs+wypGPXXiRmx2Y2qLPb/UOm+nZ4vWjI0nAZ4waFGpTkd8SdRk
zdiV5k2hlCFfynDVdw5L0Ili0axww4urIWcLP8itFAtXctpug2PZYAjc94zCh5yH
+FpPrc5mzQ6x0bnJ/PVYHBCT7RrsKZ53O+/opoBfFOpyPAiGMx+s97YbWb6cloZ4
xc8XWQTLtp9bpLjiQHoqTFpoc/og3DOaxUKn/tWULODWaPV51EYMd9TYFGefMfRx
9WLTw0YSURBeTQKjcxh4KKYWUiM8/AlH9i6kKeGgC9X0L4KGfLjDikxzse/3NC4y
doF7yIj0NmdVqAXPoU6Kq0NoP9ha5MNp3wyoS0x7r2at5gG+4ysFoi5iWitK2DhG
1B2MME2TE53xpoTa8//VAQgtVZ4IEvATGB/l7b4lOvcvg4KaqLSXL0uvRjDEdfxI
SJFb5plQjBDVLdhOLRXpHzCVh/V478StPLAcBZ6xwakG7cL2jQOB6scxSQK/WtSE
ElcSajOCdz58EeeXu+gabtO38tgJU//rTrcMxt6FTJcm2P6V8KpBgnO63HX2xJYd
iS5Em/2lHFeEPZ2q6rpaCQy9Xd3iMtToW6BRgc/zLP2PGj1HVD3BKQ7nEFKhJ9ZX
pLthFO4PLpEDVTCYJTBdclHXwE2q1IaAsqyd1t6JDrShaTZxC04NYzFusCxD8JZW
PJx+TyuZPWob4GCpb5NDDc0ykQukokHcNfgJcbCkevyfbwjw3F/b+c2klxajvfkw
0eXh7qK4oSBWzUkpyi2B0SgGE7ZoLGBIp6zSO2F1fcmZq8EBzyCfPNrdxxWt6sP7
1rwjJpNRZ5fXPIbp6uyC3oiiVV1iLu35hNWwNWmlM/NipS+344tLcp4xT+OvuSYo
7AMjew54Yi3fG1jCuDSOLmWyV11XO1O9EhiRHbWBDtdy5eCptwEhXu+2cLZiwPPo
VpsmkMGIteMs4BRb15FuTXEI1ligLjvlbj+4i5h0sTJD1DkgMxfxUr814CJS/hUd
1Jjvu8m3/GHjjRPDBLlVbs4nwjNRzk72ggICuJRqifFr1F6uxkXKhzgU513WiA7F
jz7lS/M5nURJPade8MRYMmUVGQXuzq1/QfMDGyB+wT4oHkHLo4kQEkonvLmu1r5b
SyOA86kZOWAicQAwfibJ8g8HTdS9nR9DKqZBb7c3jAbAPBh17fSHCVsWOJR0xrcS
b+lMAJcleBl+ezEAmL4Zw1PkIOGaMC+qpWtYkXdclknEopqSxGHSbKJ3lcvFiK3B
Y5kZP+V80mzIhYO3+zYIs/D5v5+BiVuXmJgjxeMSqW0DqD+kIF6/dZ3WuAwEgfWr
nv4h2MgflKVnF1unrTMfiPFTdzW08DqgRQ7R59Keg9UYZkrACDgiiVXAUiHIdh3Z
yC7lZtMIvjOBu/XWaRpneMpzWZUnjj/pWVD+D2g8yhOIQAMPSn4noL7UWJSCO7Za
xe1vbiWWYY4fnjxGGvUo1slFdbZdeEgsgGGAfRd7kbeIXiDLydn0TvWWLna5co8E
fdpmr0edtE0ZfJPHVQ8XXfkaHii03/tkocoQAG5ytlu3w8/nhmeJ1O0GiEztSDtJ
VDLF4RYGcX4YvxO3+WkF2ULBtMgavTkBnnpmTK4IKfnucWE0y7CMJGzEqlNYor1t
y6nK4kXyClh+1/GKEAdfhkYMxNTXJ62MAAhdaTq+6KJczjuUAEVNHlFuI7WJ4I0W
PWptZkggQo9h3/QcjZvfCoFMRRZ9Ybiel4DUapHnVZyQwS02IEBB5y4n6V1HGDpP
/N2O5IQ8YxH7stbRzqi3mv2lJGfay5Qei9x2nQJNFNjR53RaOtP86iXDV7InCfiW
Jtjsu6vo7h4sdxbIbz9Mk7rUbJ9kRyJjLlsoVzRHC1WOV/+5CbQQkFLK/i2FWpHr
mm3xUpfXoGu0PmmXUNS39DKyPG4fRZV3y8DBLHJgpOQxPVl6kQTdvYsQVcx0XXCT
JRUsZLRXNR4IjpnAbAwAssM8TZC7z+LhWDEzwykhl6yJ8YvOlaAquVwvLuq2hwxE
eeknlfjX9ENf+ZS4FHAdazwY+J1YOXXoApCvgMPRFyLX3bDp8reNX7Qudsy0JD93
nQ0abpr49Yi22qU9ilR5umiUBPzRllCrtxnP/6G5U6SAy/su7ssljggO2W7miYfK
J206ZeECm9YVCtqMglYs2Kj9Fsfy4EE1rQZB4mviUgt8vmS23oHJ9vBPMDK7m7+b
6Ft9j+LCeRk3odITq5jbUaWbdY8r/wdlBNkx6NMolugRHUgcMpwNuVzknM4pcT7g
uZCRxNF24fpMjB8dBIR9nm3263dflPKFNcAVvg4XTED/RiFlSxFzt9Du47uUI4B+
d6FLEqu6gJVfxCoIV4380kosPrcWHH/kNTNO4twYstBIoHDi1CkvfThR6HieX+z0
WZ3F8RVEtFUdrOU48JHcdW8x5FaIxHeLyGqk9Fd6VwrY8lBM1xqLA0AJRjqrdys0
esVLDPXRkititlAAainDD5gmXtXb/CTUCMMqXs0cOT2O/2j2EULTpObUmJU21cQT
1TMgjX41uhCSFVmle9PnEvT0BXYgZ5M1XTZQAb0SyLw6Zx5/GDt19pFbm9VH/IbW
bCrg3p/ilttFepWY/2Hq6FAldhNwTWLvkId88jBPLDZHH2MGAJwhoRT8Py3CO3qK
LVn6xr8eVy6IgOwzM44AjkzUyCQW2o/UwXX3+xYczjSFKS5RefsUC3SRgW1X8CBo
MtGCypgA0uJXFpD6LOIi8ZvxMxvLssGVY73QX/j78Ndnl4SevR3DnSyhpobyXtKR
ubzbMd0noIpkhw8DXmYM051arFHn2sHYApF0JvTyAwnmeLP2LSzXAe7c0hDg3hCp
fm2D85jzD7Z2cOkEYVo/gEtI3RVJPjk5xpBP1py2pok1l8PF0+LYZQ0f15InMs2m
FSKgDq4/7c6UZe8yXB0NjSAGhCWELkGrvohpRVKzkrMT4+t9KBpUiot6wSy3Z7F2
QTT6+djdlWMxJGKEHbHZ5Ncvzc1timPf+i/qerYjoDbnwTl1Pu9SciCsAledRrkz
hozK5KXnbvS9AW/1uq0ud/zXKDQTlh5dgmNiHFv9dvmCfeDmkO1QwGULBZzmye5x
S9F8NwfPWB69HMhkQTpw0cjiOgLsVaQUkQRW36pUcVg5Dj8OKqUHRvbPMrJuGFqR
3UA6WXbk783zJ0puFqWY+hx0VIgoYYxa5rRAGkZ/PGvvV+dXe5aFPB3qLG33tQZw
Aa1pkKxL3GGhpsgU1WNDJxgLeRZ0v/6Cf4IbhXZ+GierPH4czW+CDNQbbEs/Mju9
rgD0GkmJhf0cA1gaiCYAKqQsaqzIoJ1EXw99rlnG2Gd37DnvEtFpXP/geJyRLKqj
W1T6xxPWxM9BwRpXI9ati/Enwa75vKJ1olhvDmecX2Z5dicQhrZnhkm8wbOWO+rp
IDGkz/D1sHFpi8wg/YB4KkxnrxVGuBpUI0GINVdGRD/S4MYQjD5Jlx4VpyCXMUxV
d7UXglu1TR0wZj/G2NhAANZfDRb6T4poPwP833uDRx0FLDMsq9Ck1rx+lNNUBEli
iT45JsiAEdVkwnNJ2nAsEX/BfiGHtdtOlS9tuu1sVsJTnZnCYFTSUF6l1xsby2sv
F712qLBQFqRrr+JK5mxzz0Mlm32/2WDeWOvE9JL12PHce3jwpdM8v6A87uKjqPhR
uqNo0y7lmxm3NAfujsypmFoes9daClraHqKQER7xwvKRMq8QfhCaNY8LRIDyFEJF
L2YBFW8VVNDB/ibICxRpwfTxGabM8HbiDdFfGKx3nvj63lyXudHENkPDjj46P4PE
vWAcC4UoY1hAMgBUS4wGlfzibx41zKRxFYziYELw5BtewZ01ymj2U4kG/TbqqW/D
rgXX+QoEA7x4VX3Xob4C2uHeqPxjk6Luot4mvb8UN/kMMgDJ6x5oQEtkuZok0Dub
1vAexLGoEfSheFCD+ppMDnkpxZxmuuWlkkKmRIDPjw5yShSJ8HcJtfkCDSwhYg4l
WqYqb0wrrMhOkaayTSkRery2WzYiSCTySxXx9XYpI+jhvjU0LY5mdGyy60Fy1lCh
QHZ5sG3bqnTFYPYIaUPhjxprDPjNxQQdjqBOibD0I6OH55l7E9gvV31t0DWwg0lI
A15g0Vn3PpaoPY0aAPHwbxt6OUzd1/gYX55WpOOP3z+hZW7XltZdOAIOQSu2rz99
99Hd/+4DGQE7zcXYF6oS+y4KdJjAAswfB2VNIafhbKBY+uhsw9apfuFjcl2nCYzj
cgnr3Egkm50cF+lUlrK/SzrHAa3aWMmxP5fHu1byYMjWRy70dQTlz9CH2mHlPUXz
zhffp3G6CFHNi/Ci+V+SU5CfbmIkaV0+FRsmR2enFqlAdcbYDP+wZXzRdPtS6CkD
AgyGTPq/esgDfVln5v1qqzrRlnT34NB3B4Hw2g55HINhWpyDX+MBz87gX/7kAJZD
JDgsqKZum28gyKtKXIxq2eWOspJv6Z6zToN42GxrLJu86JDZptSyqHZ0oYIxMMd2
PSDHx+CC2+OMPVNj+btSt3SxH7XJLoh32DSczJMQFaOX7BsZF7LueI6N2xCZVkGP
VnGDIxexIQVVmZvjseydTBevr4q0yX3t6d7dZMFFdbfuNZfZDw8Q4RyvbdMt79Sc
kUZc0mXGkypKzJsW1OuuzLd5xzJ5PoEYhCZFvXjyfqKMtMFstPbWU5/XaHbCqk+A
u60y3Y+VYJkGzIpwK5ZiE7wSYS/brjJGhMLyBycwlOg6CEaSGpjv+GuF/hRhnUBy
TmQorsZFdAc5s9T9gSaSRf5Ekr6KTcFZPm6Op9tDm7gF5O/tq76KteZy7inFuzG1
ktsdRv3MvyQMA/t7ui+76D80leIeQ94eZpwjAUPp29ETGDMgJealpPzVSwQGRgRQ
3Oi9XVTEVuzTbcA046UAvT02YryOWFsYKQzbBkioeiEB8+YV7VOIfuQw41KyXHcU
Pl+w57lxTRJUtjh19G+D5jre0pUfNCj/rz0/CdQjCclhQdxg9+iN/ognJMySKE+6
53nQ2dxJthRKZjtgLDFnv92Ng8GkcMSXu8mP9eMsyeWndAkbOj8X9euFutkfwyVL
c1+DnUigR06t0RoD8Isqftbv3OFyTuUzAFFjmeF/ya8SNZYMS4qS/b74LFdjZlrq
b0GPm4sqbel7TNmpi2is7aObqjj6HlpKhilDk32JVWYvXwmCAJBem4R9+CDPgqAj
mhBQqwiKKhEJq1dt4m2dFr9n4oa/uqd/zjZPyINaz2I5GdNLviyaPb64RF1Hdaca
KynbjsCWlmJfRLaBOmVijAGcTSTgr3yG91Kg/BnvQ7ben8BtZJTslopWi49XsmZY
gzOUkXLG2hJzJ2IBTpkgt/2+KhoaIR+rrbRa39LMG7v30T5Z0MRA+7baVmxlKKTh
Il3O+k74Z2dmF1io0iCZiaGu70F92senqCFBr51E5ckbUZkAssVAtfYW8kLI/N7A
Pe6myPkKvez46uBv++SZXgfsHSohFB+3cBZ7ZvKp6cfoavV5SHEsDvMvuTiQg2Pp
nCY6p3mMPg7HU1rVFZRsshyh55y/23oHiL2Ay+bfc6XKaXdS18z09YVIuDgGn4ki
iVcXLUqrS0s3lAPML02XVWxlkhT37Fxg2LyC/I9wWBGN3AQOZYQWC8hKxbpKpT/M
SbVnrNuktnE2x4xUzPMJNn8hbY1J8toFPVYmaJeCOlNwEdoHTzXGU9lZk7r/yJfg
YL2Kl4DIuXu2+D3/MmsbU1z4CQ4hAKLooLFCMmc47MwdTCvr4dXDkhjEp/NInPdj
NkO6OI+n+xcXgX3b9dYfCw0Q+uSNNFpDE3aaOI4fjJCIstq5qS7TpQ8UfA7BWoRy
QbCloHJeSQzCt8NhUu4Y3eVrTy5TgXYpAoBX5cK7SLPEpO/qPafAQJQBhAkNiQJn
epWC6oKNOp+y4L7sW07WBFebzAjhN/Jm0LyS66O9Ac73tQVi6GeZhuWU7UHY5TeV
ePOdvPUpOumAIXZxjWaelvZT1OCwY4b8jKiWsk07ewH7YHatDRV+ov2pU4ySask/
Is3A5WUFUUabvCBS6X1YdHJls2/t/KDc7wcsHTDiews3n0oMLFkxcET5Hp5P5J0k
3qlo4lodRDrpRVoNEEcqPVelxoXycCRmiYXFKj3GTuDO/kgLlN/7Z0unUuQTt8UG
UuCQ2/Dg47VBKfnCICtr+0AT6hHS28ERWVwgjF/PGBwA64oBa/8fZybQwAHI91FL
2HnA0FQuUJbfVeXJZq03eOh92izgrtyXJNSDPJjjTHETomRq0MjsD3xaNfJrLbEQ
CQ3ddJWm3BNQt91viuN8D61YrtH6Q4AOC8QiFLJb5blF89WIC9+Wrf9zIrcyiNLn
RQDuzLWXP4E9h7VwDBYpm0iX+AwWRK7yM8tfUplTxuTj84xjHfCtpJ9uD+xFonR5
sG87jy1E27/kGTeLeXrXkz+gswNgM8NNoa2BXG4pAkLAPUF2qnRMP9VIUEVxYNN7
xl0wjcmeCBynHkN5PvmOIx39dc8D0MAMYR8O21UMQF+2zszKH6qP9IRRCJ4aPVSs
BjgGQVJjfW7GnT01bEDpLsaBH0mvaszZtIfMMDdbIkLm+Y5BLwFj5ylNHFOVCNDm
q2RydnL58n4Iaum9Ck7699+ysGgRheA1nLWWSdoWOWbwzwgS0CXey9AATQnYByJs
ZtYw11vmXHcbYs0JvZC/ztflo1IHGGE0oJtbsKsCXRrdLVAMrG/JLqwq6I9Ei6mp
DJRKT+0dzTdmFSlOjzSAIhcvwqA+Oa4mV6cDaQAQsnkBTgIqhHvqXhQ1SKT70b3u
6BQGilzvpaPDt6Oo+JOLkXWqLhuq1751AWPE6LHFik1at+WNxTW8Ph0h5G1ENs7n
1efOrPZH5HUne49bD3aeVHOCvxyAjsK/C0GcXphvM8qm41DLU7OrSiFu4I0mnUOS
oXupYKqlo/rwl+HSH4mizlZEJqyPQzjzrOwnX+FMxMaOH1CpQGnqu7As/C+vq/+5
4owRVVus4wDcBaDYIiHRqXS22Q9wCoJZxaOwcSt5keE77iJGHVwb9xqyxtLN2cXA
153kOgogBzoiCvGUXoYo2w84z/XjaKKaPkooFwH3TceGgZ6sd2BV62kiyE8X9ZHe
/aMtaFNUAjdvZwMXApM/cINq12ifOipx1Ve20Xwq9pnjOfw6DBVzJdlekTJdvQmi
4QfQBMyAc/NW62VSuLyHP2/QnTt9Oqw8iuPtalur8Zkr6iKFxGNfKekw3659cCnk
Cgb1rIetIw7GMf37rjV76ArQiWay06eIfca7zARrutL5zsQ+j8cZCaKJh+9QYAd8
ybIsknnCBWWKudgNkzh9Ophqbql2YwWfber2TaVoLlyrO76IHwkZM/CMOEOCWaJO
ZKKdXZdtVU1KEqJeOXnqLHZ+69+YsgZlSvU/VDA+doWWvUzpIKZrzy61YrCVy46j
xjpNaUMaVeaU6XHnKtohJ+tCAw0clG77Hl2BEppqQ0M8LIQXTYyybZoE8tkV/zvm
1TKD1E06AVBLnI+6vo6k03c0iN/g5WdrjgCygN1vXtVa/g+WWSplvccdfkMrHgmV
801NfDgyLkP8jPt5/L0v6hCCROQBXnVV47QnxLOiJ4zxV5DkNvHWiESSRyJytzFu
8ZoI9TpyQzTrC3hbZb1k10QutAVzITXU9NWNtGR9rG0mKDVwVdvjCSTyZlXbw0UB
/1rmTmbp6UzxidjfbpZFD4+AXyXtTe5cM/WAb83jOAQkCA+Qt8/TnBcVkLvsGCUO
aVry1d6h9l0bo4Lb2lzUDBrR2RTDC2Mn+4dpJyKWkD3W7fha2PrKJPIFZRNuPJLL
q37neyTA/QQgCJtlYNtu7pxIDk9etEKWMlZNz1qMNKQS9vgKRlhZwiyTjRjWfqa1
lu5w8LPmReb60ujtAuYA9abbtmxufGQ3qryCe4lpG2fZX1VSHw6H04W4198ommyW
KQ000GPfjb/Yl/yjl1P7GNo/EUEk8XrY2pT6Z6ZJurqdmrfTTOk2lHJ+GFYuF0If
JobqehlpB4PjuKf9uniz4hbegJEtURrrTm/k44llVr/yqDygRAUU42Cg437Txa6S
P5Z2CU3odOb5lzdulA8NHSrSmr2znCcBn1UK1+6cOlcas45EHTS6Mlx2e3kuVeox
TxpurQf+L2sZAJClxrmHQA0uGAiIrZaiLzRmevRoZwYumlCxki/MVJ+tB6eRajY5
DEfZJce0ve1jOm6XHwKb1Ejps/0m1t1wNcKqcE+Q2VP7dpDFJ8pm4vOV8+ds9sog
iIzkFIiEQa8kjAbToWlgKLsLPIWS8EH08f5zkRBdGzI58pRm7WSAADt35/1AiApY
HxTDzwTEgt/XQQpwxR9LidpJla2yh39UEJzhLY8uGZqyki2RuqHFJX/1fzoo9vQd
ddea5s4XcJVxQZuZRBvdZPw7Dtq+WfuyKzWtvrypXTxBy7IKufyeXzV3sKcv4m9c
89dTBiDSqciBBgVYmOSUE53XUwxHMw5TpBV6Q5NL0mW+WORtSepoV8XvyaATxVYN
z5Yib0kdnWD4SxMZlmCavCDJjP0oLIQoakSlZsRmThQe0SIgO52J0BwasaaS7Czt
TR3j2w0k5n3NHBlSTdhJ0mgwH+KuxXQ085kxLKFGBwsJyiIUN4QHy/wDVymJSZh6
sYUzvI8pVpRdKNNXL1A2ENaN0c9M3AtJF7dDHdV654Gv/sfMQvkgPiL2dwaKcx+N
uh7xjS8evQZyMlpb780Au0cG0VqaFwWDvxm/TDbM+8Gz1gJDM6yoxeC26227BBJm
fZZMFHrZ1Yj0ojaMVgguwqm5+1BBjx6OdTuDyK14dUc+HkswWrp69eSxULYmD95w
pCIg4z2FP0C/4Jwu9eGckfcof/cDpgbY/NLt3CuYtuj8OciNSsHIRIWHqkc+9Qwz
1YZjyJXS9MIT65aiQ7l29OjbHy5AqpHl+Tliq5Zfi726YNUU4xfpWK/0LAYjpbJr
CNb/GFRxOKXkVInpUK/KBgsrjXNyF6F4uatYq/npogg0nQqH0KSNHsylpMcwcN6v
1ha7owhwbI52GDUD1FHpsMi5GngEOnk6mw5mM4faJ+ZyGHUep08k421Fhdy+Vej6
8S3o9G8Yb7ZxSflAhlCeTN3a65bIPBtiI7Q28OuTbkTEPmnfAAl0HW6E/o7QTmXm
D0QKPLj2D5bxj7wRHvbhm30ekoXsZLWxNa1TRjMZFSHEQ4BO5YEc9c/ve5bkbi9y
hiM9jh6/fZOj6pnoNMuVUxVW7uxYaZosOhAMISmpE38p4ZnXgxpb9pFi3su6Hcdv
fun4AIAQhAI75Q7BUhnHbJh9N5Rb2laLN/WSeFZCiHkj+2L9d460JzKx2JDV6Jw7
9fI0eIJIe3eQtMjLYUioFyzu6GFhnU82KRTrSMd4ZrN3MWjlnP7tJnTN8LSe7wVO
2nLDTSG+jODq06LaFrypDPfA3iIIcKslfx+Keo49VrJ6g7qOWvB2hgawUyK9Ght8
JAJquUviRWuqLxgGcs4eFyzGiUz/p5D33gpUBW+UaiS0tgOjStnQHsEcdqxQA1fh
mwnPmG2xS94hRj5pL0MpB/j5RxF0Tjr9kgxJb1YrQclmFn+/gttV19fT+KeOZ4XV
Q8zblTSPuD11WnkxPkdQ4IloCYPNjmA1XUjv37HJd2cYWwjviotQ+zuJckUAmfIU
ktiLsXXIgloBOl/4o2aghR/meeD58pbnMGk061rti4jU69DP6tY1LiAFJZ/IzOnx
9joEQB9Eb79vRbrAMwmklzBTC5/6GkcKUiieUleioM+6V4ZrMRPzEk/tHaVVfdqT
S+Ehsmqaj9gAB0evJTrwKE1zNBSfBxhELRn5d+tu1kaMTnge89vi59RGZO3+uqsH
7S4XNvynGDbyRVlA12+rOAOCosPoKaICyQpKuveA42trYJiGUpFN1Lgmq5ww8nbm
vnVIF8FmjuVXDfClSamuHr/Pjk26By6Cn61w346qpCzC2Tk6OfL9teQVxn1dXoqN
nZnnYVzB9LNb4NDlku1LePnLmBuaeca3Q3KUeYb/+3CeTvMHlsDGkawOx93R7a9Z
Kbz6IgwTLHmAQHXMrQA/NCNQDFtyMXOaL111IXYfruvs89FfwbeTS6b/+Kqa7Srr
ci0hWnh630AyHYvlRwehmd424fFf7Vh9S0DKKWAnkiDa91ZDTmShQzYcim3eD2rB
TWkszYr03IVAiLLPuWcanPruifZokfBETedi1xTQclDvESeOn7kqDZHti8G+m6CK
pyUowvjJ4jDmcDkYcy/02u30jk0zCdWvzC0cn0UZzv9anCjIFkKEMZcRS5feCaBK
k1Bc9TNzNSy86AYQsAOJmp4cWfjWtJ0SYMJu7ErQv9DhFeix5lwotkhIj69RlxvA
cW1Tf1TSBhT45QtLxRh0cUhOL5wFL2xm39z2cCmK1uI2iiGBGD8jwETmwEQBCD/3
cwGgBa/D65FK0NrUdr0o0S9ksK+4QhVxDQNeOBgBeRVzWLLxhZeZkF7VrHDFVSg4
tPsY5cAdzyGh3Dr7CZUCanfjyiAG+7UjG+3a1FcyRQtor4ApzuqZuJLq/RfusDb6
m9YHD+5NrT3I/GbkikFRUtOqTfqzzMrGlzdqmXC9ZD4JaBroLcRHNS7ToLDBJZkf
GRYWJDbemP62bCuKkYPL4jxPhplIGyjtRj0jNBNcfHJVe/uXrY8UIrlE7Uuxb/le
w/MRwCVJBVQ/P4mbJ4uiASvU+E6AAFCxrxv9Ua7vEZOYFIs2QFMj9P/kWNw/Bpu9
khEPW9CbKDQj+LKRcm5T8EqYnUCSv2xTZjYHuzUBBlM3iG2AeyuwlnT3xopGOPWh
U+Gdy23ESlZpFPtra6CNnFpIB9ogDBkZ2RhwOjVgw3Gxr3B7RwC8r0OOFPLGTCYF
1lkVtosJ1fkl/HPAhAWTenbDLFI4j14PcYBvRep7zRACGSblorOlJCMWcCOiqgzY
RGE1CyvSib0aeIJ3LQJZ23G9Zo/pdTc38qm3qKs5sE6JKzPY/Cdv6hM300kJ7OrK
8QmEDOcTgxMnKXe0FglEfoT3lByLmBcOFgb7vlHd2MiN4XjgDonqmsbRQS0ZQiRi
EF4nAm7W17X3l9uhyMSpShJH/Gt5A7V08Y6wHCTIgObFLyVJ6pGDVhfFFT9gSHL3
QihAufP7obgR1cx+GVIIZ6PIF6ryw3t8rt1stfhlPu4iHdfCfjSOjiBQEMu7+R5K
q6sg+b+xaYu1IlTsrtbvrdYIhgfqUQ6dJThS/2hrzwcNYbphIcQ4h8gZuOCCvwLr
ZTrsjRHGElxz9TN/VPtLTstDCRczy/DTCf8UlLx+TOex7cEWJ/CLsXbbX2AwdyNW
D+3QZ6UP+F5QpkDcBtkTbY/SE5NNLreTIgjTzQyhs7HXklxW9vd/R+R+EM7EL337
J4b9J0sERyRFPoBF3Ow2QneVs2rziayLGskdG//CmYkJXIJUNmKCFD8wNGuSXLk5
0uJ4+TWZ19C+EkMX583zr+8DkOnXR4XeQzFVLaWBOaOFW99+Z0P7vVvA6Ot5LgsB
fkPNp0KxjZ09rIh334Zfmgn8v07+uzMDDbSkjRviZRFu31DGu6LMp4mOwLrFjEVb
BRJzUGa9oZzcMfxYAZTL7hIi6V70CaNdhnSCx5iA3gQJ8bRjJCp4qxZ1dwObzoSw
KkojrBB6jeSJkzWgglZ+l3m9AL2d5oVTUjAdWdyrOorUMLxC5TsS6+EPJyj+WHw3
io85+V0EQwiwNZXCDSHJql6vlHGvoHmFv6yslFBbZF1v0yy6JjotUaxcJlTqyKUb
Taye0W0lDkOadzLe2dSy5C7Q6X8+i/FBaG31QRghgNInehiN5vWlUSLFxTE9sx5i
kM7OyYW0dtzICK2quD9HUV+NKOQZCSxfQFmG4vIoQQbUKlSLDaulLBQY5wkLN7WU
yqqqtydRaKdkCEnYs0wY4HK3Hbq36e5abVFaWUKht4HNo17ItLzM7xtBw1KEGbGa
2tybYPDPGYMtgQ9HcfUlMJhbs2fllvlvAeM64xNJw0LHEtGZBBZZVnVhBVQr/UiG
ofVJs17clPZnMJ5EjAcGwfuHY5j+YyVNaXPoHEXe3Fl27bv1olc5JYAd0IrAWvZY
wx85EH8RqVylY4X77Q00JtFjMYLtWYh1eVR31jHaKyvAPRMqvXqEuuMLI9vHuT6i
qcVguM7l0CwauCNRSeylvGa8o2mOol5EVf0NE4G7OujMPFopp6QJ1MsIxNVbzque
NdEJhQoqtpwkoOu1iVDOlPlKXTPT05oUsUfa9dK9ohr/ClxN+DDpcKA7OWVYllRD
V7FJ04KjnibUhEl89/zptJbxLMsv/9LPnTRr1o53mIfT0dh2Rt3XBtu1CiDAdO7c
tYlIk57jfRdkG4GHJ4g2cOMjA6rJX5SPazezp5SKBkHoZQinjqgGC2hNZoSwH9yU
+2VUNBbbySGN7brFPloC5DisP9npYxrBx+ZCGIJOgYDX0FpfXuD3QN2zWDDnYblT
jYFr5rCW7/ijuFEo7PmdrterY/A36QcO86XhAGaXJ7jhvcD2knCF+Q4f1x2Y0vyR
ql8rSsprwMmOtXrBWjqpW8tT9QqVCf0tZ1HD80wI/+OQ44Gxo6ky9edg9+BuRW1v
g7RItbdRmjIgQmiWNxR6811YFftcpsJ5pQ8ctqtr49Y4wXyIZq43Gl3lCdrgjmRz
Tgp+LIMQP9f36Evd9UKztyA1/7hpQXEAYrLlfnl7vDlyVr13eBPir6LM7dUpPNmW
pfnepKBnzMJAU1shTodNFPiHqG6voENTDaukFZPTYSDQraFCm96YD0xwt06Ra2sg
tcpVTkyIOUM6ldD1O4wYVKg6YMHnODVH7VOpDGhUFC7gCHDrokzeEiHdmIAoG85q
tGdTpeEFfWsuA2oYC+CwtT5wGgObLc9CbMF07iAfxM/kgTx6I11VHq6waQ7mmsQR
sD1rNfssKlqXSutn5+erlX+3qeAcn/eJ+1UpVyXLpxEfsluWIRt0bIE2kR4nAEI2
PSxSm9kxfFl7XEHXx5oysnLZnnUftV9mbCqe3G1VAMJjRzBOh/AcsITA79IAqmda
/PGhFGr3Ty+BBkxmJ4a2jXWHOCmwAkWI7aI/jSXphKiTd6HgNLYQpxm6+exaZQZ9
eqVa1wVvZEEBGjToDiTl2J33QEaFvAJhkmgBQhEuq2P4cwk7WYfEqY/emdhntpyK
0xafhgjPtiMeYBm5A/b2oAa682IC+FpBzw5Cvu6pmFLym8GZ/YymTvxZVlbGv6PY
e1t7Tvb09m/Vysg8eXllqc7CmLQGQVkiJUGeY6W1XgzSUC/+WvQxzImL1NDJY3AL
NO6zR78eYYHrH6uKR9g+g6zACrJV8Iw+Xqx4D0mTRyC3DPKYH2BpDnhhnahnSfJ1
D95QYCbl0xHOVIkGQNlxSuWA0Lej/FwV9FV/9FquEsjeusez0C5LxFPwfJwcZzug
PHc+gzTEFh5Y9dedPQkxOGjKByXpi0NNm31gFK7wTq87YMVmbsalhpTCpF5Ye7d4
ExgAVewKuYIYegIvtTf+W6SXvV6iwy8koYkt45kZy6m9n9Mc3ekpkKhOEbou/NS7
+yRBVx7fV8BA3jbQGUwPczpqOmx1L7R1Ls8OfyR7mOgLFKDiedrGyfFae0hVEmXL
CWNrlTzvhuVlsB1bTRGe+eFhdmCrGyHcQhKhFnKUJd4Dho/QA2omW2pan0MDVupb
cxp6TKl2gC0gG1RCXdgNgVkGyttM5gRJxXNTgLi2x3GYBpksgTa8TIW4J5UI/zbI
Le9FvT3j0MRT9wy8gBQS+US1GNCWLikLHKpLrC9tfLI7Hzx45tnfWTn1KCi/2oSD
QlebYgAuTopffxHdFQ7Fbz95ZGVCwMCtCNoLzmZoPua6EG0J1/IFMHMPAmepWASH
DLT0X+5KXkBrhM4xDeyXd5aSXgkjMNAMAxvcP6/xHkNAQu5vRn3DHnFAGIOA7Z4c
lnRH+hAGS6KQ9lPbG5vdKfXUAMLa2SVRjlLLaUe6WB5Xx6On4G+piXyAYJr3rK1y
6kL2JihORMWFsIpeuj4sobByNRVr0NUfibpHCM8jXMen7PImo02k2NmaMIuEAuj+
O7dgXxUXWUAhvLTXsPkwTc+lrjEZzpnnSBgKaC7C3rzrijUmgK4TlFlIfjsues5s
H+fFQ3ZI2HehfCN8nXkq+43u0T3xt8SizpBM4+PDD9BQzWLXqTl3f2FniAoMdL4i
yIlD3wLzlifztbaOC+ESyrG2s2BhQ/YPAITDfHJXQ3++tE31xFvXiNwt2W8zmYKU
aAduwJBC+e6UhILd4pku2IQvB9pS4Mv5A21jOLomGnJC+K/tL01CRH0MGwKjw3tM
m3Rrn7j/Z0scqsLaSbyQvR7XIsBy85ZqIkl3/MH0mAAONw2dkx8SKGHV9XR7jHEy
6ehmtJAK3kMZVBDq++356rWyaXiRpwdS/XybLJ84943tjEHn2jhMBM6ooo3Ltj/d
CQIOcUGwXnxabnB/Uo3Wsws+BbgfEF0ClLXy3ZvguyFxV/hk9jvnlbUnRa7G3oUU
DPiKeqwWTmmBZeNYTLZs4VX0gZoKLFX9Y91UaF/Uw9DsGU95lm4CDKeBgB0Mcxox
rZgHvTqWQGcFNaUru1TLGmHjjbA6qSWQs2wzmjDZ3Uanl6CSbCKk1MdGisoZyHOi
397o51JlKp8fxtnDCVAJ4lLnv/ivRXA0tLfqb7aleQsYO0PewNqtOm/fzRcecTXL
whdBR93f5WDQj+PTL4HsB+JqqCTSYZhzwWPiG5vvMTSU1rdETtK7mxxRN2536fUx
zoekHcP+mYP/rANx3CFyBkdYfALYOEITwI0ueNHBIfEX1/OwEENGP+MRG034oKD0
vJpQiffkSFjlR0wAskgAm58jgTHIuMSnu9/Lq/VEQr1OVKnQ9io2THZu1THvRsIY
spm4UG5Uj9Y2dsbfO5LgkwbIlbOthl0/x2hMvemsiYaYsUcuigRo1l90xRS8Sne6
SYpaddovSTnlJ/XewMuZk/c8VXD2b2uvNTJMGnaAdRTOo0HWlJfYn3ZfXprTH1yX
0f2VzYtWnSv/nxcFkNh+W7SaPDNu8GblXUatjXR7rYyL7TICIBpLcqa3SLLBTDde
tUXfU7scgbE67LC8Xmh5THP1Iunlxv9uRtlvrQl7cElTo43CrgLyuTW1BQMt3Bts
FDaej0ttU5QxvWqRD0OksitJ+4yvJsC+MAdCx+8+zVi5Lq3+B/XaXyOeJgaHU6Il
XVQDnNZe/amNztzFW43folUVK5UlJ5fRfRN8WimTsLj3gcxeN4xFG29Y7N83iLr9
dLvvyr4djkZqwnBmDoF/6piJrnf7ltfkGti0eUgabw9qaO/Te1atwgHqgTM9facD
dNCCmiiOyBm9jErjl7jVcP9wDhboK2y7E49vZtqxYdmkPlkJpQMHoJ5b9aWV/rpI
ZuVZX9CrXvzthANVuz711x3ppNB54ikIc4RGMnT1TnYSNhoa0U4Ds9r2y3iMZ+ju
McRqQbz2nXcEQGQgQm021QWUf50IiXUQDxwJsy4ZiCH5Ex3DkL58tsTRKx4j5XZh
2VoRorZGMROMKnwxKtPdD6ZzZZ0cYmoog8V0Doq3gsKH2HYNHoxIXkkaCuK1y70s
5gx9miZovANdbCKgph8bCv76mewaCp06U6ysaBv2xgfKVMFlOBzXTUXR4og41+BF
lQ3YDc5OMOCIsFkExdc8qronacUvKoSE3+MSZNzhWUqiacBVU0KksSgpxuh7phjv
8VUOwg4aITkyB0c55tn5PzoWJe3ghzb9K+KJMlIIB+EkuCZPW5saGP2qrZTXQV7I
tXwaMX3lVMF5TvRaq/MtVECyiojKEw9xTww+91LrqpsZzaazVKErbxUoWCqLYhzm
9/l5mzcxZ2kdI6PdaBvZNx/ykNz3Eu3F+rKFzSbLUkSdLT+WyBMq29ehxaTeKu3G
kpJTfSw1Yj+OnaouC2XH/+WefPxoCQLF1uOZtVlXXhGyCC5bPqWg7etgnC58Q2zN
FGPO9I6WSsqzOWX8N27IRVb+cPmx4P8CUFO/lwasN6R4h4nNMfWoa/lpSGe0t9y3
l35oKwAfRZkp2iL15Buy0pxmJdaeisuYqCnWdVryafyncA8+S4GCiGr+adpn3iUF
yPpWisWiapMhsZn3HXgLCRMehwfx32q+pD2FUrvroYZKqTh3A9loVTB1YJbhCE+Q
PEN+3gzCvPCpUh6T96Q/T/GPTJz1Y+k1PhNLPjG7AdOI86FwaoqKeTyZrUf6FNuF
BRnjaVmf9rNOtXFabWv/Juwre83vbewAfbU+O8+M8+JigRR5gNd3NZGBEI1yLyD5
T1Uuxpuz8nmEubFe6MBgquCXmOoG/EYMyTlGrXuOjEyXNuit6SZzonp0ubEiT+yC
JYaUPHdWcNdR1r/zj14erve3Q3yIgfWvXU77kgawAOmepqAr45qU/jBudr9fcnCi
xaJM8pgRlB3aQdSJxVxUUcARIYhDJjob0IbdP1YdqHOpPiqCyN7o+CsW/Ub8JG3L
9Nye79uQ6EvaVYt3GImnZGBvxG1krNVP/l5JJDuJkk6AFIg39tucwWcneR0aAT4B
3hku67nzhWR2CxAsK+OKgNGWyPA42NEH9KQ54HccNHjSVBhoKk9upB1kpHZKTYQG
o4sagF40sabpik3ZOvP54BdVDv7V4ndhTXB2WODBudvBX9OjM7W7Y0Xm6ScEIXjl
Yzf5vYpQD9iStqQYSHzoebF5TETPhbrbkqe38tp/NbfLmkf0+lppjSbxLdvs/p4g
kSN9MNkPVNZGXkZLyHN5b1zdsuaqWgC7dzqbIjeOMned6VkKUCpq3JG8lOgsLMc8
kSErwRR7YIAAlryEb1hQsJCbGhP9CzHRA7k+NUI7M7v9DhH3WnyGSYXqEEgseWud
MUWfumg6uT6DUvyN0DBu9YoRcJeLLBrfhcSg0PdPrIQRV2Xp1qukgiGfB4N9fqDI
pBQm6/jtSzRJxo2h2pFIbSd4JWQP8G1F45jq8PDFAXADbc1Y4VnLNdU7hcOeilIY
HV9Rbzslc2ePW7KQtuJ498QzdeBcGHlKgJM0rQk4GAn5/ZPYysaVpIpeaOHrErRN
5fzXHnxxq2HqexjH9ro3QV6Xx4jlm+FtKo0n8CSdtYu4HHnG5TJPQDEQ47+ZBsdH
F7iM9IKHCrUHzvWM4LV6SSy0R471nedFHDkES8smZz7ftzOqkmzPBetdptNpIQeO
HrYSo4q0N3qXidwD5ROZHdLdnMQlf5122sdz5WPV5FqD5UcQf137sWxVm0Sok6/5
CM0BxoshvLPm1Or9nnLcGIyZ4esmCa+S3HsSqE0HaiV85jXtVLMmZFzGXK9+lI8Y
HPJA8mChSOMLpt85SsF+Mk4or7uri/YT8x7mYpWEsYkPAisu22ouFbC8pNl9aWzB
gsunrdesKcXHcSgoijUygcpDogidRujfUawctNX86NiX0AhufHppbROutBQDg9J5
AAkPO4AiJk1nQQt9hlZIMAKzS6qLsm1VivKlkFSq9mjsIRMJEnGu7RXACMJTxM1F
Uf73ScD/4O2yg+2dA3/FYvgXZnglfBVZkis7kXytb3a6xbyu0iiwQbwbsJqC2rLB
j2AgnPM+YVzc6bjVFNnZ6NbtpI4kzjEeRYj73989PYnz6xl84PHHpfdolMT/8/6d
yHoVQx0s2a3ltUXVSBInOUtwCZ0fCePRdQXYXqCOnTRWIgP7+bKDEp7ymHXmxCrA
FIk/6aMmA2yhycntDxrONCJKUfZ51UuAU+mEJTChbCz068axTijj2HHzUpa+wiI6
FD4whrQPzzzUHMUrRop/P/fF2QBRyTCcihsNof4Sw19NRnD0itdnFiUN8ZTRhi5d
Y5M6hkxX87ki+k4FRej7lrlx23c0Fowkz9KgFS85Tex5yUAsrE2BvhVIeYxYjcbi
B+Azohi5Io0PdH9WZmkkwsVyrWOEp+IAFmtOeIE4/+sUl4KwHMe1ejk3QDPIphi/
H0VFeeSZebtEfstl5Pyq+VlMFL1EJFijqkRnJdPyyGvcXqCFtcoyq5j10tOivbqn
euNGrt8Tm9u0XoBF354N/mf8fYTNMjmXflvuA/BrGSuEqO/y+e/orpAbfXZKrOnz
Cn1ZHTpn6dUJb/RPq4Yeo+gNzab2qCXNumRKGFx6g6G0qK0Jzj0SjAJZdUMk1erO
7HO3+XcbXZEYDopPQsmh/69wh3wqZtXYgDiAiCdjP3SOBfKmWHdkvUgF1b3c5LBC
FSC9HwhnEgtoTxCMtnJZvVP1c95SbGOhjSRv1TJIsA4C53KYRSXk5HSyuWsYffCi
bL6pvPtgmOn3pIs4AylgKQd3q9aLkXu5aN23pXIuP0NAua0tMlbHgd0lgJYsfzJc
t45k9KeY8zrqb6xn3PHv+5MEgeqJAV4w2w5WqXWLDm3DkZP/ySt7stOUneMqnTlo
FV95g1i3+zSTa7+xfmELPhAJ8Jokqy5+4IGJPBsVqQ9xOuMTwNStLI8rbwZtv8Su
3PZ591qJm9dH3nR+P4CTlhkRJSgg9iVETfnsO2yfAfCOT9pCFm/XxKruL+1PRP4e
24ePN/SLSvtrY3LLJfTr5tt9jfV0cjfPNYLrocQpOtAboxHHQlQB7nzh51X8by8o
p4sTyUxPOf/mDHIsgUMRVjlancqutPbm0dHqSWpJO4dLhEt4KqM1aQBfjcB6LbGx
+2HpvqZ9FZMfRDJ6W9xTsgGKNA/3tKbzLASb0NDe1AMU7SHcgEi+Hz4H99EY8jn9
8CXvev6OifLrRqr8vVa1JVJKSsK5Fr9OkjPQJl3F+FOOUi23hzG9cyBT6XVWLUTT
0GoG6fr2W8SPrwI62a3g43bu6yCOMhb9zpFCVpMQBB4PQumC/yWBUF7CyhX+cEq3
+WwHhopbmd5h5gnStRh2XQg19NmqrgA2dexs51rstrGvC8wPckE3hHdVKIPOipyQ
YY2it+9HQ4PueJc/8hrs5OoHgNX7sMTlLvVdcy8uSE1d1ny4U9vnlE22QPwTmtJ0
Bis1iJ2Evh9UJfMO6+jdR5n4nwbUZguSY6TSE7aO+Uu+734S1XoYkk2c2Q4g3KL+
Lz/oqK+q8gfP01EuoMuhvyxOCQTD8lGHhCg0yvBLXUScQjYfZBZYMIyOlSHf0hCz
E2J3NQQcLIrS6aoJSFw/XLl5tvrKgmqOjlbHsC4RornmcaKzGwDfOWGuNkZN8xE7
oy/f2LKyt7dJWwt9mB19PkBd8cRf7un2y+Liyau9ywTaaMwOMwn1vcE9/Q2eQ8TJ
7sVO599Y5NuMVW2Nh2C+uKyn5uacRnEYufx0neH3OpqqsXkdHgvSpOhMH5BawbGP
iLaJO8o0ww44SxJxKLKbA/U+uLyyNwqkkPzwedqfTNRI1jj+FpQLiqGSdUR4/GPk
+/ta1FNmJiNtja+S1kH1nMyfC9c8SAJRBxKvvCtu6ZYf42Gm7489QIUFOIeM/gnj
2NmlnDfICjMbT/MEL9z5UwK2RCOD5YqC70qSaGBuNToZNtCMn6VNBR/swhr00ES7
s+/Tgubt2Jy26+M0KiIjrmdcMJK8GRqXz1KfPynlCuBGg5Y4sVIwQ/PbVzId6327
Hi2ldpZE4CdzHT8Rn83k6fdvxsmyp0a8e/zEoTZHBq+as+8vdQgGAchXRkaXAO/n
n4Y7Z7LgEUK8dDy2MXiaEKa/ZJg3Ue9lDJHwtyyiikPKTFg8gLSVPxhf4SJAi4DW
aQGzAvOp4Q6T1vOS5Uwd8h0Qs5qM4CrIri8rZ2A3aVUMcacTC4KdMqk0OYej44dJ
uqnYJyawl0aYOhBqNJLkW47ZdS+zqih3VeLHurS4zHdAPxrqKJIoJZvhvRcZMdg8
tMjA23r0ShAWYoSKy6SYkPVv+PPgu5EE2UmAPmWJnPFjj3/ny5m+BnDhEJFw6EWJ
YCB7ytbYGW/afhcLRyh0MVhINTZHNG/ootbKio917PEmOHkcrH5Fwh6FX0CmTzWA
1ys48l/HqHfQq6ih8Nyqev3zoQS1gR53ISlD9L1izC72iTS2M6TDSFCapKHELsTh
nUj2+r3PZTzcV/e3F2bjz7j62FvhcKpkTw5vdQco8miCoo2cfGRtoNg+8xFFsHlx
/JKQCBJ5XYwJkza5bDXq4IAxCLDODfp4kHMm6+Pzi4447mREDIpOhKGVf2BXnwz/
bmtS4xIebD6oswi6FqfbJmbL+MQUJF7kh55Ga5+qcdC0asp1TC74yo2UzF5kJNh2
3syINJ72S1vWobrQtrRiEMp5SW3BfegH0JlT1Hz8ZmxQTaTxmri7IW49caWapwvI
5AeoILM1ctVJph5GJe+RD4tG3J3VT4QyJwOLybubaYYaLVYHY/DgrLvYzwwT9ja2
+Ar4rXDjJluoeovRzoJgFZoL2PUCVn11p4yT/WqTPAaFOrTMhpgrJQ7YXGA8wVhF
bV1+jGKjl737XDJafg8g6uJxXyNXW8e2QXqOVMabO1LXz1l5bNBcleGRBkGeIhF1
b7qTAwRZgpwCn5uwbFJlQc1BUwjCb/yt5/rPOirz0N7NV8bYhRsmPxst7Zx6lnwJ
PKb2VHBCl46DtIA05xq5PP9ehzuSfk+oBB/yVG+q+L0fIEBRK+xdmf2dAVYkf/4d
tsu8iRwTqSceNu4Dr87HgY6At5t3w2/g7qRQK/AdlVI17CO6/bCVURJffXFug9Lx
rPo3Ri0BFNBeNvmXkip78a7crspf8BDvtG/gH8bDFsUYn98Y1tvAXf6nCbLZmUBm
ztrCfBWs5R2Se4uLR6aZ3vK/qhl2iUTqaOfp32wJSD7J0h+3+00MmCQCUDUQ6Eck
FBYM9vuleo0UZABHsTW/aPLkon8W0pVVu6Qva1PhaLQ9S+Nwphd7voB+nWX+42ZT
O/fPPL3ttN9ctbEdKx4WWiLhEzoJipMI9iCoVf81a7C5zXk7Z1Ps6IkvIbX03IWn
5XRP5UDrzwVGX+LPcVV8ptYBXWbE7CGlfFwVrTsLjWRVMYs58q7l+R754XzpByth
oUX4+L21V4CkphYE26jwbp0EwUpjR3GE5xr6H+JzqzU8QfB2xvlvh1nPWMs91ZNq
pXNiVJyc7DA1/cLl6RajuCNZMqbsMrK6nEjtS6qQgA3i8b6PVYSTxMWUPdEFoeTT
ABmbl36U76KoesWPvrfTDmdGN9ZYh1kJYrvwoFdv0VbeU7sgV1FziL6wSn+b9qIW
cdICvDCJQOne9Y9mSPNJrOIVGwuf/fPcDr1rgo/52taxmaL782SmgrxH1T2Cg0Dv
s6M2vJUKko4sCNF/Z6TjT7BpMDElRIUS5M/90MxUzwd7BhOYNASrVTJ4Qbqvwakk
V0xaBrfU0ClocMm3Z1YniKLxJXol6/Ca0/ck6Y1xvCxeTafq7MdWOeDOcunHrgzV
Ojqf2/1AS8Q0FCyT1i6DhHF5plB1diw0G+2I4PkC16b1VkPB9/gA46aS7pOyaKG7
1OT4u1D3QilGm49dIl6YA7Zvsr+Xq4EF+k8airjbvprBOoU+Cfkcn1HjQ7B3xhPD
BV2zdUnnPcCqPZ6c/futc9Sry/tpvq6oZ/mXJM4D/Y0XykK2ICtAJb93zzIOZqSK
VTogjD6iRTgsyjjErFkfDeoj28aHU/8blAuJqtGwyTnw4rscDK4WEr7wCOciNdUj
qlgLyIN35cn/7uyxa/VdgKP85VxOgUtFyLPbkCOoVsJjN33YGxBrI6O4P2HuNCuU
1WBa87mKkRQSMVM9r0fSeDxuA9ck6AxbvZ+iFJZ0fTYH6dR82SUOc7WKsvTONGkl
HTsF1Qlwbs/J0KTwJggJ8bEZKjT4ZnBhI6yUjY8fsHeEWwBjaQDJoje2ZO310Gig
uCo2hs2g2EwrDMXfUjna7pU7BG2c+O5nhDzm0KLcIfIl2If0vNaeEGc7NO2rTP32
fXP22raDOs8nQ1Hc1YSCmIBpmqWRaCbXoadYJkcLMor/8J/BT3T1U4iTDHOAkik3
Ud9zhs6T5OZV1SEoBaxNvFviyTUL+HhLsQfoQ63R+9UU5FPMX+QrkRwCETE/mCEH
fsd1y5uDoNG5Sx+mRPvJrcekSgCIZN3VJtwe80+X7BumA+AkWQ3ardf/KfPpWChE
rdFaZZ6YxxqQf/Lrlze0UObasukNywjLwWPk5qzqo7qEdedtVlcpIy9QYX+9ERyH
gZgOdenT/0FxAO8lZ6zDbCmQ5dgIUxgMVhTkjZBZQvarm3horXrSP0ZXxEK9VKup
O/ax0+sLUZrUE0l8yvSFNwAYMRdT8FmDFK3bdOQv4dSQ2dyyh/oULPduMcfQZi9O
LkgvXTgeC0/Un9Svu1ySmULn/5gLhNAhwchePXB0wQyItlql4/tZ1z0rGJ6kVrlj
h+TdL5+kF9rB841dH0iG3GvzbOuwlZHwYm8qLaOWTDBcYB9FdEDU6M49SCWUk3Hb
FM7E/beZJxnMNzcCHhJy6LX6xHA4RUbaAXYyTaWrBf+3PB6fq5EYfBnMi+uj/N7i
YpPvzamPZNwsFaxWbU7NcswIuTiufEihlXd37NWlrH7W6KjjnZwR7Nq1OU0mqYGP
D50UHCexAb9mujNt+Rhg7eJq+6v6/8YZXG7p/fRXqEDjZinVrKv0FVt9XpKOKG/6
nrjlN+G+7V8EReO2O0D+Eub14EnmrEHBdrW7Mhy9+mr6mL7320cmVcWTs7QBnYV9
vGSB9qpk+pqr3aoSiFFO9m6+mRocz1orVXw2/oy5baraFbCUNy5175x8QPuggSEL
WgGIm6vNp4A8S4B2ehimD6te2A2POvlYjZt4CTVPend//147QzJQHOk2AX4IT/Bo
JIM3vjKfpxgTMmUjCD27Avc0fE1uJ76LPBX6UOpmygsoi2/EDsUgi7pj9UvUXNkS
HWGXFYmkJzaVnrgkAIeqdcPLdquBosahpz5J6WRBljCuMgUGNRuL1jGXio3HoF4Q
YIGPtzfWxGPX1gsGhd8B8Lq0ny5CF+XyEJLe7N3u+fUMBvw86jcmBH6/ObkoZBDn
ec+KNai9GwxcNoGKfFqLPNZsR61IOOL2c0pp7qMGY3IcNSck8zYbJIBojW64eh+A
g0dvoa3DmWw1IwudeMQO6aKH8x+wxmJuhTzWnO8oSRAbt1pMxBOkiTT4Z5RC71uU
/7PS8luNJ2QQhKXK8SmIRU8AS0bgcZE6NBT+GOjdBeBd12S8VSAvsXtiM2F5zzXY
hXFjY0lW7ai150CXYiZyk9VDK8B8GgH32dGHxb3Pl2QwT8/1EY4ArYbB3QCLfgzs
0HpGfGsxOQkjwhQm62I4uveRp6pDn3fpgmQLWNsvK662VcdSZoWl4m9AHkSTpwOQ
FJJFdhWdsj9rjn9IYkXjT+lQoLmvsko77bngiGkrSQf0azhWuvA5KrmNzRUe7SKw
weCDXSFpFMtjmmYMTS9xxI+ajOr744hCMteA3wp4rAzpR+Bi5WORmzcghsACHfa6
O2mCnUEf1kZ1XXuFTGKEWnirrAAMGt1sbg15mKZYTD4yUweACbYLqT0KeFKIDsf3
PMuUF8WPnp9mlvLal5BCz7xi2SAfcuqTp1tHkKY8Ef7XLFK/xvNzRJakGyqqw1sL
n31zwqWJ+WshVV9nHDU9OAUdn77tU2R/GFIo4mhAVqnUUoRlKfq1/TZo6Lvd4BMf
US8MOugXKFf8wT2tcLOVDx7aGSUjeQ3PvBbGAQMvKjFZbQRI1I9NRiBRn1MhHKJK
1UBSZ2S6ZbsidZP8/0meqH/hRIGb+NIH6KhDJLBCTyr5mxnvwbMt9cYK/zcvopUA
LwZnBokhctgd4nM+cEZLJMOdqnbiZqeaHOjOe5V6s+m9cf6ZxqZNv0DZswl69iCa
CGijeCxO3ooYH9QtOLBjz16UvdiSENHVIa3UVGJhezDmhwkB7CDdCQj9tRTaLOzp
WckJzJ/v5MsCHjYYXJ30L2DHc5/wgZERvQL7UMhZ9zTPJZwpW2A5gwcL5c6x48IF
+xp3EYgJPewpt3g9F9NXwRslj7ZB3kP8fWoF8IDKVtJtXk9/pMmz/bpgotMM5d6+
gXzZUVw3Cd6Rg1JbGlSaIINoxlksqbxKQjpsf0d7z1z6pXzKIyWWdUErK8tSDz7j
yrhIWcr2JEJziC16+ykhO3hkXaxzgEkjMgaCAy+GOnyjMm3z/bXF7Mp6ab00AQOQ
JMRXOLhY8prCAe8Naeu0ORpuTBL2JlPC9i14S+3u5J53XW086LBmI12GHXK43TCP
UDyt4eA20ETW9CPqztPcSINhwjFXrsp84xBaXbfPhTZSUVh+54c4L1E4kwVnWt6j
4MC1G1bPN8VgskEEwQLifjSEwlsM3AYEm21ahc1XG7Y1aMrk+AIB6fD6aKparU3U
jslLyIp2UIxq5gmJMwX1gaxnirLxTRG+eDtazIvYwdToWhIAggDm94aibnI2bBYE
A3ZVN4sz4ZUp0Ilq660X2zt/SahycbSvufKSdRP+pee9SQJSawEReN6uyPnURNkv
NNrKMzJRCYNZcI7hyVk5Hz4chFS7qetCcgqqmo9X+QqFO+O6wANkUDhqp5Xyqn2I
S+lh85n1JmvWQruloLzZTylrFiJaWrebrvqJaz3fMOym2iFKsPexytM+rgdUNLcW
XbBh6JAQrHmG9LDUC7ekadsWrI7NdgGgGU+3RtSODVAZ5Bek+OG9xYpfPYK+WnWb
T9HXLI44MI1QdHEO0PiQrDM/qYqRjE0/MDXI9XKGMI/NHCWElI9TiMU2uIIEArXu
3dbyjisfq1QR21mfWS/t4aH1cQAQ5cemmKJXiFcQkX9oG+BapxGiViJvXwXvPuUU
iJsbedXRgAxLT7t+PHfxZsE7mv2jEmyeOVbmZdZT91UyaUhCRSmX+B0PUyAlofK6
Mv1Imb8t17uhP1BMDjWZOjlmJwaTj4zejFxO9kYJl0rVJvAl2G7zAJDJc260ix8B
DE8p3PAyq+ewo/QSVtZ9SEchxxj57LA+KJEsNxfJsq0TDmNv8za1mSF6Dm0+RC1K
lkgl55BlJuk6+hHg0qJkIFnq2A4vht7CYcdrv8opkO/DWs3oa0JGdJ0rWdpf0Wp/
2z0K8T5H6KtRrI4rc4q9SxaGtSdXKneHRQEtlOMxRkA2g8j9ZDDw6UkOPsMyY2Wd
apQd1dfQbGfu3LiM9i382JjOHd2Hjyj0/WFupN+qFm2lngAoTQxEBEVK35vS+Vlf
MO9uRe/PD1yKH/XekCw5D7nmt1kXrgI/q4HpEUQDSo3wNF6sxk8x/mLfA37nU8qd
PDQg5kiD9TwdqqKmwvn4EPHhdAqB0ukDyILTC2AHRaVE/Ozo7Zu/q0Iw8zt3kkEN
l13U+Kpe2u+hXt246Hle7ffQglkrhKB05g1V9mCOhFhVeHXBqY3cuhOzT4e8VnFZ
hj9pVAW+wpXQGFJuRfhK8n2AGysI4hjP/u7myFUFliHwhv94QkV6SU2pEiSL1htV
VJf2mvvCvTFDk/ea+LaP6YsR//SOohwut8Gr8a/OUnRaFyUyg8UHcHYC/aELH5Wg
uDJM2uZO0TS6ZAF1LnVFjOfBer34c0TM2TGQyv2HB5YD7oCkKLcsro+0BuHZvzqg
Rm5uxmg5x2xYct4b5qfIJhgLdV64cbW9XOFxhnJyhbVczpVPIclFDQox9aso396N
/ngaedRUoj4GM4RvchgPtJv6CkeLnI2a9VnhtLHv4vp8qUvcphb6p2cwtaloWX8D
kWaM9uGyy2atA0Xgk/VLGM3BMl5GPx4CEKPGkdJSWzLNQXm6QQVFweKbHBW9IMH2
jY8bNHsVLLDptgDTt8JKNZGSP2rBwnj9qJNfWIHIC14R72JOq0NWiZ1duR/cnVeC
avD39Jby6t3TGq/UR3836MCEL/jI26V/nznS/AOYLoEOpV2LxQ26+wR8k7Ai2rKa
PRhnvalk/rXqQNuil9hR8+NmiD2jFtEzauCe8qTXG/+WcaUlHi7RBiOXH8c6qs35
VobzlAZjpe6+ZIzsZydB0PpDZr6d1ulDlSXzUIJ1ed/5tMyJNDJCRyEE1Nf59Orc
1JN6N5ulBeXtSDNK6m54XwSk4KrEUdhIMb5LTcW1j9eqnJAacIs1IWcTCLxLfdrU
AUfAnjYB3ePqlrjSudAZe24C1DQMMIaGfZRrIF6qwd85ZEsQY1Xdrdr9WUY9zTnx
j1XXDxEGriid5GKNbckGfcVeigBD91hQPk/J1HzkncHYLOLFmEIj6ISn+tg//Jus
luu6A42QVif1UMy8p2kRr+Nia9PZ5LRfSOHMHr+p/Qj1+YdIxrLfKqjAiY2fgJUF
ie0vRVGvU+o0K433dvvlvYBpAbWhwIcYLuG0AgMA1a7mtuC70Y3tOSWiTn3Wm13r
betQk0+Q81Qk+RDsuWAO6vHOBRPe7K47SQswLoGeR7mG//mL5lDa1uHkghaA/RpJ
USoADOHJhQFZpw1Ktsqhv72wh/W37MKnKzUdmhaqBcPI2Vvg+giik9AwS9vkslzG
0PqwFDVq47q1KMbo1yjLYL5h2SgvPHgQyQGgjft9ReITOeuuMF9iwk+Jbu2jv0Kj
coThhTaFA6R6FtzxFBdGUQQqGsQkkjTIGixUvbZGDQN9Ovqyvy+fIcC1pzT4t2rW
pMwKIfOd0i44VYELgeyCzPD0+Aop4djRsD+Nzr5N7VBtfzSz9MK2QMai+Cek6ztK
lnDzX4+axmwRgag3RVRyHGb4vqhsNiVSszjPdxZIloMVfeR/gYIegWwDwMKFa+Uj
ixsuRxD6pIZQ0bI5Ovm0CBdFtsXW99iU8qBbR6RAHLR3mWCif4KxM+XXu3gtQESu
dENHfkUqA8t+updB1g0mHIytsn8WQW48bDyEV74PaV4FScqeJ19Zat8tSvVUe6v9
IrljHldloE+uWjierrs6Ezkza/9LbopFL89IeuHTyUaRmxnzn6kVQao9gxl0kJNx
/n5cCElJcMZYK0/ztEgB+QTlX9+/qqzSwH1CPKZHk50FzmunnyiBgilNkPxcZ6Pw
1GaGdZS7kr4V/Arn0zSYNHCWoVzkQLxbC2++I496MYmVO6xMbRweY3+TPw8+xpwq
FcUPOYbIENaWrSsFl3xVyVUU3infekDVmNg8NtK5MBeY3p+Hvzn9cG6IuUNOv0qH
maT6LxhCgng0e3lICy1jIRGBAS0NXAXBSFMe1SNxzT5JOuxv9gB6ZOKlURbRWY6b
1l3/s/xrQaBwxCdRHAVmH23/20VELN+xF7dNs+z4c/ODjzhOiC1ENf9/sD6hMQuN
H1OrtgQ4JCFqf4rM5qGDG63PNLeA73VUkv2FEpSOCGQXfqmApa1WKXWk1qAphqfe
G8Nn9wUn1yqQeB8ZLnW33Y7sXskB581GQ/xxneIykZ3nY3AZaeEdE8sC4MDsOUVu
9TPwyYjE3bnCpk/Zet6CndZkQHLjJX9MQUkfNpwDZ04ujOAysKxvmeETAGMm9Lxq
/2lKk19pn5kUv89b11aOHZqsfatoofXW9/2Y92uHYYINafJ2REdkRRnYQH9pDsPh
XNJigFdfwbSveLcNc9p3VSdnOH2+emzxYVjDtLI0Df62osyd+C6oNjB5s6hJEs8Y
zkEXMGdegL14HuAicC7fBRIU1p2uRXEEF8Gei6TguNv4M0wh5CY+hRcA7iQTk2iO
0xqUlDx34xdWczcRRN45RYZLaDYRhDR0dDau5YkL42VLebyAhODDuX0tcKfRVtQ+
/4LUYnaXWgT8/O5nCse+wAUWakcgy10hqZi62Yy+MuLuJgoAZt4jBIWSSZ4BMBZ7
BO8h4c3fN2yog7uzcWpAJHnIzpCMuLzZN14K7pdxpNOMByYs4RpjT09AXbxbNM/K
8xNUP1B5pGlYq3YYllAEDzHMdhIcqhhDq2YCGigoWzje8t6acU/SRaOxb08A7I4h
/WDuSH16lxT+zFVq9hI4RaDPD1PuuLxFKyxjFYA9wJUwxdPCOiiRE7hE7ERYqlZf
eQXWn4oGf7EVmGJpEmOCWjRkyyO9+w6IA2oZ7XMQfC+SWvr2+Pn8s11kfAizeDcK
SLMG4fJbCN8N+2PpocQYeO2dfqwFc/UJ/ZA5KvkaLxutmCQuvwxWMnYIJIOIqpLW
o+fj9KA1zQM5HyfvZD6XUFo3kk4m4DAfT3IrFMlSZPpQbMJRgE+K0ZrW+neu6z0h
Rx0LPh8BVPOLmLxKaeKsbMjJDkmapPPEUpfldYAQXpBqNZxBigdD7bCY7SZhE3UU
Aona7fFTxbZa6wXnHYLxJRmK6wLlVcnjpRv6cqdvN1C54k/+7yif36ReDwWckE4y
kQqTg5mbbQaiguUF13/61bgC2NKLBX19CRMFU5xey+sw9nP3Cecc+o9LxyXeHUqG
xRGYe3X3i7i9M9QWks+kxGv2myimStZqKEM2VQn4dB19YDcgxP/fKQgsSgxt/Fe+
ObJjUhIGDEnao3EC050+7HURz+/CNSF0h7X/vjMmlXB01fA9WOJVpmeazvyPUd2w
FnfRPsGkadejffHgqFbkD6LhjNitynqlyYp+3CP/v9k3e9i7azc7Qk0jHarAxIVP
VvIsqh50JUjLpLgdyOn9m9UtTzg6cf+cxb6NTvNFKHw4PzKp2bOQbSwaC3Ih/3PE
H5FHnaS8P2pGBu2zw9DAttZltFsDjCOdotmXB/xjHKb+k0miuUSNvcbD1upcGioR
FK5UY+nWWx0Ehxwvw4ImsLpgdB5Mc39kyGteIy9nxk/O8k94yUIHDn97HuHcbL5z
y1/lU0M2dwLReV6fCrJ3M+eGvKRtbirkoR7q7MCt9Qr9HU06RqV8k0tPXm87VIGR
MNI2nhP0i5H5ROBtSXC7wmOVEXxnBTh9ajBsn3hmQGRc+aoeB4I8yCjk3vqa4Asg
aZffYpYY/INHS6aI43j8fnU3TBpskYtlI22KLsTb5nFEX5vGq48oI4+UE17ImkRK
gt/wJm7rwcZ4gOfAKw0BAVzYGZPyVShKop0aiPoYYU/GI4hKMBHJGClnaKzB29Av
CH65HHd0FcmNH2bz2rdCEHiVK65himy/mlzcqErKS9zl/PBSMxav1lD5nIVbazpV
JcCAVrqDRoWRuDB+GSJdR9ydP7pBd6ViVQOTA9cKVrpeQcJXuDtEzUod6Lu50osS
uxYzDVNXmffbhLuFRgn+MsIBstYvaN7ngXdcHXdraPAOXYe8W4CfgW1NPhaedhdW
Mi/8kBInnVR92k1I5CGjtdalmrUdXStV3lKehCOCV4ZSWTITtD8Zg2Z7Bg8pnPxd
xiAQwck6tZEiTO7oS72B+hfxUOymGAZ6XlVAvPjLNxBNJ7OW9xoQDZQh7eeYcNB9
5O4iztTOtEdajb1zXyWggATp6U+gwnmvSeLJ30E5IQQs/Sely+fNUxTlqUM6bwGl
7HKe0gGEsAKME0Q3OlgNkzY3o/NWaf6sCJI++pa0RQGsjuE0+XfPnmI2Iqm47ZT5
lN34AWm2lGC/5/i2sVoekmPX9mMR755H310CTB2mZHkyejWB9//fulw0Q1LzPVTS
M5cl07xOUrGZYea1Qp4ZodcKl8mogfFLmnHw6eVZxy+b8E2CzOd2etwZPPz8kp5p
K4YIfHel9YYc4G3YlJIex4zcD/swI/p249yyVrAWNLqK3JvdXiQSkXulXMWQZBnw
Ok9hpAkwHtfIXdoA7yR2ypvbmeIrCTcqnUa1kmmWMG54dLKOEn8QHAeOtr+dMg5n
xmRDfh4gGjPgtmvcOBs5Brd5mOZTzYso/LU8JdE/fmXA5Y4NiesyNgS5VWc4REd/
RQRjzioYQPq0IHO2myMVaAL2WVE9JZalDpygJxVYQjRQl62Qk7KkdqCnTJ32CXs1
yBSgCRl9UDtViRfPyHod7wL423MXqCLKoGnmMi7P4npH3ldnHCzRyk3H91Fey0Yp
i69drveZfbSHtI7Nvcvhz1LBlgFhuHVZ+d4JyQAb3SKjQF4KAJvylgtELDpKyHqm
eAXJAiK/teCwdlsot0lApNdeZJU4KwpVzMGhs/Rcw3vtyzNUKGXaLHo1KE9BTn6v
hlFTMFV4KTOjSPwugP/SjjSQtgFEjX1FbsHic/e7LWQ7RL+s1hnsPPe7XLxMS3nz
9NfutktfMQKQCoDW+Fc/53EJIAYMXNaWNZ4xnBk6rxNrmBZPw+gg/XX4my2cHYIh
R7bOJqL/jylO/QOHFnXretB3n847tYWMgCK/4qE4xAJPbXMsklhAxTj+agIOYf3O
ckRw4yGn+Aa7kItPSESOO2Pcf9pxICoxjmBopG2OB/6TY1Q2o1iZ+EE4MR79xHND
ixgfX1zZdREQ9HHsO9qGHR5hLRvutrKk+kf0NadwBYo/vA5HGGIxVbgpJzFz0XY0
1xoN0Y7j1IQztCPzN0xsvrIgGjv7rS0TdrT/zSgeMSRCUCOM4fQ7IB5XjVGqZ+SJ
W58braj1KTqT7jO32jBwXHjjHXibiml0PqZ4BY9bj05/KR0igagoZdFF/R9W42G5
pSr3//FeDXmq/Oi0oRUwEQSPtpd91ukv7HXUuK3lI567DRRqoJCro6vpU49ZH4Cj
kFtJiaka1PHiZah2WNyj5xH34OWwnMhyQbAbYS6tGhdNuye/nUJPfBY3lX+BxTdh
QiV57E8wMmIQD29Ks3WHqYakPQnZYsylgVncgvWR5eXsRZllVyPt7k1lZE4xlwq/
/nIFOybXOCidxrZ0n7deywDx74KQ3FHJk0qLu5U9tuuqhc5Ll00aD5FkO0dHJV7n
HObdvkVyDnef3K9En7IdF46Wh7XXgAmC4aWRIqgBZr+hBTc5/TTMKmRBK+v/jsC0
MtHyBCFsSbJ0o+2MXo518Fsb47CaQNqaQac6x6gqDv5rRi7LRDYG6TrppSYfZh1A
EQ7l0xyhk8k7kIgpB/3z7rfdIoC+C2GpE9mQgITjlF0oB+2o1KjP3DswPTM82Q93
pKvSwbcttQP4UejmsbH18I93e/ZtaScHcdJtWSj+2oCFJfAynrMpdEY3Jv+e0Otm
/3sgeimi0BogBmDN4b8fZiXKwzgvz7CL0fZyUT/WXVg+/LK25KIAFGw8/syqCzrM
yUsvgKtvNJ1Fk7hr+DTaAZpIiSsdYQr8dJ4+9Z946AHdihcajmwse+CBhbKpFStL
N+sgdcNbr3EII7/9LnzSA64dY32kQt8/AHp++7d402FaI3bHscX6nsacMA13pPzK
9Y/unGMLHFGxjiUDPGMnPdLOZ9V7y7qz4pdUTHrcnqJFu7g/FFDQHLAifg8uS9Lp
YGm+2MxacE0OgztYfDo3cZ/lZPZh85SgjPrKxDcfTvUub5hEaWX2oTGRTDAZvaEL
hA2V7dAHuii22lJ5+pHIYBg/r+A0f734mTNulm2ceUVq7L1ruFP3r+ZmBvEmauV/
jy5IKCYiYa1g7Q5gZ383n/EmWKt+wj7Y4pECoV2GDquZNDKHOhn9R9771v8hPynS
+osRG0i57UT4/VZEqA2KJ5jCQGSSBI7Bievj4Zcj+lxUgd7nwVLr7CzXm18YwLEA
XpAg3USDeSm28jNe8mQ21EicjdB+6IZfNqpHhZeUIFMsoouMsqxLwJ0e/glfmVnJ
7zSYXjUIsKLdK5xqLXDDDi1Ts/gMDQzMpqrMINdqp2pBlvqqHTEwX27ti1c77cAh
T0ziSz8hsU/m72c/3bDpc76xmRNOm10vDpAkmgfPJNGVFYwhrZsHm2RhaRBEYftT
z3qq7gp7SPbuS/Tm/CadKoC85Tj0CiDb4HyLgEywkkFjpZxXLbYqcHmnhTaIiwhY
Fqh/DD5U/cYyA3LKTqTKS6fHkwcNzvNV7Y3Cb8/kMAJLV4DBOrKGHLWbiK7BQJS8
tCeTjUQkTS/HrACSPMNd9o4DBSIFL86uL/8hXbdbfjfvcdDZXq/bPLNZ5rkBGPmt
GLbYh7OmAwLUF2P8kmJ8jlBm7v18bxNTGJhdFD/N+pWoCgqw87A6ql/LeqJZbOGS
U38PHg+We9LH4gZZZmz9W1kVzMErMjEvykyLO7OI67M31349QKTd+E27VXcsUyIk
lixsYM/EFjXpath7mb0v28PEGGifFld3CDgSO5ZYiZgPMi21zn5zpcqSoVTQKIck
cYnXxc63VmAzEMb/X1/QB63yPxwg1QUAP102th/EQU8LXO5mgUrEyQ2GILhNker7
Lln1HTnCom7BVLAVcDLOTHQ9ZtbJ5K1mXcB4teBnCxpsiSYVi5Fmf4iqwmS+Vk7I
XD4BqiFgdONlpPO3MSNztDard7fqSk+Xb1e7IpJJP6cH0QV51nL055Mr3+PtFJti
0HCCykmXgodXgKEHe2xbhVCH+2cRRm214n40NxMmRdLJnINvtTjQoXzXleF/u2EZ
GzjzBZQ+2ShvZKXYX1njkKg02QCiBEK7iP6+jpfDcLJjoo9JE4qQSlHWT2G1EHwL
H41QbCCJJg8XZZVNwg2zLGBfQgrDmRjJ5RJ9ZHPLxKL6aW9EA5aUZPR1Gyl4XxN/
VfLdF6evbrlHSKcKQtBNBNhFPO1x8wp5d0xoRP+aaJ/SQPyZpzM2qHF7KPpyKJk4
yaAVeVlziidITsEJcVC8b9CezcH4MgQieZVXG1XGVwUgDrqZIW002YtQFKSim+Z6
8IRlbFMKdpCP2k2uAJ4qlzSmpTpH3TPLenz7dzlSHXv6057kmS8C2zOSd7+gT3KK
oZTNr87OfK1wHTNMBm0Q3bVFEcOjc1p7Bqd6Gi8bjcdMyeKZyG5WcYhQSEmv8oXc
yR9wN9q6TTmEiKTrU5IJAo74JWhDO+N+jdOgvtLg6+l2KBfsSAJ+ApkcavpSsILh
W/I92WZ4qrwGvq88BH1ViKDS271th1pzct549LNpDLl0Ts0quLIU5t3ntvzndlQF
6qZx+YWQ0wT3YODzKzbHmB/5hMxNVEJ1ODHpKmieXR8vNayrb4Au7Z/fX+6GQcVp
HrImvok8vfORppy9DUST54BNGDZcsPhmh2Nuh9r/Ve2sMvQwn3cEUf0eAe/0Pt2Q
FnPYLDmuOcBVwQmU0/SycOaAgsHQVHd/hOziiKoRu4BjgYtmmAnwopBS4q5Xkyji
O3MjHrQaDCLQqF0T07jHeppHOiw43U5JTG9q41BxqCFlAggSQKcEKbeHgMFSRgU1
7pLuH/Z50eoK870PHxzc4dqgK852JHVlaVlaNMdWvjUL9DGIaRe5PMRQUOXjUYag
JTUb/jBoBrdZB2igDFv8vKF9KtDY9/Eu6BRgAd0RvvOVyOlvMl9jhmFdKqdC9t5Y
KjowQjQnhqX3i/+2b4jG6FTr5mthROsQ6KP81dxgz6LUKteNo3tAHNO++py8fQwb
9iipR4+bmjjTPInCf9P0lc1aMakpKi1e6QUS3KCdOLZ1Qf3ktI6bl2BXN0uGT7H+
t+OXzP9FhEbplwvL5FIeSMVRXJlxBh0JtKNfmal8tMQ9AYu2Son94X+hf/PQ3D9d
wonVip6TTT038bW5Ftoad1x+DgqqO0KnsJnfRPAh1Ac782EbUn7I4rLC9gpm9A3b
JFhTnSivsAFk6laMqwSsLSftgPXaqIpYjig39u37wF3njIreLVaWDFG2XnsiAAy+
kYH27F2d4lBtiVRdBTFFh/Wy9gGKTsa0pZyQ1v5dSUCDjSlJG8cA+D6q4zU5Z/5R
B5OU3iio0mjy8xJpAr0N/wUxOn5fBJB05zKZQfJcvAu3QleEH6ttIrTyK0UhX0Pd
fFuXPNzuddEnQkBzc6ni1SChIWaNtcHN1MDLqaTgAZjp0ZydmhKGH33VYQUliP6r
gmgQRaGaRROhX48qgPmYKU5k3wClD/Vgu9rzOxKvAgEizpsnAJ+rx+zPj7TOLmoV
DH5WYlN3fUuxfZdxhF9cH9Wzhlv5HAhLylC9ppNBQ1ghtEoMwQncv7L4H5zr6Qcd
HJSgrEXrbygZ51gvLz4j/uMN3blevU6gEAJ92DFWUKxfCG+nIQ+LCh/c/2ZlRt7A
aMiz9pWcMTdLSPXOX7GhKXD3tcYi67whqBri/vdTgpUBKfvRJot5NH6pQ7L6uYws
v2fJ2a/DwOpB4lBKvzzbsk+R05VksrredU80SN8pRWSlqBnVmHyzWBkwB4rrtX41
sUvTXdhNZCmv7Mrx+zsk4+LRzf2sbTSIlBPGEX81SS+x4zUe0uz/ygP8Hl2XH3tj
KKWHmZZ98bOjSWTAGEHLih7YF+ewNGhNdX19IcYyxVcSwGcAnm8pzWw+T/r18zeq
gzqu/kkq0UQnqpHHxVSeq+cCTKcqKSpRhRM5AMOJu+1r751gJHMAMEMZ4VdCTCwV
W3bTRtgGAEMgy2rKip5lylhYu/uze8ol6vbZZPxqdd1+DaYVpbQHhSrrkBMQkivP
fxPD8mm7OUM//BRExq/bVgODg8Dr9+V6HlEdLhwaZnmNDyslKYrwqkql0dIea5xo
89g61qvLHJOhRvHF5VAnWqOzGS7ZjEy98HliYvSt6n9utQ/zEOuYX8F2mzFYlcHP
Xp69/fW7PwhXUhTWRVUS7iWyyhYEV1hKLEG2odKY50O8eVmmi648sURwIcDNfzum
bW7NlWG+pNgBWzK7YB8MexZ0vZAOMPUZFuAlL75J3pfY9c0yfqGTWjHzS6wOS4ev
BTjYedPHvK/8PQaWz/KddtiMaWE0FtagGeA3pnLt0AwZOFj8viFRIfbYsKxjWcT/
0JoRKb6lMgWht3CN+Ou7IBYODd1hU8N5ziahwUaNLQUpYHJ7j0hM+al0UwOng5FD
Zl+RvARR2Bfwu+qzr2HGfJG2zc41xfZjsKHkWgQQEaB4xjAygw0Rsu89E1/IBxo1
cv1j72ExHuj8I8SVBHLU59rSPZttp3eHqw1SlZpaiBOLz90XkC9mvK1aHvJ9Z68s
DYnfa6Lu3VZaZQG03wT8hY3U979Spnr14QDV6YTs4WnP+oLvrZQluXNdMNQ+Zjk6
8h7fnk6EZ8dYv6V3fi+SUkqjBQGzN+FOJ0y89JB2wRv63iZhTeMAaW4rrzvmwK63
PRnJxqWE32tQPk65RcJfdQFIQ1bSgFQC+cdOPAb7rgSsz8fJBSPTY35YMLhn490X
nJmzGthJi7AIwL1X0sp460yLBbV3/N00XX+2QlqPHWVH3TgIP/G95Su80lyk6yXn
1VChrcQ9xEZFpqeCNcG97/rGkLadI92Q+1F+jIRJtf+vW0nNSR6+juXm/EViBdZI
V1P2suVNrzGX4SW0naXiMsWiSWZaLfZ6X8SJIakuZtUOvdtcsViFcL6WkIE8CHpP
QVWOu+ScFb7wyYr9kBK3AV5hDNCF+Q36eeVkQjQGRsXd2EhC5O1UyLxB1FgBJUsZ
NlxSrZ5IKV7uWszNER39wb0132PQwVZ+2M04bXfbwj4+/9Mbi2HHeJBrsc3w1V+f
u5WvVuzh8vhUHna09Lj+YQscSdp0Qdu90aExVBBlH33ArSo+fNiWsOGJSlawjssO
OmGrHEf1ctBDKGCgYub03aIAL2s2L0pGLNdRubefUDXY5PY3YOmOfxNJ4VyM5BnS
T37tM1iF4jnCBym9mW9PgOlfImJ3xD4uEeNZTEQ/7fG39AW6JrmKy7DskIk4XsJu
cjb/LlBSFdxaizh6YD0pBWx2zbp0Nr9s28cZUIUhIN1mMyqn6Gb2V3sXw/pukPtK
J/g6PKpBWrDMjlBWDzUAIgO9bbdPczsPuziE4efysH2s67bwVEF1MO58dCXPJtQB
CdVvF9iBcJUA9hwbjm632Esi7Qy5W9gs0RS0m7z6q91WcMfRqN6YFlCgSy9BgAb/
PvuWJAdYrZdM0N1oOVrThhtyoD9mqzD9bX/2RDSx2674VVdrB4snvDqFbTy6muCg
9T8qymJYeEaYCdTch4B01oJLTCuc+T4/+sx4IiKd3J7i7cKmGqv3LA0GeGSUbPKa
pEZDkrhANUclMVja/iGhuWjeICU9FTjBmBttZI/FNNZcnff1s5gch506lceyZijd
15vS/6ZbrxP3gBMkSE4olTCWovF/ByeOnkYnia92k2vgx7z5kEpVkRW5MDjs2Ls+
TzKRHF1BxhoCj1tCWAKUaQyKh7gIjntyll936F9wlJ9oTUt7vt1RBsfducPTgTU2
W5kA0cV+/HRnhIBLqTubZkyazkkzvjFd9zUlW286UmWowDoBzLCFFq4p/L0tQWc/
AgMbbCuLbacdhGep3Bz6NOqo1UxUNs4g0U7AwUy2bgYBHAAs9go0B3+fA+EyDDd+
MDsvdehbOYJ9Ox6YdOB5UAIGJK+06ECMBoTPZ8msxOHxtY5BjnV5XUhSJMS7YNC/
i0Yn3QPlyI8Gw/Nu98T/FDCshXL44kKRXrwgbEN8tfyU9p2uoR2qGAYiTVeVHG8H
t4KUA60OKd3nxUpocGHyz0m8wQKBeF+J0sNoyLa4d6ekLOJ73lAfOtVEChKsQXjX
RANI77MwVPZZRuBntYWSY/XVEhWsYBYIQy+uMGhB2w9zKDj5aqntfCEYmBF97MtL
Zk0JYkOiiEvq0qSme7B3+2WALQUF8ScF9GqdkpzT/O2dn91eKhaEJR7R4sIzeA0u
trxFIX5ezNL1qJBKhdZTouRdnGa9y5yaxcR4PmNNDNeclSt6bviV32hFJO1QpU/T
luINIKxMXu9hjXKGJWIv38AraB6TD4kEUbc3p5koJrTt1+OQoHkQEpIlt2ue0QPS
ikXjCfH7XWrvDFyK4LtUzRvN4bAFNUzkBxSTEZFkb6m/GGFsJIRjH10TO2ObHWLc
L4ACvB2qYqXRG525U1kNulhQX6umNPJoYsJCAUUPXsdgSAr9CAbVmK3rR6IcX6j6
RrOlMvKcYMkKbeept/IRy5kq3TzIaRoejbt843K9xBCLvbbOCzs9m+Y2z26shy4y
RyU8zboGAFEPw9NjvAnpAMgoTOxQW2MWRw5VyTWlDBJDpDmCzqxXgPalcl+EW1fq
epghyDNJnhmt9e83yunB/tcpGUrzMhD1gT2Lwlo+dMbgB/WKmxEvCM80coziOCg1
u2Ue+92DP2eZRC0zt+0JNiVUaFwvCWwM1lB/i5oLiFLxekkosG4kkfgf4pCC8H1P
aAzCImUErkpIZE6IU0WkostU520jg4SaXGEkKe0XijF240/OLnEWRNwH5e3Esc3w
+GOr2cSx1mdL+G5JbsyTyLNOnXaiUOw/lvdIK/yte+AB3Z5C+9IaVISojN4wrSYU
RL7o8IwqL1SyAW7GAPXY8Sh8Cpysb43ktDbAuL0sVaALx4pUy/oGLFA4LTahLvT5
IVutFusPCP/rtgKiywrddhIaKx8ZCJ4VSt/hFNoPBToTSPS6Pl2nVmYmi/Arqe9D
23ZxejjuutthIonCwR19TLjgQLPpJ1JmpuRpWIjtGnU6pk7mBexSLazsbb0BnOY0
yVxv3JcWpeFOgeIuwXF4tk3LxcaKlja99n3fmKVk28WZgFmaxbkyR4CjEWSwOT6o
IbPAEdrmPLSTrZ/yWtxgu+yyTWuiQ9MMlqQRzdQJ0NU5hdwL1R4tq/M6L7Nf/xc+
Dh7+ZmFvC6Lm+VOHl5vufd6xoBZ5t7IrpS15OLJvkbnhnHgo+mm+mfYwdbo5h8OM
qrr5kuRPN+Nsz63XZqRgWMQLDLjrfSAYbfo0h5qv/qayAd06zMGe29OmvbZTdaoV
gGp7Z89D8KGQ0KOxzhRvkyPRYXOGZxT4n4h+sixDllJ7FNgXw7u3yhIRGcXX/gEx
oKy5jBArNQa5qfPhiRbFhE22Xauc4Fclam+Wyrtr0r3Nf7cHZcj8OHgQvGw+wDmS
51CqOqjpoDwRS4OoP+qPdn0NmS7eGehxMT0WOIxa7UjUMU+6ON0A7lw3wcVD6RJS
+hoa6p8ILm7PcDGj/ah6JGyTy0dYvakvzW0bnC7uFG8qevyzfkcaFggQ+sJSLYva
qItO35MNClFy+1D/H2THFlhH6Z40j9JgLhPJbUT278nBKVNJKe5i22j9nx12eqKc
lvLmo27VU9g0T8PFbODTaYeIqqi4KRcSwc7o8Qtidd8VM6Vr8hXZaeK6dAUqec7B
44XFXxzAcpYwLYDD7NxSChSqdz+3/gTapnwPsUhZfhoxad4JPDQgmOFNFqrNr3oz
fwcPEn++GBJVUbXYBf/vnjJq0COOkgwJaESRwnIbs8Kx4GxVFDhQoOreuKe8BqXZ
PWANXQtrmKZ9IK2VEFQTjJKvVcfQx8+JH9M7XCFAexQrK06uk52ZbF2ky/8ZGKvr
MbV4NuUaCKPMEnPWL/DTuj8z7jCRgY5Ys7f91S2YSzkDSJkC70i38Vu+n39NjfPw
v5Zts41Wi7qZOQ1CvTHXSFkehZuYJclero4No6kCWlNWUL02YLbyw3rUFBzXHWJn
JbOSprpXprctASpI9mdd6DRq7NEoYMWU/96w56HfT4SuTDM7G7r/JBe+h1EVeZyZ
7zB86tR+l1TbJ7QQhp7RFdNT6vKWwllwfiwN6WwJUY2GttU38RBJCeCS4HXt5n/1
Q9HRJl1x9OQ+yb18xha12cyShgJwa6S+ypkWr9Oh31MgdPEPVuqp7N4HfZoKErYy
niRfzVRkZauiOxu9YrR5Nziogh9c3DU3bFWRckn2iezTh7eLadpnhb6MKn4sINJt
W5pi2Qz/0L+K4lBL7AaEC7mkaM2DUmqJWQk0ELQkQ1m7WF0ZNUhBoCXCoSh1Wy/D
8XaSRjkLY5UuEVke0hAN1LtlyLwmqliOOLAP9CE+rNhV3/KMucd3aCwMlevexhRA
L7j2Mf46ZHesgxi4z9YmNm3k1Wja2+JGU5TZe0hVcCIxQvSXaT+gjGkdCv2fHaE4
lNDhmJt/APMhnIwmgBQvt2UtpTn6LzPwoK2qRmGa5WkrUXpgPQXE3AY9fQlgGZ0z
TldSOFQkMtxywofgnVlpN+zxAomReb7rXFF5eT8XdqysAChSVwTEjzLoZnWLDSaG
eJdzj1EqGpDoj/WRmEG/VASZFe7YpzRyzQNOBlF/jfViGHL3kfkTu3QlAnk3Tv8i
gZJngeR8SNFpmPTpSlxSMIXtaoH3tLewu28KZ0cQYonSI1eJXijCPHWav8KpnJfh
p46NVkatLtki6P136gQBYbXiz6iuYkiyHsiQWLEe8j8U0ObSGMRRL/jxMKZyoEhz
anD+WA+5jM3STjzJ69pE5iSYf4lBZc913ojc3Dpg/PGii/KqH2x6ZA00OF7thBCf
vHaeB/qWbreQR/HqlBrOAynKbB7KFos7iSHrRThP1QUW6FlNkG5tdjBwARibWQef
14kFP/ZdPJMv8RFQNxT5chCQhUiTB8LsYYvY1qGCzNiz4a9ORkV9xC9KFGVCBpnm
Rk6kzUbpXmQRVwODP4c2CU6krZ5JWpFcR8mTLO6xSIghsxCtbRYldlyINoVpfhev
GqrAEdrCdpEL45bqoOlTvFutPs9O3iAgzlMtUSBBn4vNUhZb+BYE9z0sW4JpHB9j
ynLJ2Dbn7t7yrQtR0UBtd/Z9rKdYXipieSGfMAeHwo/i7C8TAEIm7AVxeMGTmR+1
Rs3ka7cv6kQnTuf0rtsPu6SUZEb//KW4iyxLYwaKnGyuiLTbGNxmfbifHjOp0X3C
J86PNH+42cpbI5ZfORdep6VZZ9YTDOWLmoQNPhOIFNavnucYRLPD8P3Pe3Y+5X4a
YgtBURIIsV2ZZ8voFmxsVhhcf/p94dTwtcyqMUYpsF6Ovwgc0QC7pw2axcXteXrG
xu12mydGjnPtKJCvxOahwPItnQTRyM/jY7UyLdc7f7K4pllMdWZXJ9jWQS1g3syK
N0xdTj2WwLN35FKqrGGJBqa4PQAO6g/G2yo8ymbjuQzxrzL/DbbnlaJuIHKLmCxY
bcOLLZbWIyzCT5stXgtrsTivvXCqTkbjjpbVR4icB7LQEK8y2v7P9OIRhvyKsXiu
6gjVIT/VUHz/5sCmgNTfZAat9VRH6mnhIea/jiL362zF6TCAoxDhHNESO4KyDhSd
3CVxXOb4c8SE9ntgrebrWrEV46ytoJM9tISpXcDmvvuwog+YgtAZKAB0MuAOEN7V
Ho2ADcLjnpxP23U8+UYTAJ/Z7VSeZJ82haV5otJLrTtMnGg7/aCNHUOOdO/pUcAy
w+RELSCFj1AR2RsPU/J/yJNDwpPnTEyRcY2YknKt2sFAvx8eNpj+hSeaz0H6nTi7
HiI/rhxEE6W/eCKq505Z+8LN8Ewl/jfljN3ZTQGaFkg+FB/oRDZBSDel2yPKgsvz
jbie7tM/ALBXHCs9MPCM+hXlXndHofRBFH0C210AlmKehYcjPJxrhwJjiQRPCbhv
USylAbT+ixA9BZs7tAt4SWADVe6HqvczJ6ho/zEdlSGGiC4ph9j6evUwbezZHj6T
iDOvBGqrD2g3i9Am0Qe69W5Bfme5CXgRBX+naUEwMyAcCIKyvp4i7UkbAGxeEkJh
L4cuXMKoYKKLqo9C8eMAaNXNFrtBbPwyW8HssULg0ysvjUPamedEoZlBMm9vQtzp
4mUYLQE610hBQWZgdZlOCvQNZr8RgPNFTNedLQ/yo1rGow8yMdvkKG3dITU8dXrw
H80m3bSVEtKx5Q42F1ioH7SslnVzLB+KgT+R6F/xN+Xrp/fuQEIqRg1IYilSN6kB
A3v4QEbdby4sfRpVzx84Cr4YIEFP5pVIaH87WTRB8tbe8F71Gm+VIXqBUD1s+/95
xH+1bpTxbUeIM0io74mBUsWSfmN9xjaawxcV6Dx1MJrl6ISXur3jNs2LnzYja4el
1nlTxx1JSE2i8+vWucRZVL0ktBvensiR0d9bD8T+zYDCuW7YlFUWFLvn1iu+KnmH
PnV1mOIgcdE8h7PHr1r3mgOhoDrSIDv8nziPQqGAZhk8XUd5Tin2BM7X2x6PaS+u
QjvmyX7iSEjNve8on7nvbEypwRQgokzCZC9Vj8nlAzgn/tnM4oTF22NTG9ng+6qn
6t8O5t74fT5Vzjl+9AaYndeVQmqcYYGsUR+pUt5DpTwyohKrm67qau/Qe57jHbSn
h2VeCidaZa0iEk/WY1z7aZzSAQoVLIW0bgVvzOAlAqXXL2jYDOSV/lO5BENARbCL
iRzKsTKFlh0Ix3WX6cukclpPk/s2nLLBnPlNHi4lFKJv3gMCjUzy8a6upouaXnmp
7HKxpYbhsydSZY0kv7vKBUohC85oXtifK0eFp+wTNHqgf4xMXW/cQ2r6Pv5roRBS
mt6m7Su2eZl+vlVrvHUSbkf3AI1h8ce9p4yx3TCpcORQpqICD1pcpmgMtENA/Bdr
n8poaza13PIAVMJW0b8zwByjfGtQLvb0kPDvUjHziKJAMfdOwdZPsDVWor0K/Jb2
XLGUIWGRFywcW5W5wPDEDR0XjZ/PM/CNQlujsuBKzoAkyGFYHf+LfUx44rftZO6+
1V2W3PU/4tuszPrANWeThKdRtGepfV2p8tWpw52qXJDh6CxQYkLJZnOxfwW6dxeD
IQZDfsJ8hA057ZXzfNzEDb34o4xh6p6YjW96zZYqH/lYHVW7qkLLoVOaLYWDDjJj
d0Mxdt7vTM8Wbs3E15pfwn83UZpxOryDvsZo+W78TvlyikvFe3NI1gGzYDQZqUAm
NHwFxPEJrR8jLIR3KO1pWtA72zPT5hbgCAF8TIA17MpnsPlcEhLu8T2d7pF3ci3V
g5qwLXbfMgZOb6MAGhgJXaRPpWVkLFg4FWPGvCXjNRmMIf2CxIWZQsVecxO4lcfA
wm5X9NjYe0/SGZWqXurqOtFtuv0nwxxNJfqB5azEn8Gwlr3+I8uNwGjl1ADhxAW5
ZToldNEtds1/T+GEZ54MHnyGvh60xbhjCZkhj6q3i07qKSzBuOAWea9R0hso32I3
rT+yQQrxq8cnYetRi/wKSlpCzj8GTYzgNjeaDkcIot3Ewfx/vUTnza+kFLJ7RYjK
V3I51lcrzRKDbCPHZFBONUv/LZk54qNbjF/aLYh6pqZHnsK3KfahZbVo+igO5Nd0
eLLpm4ThWb9d+eV2lhL16he0CpF0XDCGKiTEohPypuUlAJwK6HO66C94zTXWyKaQ
ZwgkIqeSJTtpjSDP6ti2jVgDb8S5za3qz3mydD7daqhFS7dsL+n3PhB7qlwg/iO7
Vni+OJ02nA7vWXwRKOpGbNTtq0BVidwflnlXcyBAktoG3kTwPEA+IAog1ewTO/tZ
+kPVt30BEsqHa2J26/v7tWk7uzoN8QoOS06I77IfKBxWJPFL5LyIjwMeV6/3v0um
XNeflQRUOP/qllF4VbAnBJ7Rb6Kweevbemzyu2j2QOlyfb0sdiFyAVH6EGnyiNdS
Qw1afto1zBe5VjmQgUq5eN3pcd2kQ2Lc53hXKCPG0hR5jOHHBh2Tzov1+p3b+1eI
/HeG3fNQ2XnafGC6DpS973EbE7ySGBFaFzRanmB8vSvvxbV7PbFnUBgKsezPc2fw
cLc1nYZOA/u3HOwjc6gOMfOcmR5oBjbHg5bBtDXN3LAxnXMwaRqDXYb4nOV+g7uz
QEabGl1H0TBxYRHm9OYusDlDSJ8mhiy/gzGKRghvbq5L6H3XYee8OBoOydFizIu+
3UumKrIseVv1eMBnDsBZznQtcKRodOpIbF8ZDkYzT3l8noTBBVR4jcefyZVmCIm6
lo8K6VNdSxcPDMXtYWMJ4FCkI4yiJtq/TNFtCd9KDUw+X8EdEAGibxNvyje66BmK
MCfcLKI3iDET74RcwlA6mr0VjSwIAmZvNSP4ApRdGdLFL0XJaiiyStzLMYzrEeau
XxG6kRqkBlPUtMtwPyBLVtd/HrJsXejism+5Was4qj92RCDI5X/yMZyUdjuyNfzS
JXAZRMPy/O0sgvQLhTbF9+IeQ1Gca8gwyDn9PPi1NEZVgiXIN3sc90iiVnllHLiY
DESik1/8YwFaCfUTM33gazgOobjGAH4ZKvF9bPcithmPC5EDH/LsIMlJo5H+vJFL
0oFv9ZuIYrRj5wwHpCxXuiXx+XigD8bxRANyULUrgzFquOBON7f+h957hATr2dJT
SBmyVIcIJAd87QzvS7CO2cIbLtjMMATbw6Qm14tiQ9/yJvBSRY7OsWrXbOeaRz+L
/ugP4QyA4phBGRFZz65fkFqY9nrZRtbRCxWe5b2k5rW4icDF+9gbu3C+hIoLHyyq
/n+Uec0qnvFhbzJEMpG2U27FG22650lbz6CASJkO/fvHV9frjQb0ioDP8uB2SI+X
eT6LWQPtNi0B/UeKhnnD+WnQqyTpGQWJKDbhgJEelUXszCxTfzVWAmUoUmaLdkNF
cbGxxTGBlFKSVH6q8Xtwd/IqLSEeozFQNEAqQ+qljNRiYSe/13uYFYaH23ZmbOVt
OYG1v8mPTutraOAy86SfibMIZ6uyqGOixZE8lHq+4hBPJ+ds1uo3uwUNiFm/vJPl
5ytYnO1wbyq0OxnfDNQO1ouLRlAEQiVW4WKSwj0ZlMg2EnJBK5uf02eX0pmF3VNq
b0nxTCLMS24of86ebXxJy/hYVS/y51q+IbI/Nl+4BhW5UbdxUXvwRlZpizvxFqLK
OiBIVpoOaFnsjDetJMgtpe74UakLWKjEXwvi0xoLcn66Gzxm8evzK8drAgF39ujq
2PgmqimVEPLXHicbW48LkTN43RQo6FaSQN26SUEVFi6XKBQ4JAjeHD8l849eDtZ7
/reG+d9kT3uWBuDcy+mlK+H9kZJKaEjwDXP7ZEhLn0cHZwJlm2da1Mkh0wk5rT9s
IRTpb2nUZHpQ9nfx+FAbUbXYkEcvQJrSaPV/79MSKGaeY3Rb/RLCUUqOG8dgg+Wc
XSJ5RIMuPO14rUac1C06Fbw38YG5U7ooiDJtadNf7QKT0vFdpmU6P9hg71BsHbPc
ic1d3HsZ7BNt5Pldb3is1O0WbZsXiE6mRy30Gn5smPEg7VvQxlmxM4cGDlyGMjgK
yge+AKGuF9xumQbjEEnWfYkCFUoFGBKZlXiqdTyIGur07kQFT0lrEtIsikel4cmF
mi016hHt/fKxdrwlj9gIoo5tcXgX5DXDjVneZGT14pYxOfhvLyYtWR97TEjVlEMT
xfRD9SoH6fBTDzSmc8nnLLklo0P+QqvbMFAduiW3eduWMIE7ADVWCnOEi98ME4o2
JUGdxAq1yJp/+DHXeqONKw59lNRCtUK17xby7XtJqEkjZ4qNjWGntRu1VRY5ANKj
dJu0r8sAkSzZj9uspk/w74DklgQ9on4Fmx0y0jverPjFOay4HAFUMd2iV1ilr/O4
Cuif5DKE3qWw13dqbuL9wLxBFmGjazZ64PuMsQiwuYfJOAE8IvDiwJ+2G5C4PwzS
VQTaGKnFXGaHOqUea1f9loMM90wklwvNKV4FQLbRLXCDUigiCTANY5ppPelSSogT
zZfKZHq4PzoLP9sD/9Wo076GMay3a6EBFhG7+Qohzybkt1LRWCKmZwTCjgBsCIPS
q6Lj88RiUZmZILpHfjQ29NHMULX0mbVJjq2Ci6/kTjIIz7e1+qb3R0hXEZxwZINV
y36cIH7sdD6d7PA5KW0tBR8cm1VErOzXGsiZeI6uKK+OvBy59umDj0kKLu37m9nq
54LVRGxsXngJqu87BG5yXxlZcpDcBBWvJZQqckeDR/KMAb/bE0IIPQ4ikbIuq7JP
nubPN24DXRC2JLHbYfCdnvn4+fGjoq2y2ODgR7uepZOHoNa2FA8JAFNFkixa7e+A
S4dxqkkGf3QPbGyY9/UZuClgcYhAC3L/407QV1f53CeWg8E53Ef+kQZLt7PARVY3
uavsNxc1qB8RUilpFqnECAcvoB/8EyKMA2GJ1J7P8+iFsTskGBIMDoXFVUJFHXVW
bqSmR9QZ8EbRe9UCq8HHzfDwpD9elZi8VZSr4dyZ7/F3CKPPzEGbcqdaXQ49zuaZ
Av6mzpcmxP6B5338a7cHK4GBbsdfPh7/vZy5IIeeM/rGTXj1zdqNKuqQ1s+RNKKF
e8xAyt5Rwlb4jZjdhoa4dcp1uXB+mFcH4hJDhO46Dz8eLPL/NVJhpdhgHCFsutmr
YtNSxjqz/iew8ox9IAKad+dqjdH863atd6ZHvhouf5Bm/T9gD/Qzb6JSUReAPH/n
QiHqeN0EwBV+7aknpoX9m6Ho4R8iXlDKbYWeZ6hUeI9UOimOVRCvKFxJEFiwZzJe
B0S9SvnizAwdZKjwgYPsdQsK7ocMghQuQO3mJYvrPeiBZgBwD9Admjtr+RmOI1h9
gDj0+rs/PqBBmjYrsJ32hr/+4PTCwYHKXp5p4ZnMx2DHZe2gwoUhSHvyhrr/M0nP
sHd1UvVLd1OKON35MICkc/Gcc7gCk7LKt2BhoX+6q6HgMOUZPgCEvivWMma3Vh5k
ku1swevwY31whlSSlT4v7lIA4kXisDsJfsfC7XdwyV0q5T4VOqY0WK0MRw7tp9r5
2c+NWftmqbexC0JQvuMkKoj7eX2dvooo1Vs4WGrAwrhoGGB2zJYtzp7Qk/ihZY5h
AbGArWQigrEivHk/PEW2Cq0k9HPMs/8MPynQizB7FCp2ApUMqlnKEM1ckdGzcMnQ
Vs+biRbYqB7vup51xm1/vbzG//537qol2Y39MGX2Z3PbCrYkrFPbQtctOT6WaQ3B
3ANj8/Hn304FrIyBGaY3p4aXKBxianwMB9vNvXJAxhmeuzYEVbo+JO+eXFKgwQ9v
7VH+BPVpn46adM01Q6B4Q5F3KAZGfXVUCxQRSsGdUrPctLVbwGFIRTXNR97C5Jc0
l2lxtgFDjL0EbgUhHfqgsU093UX3LT1lZF13WM0YGXhszodtmrpXv57481mPaZv/
nD5+cj4VRGl1216vFNPPTE02oKFJ27NFCHt5Qxwk/nwqsyqLTA5pq4EjYeskfwcW
pd8CSXvivLqwXXf7Y0maJkYrRBGS9h5TzVnGJsXFxMX307147MhIhbpxnDOj+CP0
kbY4wrThVdeC/wBAYCHdFtbBL5M+ZkZ0ER7oMJ18VLBWYlUrRjD1kjIWnFbQd1RI
xg8lQy3zvjCgXfjxTGMB8SpmvXHofkKDSb2z2SdhKJ+TiRyt1iBed7Ihicw+PGMG
oBOHfkEhfNGrRcBNbjdUXBNR2lr8HPCeUqrqRVNB2RRTHEWD6wgxe0xZ+VxwV2/F
tivNLu6CmeLT97hUOvE1yG4i1kEEVyd3xeMRj8nStoTJPLt7A5aDE755qZv2Zh2Z
0hMtXYMJTJ7bqwAKA4u75rwvafn4VWU23I7R8oWbAKNmJzEOq4nj1nRKU8YeixTx
aF0+3OkQCY40wRQpQ9FAJ1+Wvsx36f6dfeFlDdugijdk1qs9kgFF8LFkQiFW1t5M
jW1XRdamPt1IiBKpHIPFp9AHw9iHRF589uSw/UUZc3UPFGQONpTLL7jrGLXMc/gh
5Nt3M+tGWq9p2yHJQk140ALwMZvMDsA7wtyIbzcrdL57HyyAeSjw3HrsXZS2OOWR
CN0hj4tNkUp01dd7BmxsWcvVSuApHyy/tUHY2hlndLqsUJnpxnv8sdJAk/YKxn0u
MRlnKuwTs4Xv8E+04E5CaqUgvM8xbX8u3jiEVuI3b9Xm6+T5o/yaKbXClcUBsWeQ
AAiH83DfpSS9YiAhOFttkAfy2Bw+hj0b8Sase9F/RCCaJcD+CYESPyXOzY8c+RfQ
xMs9iL/BZkmV+lZ8pt9/IFxvxS8CEM2vaZFdBODsKKq2qDG0zgm7tflFbY7T7hTy
Kis+Kp0wXZCqmCX/wgFnPxyv/Wr9mY69nwb758yJZG/d5Qf2XgBWKFCp7zWkwLlm
949JbcmS8LIGzjJUkuupXCzDQlxEXtROpwz2NYZ3JiVNvKaQKKsvW+2muO+emjn9
bovouWAdHu4qpDswqX8Nc+cWTTu4/R4qUvyLP7Lvt10OGLOivHpMqOK/5jMWi/z0
pIW368EvJvzEhIYxvkDTLq7Gugzj6s9UQVAHKV8MOFt5UvmYTn2HLanoQOEUs/04
L9aPeRdkvNU03cZ1AW3ICYanR9nozw0U4ITFnm1erOU+3MYlGFXj4H2PvehH52y5
62sBq+VSiRnOYggaNsrUAoAgQWpXb9DhfQKb+uia6YSQaDwmxhSAFgcXMtVpEr59
uH1eY26Cl7dXIJENVhuWGlf7S6SrJf6Fd3iGtns4a3mEsmHrULjnKwfig0MCJl3b
nVXeoy6KJdMzqfridzX+qRglByuB30PPjb5M3UhI5w60v8yuZnqNOI1QAB8lAfyn
f2F5CcsrJuopmSIqk3lkNIT4XEyE8Tz3CTx1sKWjsh/6TNrBdiHjLk8Zg6XwlBNk
cYYm0IJySIsJA3ylTebcgWSodtMrOBvLICQpZdUU6kDt87n0Gm0rOkVFugz3UhLd
+oB7f+8Oucvdp4mLgc6sT2t47f+lK4nKPrHuvoTOtkS9xIO3ZJ448kah5aMwZZgk
qcfBw//h1JCUssqFjZ8UqXSVJnwE6hyGkJldKM0VrQLFT+e9AsBBcK+Ag41uTpde
ezyyGVQFI6NU+VHFFgUMhq5uAq5XeAaxBgpLzPuJi4yW0RLWbywg4FjepzCRblMH
fOcNAN5tTtxK2Zq5mJrewf4H96uZaD7uz5BdFkztqhEJATiLp3NMSx7ofvhOSst1
feOGmNRvu8SOm4n3tCVcO+yavzqDneOGkp3vLE6yjNEQyhV2xYXk9LifcnhVpeiH
wbvNcCBsAeE5OfgTEosF9rIL81KAfoY9HavoYQonsWVPRu3avY3ElzzEjPs6rwFq
X13Y/bWjfC81rII3pNlBf1URFavjdDJyO9s+KUjH4ZzQbKnPl346Dun7iRdcu7SW
/BWNEOvsgw/PbjQw8dnz3qz/BQg5g+vww4zXRGwhx7rPIcQJQuJlw67WYSmEFaVJ
zZPlMuWGsYbQgdy8JPEtCIpoK1T/S5H7P9Mgmj/NhY52z4wIBALLxkMvqwjOxVgs
opS63HcfLvy/6PxraF3lTKx8pWcnbvqWgx9wez5HgMN4X3i49IsP423iW5pKzknJ
/SxndRKCXPvoMZSomoSVsgaGl74glPuE5eAsBArGKfW/vr/SsgueBkT7HHQA1OGP
fMdq0CFhbCTZMnDLGlUBHqLiMUzWPnZH+z/lYOPXsAD5YigF7VuH9hzhOBL0w1Gl
kPGqf2HsEWLhyAx+M+hxnpE5Aa+iMxaBcdCzKFInSq/ZbtO1m8YmRI10rO25z2sZ
ZNO4wx1IFcX5jhhhAlk7cOOWQVLZjh2GKXujDOs4df8oHEhJ45FqGz03p1Okoqpq
CNWIO1AObA0AKw9DOb8b6ty9Fg/tbYx2ly/yOS4a7bnESqonrGoWlQvJN9DlTznK
Dbhoz/IrcthJmPCo+FJlgUDvmOAkp9TUuF6JhVXjkg65DlHM9uYH9N+DI2QlEv1l
jTdNYk0Q6ooYX6A2SYa3zIhiaGk1fG6J5zONdVjvkzQi/HstrbE47gYWkjI9NB6b
Z0Lb2NseZHy6akqUOHNa9yM+rIf4xh/+9lOKuKJdUgTfcl20q4lwA2Q2eX+yNhCA
IcVSM6R3nwfN8onXI5PA3M0Kr1K7LYd6fZVorLyBsSuVMkLXlivYHufQWrFfRiTt
Ugu3WTK0MkAQFXLqNUwf09vay6D/trIHCa8ifbwqgZwQAuVG/S4YRF3DvV5t2+Ga
6ESH61TdkeTecTMxldErNzg8/nHqo0cRNCqmW4hoebCOsmXze5qa9FDG6/d4TokS
7NzFoohp3a7BBw/tSTuRRtRRmTcdz2/ko/Wd+D45WO7VG81iroZjBeCWA0qEWCJc
fo/AryPkfgwuz6GvRfSigBMsrWxkcJg29n2XOjRvV1xHSGxJHnFSoR0fgZ80PcC5
sKHbrTfUuq6GBVRBwhqAM2tY4FMXlU5Yd4rDjcWL2UHzVrI0TrK0wi3wJ2VVeBJq
iRDLeRR/tOJ5QGI1jr+v1QjcriyMWYkSId5zMThgvfp4EJ7EQQjRY8NY3f314RqT
ovShWKudC+iauj78oy7KadDl7CE6PGw/uq68J+cVPaT2SlySbyA2chu/a76vMh+9
pgYgWxXC8w8/D4Byw3wZTbt7ksJL1vrDh3+CKxe+xp/RJabAF0zG7TheMz8lNc8b
5Z7MWJlq1Ua51SaLlSGBxMsTPzfoH2Jdk+OISKrKm42iXHGz5FYtbyBLvDAo1WsG
6yhBZoZn5jFV0uydjntmbyyUQkiQQyYyKTwffNWFN5u6ohOhncLQSSH6rf2cG5bK
DzuJJjb/hQuJKX+GnbqFTmDPvzCZYx4vzt7HDzCuji0L/keA/f6FTxW2dS4BXHKE
yvaozB1m3kZNW5o+5QTEu/zwW3BEaeda+G0hJBbkgxRDuGq4PnbY/HfBH6Rkqt1B
Rr/fYCsutAQ4Uxpd7N1ILl5Bgm8U/9ZaV1uLyfzKJzHLWV5lwWsGxnc/iIhh2xzx
RsIj7n/ChyQ8VHKJRF+0SJposKmm9zE2b3960AukJgF6NFXDRruelosr4UakVQ/S
bW1RDiKPWzRMuPwKAHsx4PB5xsWUP3N5cIdl1F13UieAR94Sn09XTpbiL+kKrziG
fwFt2zeFVFB4yO1r/ZkyeLquKggXO4lQJNBrjDHZUYaX34iHQwZha0IzLzOsN+Sl
unADK9s7n7uUQnsevZw1ViqFeiDCM8JTzxewDU6zIIF+pFLduenpaX1FnDdqAQXn
t3xWDK0OPFVVk3Hv5norlcJot8ZkRKcY1JPtY7+gQe1NNvaTZ9L3/ERJkrX7osMQ
n2jk+rgI3yn7HDvJphB/aCQSEsrZshgSVEdYRL/oz9A8cvxvaVRbpVRUMBG0s3rS
9YOHmS6kCGlsGuLvza7iPZ351cJ037hTYv8eK/DS3wctM7qSlcZSdVk76HE5VL0t
p5Lw2/ogRKZNQQedINL7ixBX0PGMg3lBS4igVtPYuE4XaTKWe9WR83+rVKJa6k4u
J5+UeDHxYiMq0bXSGGPnGUoGNKygOlGMqMAz1cWMISHgqQt2Fkj0hkGPotBtJALe
UmR+DYTph6KIWstJoEqz+6cTMrHWD+soQj/KWMUFEXA01mDO0i56g2ierc1Qn3Uf
N5fC57+Y+DVELZc9gv7YrtVRbWnOO12iLUaYIE1hweRF0XqAcbAqDCb5lSSVGYc8
8SK4QBRMPiPAWMrSh4NdtB+mzrozI4tx36TO6ZqHX29XlIbfiHlqF2oFj0oB2t3P
0sYTUBSL05wuFmKU2DVjpQCStIwAXXc5MvOsCxciFWIalErQEaMaan2uC2O/5eMj
wIKEoPCVfmcVxLLy8nPUi4IPuZS1Xgp3zd+opzTVMfVYaPM/j7e+c7bCdgSbOxIs
cin/6/lDQ+iJguN/mTnw3fvZxaK59uWxTiaaR2JyT3b1TSumbYxrU6W1S+aCpFTo
LtS0O2mJA1a9A6mSGuU0RCJ6AndvJfruNu6QdqTlKQ+CLcAN+2lpdebM3hwJvPBd
nmo3HST5RyTMKtpkg610nT3b5Axr3IHNlrwbe/B2O6M9wskxwjH3YcMEjOvCtXF/
5BM82HeIX6iJxFR5hPLdHGKukSC5uXooNDFwDp0mVhvsh3HviNXDhXNccO/P2ki9
O+DMJFLr9Q4YKn5YxOKM16Eugge360aWR+WgAuuC5yNdZR9z2D8ZgUdb8iOScFQ+
U8AW798PAI/xYh9eHLqoKpgpJbczrNAHjQwfJrANsqDbOOYwXYcCkR/41Lo1CCrc
LpeoSGUNrv4jEOxFYWOYcwve2UC+0/9hGlcgnolGy+TQV+PE3UwcZ9NyV7M2mbsh
N+0yMuvYxcB9upRCHB0HKEQ9jybK+HDWYTnAV+M4qgOK7ZGSclf0yQljxYF4OAtI
mndo+KZ9PHbMz3WkC7miN6/lqqw4bBWgGTeEs9XKk+OaCtXtgA6Tyke/7Q+v6Vzn
MzKMyc4R05YqBvzczuj8rd4UGa94VteghkfyScLSuW7JceHKEeOwPye8Hwwy5lJz
kQwty4m/Z+GaMNXbI54mk8w9notgcd7DTEveS8QzpuEi9YchfXgpNEIo44W+4sPb
NG/rnii6ZBX3cev6Bhe2eCql1LKQpqhbzw66ljjv2A5BLLW1A7+rQSAGlPHwNsNV
WZtE1JaYEkgNelBZhCGCieDpb3zbCv4Cwc4rZlEezYkaIUyQLd1W8WIqWPiAzJaB
OGMmjkYne2s7Rwo0GI8jkiCtg3szhOG6DiK5ZEeeYS//F+wNYwy8OyYmM6GCuII7
zqirSi5QtVAkMlLdaceigtIKNl70yFuCYg+Q5lsuk1jQxTqG5e9YvqohzzkPvXdi
EiEmAGwuNL8tandZOteWpu+9wlmf6AgztJzFAL5AG6gRc4Gr7NCoL4Ij4dbwJRH1
X/6/wyN/dLariC+LLfke2xS7okZM+grIZ+arKSflSPcdUNVbl53bdXonuNe3a+OL
HBhqFzpLbw+P/eqMVRdugDQSlkuAAklPeH+rjDRkpPYJq3q9Z5zmyXPEhWdIkwSQ
5Dgu35w5guAqzH/RmbE+fEaivuesgCusg743UXgdCMUCYa0J56dIazvGxDKoFAAp
edRhU8c8CSoNXJYqBNdDSvrlYq/jdHaRI2hcdfQGNxCszdn6oRjVtSkA5I6xbl5l
6ORvtjriWX9Nv3qKS3w5lx6mX1QHKfYD9yL2zS/wNeLMMRJROZNy5byLTMLth+is
yo/WXrg9Q2ojdjfR4g4q+jcd7UEBRTxGWKi47NzJwVZ+9Yiqab6o+woSD/VXiaB5
vtdwyZbRaUAYcxmIjnkwxiIk+H5kgPwQl/QuH2MMLcXvnBj/JV6R9juCYSqGHh6O
V1LKewHPheDTjf98X2rtCi4MGFTxbmChi+3Xa1AT1HYscXlty+RYgi3Z6zyBL260
+RXuczGK+tBRx2YYZrfyqjvAP2VSBf70NygL9wJjxpBj+anEP8hsEIW5/hSBFuQV
v1P4SQqi27GnaOGaHAnJ2IGqUTuC+iPiLFbxK3iYfLJXSjYZsPOkTzDnL+VWBpcZ
o6RV/WJ+Os7RrtV4GEcwoNDQ4uQYVlEBhe5m5V+x2W88kOYrI7EYnltpxlUOvdIo
pcddQsIF1KydOZWSykZtVmDqCPeY2dq4ea6JesSuPjoQ7pT/Oh7vW2/X9BKkNvwK
reqm3Ug9SL6j0RWwAbmtEqVkNGla1XeRvcfFXqbgvgEDEN3M2vqMkPN4Js+M49On
Q15VCCNlhMwQeKJTNjUvg7VP/Y5oYg7yTiIZwkpifO0NIW7JtesGV+m0K1jEKgR4
g6Oux/tFJHnczErRYJMwn6w7HGvu6SGq1KgPGCtWO3oL4pD/XZ3ED5ITDrUueqin
7CUxCFOHVYxg8Ehax0XYYt4KTSn2be6RAL/NySPZ82K1ArQz9lkzuxeQfY1npDzX
4plmPEMl0GxL3rK3ps3IoAtUnaS+R+aLf1e1Jbsdx2Gxvhe1C2Jx+zKa2AjuvBdN
F0mZ3w4QkuBilSqH0klQu/2+FNUh+xZ1YR0w9dW0MW/vC912/tKSLkf8nYhEzsMn
SwnqJcRssQaKpGtFJxCHPa/+cJegTLJA0HfKca12vNi5p3+WZyYC4GPVPhFE1Kaa
B7fadhp2hSTH62x1XPd1tWJ95pBr1JvkowfQ2aEAaLuMNIVbZo/lM9mwJTSx+tHt
FQedo+OKTd7weOJq7zsU2+Y+w4BvQKfPLPvAgGOHbi8/3HSckrUeu7HwqWZcVTEr
BqY42Xwq3JUYbbm1OcY0kVpDAQs0xu5iL1gnJJwrJvPla5IYdYajZA1k9buZ8jM4
rEiA9MbK8gScMJm8jCiIWGddbINAWQ/vH5MSBCbNWZMWDzS5tJ4Osy0WJWQZjQL8
B+U9hj4u5fYjkujZ5fHSSdXRrwNPTNc8YzUgFnOsZmuS2wmOwD0QgDcsO2wY+Iru
psrQ2TKH8Mz4oPP/JgZmSUHK4/R+hnA+qarG9oAhkK4t4fimw0Hiz9P/I5eSueTw
Trh28PYprBO3VUeV8TtWc589z4CKz+3J07p7cGNFL6rumFS4ziP7XCFlp0GhsLK3
OaHwMGe69WW2znuA1CTKnnEFT7eW1IH+Tbd7g5F80Qxib9T1IIMxMhX7s+bqBb6d
Llkih9q5gHQTtc4ErbuiovZZJ7UESvm0aNRLnDBay03wJlCJ/kBWZlaKsvdUkA5Q
uuxlNL2Ao6etDkzjSYt1CjFSwFAJcYV8SGON35CBjdGPWcVfgV7zr9HoB63cOHOz
3saoXY0/1RlNVpO1fCgSA+ziecZyPMJDLXnQ0/dKn+zKDjpHDpFAi3uFkdrNJ+6y
0xIwwldIgbyZaOxfof3tAuHAlOxiryk7PdIQi8Q7Nt+YPjoAMwdey7PSxiQmoaOe
Oel8kw+v2RE6HSP1qCNWJ1wSGQvZgiaT1hf+TpsMa3xHdn2yK/NAGpFAuyeHVxiz
77RZ/FMqWlE7rv56/wmddiUP0MEsX8xDi915xDn5DcO0jlBrepSTOHVqt60G+VIj
djdLdmQyHjyh0t9HobGk7TFkv1jP1PO+2mMXBbNK5Z26jHWZg2ocnBkbmi9Wu8mg
ndEhckX66CDTNqkjUIO9x/li1LCDcYZWQ6U7fnofq8ImQc8WFC3T3VuvsU2v4NXJ
OGBwlST5p0zplYDzVadHEhjDd5SslUHU5m9jfqSOABOS6UpDhexR/6vXW/fy6nLV
3Nc8iSSk1+IDOcxl8DoUJpIWu0GLnSkRtCqcmRosnuKB9pKMTg9I8EpSouksyOQQ
CPOCfwbCG5BIczs8d9hCfb9MsMeeUL34wGB9QMTOoopBDVsBgp5c1OyrqFDXXMNZ
62tO2j9UfbmwQrwBqvLveNShz2GkjabxadpcrxkXUvXsq25UaQseaBYUk8E/Rq/9
h9ctQZQsbXpHdv87rtv9+rnDUBaKEVY1lpDEwSr5MdMFHYwF82JNqEVt4259oEfo
re/f867Q5j73e8oZrsB2P81+WbiXvXRmxCkkU0PFzDGSTa/E+1wWhio4zkB+68YH
4Hc7qFuIYVgGOgX5vSCWX89QNQWLd5mDxuYAkFnVwe2lNKfMWB9r7xP0crQNLUB3
QTc9/vYM3WtX3GzpGIHG4g4OfbCizM50/g/bDZWLbRBnThDq0TEFKX8DIoAkr9kQ
boDakLmKfasfLPH/8s45ZZsXzJ7FvQ7ejFG2xZ+ps2P/P9Q4Al2f4su/Cds5gg7w
jS+KtnSIATER2aeC6ggOpLFsUgC7bOd9iYNziXhZguCdZkOBdzFfiNKiVqwRZ8xP
obRf7ISmQfJ/UEzYUEg8ztmzw0hskdRu1PIjsnxLQxj08ZnEvs+SpE5zJbo8fTeJ
AveBfPOIx5UFlBgUqnS7Wj7nyBTecAehfDoPnWinPxDq7bIdBCm58QPABXQs1GrE
dPgzSQqV37fzg+8QGNMqEfomZl3p+YrmYfehTjACO4+vhkGOG/+lBM/EEt+wv6e1
cape5NUEIpbC3IXP92aczTbu+jdmsuj71z+csy7Sj/4QU9i7Aid2pDPcrXFlhl40
Sf2DoDPF53Hk57Fj9sNqfT0rOs/NuRc2Qx5lKL2Ly3mMPKtU+w709gIyfEfK6gnp
D4irOR7DwGN6LdGYORNBw+L5LrHO3YQrZUE9lHAkuUFMLrrfg0bphfK1GylnhRMa
S0MUTy5+YOnQsWluelzOhWwwRxJkfqTyHbSg86r48ma0t6EmtB4sugrnAjyPWNfe
hheSe1RsVEcE7bvFUzxIUQloKQVoPtBtZYkwN82Xo8CIU5H8JeBh27X8Qr7/fVHJ
3XfxPwpfvQFQICINeoONHBjc7jt3aQxK4siTMXUtZrEzvLOduXS11WZJDOw9RBi7
TGn4PutzfoCVbEdvtwtA3fkLcKNNJOqxX/gzTnfnjxORVraPlw9FFosKLwMzA2+C
kL0nZ5WMx/qsRxFNmxdDJt+Ss1gJY9LmXuxpIIsTOdunihdWoWAIZPZxSVlJ2iED
9QVE9idpcG9DJvsvb2xIDfB1B1OdL9arlUqskxK08R7ckhoLqLuNXOZhdvrVJQpj
L74nuj1oleNPLBJv10cgBTZvkcD5GagnviannNsibLuGp4dZaAziUIBDEJiZ53aI
yCu534wnJ82DjkJr+k5gzNqQvLF6VmxEIzzSCyuqUMBrhL1bfwA3fOMJrfi1n2YB
CnhOBfghupocsIpod5hHncjHPBzVjG2gW+50DCbnyRxcwORKFSZwRVTYDDnnDWrQ
kCVT/q8dyjNDz/Ff9Bp9WM1xmwGk5Ubw4oZB9DvJIJLMcdSaCGeg8vR8OW1EeYLc
KqixHR7hSr5ukQgB8uoUozNSphHz1mnXQIuJD7r9Z8pQRnQ9rEhsNJ5DL9EoJTDZ
AiALxNvGspKE8DegEP/qrtMyHyZjjO7nWwNiXd0bWCqxWsAl7kbx8eoVCetrsRuU
pM0jfRjvecBvuJplbO85jte0iyPzhXfR1vo9HhOLMO0MnPiad2tM/ZvtQ786tOyP
wutRkZKxSSbBk6wKnEvf9/qu/7B2ZuazGLpH1MSCHMtJc8x29sGWwO/fOzyZyGt3
Owug29BU+xuzOhX2XRBxfad5KbNWxcCQEI2QB0GMay+1fJHsp7pF2uAgGydk8Swc
JOm6x6XWpzrPvjM1JyKbNlIn1pXo8GG1wpQ6Mru8O+Z+PgF3kKHQY3YApMyClfJl
QoNxXEUuzcWrxVteXapYgwCvURb2qJvs7hbSa0lVc+3dP719fr/2FzTlzT6vVfX5
LP9XPXUqIBMwouhNvGYbAIxrsc0yRlLdUdIBSa+zGgeHMyOlX7MCVNZKTN8wHX+X
enbsxhOUX0bLRUeGV5gnzdU6hwUy2jl2/OtaAvY3f70iThsMqdfcLxZPD9d6TlHR
kRLCzD+31g23ll2VvYNTLNm4vtAT9EhRgmKfzqO8bF5Qg3fpkPMnAPQRGdNGWnM8
QhyM7USCJuYJ9R94ed4Y/fxGjEMuXS+ecEkqyOsXw9DKPrujUZjaGIzLkMvBS3gd
pD1knxuOqHjQ8zbPfJhpQFA/+q75lnJFl8kUiaI+GpqRWZpJiSzPOL200dFVgsHh
MTR65VNaKfXvtOWsHOUHvagMpm9HM9L6H/xHGU991K/AM2LWE8M/Xh2qSkbgrVeI
e/C6PVcMNL+txHoTXFzbyjgTdQF/bfpc5znGVhokKW6oNUe/Q7sGWnK8emvnc5/S
J/M4yZ6X82Ozh/9aLE7h4aWedM2SWBrIGHKluHsen3Hnbb038K9mACYX5rIzT3rj
EwRqadlQIInz5GfHjND2ICM4ENKWvKal8F4qiyrZ60Wyir+9McqqyQNAdRrJuWXo
MMRXLZpLmO2B9tHKRfqEt7uCr7dvzb3D7PbgEQF79hRK6bXbbBiwEP9lK+5YDphL
dY0rdI4BStSZ/AyklSdVl1Vs0/7so1s4dXvnENtZX988gD5xkbz+EDJFWXL3G0QY
9stQ/YacY8USIb/8V3/dTTPtNhAn1oGKu7MfYCCmPuQWmYd3Y3ApIiwlzqp31lV0
rpwmAnOhzkFUoRkZ8/tH3TGUTKCpOCTwdNVg/59Bb4U60V9n+ybd3l9twa26Yp4r
BXA3G9u0ajKXFrjNjFn7EJML4gdpdXI3ktWHB+Xau5bUKL9ymM/D4oSqVUKSrqIZ
P+vGdMrlGpGcw0himWH+QKCsEu1nXvQAw9cC30HPeoekkVUlIH328XvLmQdRk2Xy
VBWfS6/DDdagNpAbcBRXAF0SCpbJk980Fff+dUam5ijVeDvDjHRE+jNf7h/1LWqm
qic1mEMAD4RBjXyQA+rUfyOubJXF+VpJuyUIsCYC48fOA+epIbMiuCRIla2eJyXm
6NAsQSctAT/UNhxyWQgU0HgcPSPVtHuyql+tL8X5bE5xyTCQ9lpAQWoAdDh4QT80
vzVryXaC3XWh2Ir2iiEvmyiL4aePshWJ3WWOGygStiD/l7AKtTMB2Cp5qD81mL90
2eyOk6T5FmN6ogaCqZ8b7y3KQ2A+vgrusuXCvYJcqopQjTa7iWljSzi4fuxoxuXz
PcWJxFUkxvcbzOh4C2DV06mVVeBwH9cjp34Md+pS0eKGpnsV0KSGMz9QLtdE8cAt
VEFd74pyNwOsxPFZbr7ggiXt4JLwTO2va3GfPFN3yCu9F0CdKfCUDaJ1KPosbkil
yfZ8y9hZu/To3E/GY7dFAC2np/8Nv75I59aIu1IQbDI5bJwAKnaKsQCtiQeOd7FF
vCMRT4+Pz5bfcFBf2X0oJ7U77zvqUKg92kywFoKKbJjptnKz2jmW9dQvAHsRM4lS
LC+WfzsbdOGQyjjPXfIutE4fEDXDD/RbmCWx8fn2ugbGk+w5dVZ1UQgpDW74UOlA
ZyL6Ye1hDunc2IfiLkUrDeCp3cK9IR2/e+47pI4sowLD3EXka5/i/Dfm/zTw05Ym
PVzUsMVUnCijv1nFl3sKevfmDLlLZ+WBj7SRmsc2Uqx6j7fFwkowsoJTVz85ZuQY
oHS6T2Ck8m4puzDV/2CYnygJXuAFUoHxbhWeaRk77bW5rIC7MJghz58Db/aEqY0E
DKciVS4xaaJjG8n/7iP5n/mBejPeYvVcI/cLT+WLaQbRzfn5CDh3kxsVxH8xQ3U/
lCXLWs/V9OEL6LwkIk2K9OKXNihY7XRDDdfxbIZ+DeJQrnbxILeFlNi9tFnSzKJq
lQ0FJiRic67ondPhSROsLhMtMqyqywoFpmssya/PpRuT2DP9ZVCpoA27ZuQef0Ec
o9YfjqHLWp7hIqnxQlet6fMjZ2Fv/UQhEQy3vXBGZmrm12ZQhgE17WRJCPqMVCw3
qInO+B/XITNMMp4xmhdYl4PjnMjaey5IcYalI43wdsxSdJpyBANgbIFus0yW7tHE
AdU1cpDrk5D9FTf/kXodrokGVko8yU9yGbPOsopAQi9gv4FfLzThj7MUXXOsGOVf
6rUVNcwUBlpdpqL2u8Gzozi3T0lbULFDTC1/A6y85QNCtd4BIFwmF+3DmDBB+Glu
4rsfomQAMyUMfePGayK4rU4lYR1tAWtTPx9U6GPMXnUC077igQCU/l3zLlzclLge
lC8SxU0KSGf96JgMP8SNYUJIha9Yw5OHyQ8oHC82Tiz1yyNpd8cqtBI7ytsqK0ds
w81bGHDVVtsCuuCvQO90VjUfHUh3Y9Jvpx/4/94hlfGQj5WQ64dOXQxSfOAbXr1x
Hoof15GJVzYzRER/XVuUi0rpaU3nBQP7RM3xqRTmFlHkyNxkME8+z5N8EBRm4mNz
vaR486RSffifDdhb7CR45MMnwxfcXi4g7UEelVolYxGV/QwZJq1vKoOvLMttVn2u
2SUe62+EsBNl4B2RQm/awsKd5doPkCkM1KzNnfXUIoibYEY6EKXBT3+w3tLPDdpl
bFCyDaWSWeHpGs7Y2M210ATq12qJTgG7bM5lvkVtvTonkdgp6mIjG6R/Pzc5Bksi
LpCC1aISZTYqeg37PA6TixXxdejNALGLTjdaf18ppa09MUPTtup5IV1VYDpoHHdT
8owonsY8HwaBPU3qBZmys5VdWMdHnFc/XUK6AwiqJJ7avdoY9HpYe8W+j+6jLmhu
09jtPGN8OZY5x0CFK40P/yVdGA72JVTwOUY/cVlQgJf8GLE1ZrBKoAwOL4ZHzjtO
kZY93bBq6yMd6mK1W3PTmHVo73SdV3Q/BO94PWewFhbf2+DLLmVQM+lYefDcuEgg
7dTD9Q2t8vLARLP3QYa3EwxCMd9aP9RpZgTwG6JoSRZCjSoWp30mFCb4v70B8elk
jkMmqBXy3PzvKm+MapnHvwIBD/6j4IquqdzvHu11sqDrC8XIyk/cNzt5WyHbW3sr
FN+NEZMfLp1jmHQf2mRBYVJ45nnobsQoQTm5ZCGEulotzNa0nHUS1blw01UIBCHR
4zWTSlT/1bE3k0JR7ndccWqNKK03dTWpuUvxo1x9xzsUMKEKOI5/VUC8muh26wCG
9fVJ5Jrl+BfJSHzCnoPqrkDnQYUXStQoDgJrZ9EZqUFGslzXKz5zw6XBbYLrq8R1
W38MqkvqvG0bJQBv0tczqyE/xQwNubTPP2Kry3iqIb3tLSoasqtph6urDM1gwtIu
fUKQU5XIrsT4fylTZzilMaw3a1W4UUwEu2A0HBRy1ny7X1tnIxZgBV/xvBC4ZTpM
Ur6RfL6mPlX2+tmoPpWlazWE5vHpfTpGXsAklwuVh1OfeHpd2Pag7aPc/jXxvTAB
JSO77iJdjFblP4DihZ/R4XgNLkyNQLZMBCrI8G3LTIiUGUAupR7EuALEkgKh0KWO
9Z65Dw0OVJ7F1wtpzXupo2YNl9veJOQ+XCws0C1bkp+o2jmAoEhjndG02pus1Bbl
qkG90WSgiBcSJEyF6liOV5I//5pcF4HqYs3LABxB5+mbjOduL77LBAcPz3lJ6a8f
fUKguqqqcPaZEVBMzmVsnczSfOrnn9vAoISwzy2bV2zhkmsVO0rem21203LkKBQ5
d8Q50UvQCjGtw/F/SK1Zjml8cexgDIcQNRYnBIiLYJtpvr7bgUtZH+PDFblJ/z5S
2wADAAPl/sddKr0tZ7Y8xxdd6toPCgIBfvCs2QyJeaRxBu/OYvSQ8CM180d57arE
I+GlftEats9doaBsnbnw0rYQ3rFH+8HHjaF+XbXGGDOefyOCXuWDtlTa+/mVWBjk
j+6v26SONKYIxyH6RWd08KpVix6tbAL1fRgJDRKF4Uc0f1mNSTaqow9S4wNniQdt
OZeGPuatcv/BCjiyKMcwptrz+1HUQCBMTgJbNO/N2ROLplUukQggGQxxWCR18meh
X7Ak6Mfy17VPYjYksVPHuy/xNXRhH/vQtgd3BFAhxDvxJEM8BrtKgqQRMjatpaFj
IwAzUAZsdPBrOvSzz6ItyjXvrFVgIHHcsDIloOSFL+aSZPBogujifC2dqKSTunzH
xoPf1gQ4UxtLsh8ux9z1HNnF9FXSMkvzLKwROV6MylrirUQzY5kcwdSmmDdHhTpb
6PPrqc/zbXrp7ogiT4ycudVEqBIdkVeWWk39VIf4sZbmzjGGBe1rUgrlG2vG7bvz
KQqbH8IElpFyFXqQUP7vLnUIVV19mNusmz4USNgS2gq87A1bmrU37dNGoAIYcvEr
vb8M0PBiICxsVsSTvsPOVbycn6aTskzD/0EhokmjCgtkS/TVdwLkvnSVEgAjBbU5
Jh16bxCG/WOOtOMXLCbpR0ozYQnZpNDaAhf26hyAug+KbHq3Ba6VriolPq1Gg3h4
02rpZ3wHry56XkGRUU6lZ++UPTlJNliCfTI4ZeaPx+MyT+J6ffNsNRJmYGD7mon6
N69zD3EIW0xCNygyHHw9pjqMEryVa9OpQx18J5rzKfFqJnr4wISF6TKkRjqKJTrT
kjy4FEFvdqlEwdL8J+zCBKIDVO19Vf68UzO/9zI06MxUETDwjD4eS3fBXuJs3d5b
RfwbAh1IK4KsbZVhbnd73IN6LGsBzORmaraj5Cs7OxpzSBed5G8puLL+UgGvrHtv
pLuwBegeGXQK483rkVBICCWJ5J5h2NXeysgxZoKADbd9WPKpOmYty9gwcxUYFGbf
azybewtjKI8IxkBwJJU0wWPDBM157J5IpCalcojUqZv+DojTI2+7CpOAE9LCSsoh
cM+4lTIyc3KDTXVTq8OchTQp9SG41IJ+xtZucNmxtJCRvY24s6kVBdb4Fs3AkO/U
7soR2BXf8/YtTRV5wSPGjRSAJEJPHz8cRa1yW7B3y0lA2DDj2dEouSxqfiKnNAI/
TN6ERYNlz0PSTUemc4eUCb3ToVlX/tNziO2Xv9TVaISpcPSC2Q53hP34OLp0BOV4
jARfiphsQI9ohBOfb8sF2q/CBW8XT3lkxZoQO4F7dWVwI/Or9AR4fyktfldK88N2
6xf3vojSFUPBq7tzQ17LHOWrsjJVVlko95W98l6iSGHHxjm8H2AdSnppQO+4U43O
XxVmy7Wj3EDKdd3JyAvUrLIVmjUooHq6Bu4eYEwc+oiJmj4vmgkOC8/e7oJ2FU8d
rSGjAOWcPDIvyQEMHdlMaNvgdr5HeqJlONn1QPrCUvd2AiWagJVcTAUjdpUA9+rO
uGWJbHkaWX2fGLgHvV51A/JO01tkpkeXX4orqi6eo1VzD/6eYuL9UG+VPyaZ/V/O
fRh3sSQK1dWeUGxJgm6TH9urIu5KgTbfzNxMqVtbu1FRCpTl4iFZnOBv9xLMHaUV
iLGCzWd4Y35sDtMSv1irliklEPxgodZq81MMQBbVAckQQ+GLnUWYL66dnfarwqxJ
GsJoAvBmZO0Rx8S7z4Exb3HQ5WT49fTRgGrKkN5Y30bUdL0ZjoKlb6K5RrYNjmy4
mTPMX8xNg70wqKABO9FCywVwjCB4LWz1/ZQyZWL7jr1j2hInTQApsp7yvoT5Ne6w
yMkv1WMaMRfNtSbAB6ZarGplJEQlUf10lRwg3O0EW0mpDSMha9RZrV1H/uYCBUu2
V4YpHMlqI2CU6tGX4vjyNBvCIJ2UYhNZ6F7lrXG4gvsfsvr0Mr+5+amz7vKJpQLI
RiwWY0NtuQonJOuc4ChYfkR/QyXGZFYMvUWNRGBBA1ui1JfFQ9WgxoPHjmi6mIxB
7lp2NbBKt3kZ2mfrSBagEiaaeccbjdCmBZhDZo7jdT27+5eiV8fTrat3DytSZOHd
ituH8EHdTE8Gz40ND3fJmhnMhCwyH0XwGYqC/j1qgUrXTHcHDLsnZ6WsqrsS0S7n
fGe+Aj57SUJwShIxLxF7QmRb+oSx9vUnmvd08G2WuYEGDRlph4EdWOycB1mdEjzc
lVH0BRAInNZFdPcDAh0DiFfGsO3zjJJk/o/1Y4ygVHTa/pWzHW5VEpwX44dJAAQ5
Bw+wjFGkOtNt66Ymd5COhh4lyiCwm3N5nLRRAd7ARsC8/RV+iRi+V1daz0AIMPob
xrTkznXTYsAPaUYuArFXATTdpTuaR+IgasrTyfahyWqwqzmUGRxMJ3rd8V1S4tJq
nZMj5SSyMsA3myoxo2t5V2NQa0I240K7+BDiZoao+SSrYi9t0/7dx6ot1ZVCiSQ9
ehfc8vgEmEtLD+82G7Bdeq9L0LYkgjVY36K58ANnCfGVjne9MyeoDPFkF0uD7cqM
r59shWyHo5jdBt4JJEvHHly8R3XpHJUKGad1weBFpK24YnKxrlMjeabZHjRMt10I
cVhcUp9/BdHuek4EervtqMuRyWRu+o9/7g3zt/XBrznl3pJdloyRQc6u9AyxyiXG
q6APNmRuMH8MgQGxCjDTUHWg200Am8hjjYcee0DMXNs6ZFnK0Vnn4EL8fAFhmiMH
ovidxm+JdcUZcD3SgL+bjQWJojnLt+/82dMro8XOnfMquHDgq2yxUjIPxhg3F3NC
8DsjKjCtxiwbEw1NBisX685/mNejgB5UoXYPS0v91IjvmRma66Jo3uAKqTdFsX9F
rEOkqzERQWnqsSuTZQGM9yJditMzHNePs+ASnG8B0NcYQqR+UcDgbtBJoz4QgFtt
ioDk/bN7eteQBu7yw5QWvt37KEdVtcwwpvT/pROTspoTM1bDaJS+73/CZJe9rWem
BqRtz+DuT4cEFi3zSERNNQZopkWLq7zVWZTSDlNTdu1zVMeqcE4AJHXJWTlQzm3B
Fy1G4VHXo6OTcPLKkqj2D5zUGQLTL3FXXu4QU4cBV4n2cZRlQXDlpLPDZTHZU4Ws
Ruw0bOaQOVikxu0W1Z+DbsXeJz0XBHTdJf+hnFyxVOTTYvQeU4gjlZ3nIkHfBqHI
8KZDsoI+2vB+m1Sxeh76rAWKk2MYcjtoxp02kRRjjtAG5RDQQGBgUz9g/EZNtGFz
lo7z7g/02dUvN4GVI2z7JoILBOKz+DjjzGjjwGmJr0Rug09+6JdpIUStc935yWVn
/z+9Wz+7m+VgMuVmzgO7ENnNVKdsFFR4CKIukKxLyuPrmCq5YsVm6dqPYXVoub3H
ME2aoG3t9oxgTZfuHvHcWWUntFLJNjyIQGHjP4fYmDWS/Nreb5M4bWLYQUCS7bPl
VZ6BOB1ipdqPRMY/6mLDhKoUYtiWnUt3NgbCrehM+6SnGkBL9wlQqEnxGL5Gm1J6
rsz3bSvElKS4deEobHCL7LYEQZwYEF4YVqOFjjKSf8kBtvoyGiqW9MPGzk+mqRgM
tNGBNAczLCZFWT0smRJa0ekJ4xYNyPu8suF6kMRu2/AopJ9v4PzrO1Gkv1XLEfuF
mN+J1qgPWrC0vS+qEHOqYkqaW5tdLOp7O4ZUeq7y6WeL95WA1M//saudKrOu2554
IabB9DNaLBFRN2jLA5sMHlslJUX4jt4coGyGWNfhz4LoeFvhOKPCP0Fl9Be+xUsr
s5fE4OZd23KGS+m8LDf/iUTv0KyVspcF5gMiOOMOOnqeAdzV6XasrB5If1Ej4dL1
+m3VCccxcAtZvycoP1M4skDBx+5Jih4uJkeuyrFOSjne1e9Zao18UIoH8WlYdm4G
8Spz5b3KaFrYqjinZuNERlDQwkmifRudYCxKXtqZlaOxBv8rlNgHB7kF4d/1sRKj
GObAexDv/o/jGuI4s7Fh0ep78o7Fin5NVlW6ueyu1U2UZPS9idMAefeKFU+THd81
kTVqkZTZn1meOyrHpoGIlt355WKZKKmuooLi0z1XpWCZ307WRjFURPW8bXxDchPn
H1bPCSwgiaSJB8S2C2Tw5B2vgW3/j0O6h5YHrC1AXY7iEX/7puPTw9A6ynmx+KH+
OMsBDHHtHjzb52VZjW7DkeGwM2v/vvL15fIuj8VHHWLqpJQJLrWLLe29KWZm7Fq0
ZCrPVcCcIaVJEvoBmvbAY9C4HsO4Ls/adwUBUl12D2jGM/xeRVhABvsAnmGbsJJm
NJ9yd39SGAKOLV860y7mFAdWxahcYBtbc/A4x9Yt8AIAegPzgTsXJKXuZCcmY/hf
xqdRAy/H+vARZ7ExHgZWAwrwyk9nTIPu37LVexnZyuqQtawIiqciUvZfn6V1CmxP
QzJAxIIR4SxislrVrIAde9//CpWj3Yv6Sa1CojMp/d+5oq783a+TkDYrspjt755m
3Rvn9NV7KPuAZxBstPbXyOJfSp9qrtnJq2df5/quAm+pHB0a+KsJaNWxr5t1prw+
XE22kgvpTM4FqB6tkc9NnaEemqq7UzEBZ8oJ84yRBqTxg+xHE+VMEbe/vHYnHwNE
nxeGZjqJcTf76pl8EEQLgHL3cnIpdVvxATLVA5NYnzuzRp3muswqHfRDoSjYV7CL
o7zzkxi3LA0kyt4xq/z4jBP/e+0F296WOPEsDE1RQM4eIeXahrlaPkwvwOxtiagL
XnQCCE32QHK0MXEKUx9rzaG7Dhu9bNpLoglmSorbhFL/NPM0B7oh9hWE/8RlJc0A
1E8f2BDY8Y6EbjcEPB1byBjncnylwIjw236T1qs0F+8+IfrNWUmE6kREl+Y6GuDy
cvKBjkK2Av2gyBcim9/ldDvLqBwiSW3LCwjP7FlTHwCJBBYvETbLpZc+GOqb48K5
k3BOPYLiw9Ems7Lw6Nub4eG7Ad2gYbPIbiKUxBSTPITxZnvfx3HFAWC5UQm+B+rK
sKWlvu+EFwXp/s8uYmeXIMe98OOo9lLdzGeSmDnlGEAE9AsQx/z+JCvauJu2DjRm
Z1eNJg96zBd6ZpmNEjYBgduxoAs8nx8AjnXiXZg8iWXwTospj4C0izteaOqUVsVn
EyXdhgNzOwRukUlDAVC1Ey0bVPWI1PsVOn1GIQdlbaXpWrj1WjRstrK1UOdhSJyJ
5knoEW/BxyI3NOPd6axft8zfa19dr2v6nntiBS2CECXcsq016ONnk6JrDYOTMFS6
BI/RaNI0iBljl3tFauQDlQMsWRegnPefGSKpjSPhzhaQNDx68/6JbUGmR/XZK+RZ
euiY5c1sEC+9nbsKFoNWUtY3JtXrStFGYlEvSnnwg/pEi6wXNaJiVK6+HY0RYZje
r2WOEsbk3Mw3YNyieGNO+lws+GwQ7pS8CPG/49z2T6Qnd8uf79rRSJAgMD9B/VHW
Gtkfv8PnXzOXZazKuqfroDSrSVxWivJcsb1wo1uyJUtsdFnw+8UKkk7186LVHooL
b3pS45x8+Fo88ijnCKjR68tOvGoaipDNc5ajqhokFaFdGY21nZf1FtGn2mFXB99h
TQ6ko/pF6KJ2bpTBRP4BQPGhNfB7VnhVhlAF9ZhpsyAjB/S2wGotZ7lzdqRPgfSQ
0aQGRQP9mcKIoqvQ+C9WP03xgmAKuo9928BEyD1gEAJ1oWhMfLmxWCVZN8jE2ESP
nL9Uw5z/W8re2HNvpwZK0WxUWPSpPnt1bcBzQeLWtzpsUltjhOizIkoET4hcOw65
oVysy6irOb/sByScU5kIlSmZgMk60WbgbgerHOdjnLoVk3gxY3hLq4mKvRCHANpY
/gcoibJDgw7EU+Un5s/9LjQtZJmo+BlXQoPCvlNbSQXfLSrURl2FcfbkBe5/K+2A
B4vuyRs2ZLIFrikuKpLsZLO//LxatydU37sonEYBR4Af2GvHRTEsWQWLnorjgyDi
j5c2vMm7nMpEB/xutjKFjEEgSmiBmIdAjNGx4WfbJ4yr1LkTXN7/yAZTbJrzuKTo
mT9MKoQt73GJzFs8B3a31CN7cHLZm2c2b2qNQTt/VQrkRany+k6JtfFvVFjI9e7b
OJpT3mDFGQLNmVwuvzuhWB5hXAbFTuEjx5EAgXsIFKDocYQfmm2vCOd6/30rEBRa
cl/eSodLk0Z3lyOJLf8PAvGgLzzlOkOBrZM2741Su/c7XgRRWkZuSMuSbtsqRV5M
vOGXwOFQF0aBAOHwkQhu1jQHhnO9s3cPUbE1OKXMU9li33G+UMrQxB2g5unibaTJ
Bs6a2Wb26CTUZ/sCnholTsoWqRV5ywgjDJ22FDgJmQU2ToCgaN7+/rX/SaY3X7lG
gib2Na6kx18ZfrrkT3FP6YksMKGqOw+NLFhU1l9Ho2MDmeW8uxz1gXcyaG+kex04
ImmHJ2Ux7lR5AtG06kdJZcv6l86xRLqg3zlxA8QqtLqOVOFhpDg6ViMkEX/q4rvZ
szg4tbJMQHCz3uhvabepnaw/wSaXwcISoS0WgYMEhOKUQ8p8TbzC53NzLZqkUcZB
vgd9p7lRJX17IcA3McAhD4MCvbsIxqz0mORIBl40S9kzXDTzRqdwIKP8LUStX1Ja
BYD7dEXcrOYc9Lv+Pvzqw/56NOwBtkRswtNKT16fWGW3wHdgbiWWSHmwmGoePN/C
cKjock0UpRtEuvlpcoazc9RtPHBCRISR8fqMMNVKz6R29t3qbtRMmZ54YBFbF/5C
4Mym71eMgGRXPr9fctzAqsTmnlGeYWTTkmA3b8sICpHRlR6mvzDRUVBShNlEz62I
8XqRVCpQJEbw3/53k+jtaUjIV/2o6THf/3uwKJgSumrqDrgSOaG06kTgeXO9unO3
/2KRy6tis8lNycyp33gepog8OVTQLArxNVyAdLd2W+d+4Wns0h0thN6/lq59E1qf
yblCuaTazfaoZEJeRCMMgBwQ8DvI2A4K4dMAtTUb38y/UgkKw1LhhCI7wNSRbC/W
w55sMcgwQlwPTn8FOfs1EGn+0+oJ+HSCMog0T9sy24X7XccZPw6Hp4R0JHd3hmN+
e5T8VxDF9WsDYEUFbVV6iCxjZsNvLPh58xrWGRhkl46t5JTiFyRzRIY8zLB/w2sl
ISQB6amKtpVcCuiCHJhZl6Bd9lupyppiLrj0XhmnVVwn2uoYQKJWOVJkh9anGZcC
3ViZC918i0AbOoB2iVEsR2aV2TForXDzU+otSkcquu9MTc8lxCFf9yCqoqM3NW0T
47ycG3wXPEspl/MhFO6PBXvI7YDqAXAQmMN5hUlE788FTDMZQtrVMuWbwSR1l+kj
0enqja1kiOTMx51dGLHMOiNAFCffebhkCE3o7wCe5C3yQeedhIzVuHdrt4zBQ7r8
gAKHC95NEPOa73zBTQDV+4gSH4sB2raE1QP399uSknp0XS8lLqsCfwJ077oYa1aI
9LwjsqR2SFmwhu8tY4y6ncs6oz6gRqAtpkV2PuRr3IYeMH7hde3ozraVnUzlVXYu
DeCFrpVR3U5xR1UxIfK9L4sQvfUpDU27shGTri4lidhUWtE9RcjN92dgyNWG4T8n
7QcsdRJcGhmVujSWFh+NkGsQNq1n5a2PtW05QTd3u2otNnI1NO8Tv+4f7GkRoppc
3GgRFwI4hdLUR3orOpqWJ2skD3EH7NwS/Bza0m28a6VNlywcyRCdTl8Fy5a801Uc
txkctL+U6GbFnPwoOSdU20DpGRXJ9JYm1ETQWypHaHgTSZdJvJAcSwZdmJrMp4EW
Y03kPW0k9/88JR+kHin4ZFrVc/lx4dcoYI9h7vQIhQHACzFsWFasJWZxKV5yrnSK
HrssVStjnIFhjAcP9qqWvQiHjKh7+Nk8Kr3ZqOfTMKiHeg4s/5jmFwUMS5+oR8KO
1Dime4de4ij9FW/acMdo4sg0cEO4TZhtj+FKnPWOOVMxBIfYQveOQcNo0vev0dd7
bLA8RIt8xb95aHg0SoNUAGtFBBn55qie+dUFXCf1A986xpAHWyQnxtuIc+Zv0Q8a
tbPUStxkWEHBQuXKR3bIFg8Hqyww40tlUTCwlF1dJjBtiWIoDI8kudG+bDKDqAo1
7xWnPS0OFqojnQXdnuvPrcJVUXAJRijaMgjsxlDgyShIVoglW5AfIdJAbkxQOVEx
l+OsqIR0/cT6C4Liu0Sqs8O5sghQNqOuWbbURgOSyVqc1868CKWXunG/zZbOsRKp
SCwHLpPyWLRnH5ivyZuEEn89124y4ZNZdcJhdfBJmRAQn8qWJwm8FhEEbD3DjIIg
6OQ13QgzixJeRlty78ygUthipQyFUdMo2/okB8+3My5lB3UUaVWZNkbZVKWMkjdR
mL059qfPznIscKIrqOFzGKIrH3OWkAb10eV6YTHkwjdrt+KsxE4R64n3x6Fy40j6
RzfBJgwns+Lhg1oBCFz1meOxekUvBI3urcm2bbpql3DWoOcJw/+cukyJzIa4wOJ/
DIUCmZCxBTUiLWftb5Iq9FwwiZy1bcby6czxxvpR4T1Z1aJt4hnpZw9jLqTL0sJJ
DF5Yr+JgYD7bWh+fLXxOrkyJk7Er3biAib/bCyJD7X8T+htx2YMoLv8ObzOtJm2B
nUoeyDdPgR0Aggohx+ZC4FFZSHcZy3DhY9yv8a8o2QG1kx86dUlrjlXaCR2c+sZU
Us5+d9fjH50ksknmOID4yXlTi9w3swKSer6/AG6espm/Efnv2/bxBnLCgZY0wmRn
G2DBcI52RViiez46S9B5xPlPsGrj14r8X6t3/B6htQ4KiYgkbaGWEkELag+s5UnN
jSLGRdt7Aa7OaTTxfavTX0LsQ2U1x3qv3R4KorDA50u0U9THojb4Ih4kE/sXLh6D
DYjQ8vw4kHyvlL7jAexOVnq2pkqJCy4dKQhUQYsHdmMvuDEXqu4haehexTB9hrzB
wKJ1jOXBz67RS7E6wCqTo8J4V4j2h0sUBH3WpnPFeqJnGWiYxmCyZksYJB9S80hk
lIzG/GFs1UAwD9kmshSsZACbq+9IJQpswcA1Xkn4aXUEqeprlpMAAbpNfyFvRNRo
HGOPxH5Oi7nBtDuYsV4BrvgmzZ2PYjhFO+u0ueGDMzbroWafozvIVA+pseJ8v0DE
nLQZSLLTHrgGz8k1L3I1aJQVvl/JPl9VLMuJsV/1COaYOmvqd9qkiNrfbqr1T2or
gxlCaEqj404SMI2+mVcyzVdyX7ZJhBffQifwdEspHxfAjK7B6zpgoyQMXy85tpiQ
Nlz0Qy65MvdCaoMwxhXu3XjfJtI7Ys9dPbuLBu15U0WDuMQKC+eoqL2T4yE/LUNK
+vE1VlgJW9ZPwcM8UCrnQxmTxl1h5l1+xnCVc+DRKYZX+gtcJBM41p0Y+mxRKyNg
S3XXDqNVkjLW2kVfzvhhIq+E1AcXsi895yccyX2vOjMHyXY+pjhppYc6HR1cwKgI
Gt0BP2Mk9pt+uqE1w8+zGSYcHLnhfYuMy6+MWn4lk+Pnp0WB6uYuuPPvuAyK6aBd
eyZmjEO+pcAYknHFJa4tmnADvjT+PRVICKeHRwJjEA8VUqbqGZFNMgjazJOrrUgG
ZG92A8W/hs5PynJWWcdj87ktKYdlW5/Y8yadOFNUtW2Em6sZzu7xbSVXL3TVPOe4
NJYF5E2XSsBh7/WdrAxeTUhgyCtnUj2J80oA5pyvXGoFHE7n5sdU89EHSmwJ6jHq
QVlDP8PUy27EpfZ7u3+XnQYnJ1oGLnSfWtwBiicnihEsjjD7eWQ06BzhKeMRkr1Y
hbkBJ4Lprb36PYEY5dmpc2ql5lgT/xj+ofq2sG0hK/3q8Isp+zrRBFINxCYDOdDP
miejatMI6uvypSmsA9L3XH5PJsCGimC1+6axzNy/RgbwTST9GdyJlAjQHe43GmHY
8sfqS/YKToJl2aiQlp+PpWPyQhhIpB1CVtH7Qh8KL2X2wxQEWF7+EOmFP7ut9Q/T
NUk3tIDnZ3/4gGP8IydTBXDf/RkRU7sV2lydHQuR+TSi8hAya3uLnUoZRnIcfjL1
7j3k8TzipOo2EB25/mGAimJ+coe0OW0LXsS3ZhizDMtPGU7LJaiVZd28cXBuhgZQ
KiRS/bZ4/Z9U7OZ8qQnpLSXTTLqAldnDNPx4PLu6/zNpIeo6DY33QB0E0Wi77WqZ
vbdhGGNXczGFkzYFWGgdM9pPqEzJqj1elaVYflKGlI+BaArmUxCS+Irjhr5Ix5ZK
6ZkxDAWqfRKQa5EWTmH1ZNTCSmMg1vyj05UW97aTq1uLCt66JQSy9T3RnOXTXGVL
vX32CXAngRrIWkMC/+ct9HSGcz6st9G0KrgUocrOEtS1zHmjV/4dIKyfkv8RWkDO
HkWRz0wiBva8zruamEVPCzuFEnOsz6H0nBWdnLT+efCLqaPydsYxd2WULPe2GYW0
Jm8EuhVKGZBBHLV93roKiWUbOR5FmlRHRhOstu6tRhQ0NMG2EqWrPArGBY0zi0nr
nwosx6aAD+j35BMIKwYYZot0SowxZIJmjhxnw9vmeSp1oepJ5CGjesRgNcKMiLpx
v2AJ0ckUhDTFP2PZFj6hsMaxbUZ1a543jTj9Wu4ckEP4xrwr03NqnBK27J1QtJwH
t6QRXVjzk8HFmFmyrMDkAzRFc7ehibWRWVyVL7TMWYdcNqq1Jug8MwuGh7t4uFvh
q5MLJTk6X6BZwWviGjwek19LzT8z/9+acaTbT84YuAxi7nc8ifL+HgK6f1aG8l32
XcYxIkyaR9gLn0IQXDFQZeUWHyqShdot/w6RJ6ulg+J8D5JIpw0BGxqvv1+7TooE
BnpdqQTdBpjCqaffNw7WRAKLY8PbBLDeRRuBPTt4LGQKz1rX6YN9AySygJtS+giH
6QYXSmorbKoz+1tsYwvy/qdhM4wBAm5GBTsO6e8/Q/KFjkSDpVFlt2sEm7EB21oU
Apy1C3ERC1scqc27zeBpmDZDlp77ngfTx7e2SCPX410Uyk5URqQ0Mf5nA+VX5tOK
JNctBXOPt2EQ6Qtg9r/EpWgz6NKtzYSgJzIgJhHWbze3K0IylLuC0iTJ8o1hRFYt
Q9nItwNX1TsjiSAgTq03JmHi9apqsvc7DmFW8xhhczRQwMmfC3hCQ37yEEVsO95M
ex74cUh3X0op2ZlYp9q+jAhT38Gs/9L6JrqKy4b99x04gqFDvZzPQ8Lgjbml00pB
bJYZvDbuL2lJBU5TfyMItR2qVaVFQuWlrlJV7ElTyWgTizND799qU+iHYJw1mtWZ
ZadLVtLBcrEmtaWj8nFx+mgdRE1swl4qKYGVXoY2oZlEefhuT0Df5ZHdb5ssrHQm
IDaaNCddFSON2dYFZSjqW1SW0GlF9l92obbtq8WwCKWbk49m2bG0KnA18FXfpiod
cJMbdjCC5sIoXnVhodTdd0MZ8DWKBnFzK/rO4N0mMymGO7NCOuPzcSMBaij9+Hk2
dR8fk4YXeJxUg6F674MFD8E9zJL4OG/aDuBM7FeJn2LEoquCpn4sy++TYcQ3HD0Z
3dr6IV2YlcHPOZrIzl8XwkeF3JNQr6ZU+Jrt2tu5rINcVRNXVCQhhKsGt1JwIip3
A2nTAd811RK7XYvikwiar2q9eSfmML7TXeP0pYxgWto+kov4hPZRsFpXCQBoWD2n
yHFkKP3jmly2DvrrXex+Y5ssr0ph/ovGuug/ACMwAKjBnDMIo29z32W7PviMHkQ4
wWKbfnf7x6Rr+a2TkJ8xXcVzF681gwa5P9jz3L+tV1Vmz8vhbt5/W9rb6zmXrsz/
6SofHKW8qG7EAOdtYjvVRVDxENhXcbR+ZkU0I6uyc/+PwQ5GVtFC67/cbQbld3aH
W+ilFczGTddcNg8L9F2TyoRM0RA4h2bJHJeMc6GWL8fLNQlJ8D9TY7i5XDX2cjQH
2Ex4Ba3RGlMciCdfFux6nOcbswK6V07Y0oHTqsZQO7YEheZSPPkRYhmmI879Y1Xv
Znx3ynHFVYBobMzkCNlUVhoHHcJ1/pNqYjtMzzZdexAQUmL/6dsXRQDtoW2KbWRV
t66NuGAPduxj5iLmMq3x1FUNR45VXgGi7LY41Z6v4O0ROhwdcQ6v9GYzvzXZ+wZH
nHe4y56FDGy3iHD9rGbdasEJfOs16EgKm36Z5QUT17GVj4tIQ+6ILRkb7on1ZGY3
9Hkn/KTI9M3C6DY/jGZO26Vzd4WUm0kUoKW83EvnRG2mNZAplQTB5ZSK+/+KPtcQ
1LlTMwPZ1Kvag8GYw03jJ1v6R/fjft6xJsxgqmtxAsWclD8q1JPRgMAlIjz99G9q
jmSCgvCuocaTXUVenFXbbx+vBYSG/yUAcJVjs5yjtJ9iJGwUnekpmzzjH/qOgmjP
7VIrr/xxZDnIBcYY3yFAwxhMYHwdtV0nYcYO3Kmqse+sTJv/q/CpUYqPS8deNB+s
YRcB4v4oIvZsGpRaHOrbzBe22ePo8Msw8BEffaonmI1ZazPEDbo3hyrjAAZwLfNR
dUSyDcq8+hX6L+gDS2W8ixY7wcfPPZr+h0RXXAmDofe3dljst9f6ioXyZhgcGp7l
i83htn6ZxyQ3Tcgi1VcW1TGXz0VOgf4a5qpEMXC80oXRv0eOFHEidqvRn268ejq8
hwaMPJn7RUtY04vCSVanO8qdxLf8U5D2VpVYBqpZfCX3MK7ovSDoj0Ene5TIm3Vh
3GTl2VVFiKl1zViHIaiR2O8kUTJP612RMeqOht1xF62D1l0Vr41rj+UJsMa7fXCV
+3SQHJDR8wDsAK/ggwdBkIdWiNgrRzcy8cOIentHVIXyQuGC7XF11lhGrmIvSoJm
ODxhFSmwlPz2qGJmMnhfsvG5lBdqJdcR3GF8KyTdHMpqPlMOkTl8zHl6xhHDiXlY
aJS4thE3VbLnqG/lazYWLto2xojXFPtq0m9CdlwEUEjOFqstYIJ81dpAY3xTQURX
AnioCVGPXIxby1TiBM0y9xJjes0d4ThoMuEyCMLnN3o0PT03iEb7vFaqWF9Xk4cl
Ylz4oCWlnMWVruBYEebQsT/ph/atJXHr9QVXXrTuueorEDVhsy5upI3hGW8H5v6W
qTz0JzKnm4V5cbfPp4UW5AekHyyfG98TdC3r5ts1aX5xS9Fze1pg49NNgvWE6oLC
tC1E9Mjut3XjOufZyvYl7JLgdypKExXiKctHs1JyE0kpTPkOdK6jCH412gsFkvYW
n/kH9Qepc6Fen8l0mJfJEkCRTflJtaKwt7uQQ9fB1aDvp8ypdYYETdAiGiL//kad
NLGhsytIMElswNxw0a+c98066MnI6xGio2ZEtwVyx9HpeX4ahl7Jq4EPkON4KNQx
JIJg8AjOz/ZZuTWZ53rzABBXC1Dk2jRxKr3VUrXqYcUtinyWFbeuPyS5nj5vKg5/
04T7iG14KUVIxZF5k9i9Ggzn/D2pVxs8ykedWMzLseLpCePX7iVQTW2ysDa2Gyaj
GqDHx9Nb3R04D+b1FNZpKHdy1ltNw+p3iAi5sCY7Jqt0n7vu9SEsYxB1Dh4btVDb
3PDjnS+F6yK1IVt07Zz/f1kSBr34szAruczBOY7F6Mtk/p/kA4pfch9SJ7P3rWf8
zQpDmo1a3kMMmIZa2GfkMyt+60kazdeFKD1GDseAnLfB3C1QAjehwln2bq6sjL+G
vPr1a2O3vSJIaomXo90JWvVzT5C0Xdg65APY02+11FOB3y2aZFEw50xkwmdAIJvd
Jebazzl1VyuN0hHuWzN/yoFFfAg5CSLfHQvIIFiTdcKgwKu3/yuPQ4Ypuu3Bf/vD
4Et+IRKHNu04C30f27O4PW+jv2+WRVD73UerfVDOnhkETRGCNCXw161paMvCFjhW
1rWOWBbWRUM4bBeM+EYVJ6fmyQAkZz0jFgyBDYfplvgkdJbbHwjGhRulex9g0Wd2
daiHaBU+tikvXd/OFdCPgWEpRWes4NdJNf56ChlWjCGnph8JW97u2PihSWTzyCEJ
idLPOmeZ2Mv51gTU2wbbZbq/ULBSc5OP4mY5ePZUSBt9j/lDVRayQJOd4UHNMUe0
sbTQjllAXs7UDhitsfghcxl/8ikg10LoVCy4Kj7nsytRJIgUjRiqA8VI8id3afIE
CN3mCPLqmbzK5JjExAGhijr133gGDMN50DOykYuhklSMaA3dq1EI27S3H+eDbouB
FQCYqJLFryCQ0mVIPVDHRgSK9NOuaV64IzdpQO8rbYLwontnwCvZcNy2pHnD0Cgt
PaBW0VpEJoqk6VEnRFQZqKp28+a851vWmItieZph7IzHAma0QAdR4Rqa429DHonQ
pN9mybobVaTXvjditEmfz5y2rInIqO50kwcIZMX56dGTc3yVGvr3MLS5WD4lVLg4
7xkaoxivD2iULOGv+QZFGnS6vMsmaxETvMTUqfFTAqBXZ6vXBSUnCFGuLHdwr+2O
FrXZzLtKl8jFvNboCVUPnGDys6q5KQuIR1aZCMG8c0ildpqpcMCFdMd/zrA0INoS
ZV1G0ZuLoZG7eUpIVSpdzFWFqm2iBEECxasXQWR823KldMePKzMauRjvjNHifWfS
x7m8wq8gUbBwU8EDqcHMk0xJXv80CWQr592md6DfGyi3+v+nYNwhS8RiBQJAkhfF
a3u6Va64s96kKqx4MXy4W5iavNUwYzm7K3EzW+PzmUzj61OwcsYIsyFEpgN1Ht8Y
QGT62bPtGN7mi6fTge9mq9LEq/vBsqWumS/3/BfTnXZncBbu7vN773npCcJq5W/b
Ux4lbYpD9q1US7gDkTT+W2Sw3UtuUQSy0nFRfJgh51dqc5R/8OpFSZQ4lJTqyY//
mrrt6XAfpFY4s0MKAi9y/ERiMsliU4UL/5AZ1F/tnSblxWMnW7ie1hykcqbvOodl
L8zIp+tShvBTVRRYNcjT7oQsuGds6PYL3SrIe74K5elFgKs1vawbDwHY7r8c3GjS
3et92CbSSqrtp71BbvJJ+dxvnd6r52v7FCYDrhhslaDTO2l/IvgtKFlyG2uSdrTH
50S4v2KaFVbUwaPDYFJYLlqagApniv2XHjdAMfn2y6kY1JB0lvQMEHB4kvdMuqE4
FovxDA4t2g3vnEE71xCbuTLW0rVT9Zm6nZ3MarCj2t9rBDuC0wsbeBGr3b6rinWB
vFqa8Nf0aMtxtd5+w482NTe697xSa+6RJq4Lh3l8ujvTEyAw/yIECDdMBQv6D1ZF
0Wlk8Afy8X0HaY0pEMdtfluQdSpxxz+V8GYtpSic+BTTwXSjG5CMPJDRFkAiYWai
byINnboUWjuqHGNAQcdEGXmSs2VmB0yFC02Me/RdZEFcOA00BgQcWlvKDDA+DhR7
z+x04YdVDz1eYqh9ZN8uT/9xTixqUn3X3/+uwNnreQCHcqH6ra2FdzMka6EPatMu
a1aShHM3m6WB8WtcmLf0sY0yrRCxnmJh9SDYHDfHTEFAyZVSvrzWhzCN6wK3V6Su
cTO/38pEhIOffGX12zqmZKBF++WMfagF2LIBqGk7EiIRcivNvh8/axfiOazco3ox
RLW4eWj3OrSNL+yzEmqGxj3bRs8W8AFJV2bfreDCnqsbzZo0n65yypPHDeo/Xd9l
fUxzlJ2VGVSki/GECdXeUkm+dNRTbp5SMtUKeRNxchLz3PI/wvNrsGxdZDjxDzVE
sEftgBK1fhKbWTkGZeuCQEpu0t21oJ6nNb/nuOX/Zr1xp/NvMKgwTIM9glPplz13
RD8c2B3ppKMIrRlwo2BT0Q09Rk2iDKvhQfvXmQHhAVRii3IIeB7pPvfRuICCzkjJ
0p0GG5hpUxL8gtqRxqhbaFSmznbt3ixGE3j7LoDthtLI8MzivtISLtAgwDHe0qFt
mTUk0oBVd4zdWNYCwQSvHK7RxcwybrG++ISNC81XKll8XYSwt8msvhL8cAuJQJUY
SLWRho7x246PknQHWCzhnnwJbFPb/2obIQ+TmLakxZJJTShzXICzJarBcgzq4WlB
bQbdGMiYcAXJotn5C8yRJpqtCSs/un3LGVQZGx3y70twkCXbzdzLLA15L69OPP8B
l8+XBfGE4lU742ARSWZN7xg+6dKToa8Bkav5mKb3x06Zog98PORzUaclLU0tSLjO
StHCjhYXN/UkdRDyfX4n1fZ7EEUp3EJPsTGoY5oiuZaKNTs8xHnxvN+ebLEvZnlN
I+np4gj3LgmVPQzAtjCDQgylU18DgJXSRd9eQprUOIf3medkYw/wIjuN6Ijo5oMk
3ydegRAamuoToFd+IOwyOtrWDBmN2QCkSjNaeUJ37dDEQoTKFUV8sHXt3RQkD/pB
0qompWk2rXAzMT4/07nESkYtk0GSgtD/SOIdejUJ8NLvlPgwHOyR+ReKXtR3cCGw
dvP8vQr27iIiIR88KCTXgHyX/7zQQZvqCZN/IPbN98Vd4yv6opdqzDgr4SlOmfFA
pdUea5mVHG0AAoB4lgkUcV/F2oudlS/X8KSYtcd4+ngrnJNyolBcYZkZfRbdEswU
RVg/KFOoM8xIbjUnvUiT2Be3MCtxGg4tBpQ5E3nBSmJ1Zqvvxsq1jrTYp5KoJz4C
4xN8LElWn6GRXntsP77IGELoPCzc0Qaqbp/4xTWUWz3DHttOkw5687ezeDqrU3ZN
9yYlCP7KGHzmyyR68pP5UBpqSMvfktq1wBnRBag7pH3Uh/481rLLNGpwZqvIACyE
19CJI4wsyWme30sgRIgEEYP+1jMdFPQdqruYpOZ+Fyem7ERtF8Jb5Lb1WdBpCEXO
U5+pbQ2+pBzvVinL790Bs77EbXVTfAsFaQclRhoi4k/dEM1dwpYwE9LBYibhk6hO
/j7bG1kFg8F/t+zN2A+xhwVBVWdbfMpChIexK/r7r8Sletx0sI7hM1pEBnpuvnHG
GEz5dQCS0lEsetDerYgZZJ1X9/amvCgkULHlPy4lNa0ZEerL/FXlJ50Vwwfga+it
MnOFALg2RA2pC5ieeCShS5Mw9FZndJBJb6rkzUK4tFhGxK4Hq6LLYFflG0BrMipt
o2LWSH9G2kwFrogqv6GdSBygkEx2csCyZtEMiNA5CvzykafhPdtIv5c3/zJR/oFS
oMIiAmsNN6IpplW6IC9yb7Of713pSTRu3mGhQUR1TfTu+wNOlQSG2b/e7EYQ2bKi
ARKQSFYljRUqLkQTJLpa1qohYIuOD6HAaUi0KK2sFRA5aroZiEyrhyxc7gryp4VY
G9xfgBIQjfQoVOdA5eQBVg+HCoX60rbewRdly79CTN1ADL0z7ZR/msoDlqN4/vi/
NB9uCW+UJ9VlMNo3FfYGOtiEahq8+aUBNAMp+2ZAFclr/HPA7hBTCozgOGwmQafD
8T4xT+NQwURBuPy2m+LCuxY2eb0jw56edigNwUF4AT11D1PM1bkjYD5huUEWVyJy
2PCfuj/D9ZqQ+p3T+dEFGQvfNTAzxyWhep/5XZXws0mAti+i6TQZto5Z3ZaOsQ0/
3kon3I+RsBHYdAOtnInSAtkeBhr81SnmOwBGwFGhJSLkhvVAT/v5pVeV2w/EuZK2
X+otgBV41kr6tj9weKaKmwoZTvvxqW170TmMs3V2CaOysidQLNRyh4XJkDF1uKOc
7sKDsCeHRyNv40P8PwbyOfUOQg4IXoDQ8vzM1f9C584Oq/N4m6A7tvdBNOUHvbgM
avp3/qO3bEfWDLNcgVOqK42u4V/lTSy6ZbQpgC5ReI3z+iS9FPSjkubepjGUZ7PE
V8dQOHGk9XQA2PgPqXOhGqmYiSzsU/aQ9Kw++oxxF+88ogg8Hpyf297KUE2c+/mJ
+9MVfAnvhb685Y371S6Ct+bk/4Ttpd0pE3pVMcZM/XrHKCR/dJu55LrmUCrPFm19
v3OLqX2D8405BEhBKT22i5bdCLEnLLb6aMAB5a2HUcqmFPUpWnypVwCiWKN02SdP
DtSGLAwhPmTcWFqErptl4zOARLMNC0tGVe8ejDnZkWAnI977UI2wcwdkxqgkaoz8
G+lsBOY8NClNsPaPQkgP4pcMQR1pnCibeteP2C82cX6phsbN1tKt3PBqlWmUIsMq
PfWFfTezMMRAH3cuvmjHUwnBsJvQFRVjlvgwKjL65kfdKoSTZKH01i8QH/gLkZyv
KPG07fObAoP9VmD1P5AdFJ6L0tv/r0EnYJOy7fpiYnuHJ5mies0ciWNKg1CHBeXY
JmP6EVk7s7beCbpDwHz4uMdJK61fpr0dvTWyrZMplO7OI7V+eRSe8Auy4XrlxWti
7AMcP+74BLDCixBXYDo+VBXMgFxudI8a/20VGn06582Qm4hATJ3FisR1jsu6PDgo
7AnhuYwe2GKmy+la7ynO8YRsoWja271UE1w66vpekw+n31S2RVHlRbWOiOJ8r31j
p6/OCLAKulzm/CGPk4nMcFk8h1lQCA0uSyw1d2IhjRbgKEaNImVwXxzsLiT6Wqni
YRRl8L+kPDYlOni+EKi7iaL+DFQfKhU7XrzjY5h5Yru3lJMS7F1APLvdgSHHs7Hc
qWMVzBi4YES2snbQp53ocAXrBiewm4MXZbnHGibtxfcDFAcFFhGEuJA/ZlEbo4Kh
6a4euYJhA+QmFWX8S163+KJ80XUKo4v1/gqN2UEwVNdhb+WLPTwSfCjgPG8DTII2
t++zkHtNfbMUhcL7GiXDbhOhgjaHXAgUfAdP2aZAKb+06n9c8dH2RdVF8GTQ/99I
5mYbQ7ZU+oQsWt1Iw0D9sReBnKwZWBx66zFJVWreHXoBtPYMJfty8yVooAzKC6fI
g3F07cS3hwIkI7v8CvZh4jAddbUYbLFPRMrzw3MiaRlwK+TlNY5+v0YxVPGZ+775
xJhb3SN3i5HmLx/VVoECI7MdA2PBqFpWUFmrg770bpjwL+6SBW6iMuIYyMCYxaw1
hEb2az6zpYqSkpIOhtDH0wjtjZF/d9l8xN9SiBcknYC0cQDd7JXkFFUZkB7AlYED
KuxWLFBH7Mqzq2lzKL2QjYy4tSGHXryhXYqwoTfOabGR2klPQgAwx/zI2g9tThkx
C3QtkX7F4ogumSh3zIg9J+f/hoPW7rrXyBgqtLPxA7uYNMtqcAxHENVVYeIIU89t
FV/YRnzikq5DMiu5HD8u1nt7zOpjfsjKQl0Zw6tW13Y4MfXEboyE5VYoaV06ZpTi
IPBXT/dexferbB1/ecuMGNyebTrJ7iITAqxcsNK1RoVn8RHOZ5pxsqzRbu2xSCxf
ze5eRteD9ECpebrCmosDzoSHkIKPIKVX10GceAQ/KmGgfXz1TYD+dVBkJ5lPGDAY
mx6RFuq0I1Nhd9CfIKXIVGz8Mk6+Hh1NWFgtq8QyiZ/u2yIhZP1S5sSmhEaOONcj
K8B8UK/W2AJFBAIZhdHnsQlOPTqA+4OV+Fmua/fbGR8EDJfJoLKxw1VJKwY8mTZI
k4gEykIPDMjcsRrBRvMXG75Ryf3JXlQ26ruHSXJ5VUhIDGwbJiCgkUNYjo2lu3M0
TygAXMVJAJjNyoaGzPqJzza8+d2MZIJQ/wa1Pr67thK5tLA7umYIkS4cnZxUDWbY
1Z0d4VdhvKydkrUdZ5k6qOuj1l4W5SB+YJ4uCU+lU0EYtP/tOcK07nscuGCYJVog
0l3MQmibMz9yhKEdh/s63Ue3r9Rf9e6dhquxEdSBu9zjyp2nhwxl+wSJkC7q7W3O
CTrME0TrOXFjGHt53qnZ2ebdK+moWoRIRKEbm5dM3kZG2IsR7yeVrlaeNGgcjifV
7JyPryVn28oBzaPKscVLWBn+9ymPB4NHEUNJfAtT1CIKInI8SCHGYeJ+DrqW0Fi7
y3LRMXUt2ka8WeWP0iUdjs7nJCc0omhpN84QgVd60nfwRcu23Aaccin68YMkpqjv
q+Yfz0jlfvpWQA34gyzkywS2qMLmf9nQJwdllu1sPKNcuv/eof2x1QRpyF7WxQLt
KMb12+AnAMQwIp6F2Xw/LvlqSBDfm+EfOODimnicoWocsx7nfAAb0H91ES/0sCTp
2xdc9FsFAeZp3MMntmzFF8jvSvPso7kXoRYhffuQl7FvYcc23zRu9VJMwbPG01gg
agr/I1m5G/BoBt2nwEs/9mwY3rMNF84xgqhUX3J7qyUsR1CrKqzFIaI5+pHEJlKg
YvUO18NaztMGojmkEvTAKALwAm3c3j1Yv9OcskWfhDp8q054Mvm7jUyJUk8hJVvu
51MUVMS4qLUOGAVOCoJidrlXeczkh4wKWtUy7cfwG1HZ2G43EcBWZGuUoCK0SK6F
XZf/ZspA4htZVjFHH3maOOgq3ZnFH9+975w0tZ0uniF9nX0o5D1lIGqNKAeMp8bb
PPp2IizyTk+7566t1OdZiwqcFZOb/bEYk3Jxc1YoMk0phZlrdXTR1lEGUtS29K4f
Uah27jZuYKwEw13Te3u0uQygghN+3NmfjxWJBNXEY9fP/CufO3ZbSym/VA8FEmDI
A+8y7Wkqb3J7bvnKofcUUrOYBrXH7jqeqZo8G7OgCKBfgvaayNSUCIqHLavI+Z+G
3ZOJHQp+SfTkUwVn0bDUhwf6cNCkF/afGKIH4dHK47uLSIGR+wWOm/fBlQ3kSr4n
BQ0Ak8BoYVLgXVa2gsubMkrQa83+ZKwZfkV5b8sf/7u8cDRCBVMBVPKhDKT36COp
AghXdF6MHy4NsB9HrP0flVd4LguQaSWmMZrZ8gM87btPstYv1N2JcRQa4DS0oq5T
csYlt6ZPMA0gjPMrt5ONLiILPeQ/g3gm3UtkMKjLW76yo+lEoZJ3wQ9zVhLJvqTg
XxD39s+dxL0hxm1LQNadmQSqgWClhjPy5+bGQFd2CBEhsXOGt3MZmhWkt37r9qZq
e1MI2+WFF3Q2G23bQeh4dncVL7jr5G22dNvtkVEc8duC6gLwYTfrTZtV8PdMgFZL
ZaKGcLDoe+C7Q/SqRTwxfEwNsbFqneT4huIqOdpuDGFDxhtJYiVxg35zs02yjmkN
wM++8EOb4Yw4Zr03I3zlfNJUeEsn9HAbfMDQLDf8v9GmqT1gk0GPJ1csp4isCGZx
P8U4CL5y41NpIkTyB206V4ceWtPzCwkFhP0SnCsHn3VlE0Prr7oiU73MUQvOEwtb
rKXumyR/6xkloech8BpseJH3aPdKTg2n7pFJM5x1mn1E40CxsLmhdRKGtdlMwcRD
VrJjAN0o2X9C86aQ206XVCm9Ftm258crgMx1mSlngMiyjEtyizInPAcTl65v9+dl
XOV63ndqeN8qDKJaMYj11h68pJ1uBDGx+Fy2rVcz/+7ir8RRstcTeOlGx9TPp+Ea
xODPm0wjMZx5IP62G0KAhxDtjNx2WJ765u8rgD+DLnMlXxCPMoSD4WkOCaLwkxB8
MYt/cTX42d9p0oEQQSfAqZ16JnSXFsTtlaP14NL1se1C2Nu1kG30dvz8N8mOr51n
qTwA9kwclBIOVXjAvbRNgde6pxgO9J6Sj93f0osy6JeXOEEbH5jcDQctfnYX6Uox
bEnMYkC7Nxn09cra+zV1aasDsB6t1NbrYRMTbQgEAIqpo7yDz1SxGvghKOo1NGbF
ltZehhKZm01OFEo8QMohjRa7ehIrQmkrE1QVvOZujc30GHeWwYWc0sL5VcEJahpL
EVo7krLuTsxkS1eIDFZO8/4R4VsVhB0/8LUFF9kQxs84UClTzc/ruHlOLwOKJqLP
sN1Xg9yaloJlvvUXYIh6ux1Dj5DC4ptiiQdZM4amSVhTB1NdjN1Q4CHT3rkle+bx
QAQxY3N5g1/pE+gmqt2jvq3ySKric/WlQXkZJ+UYjCXw9JdbPyC3WqkibnIEWkYL
bkstKsMGHXHyWrdvnfJcFAW9pFhNoVM66263paAIqFjSHw8z3j3Y8zHcCtrxbT2o
bX0rD7p3ZxxE1WBupo6IB1iO5h6qjpaeZrwB9ExMNxDcOB/jJvabDh4amFUY4B07
gp7cJ6/kIr7+IKFh8UNzEJABygK1v05Ac2TwnZpNNSy80c9Uk9LyN2pfcsMIqkpt
qO/XroPqdmg/YKtnfoLJQf1x8RqnE//pFGdQLf8CNio8iQ/dDcJ4tJk3dZ0fmSLN
awi9wZveSmzlvFmhMuvwWs/tbyoZJ1iRXvhXT2g26ot/hJi2Ml04asJ6oPrdbThX
XuiS7H/9S12oluI6Tf7/GWdWF5mxmXU81Z15XWNZewO3kuaL7rR6S1nVjVYosONs
ZvrdujunwBAvq35ipHYubd+cND9wW1Hqg7ch+J+HoG3S29Zb0lMmBa7yLMUJvIPx
YEw7jamAu510J4H/dhjN79ZGC4GsUgGsmFPLsfAk2aCjGq2hQpej/uZ9G+IZJ8or
2YgRsTOEThFv6p1c2pP8NmfsbZTb2teBAsbAfCpTF10YZORzQSl3HJAqELlJvHKf
lkKiIkaRatNMXkDHYSAtdhe3SQwm+2HTS9qTV0OsFFnpEsalk/Dv0ghcS2oHkd+m
Ao0Q49plYIGTCUjjEjgmt+iUBy2T7hMb674v9excoZ98KgS+JZG5dUmUGU1/jiAX
6bhMNiJ4GdWZ76CSnOsGPVWutnxr7eq3hRaM4UyqhuJ8a+UsKy+UcTB0jHWqnnIm
Lm/gkYfhvCA/bHLr+TBWCr12AfPIVMZtS4WOexWGmZ39hSmJruoG/Se6O1lKMAfx
TCuVeKSMhEYH7FClQYUtcv0t2iexTl7a2Ep4Ei3LN7ncqEezJxb+7Wug2KmmBN9I
v3JGEyDXXXNoipKACwknvbKU8mVF6COj5Bqad6J9CnTHDm4bqEK00E+s/J0HSlOO
bhIoz1Kc5W9kxGwqWIkd+Wtweg1PZisimQzmUIAUTSzUjFMAARDzEVo68EgHjASe
euC/xTeOhBz4vCe8Yi8mf5pA/VMd5czKD+qPN4Y1HqXLcUk+RCojqdgil2HqDH5L
mbSbJLoc8cPnrAztcSSPcPNfML5jgeS0bLEZ83G1OSyD9pCzPX8Ub7SZkH1kUsmQ
bjruLLpzT552kwcsIN4taaC2dteWMpY/Nk8MthEIyociybXKkBb7DpbH328FgMP2
p7q566EHy64AZRQ0PIKxiWCM+bytjxKF190SenjbAntNnIDYxOiilZUsquBeVc1I
sp2Z3m8meI+DW/FZTsKE3vF97hSp8tDHIgCFJzjga7yvOhLfZZaR8YctY3Oo+UbM
Kd8P1dwNC2EGK2s4PoDurdy7lTbH+C7A+0sjbAHzegsei5X1H7G9q1U1+jNXRsAM
HGW8ArmLhscThI/suOQTUKbkhIJxKZPB+i16yxXfoVKrAvCqmqyciXkq8P4kFo/j
s/bFG3v+aKookyK+Jdi2oylqXQ9qQ36OBBneb/QhTtH05rFYPiBTK+T5CNuupJOz
e6asl2eR4GBTjjDSWQlqn6uPsEdJfVQoMHnNNHZ7J81zoOgcbjE6opbfN69Q5L/S
sTO9MpnGbRGWN5Qmn/I+niJ3Vpo0GwcUMY5Qdkaxgr4zUxBXx4t2BNBTcWr7dkGF
N2SrwIAEuz1XYa8FZvq4kiJguc8EAqqRP8cc18DAnQpimcp6HVPmh1dCIflIO8gb
mFCZB/qKT2QZa1dmxmOu0grsEfTL4qokSX+Ow4X3OKsas9tHVuh2y2M+e4faU07F
thdR2RwSK/eM9frtACUugRa6V2+mq/kon1h4Jrvk/gsvCiRjPksBZplyUof3svVn
2q99EEH8H3agCSi6cqzfsggmSEge4BBeB2ZZ6Y+uPoDKoZkSlcgsYSbkCv/oKcxb
BmEh3dccABVSRDru9HTHj3rk6eGjBwi/xQ+cTl6mv47OfMjBuSGVjYq2VT5sCJ9w
IuZprzJ883DEesqruCk2nTzhpY1orULSW3B/NVHWXT/wwPYwQXmhBK5DZL/dKDgT
thdSwaWWzAqVA31AUIRv3hlLm6N0lJ2DJW2V513Ss08rVTEk1LWGrFqKSdYAtTfk
ESG/eLn+dlEg2pH4/qd59H0e+X4TwHprxhu6nk6OR+6rySA6uo2yVa2DqPEWxE88
6IkMEGJTQsbe0cXC+Hj+AQWhKe+mVLdB2P2KalKvY2sXPymBthGUKVMEaaSob5QM
jmpZtp9IVqtXbJvMLhiVdl3KYiBnBbHLtKOjkqj4RCby/6je+/0q4GVs7lSiyYSc
1C5pa1BjnlhYEV9C4Zhgn6Zr80UmHBKWxy7kCS8PqOGZ8jd8HX5tHbczgtVkWfGm
MRN/cTDSUyIQrQliO9X9c/SqKPBZBqueluiGTY9WrnKPjQr8t0tulFI5a9m3XZWY
Rw3eO54GVvoCRvaqTMvHvoI2v0jvzNCob8FkfyOWYQ4adLNJmSak9DaT7sL+Jb3/
QlQL2ahicIV9uAa693oGwilE6jOliV987DtPUvTB6pRxmVyGYKHQ9l1/F8L8fPgX
ceQ4RYnhNX4/O4v4fctt7OAZXbTHfKoPi+ZlTPDkO6me2m3p6SuNRz5736XV+ft5
ooOSTnztH+ofkY0ZRFnVXar9EzWjhClHlSRSsAQaiODDK/qTurY/nSKEIdGL3xKn
USD4EUWQj7bLCp6wghlin8QxHevO31/d1xrqEmHK/zvqau+WW1lV7wgBFETh8WzK
JmDY9LYvVZzTM7ApXtfNwsbt7NrfkhuuCbI8+PKjKwP967qwSe+hxZptRHanVEqb
O1Q9Y2G5Okzrl6RL8NlhOv2ywffhGGAhP2H+xfkSvH8ooAhP5NGSxTpUoVVCWDy6
X++RMRVlAqBOfc348R4tWE5mBHILivD41A510gNCwZ0F7uC5G2eeh2owO+ZZSFy7
oSJYepLwMTc0BmTxnyHCzIqYHzT0jlYvrkOlin8+bcLKTkZEV2nvLvQvoyOeORrq
FLliu/LeLrZgTFJBTHTFWhxvYYaHGFass5T88FyQD9UaefkhE6aNx5ALM6YqEVMn
XRTvz4V9GqJxdgIWdrfVu5LO0ppvC5wXvFgwp5/giJktYPc7gxYicVsZVr1DLbyu
pvChzofbFuXh+FcnNLR/nYKdrKHCYGIwhWE0ZjJH1qdByJrz7nl63soSNbN1T7QQ
A1jVVmSOy7ZbolHyzW2ca/4a2Ws5uw9esCN8tCaCtjmqPirPaZ3PqNWt5gnWu3sB
iHSytIFq4j1zW/SokOK6jpS8DKPb4G9sM2Jeow1zWZVutQELifNheVx1DMb8JdQz
c2isDckqmzDvI1eP8tpa2H6l6dGOs4U99ukPamcK+3ZXS2iuH6VA5j2kXZGeruCw
eGxinQiXgyJfp8D+rsfffV6RGgKfNwh6ARQIx+TSg7lU+A8YmLqyfBh1dk6QL3Ge
zqwyYkl5mPPSCEaD4sszoz8XHVWFB66Fc9AW/zQx9t+reEgH9nDbS1FVFl362p+h
NZVuY10fAJBAltRl851Ea+TEA360nvMW0Vb0Z9WUZSnWyuqmPj1q7fi4kpb2ixRw
gA4PRlC0qk+RzuAtaTIO2gWHnw85/bzWu9+6qG0bjrrzq6Vb5pQFti77OZP4CvgR
mAVtpYY2j788j7Ugrk9VG0a/wZ0NthBT1CIgTUncamXxnf2DccLYsnXYwwkjBkZ6
wOwyfAxvNYKpZ1Vy2tMWGWyNqTjVPlvMehBymJcKWWlRcwvSk52cN51S8Ck3OHhJ
D2ASuXzT5QNgVLZVnUWhqU6Ab36RdeN37K5epF5XWWutJoDOTFAYU0o+UDlSmmtm
775vin63WvybFVusnn77pT5VA0HubPP0UcYLitumVz7/4eRDLicSV4J30fE3BGiK
KP/5jj0FuJg6/nRtgjAJwyAkU2/sI7QCoY8n4zU1ksKO7apN4S6gkSwrGTY9u8l3
J8Ww+2NGzD0t3g6tj2/3KWks4xvtr26aHPIfj2MoRs6r11vh16638yneeNy/OoHG
ib5luKx9y3GIFSoiKLG/8K7ErxAHBlbhU3fZDqo3kE6VXhQm5dg/Piwy9UKUtln6
uxTpGrZGVJG8IC0M9QVZ5dQRzSkbpcuj1f/eYaap/wAa3WnHpUMmHcQ51XJCjQ5H
9TpI58jpNo4vQAVtb/mbuFDb82RZQ7KOuGStUWkAH3TPgC30LbzA1Ewxt0Vqhzq2
WgoOTNrCzliy1dQEP/XBPWHuMU0sMZBMOtEdRBxCIG3JLS0jrgJFtbx8Tzb+Z3tk
ziBd4XjgeQqKXBgN9IC3vXFzA570s7Ufh5udW+1DTV9KxWy1Veytjt/PeF9FR5WZ
e8/ldahkhnYurf1cWmLxGOCkJloGYXYJW3RHXa2cpm3xmnLgCd/0lcKSkgTZyqIa
EgiTCy4pt/jYCmWeg0VPTz2bhWO3ZYcAYmi5VrQhB9HHPlE6zcnflGdtnArXtt97
CQqdxah3b2UJVqaidYJQwX6by5b9hSbx6/kg6/Sd+q7Mp+YN6ljwQNxJJruCWqLa
Z3lwXRlg8Z8Ci/fgiTr05fPkoXVMM8joqceNTdAdQjWpAD/Da/50IhAvEkNZULuN
GRtX7ptbOhJvTdIYKs/JRBzbSSOe1zrEU4ygEqyXOJ6Cr79haaJScF04jDPBfHqq
eAxYIGmk+WoqyQuuDnAM/q+HYusAXE6I519sNJ1c6jUXOrVpwDHYncOuw6CWskUF
A4FieFE3/PozRBR9JHPeWYTU8eWbyf6uutDz3rFLV9WmgL53fE3xtnxc5Bo+3/cR
GDuxlR8F44l162KZxnXWYs2kDZG/2KeHTdiIamJMPPGsaBvRBPkcyYFQA74TOe70
CJMZkciWnAvRwOrHHReUZ9S8XK5p4PiOzGmXJLemTbnIwxNRwOBJgu1HeqiSG6Sa
+1pc3lUtNsnT7F72YZAe+FLwk9V3wy9sIS+KqSsXHux8DxRJ6no5ccERq+ksAZUS
wffaAtAaB5xNvsFRHllncw+E3Qs5+zDimsMc2zk1iBMfsdltWEt848LznbVpm2fs
ODCAHJuwyLWlB3PYqtMHcxOK063RlB63zMneINlGpZL7cpvJHG46Uy9cvr8PILEO
AQ3A3/lzCljmBI5c86icykWkW6pq0GR7GomtFXI987NpWHYJku5dOuQKGX0PSToz
I57R9eTv4laUBAIntsi9cvlJOJ/7Rf+zCFBcwnVAWhPvXdgciOJiNGIvtxbAKTuI
WAH4TDLcqnhvOaVzWy0ApJblKdjLKkM5qx+UsnVxNhGmUeosskWFtrMjeLffrmGj
e30KpkJ9T9LGuNOc95N2IG/0RAhDlMGh7RdXknW6hoHNBQFcLqvzMzNvEONbGYzN
F5geyIsxmJZ29CLWl09kznU4/GFfCRXdZQjzvp84XRDjvyjOQpyP3LFN0dOXIGFj
NMeKnIUp0pb7LiOFhPQOFL6hl4m0U0Dk8k/pk8n9RzAddugqEkm4AYaZylv4G1Zu
mVi/gtxtmG/zJN6AE9N8p/ho7XOzGOCIpA+yFl1Jv7BYUqWFTj4BLjM2PPr5ci0u
tF3XhQG6qDcqLP4QLM0hcoD7S/Y0210NaqPbpe0PVALYUQeN+JPdgxFRyMQ1SkkG
p6DroZdbrpHN1ukC26+4diU2L0fJd59oSgIUzfZdE86ruvoad7YVKgIgpdhlMJDX
RJ/xeEbSLtaCNBckDUeL0D8FDLFs/xIVIHxZxqxXt7P0dVVUXVRDa1bLM2lk1owr
kVcP462rp65CeqswQKxwPMuysjt1EyVgE3nQRPfwBTv34AXkP83x4KIrbzBpAzMF
vk+FnDSlpvxMshb+nJZUU+9HcZfGtOxEAoxclq3hOTJZc7aAa5yPttE+rfRXn4n9
FVivnDMdwh6Xn3QcWzKlRtcdJfKD79bmTtmzbjvUilg0lh7zb6+fyUMgTAJOjd5o
2sh7PhWKZ4IeIkVrt6COsMBb7aIGbKZOmcjbvadqdO/RBK4kE/4Kzp+CqSXyiS1v
fNKNJuNb9DWHcpaikFVP/+/MTlyk3OB7Wv9RKsrfO1bd9hpRf3aq48WjQeWCCV3b
p2Sx3p0svZ4IlSsQgfxIC3uK18DzfNHRxvh9VD7gCWI2zHUGmUH8NsD/Sk6ekNSh
pfyWNTEku9l8hU8Mh2iLUY8G7BQKA3632+gBKYydA2S7qqds4Nt/OnlHPRA87AHp
Ws8Ey3GmvYzkrehMtvKGE6/gdu+Kx263afaryM/B+7qho4Am71Oy/ZZAIzetZZSD
U+7D5bbtAOytdtxi5w6hA5Ip3WkyPAWxF2oW86VKUcCFA6B11rBhdQaS1Tzy6xDQ
X6ROgSKBa2RT21qK0QXiKiBoX989ATulIIf3PYF9toEVsXFmuih3W3kP6xE4Ahne
slDYB/xZsKSEdXQ9UkU9aFiC6LoV07TEyTUs7czmDFrdc8Y1hEyQjT7F8TKPJLEW
O45R3mAZsl9HHCgJ4sIIECOpVeHvWFwGKguV9jmoOzBQUaNGS8KYOUeaa1oYwcAQ
+UGSa1741gTpTpnBcN9V8Bp2LOFixLRPhTHW8bIcI22iX0D48xWuOCvAFKKNGfim
Z0AxURLOcO9jPMYn4huw5aCu8G4aWZLK3ZmuMkiLlxlvgc6A1aziFEE47pbhLoXM
0t3xbxZHFlktri1QS6l8A/vA2fQ74uTmKr74o7ySe05LZHp+AWZKl72uYhaybAa6
LIlW4agIJxFpje2h6jXfQEVya2dtmPz7yrroqLmHYgtsm3YtgOhRsu+TYFTRUlei
zxCw5fdn8BiCM6BkDwh9N4hujYT1AzAu195s9qxoEMyWmF3/97LAHG5vkaOUCDJ+
0d+k6Re5hVmz/uE3jc/w7zE93P6LG/gcA4GVjmd/wPEDAABY3UwhWS7f5qJu0e1T
sra8BtCahXz6/r8drXzJKPWa9QcBA3YujM6Mt49hwtzAc+zNtDB54UnolEPAf1KE
epY1jzfXvJs5l98UIzJV7RVQ1jujRpqBKYgRog4vN8E+Djg+3yaFmmG57nsALT97
QO3KlXRmq8dc4+ztOP6J3S/X5/B+l5bilDCQiwIvHATnDxPSKXqPV6wN6ZPbqiwJ
cXEiI6ZRqb7QMOu9NGjluzNlgTYr5/RrHsOn63jpKRqb+K6P8usv0E+UBcAm0Oyz
S5MIAZ4pjX/aXyr5VCya6deeraC2+vMvDaOz4WnohDPLV6pRqMOoC7Aano5A4Ijs
WCTzStudSvnt3rptXujgkRtsFnTjoQ13HlMhaNEuiIeo4SsRgNQmOEKEjvwT/GZo
iMONANugmnUB8l5eXavtC0Dx5f4/VQwqVfrUeQ3aMoigl+1PT57kwSwl9AvpnPVI
0UUxTExRKjNYcnGpTeFVsitM5ZBl1lp8oHi5e+RlUwKF6PfjScZUblvhsWxkJ9E0
rubK6ECJoVtHNkxGiD5Hnvwz3EfWxAGl+TldYITOfzUBmtZLIBolW5V4C1AfNEYS
2NltoSe01D4MOc7+Vj1JlhraVDG1I4Q/64XsBPAM459606upRArSN300IGWzBx3D
LjV9g826MvnDM5f8u7VDBOJtqXrGk06Zs+fgMjw70txmcN07QL8H2+Sg0p3vr/T9
HhRRL5FjsFIDyUYUjru+4qr//bGgFA0oyJ+Af/J4PSNSt5UblwKYDWp36NiSE26s
MuEUoMWlPs7B2TEg6XxHfHQowIah18HYzc8MjQY57Zjc8QHq+E5qAGNKhQc4L96q
gZuGYud1j84SMcdnOdaK32HK+ELYeALIYLPjjftcKFyV4s3FImEVzxlKlJ268XoO
xnCO3XR1oEa5t1DyuKxDjxCsYNIg14QBu5U3UstIYdVAx+qbmOxw0nMiVdmPcb8e
Jro+ZnSoKdeGY2g+tEj8JUnyzI9l+14+6nNhxUxFj1qIF2wvBTya7W4Ua8RSX7MO
dWiSvvjFuuuNu9ksyMyv+M46KC9t+YZC5B0MTSoVmmKh5yffvcPmIsbXiUwO+f76
4R1TsCpCVK7etzN6+XdE4ezK7LGKrLPbB3ioueR1/fHTnYhEBUM9ZvwiRQAN2OlM
rhIH38FZ93bkfTFhMMP+L0C49UFt6qiU2byKwSgycele5Or5yFA8DUuVTe34zvYt
WwrMo2P8OlrUSQvcZS6DUGO5F+uxABIUZE+CiffKMd3ehDWlRjz62AivabIWuU/A
9IpQEFIrX/ZjIIpK5e6j01rgtx6+qUyRJd0B/C0b/8661bHqELmSpYuM4DaVaV6X
+gt9jLS/higgeKXjEnqKP/zpV6jRg978HkJHAJBU1SIBv7BmJKA2jKlUi21hdsF5
zLcKqCJeUx2biOAPCoI2kkCuZveKm0ZW1uTuZ5sTtFB8ZnOw8gLDXxPypDNsDxMI
VNirE104la3AOEfeT0aIfSRa8pJj0pb/qLpY02FspG2xMhSYmgtnqUZzEh88YlIY
Z9YblTQSDxQ3NqJd3aW315XynkpmXjRWBM655qW8cmM7D40IDb+kP4aowE36C5B9
wsCbXumn16gQ0Mp1wEzZ+jPcTSIPQGCr5hsdncXfTNRk8GRAliIp7jXHrYkWEZRI
Uqa2JP5nJa9K7f7DUb7gWDiqUyJjAa+aULkmPJ0YYbGCAJLuJdcPkrHnn6dgC2BB
eymJpeKxD0EFZKkUo/0j1Ih4zKeexZW6pRAqXr0eTM2pVgLYMOul8kZvbxhwvD6V
lQ471LSZUkBiQVIjQQZRhBgrtUcGwiiioyPyaOd6nw7X/uNSarLGOjoNZwEmNb4r
Ow5fAb2mDOLeY62AG0sQzLULOe/S0l9MIqfOEMP02XEM8Xp/DK2vdUMZGetOdWCL
e5GVB+F0abDg4cutZS2QJ0+IvgvUWFVdAdFYuHzQyxKk89AyXpSkic+CIBLik0gf
ubizdC1LNH/lttCzr6LobKCMe8W0h+1xpSKyF5wMHDWEpaiW0avxIN8Eg8Zz07a2
It0eXdX/J2hRJcO6pmJpw11tjTCrCgoq9XG9H+w/s8oYEO6R8OAG0HOfoV1obE49
P9nN3iAZm4BBPeOIxVWSENNBhkxI5eGXCZqoTdfx2zPbLvLt26fvcE9H+r/Y0QVl
RfjfaTmFUv+0MddSidgXi4CMYS1hO2KeBC04wxMJlN7ZzALsn0Bl/wCjSP2LSrbg
KIIz6L6Z+kj77wOQcIlt4tO9UdwzY3NaNeeXvsb1owrCYlHYUJ1AXiU4BsaOySgx
Uz875XKteib/fYKjOG0yTzWpF452eQqagsI6FhEtjWE+FzuhoUdQFdqT7LGfb4L6
Htwi/eTMgfYfohqRFpMEqF17vr62fWsleEYmTKzi0PnuFxUsqRy0FHoFeyIu4ZLI
3f0x+pQURyqMHA/UJbjrlPaToVMya1v8TGcAdmggUkJLdIIv7vBwjWW36XZpVUu9
cLe5O9J38XUAnfXRsgJloAE4YWCXLak/84bgQKfI8b9oQrMrKG4jRJ3uGlWXrct8
D0nvxx+iAyiRSdBG1dLuRy68NRMAVhDX/BMm7zr5A9LgzCmTXuf7c6xP2bFoCSRh
HHLb3nksSTrmuprPk6a6Dnr5zVizJEpstC+mgAomCO6PcERWSgrCAIHQ5GsnFdO2
xQjP+5NbJjOBMqPEnIx0ebdLbWG3xV6g9t2UgGZlkkQ+xWnhghs0Cl57c/zQiVsR
WZnYCLiZvJW+z3t9R9RffDTBSBx4T/GYIpNIgdLxSAskX06nQKw7yIrWB0htU+F2
mUw2vS4zGMjc0/RGnV//3UnDgKN6QO+F8WDxtWOa7T59LpTtrp3Assfm5FTyV/xI
1IadUDj/AmekQGqn3EO3bk1QT9R52r86vYewNEFWyzL3oRI7DJqS1OQ7jWAevEv0
Cb7+fNOt63ahOLHobipOt3z+BDPwreOsGTFx66w2v449bdGlY60j2tQQLlwZTSYd
y8cA2lSgkZG/btslpvSfXhdbg/x7ZODMKjbJHDxW6hhqkIAxLeLy0oc9voYOzC1R
wGfh+yy+purx6v0ZEolk5Z/K7d65z5WckurPxLQ9PTbx5ZtixR71ZFHnp95tAe35
Qid5MwRoDbJIHaWCQBu2/2flOJXIyukejRwYMMu3Ff8vLBZBExAuUaUw5bo0heGU
fp57Ms/kW5wd8OAU9C8t5RbjIW8Tea81KttvFHO382MFm9PKqL1b0ExKuHt2mMlJ
iP6q5LtKM01iZCnOFvuox4WdLj79kvwgSSUjETnh0t/NdejRC23406I3ovtP2vQx
awXxmacDdLgXjgE96BSQG4tZiLMeABj/azfSIaio3UBtLlYtC6t5drCavnxNa4q8
1iPj6cpENxc/cMKaedyOB9MFnOAL1QF8NpWk3HU1vhOtfXC+NrXkgSto3n8swkku
//lnvW2zYtTdaNGe7Sxl2rvWY8SKCyJ2XVh9GixRoH3ZGmntH/n0ExnDiynies+H
STFVTEuy4wiZGAhQ9i6quIpOokM9tFlZF57CXhLxgDPU++FXcbk9HNtsg6mdHVba
7sxXQ8zuZ129zAFgNhjBUrB1+5s/pHnQZZ0pXskusShTkvGe23ZW+RRQu5YGxRmd
y1UQ8de0WBLfBr1WdEsyLOJam4HhSH2G1+gUWCa+/NeU9/OBbmIXLRnC9KO0+fVv
Oo/f6ZmiTw3BDzk5vHA8jlA32AwHCO2RjONk7u+yS7AHyYlzv8OYsjSQl0L5f0Ms
+FxDuBAtZcL5Sj9Q83z/0uRT18WrnRdF/4Q9YtQ4e9HgWmMHUZRzosXHyydEPPL4
pPCmuzMvXMt37LeS9U0mDkvt1xkXqie5o1ANuuWAow0QxOrupMSJJLTJSo6CpBKj
ovGgsWp2jRrl41n5ZB1Y+RgOR3bYy7Ep7EjMhhBvTbOGxOBCzMP2TSwUa7pP9UEF
pUxIFCnrsTtNorXSt4iMoohDqphRNLw0JXVmOTQDiMFbj+OXOKJksuQgnwNRw5OL
R0fe9wp1YP2FMrdq+a/o5LpQT5xd1seJcUMAWf5kN6Q2RJ1UuAswimmpXyOuO8l3
y8pqktH0j/xh7hYLEWjUX2BZ397VzaAR1vgpaOPujSyu3HgsTlMIrraP+tgDz+oc
k8Ln+6RWbnuiFAJrgH5Re6TknpdNaiLe0gj6EuFttjY8kQ+a/U22C72OySkfvNke
2hKD5SbLWt/pdWIlNVpwGYo46udCr2R5vKKZx6byuqNxoUkwQW6YO/eBfFUqGHxC
TiuuitQBhWWEfAoPrY8NwKXx127gc9oCQlI7ss+XyAqXTfGKQKlNo53HPGV7bOgu
rrFiP8qfiDeLtbapsNdX0uUprR71k318d7l96eaivedgPTzDVwSjEpXcckiJt4Z4
phF6HFKhoszR7fYNaYmpISO/9p4Kp7GTnvxbx+ZpFRvTt2/sruo4eiuzsyfDXvw0
Kfr1jb5ufPWidI4X4+MBbCjZZLNrwX9NDoj4djdG1DZVsKLWhwWCgbuA5pHRrhMa
KMBxzdEYra/dY+Ej7FlOrOCDZ0RK3xYkq3WW7gT6dNUkrPDi67f5C89XA+X2B/sw
gAzqMupZpU1YWrJXzA2p53wZC7ZxI8pwGTAyfA2IJVT/nCHeMbHoaaE6bMh5gpep
cuTtg08tH3YHHuXQIP/jSn5qTAR28MxskahEABK3OhzmMaAH1MWUm7rmVK25GRXv
Tc6F68gp0pxlcVSLrtRwItjPmPBzbgUjT/3ixodeNgnbbitnqLOkaN45R5MPYcrX
y2U44KTgbRaASF9F9H+mZXsbTepSM8te886ljaGFSt6ZMQvw9eUd2Aed6lz304yr
JdcjuC2yw56kdJVSbjUOItXHZKEUbDPeJFtrXIOf6PII9NBHiztpdrmRk2DFYhee
8g7AXwQRQJs+PueMAEgNU9BvroaAcEbFgSvAp/rK61PQXuc+5dJbpk2e9mubExd0
N/xamY66Zo4kH5+J6XrUlI2HiQZjx97G0+4br8R0Hw0Q/LxT0l7JhnGFk7uNCfin
edUScK6cgh0KLOd1LnOSgV9FweNvHBGpl36DchR58cvRcaBUc6tZCuE89NzNL9P3
9Q/GnQ7/B23ItTZCO/8EdXGpKRIirO6DfYcpMPFyIPCUsokiqOA8J5/gUIvy8cFQ
Hi2KkHFj158KbeOFHYkOLD6DdRsu8imvuVViMSMrH1dYrFAwFupzrYYXyL8adlkl
lmhGYWjIxFd4F0zJktHhl4FugsmTMFF/sNabfjNtk8Fjxtg+6j3CqPTY3IITfJ1J
Tic+6U5/O6+k7QZV7Wcr5c0BtloULdhH4EXm7YyZJLzf80CLs7oEwAVjdbsXNqbp
htc/RdFqUsBotccGvy1whWdKld44yOsWYZSXIHr3DNu3B0v+ZzOc94jxBjz+PgZD
J7Ql4S3VOrx7mNFx5Iwyz9RPDGFW0s0TA38mHeR3arVge0j9vbVFfPG3hu0iNRvj
thyfd1/L+fG1NkJVKgbL1Yt4PZQ5EHuI8nfH4jZ277q9PfomEWszERHixV01ZqXP
O9NAYLa8sPsNcEDvMSsd3qC9gemRMbG4URExD9mh39ev0lmjOirtjTmhB+fI1bDV
JHfNiQPFDbeU0u+2kEYkMP8wf8fDfhe1jylz+SjPZpmE7h+jnhtGkfG2g6eCY/0s
rrW7b7pW1L7su9e8+ia/ekifGI5FhM0toWrP558HTUYDdzr0OuUXQ+xbNcKuV6xr
8hoOBc7uPGRXEle/bBYDGMSJBBsi/uxD/daSzD9reFowvUQhlOT/RjaADtg1cmEl
Sp+o3Gr63seNioaflGDajHcNJMZsTU+PQixvwxu9c4Q36s/gHoTQlgdye83YJiza
wrSuc7F+X1WO6HKYT40pVz3WXced7Hu24qk7ItPznRpnDsKjoCRGG8iugsmrX0bf
R91XuxWfeto0jz9ZbeSeybQV05mQemBNqmv2g0gGYIiEhs9uxwyVfp3bUbyy/xPU
RrDH+GO0dHVwSTXUk/yC7x+cbreCS3oHrjcJU06UVWfsD7FBG6aVWY17DWQAWMdI
rx2PcJ+pxDEIajeYzZrJJogEd+1LkvOlRFSC1QDvmH7UvcTp0dQejTItZrBSPM1/
Pe6T9Q+S/LUq1pHM9RgWeLtnu8leJc/iBQoIFOPFUqu+BqHyNUGrJaOCek4vi89E
I63mfJG3PjNsDOMKp3sc2qmZsmP1Jalf6Ke10DAJn9/I9sz/yAmyN8vdM/b+i+63
rSoELj2JMSCw1G7JLtMU7kDSSexw1hW10MP0RQdfjfGrN4DMz80gi0rntQP+y7aU
xRaI96KHjRuFX+myy1ymw6/ouTlpmwpx7zlPM//3b9EoHCovrcBQH6HR2ITl9OrJ
e7vE6TzRKiAkRsgoI7+EwxlfxsU/sZZ7WCDTzIi1MLfV0udxxV97Fur6j92Yx0hD
ov/KzTY4ZmX7+UNA97u4RdBsNWI8+wCEBMDVfUA2XnS+1FpUPLVY5rhDV3CzJpcO
HbCSpS02ktLDGEfuQYgn6Y1c93+f0h5+Gl4t3eu67dWto5ozJF1UR/Ma64h0Nbtt
97ylGICDxoLgy7504ZFw7h0Gv013qtQzkjuPFnwIciCk0ssxGy+FQE6HnllYVZsA
iE6u7tkb/FkZYjSFIiEvi6SCl8Pkg2AUuYRc+vx809jLLNZpO4tpL4Cr4ouVtS3W
IPViv6yRy0BtItkC4XxTh6zUvKP5o3aCPbPoP4KcSfpp1KK0BEcU2t2Vs0ujyLcS
edcEZdFn6lAy/gpiGJ0UMnzP3+GSYu5N914GPQzfAzXHAdDXrhFnv538Vq+tDAzQ
c+rDbiBQhQsaEqT33H2K7xOjh+/0BL0alWVXr1ELLwn0GU9fPF+Z+aVYX6j8HqW5
gH0veezg3pxbdrx6UNJsJg4J/IAuR9BdAUThNWqCSeBAWf/oWJNDkMffz+3wd25c
65WCZo0r01CbMtUd/VYJLI0f/cumvLMoDcAEhHUxF8VBvBDvkdPAnhRewm3gvK1Y
ygjk+yQamNKkyJaoyHAoqrlgb/7msV1SNo4N0Ei3PcUfpokCDmw65Fan3oXkYfmh
QxmkiaNAQkhASVCsvrrwZ694479BuszO+DV40HHds+1fY2bq5Zwtq5SbJknWANUn
FlQwpSRKEbIL29oKVYaWmzN6J/EIpdn26+1cO5WbWA2ID926NA8CTlMBJUY6aoV/
ie8lGOYauIZw+7JD/jlz/rNCrt4f6ZIIN58X9qJxjDRSrdG419pWK2b4TOEEt5vc
sKsIuENnjCSm6cm6tvij8FVhveUqadifFAJgkuk5VD4ampxLH0AcVS8XCpTXfyHq
2UV2+KxsgpPyc9Syx3LYUW5vaLYpr1V4LiA788Q1rmxV2fTaA3nu1krdXf0NBMQq
UXKSF0jZQ+GkrLiynxvgMbc8SNJULshuV0y4WDq+BFLR11ilj7Z4ehuIiqoTjjD4
yvwrHOxK6LfWgHQ8hXmiopKQoKUVX0U+UwvTk0pr+6gijrN8/qdS+455Kqns067F
esuclA0yKA3ArwMZnXqkkd+vTqRIQS91GObXchz+1eOf6AeOULJRL4q7CekPAd9y
agYqFziI+zd/xp2ih5W4UWAS84BbKv3v52nxfaRA7LzTQZkpcRKC40pwkJqLtGTF
nMxtoscZGfFCkW7e/3rP6sCghejZq48RD/W1zcIFpyKMFMfdtBTTdU82OHeIaqQA
YMc6zSa18yJAQHKl8aLNnHBquF2Z7qbFZamGHrmE9ePoc9Db3z+qXCEPtcm9v6X3
EU8ADI2jdVTxKTu4CDt5nvXPbBOGu6ZSczi/PBU2L0g6QOiA3gI3XiD+vUIxZ8iW
wQgPYpbFMmAsNeK5wQ2PPsnun9A+/WKkUx1W/YLd1ci8vqbotB5N76xC7/iBkZGl
+QR+Gq7FM/k8XsaLlwgmAwPV0GtQOmiLqeTjcZ2+b98HAsDtJ4ID2DBYsjnlXfng
RhZmcsQxOBkVJWU1OZZXUhHuAYO5+ZBBPZAigGS7lb+EbyzypQjDd5UfzNwEHNj0
IzXy9d0iMlC3nXBwA6qPZbaXQPWbrfzfXfihTDEwERG+iR68ZLWYBxMxq9RB/9NJ
LTuNxpIHv6F0if0QnLYyOsAAz3BV1DrJNNi7zPLscaSchdSgq8OE8zeEJydTRgK9
thse4LGqlN/5MaFkqQHI2AxgsZfIruoSQIlAvgX8ZhKXqLs0BejLyDmb0OgPzzTt
lfgdFOY6Zr0PHsarWpPdpOFz9K9gbqgUBeLH8EdWtCpI4T4+NicW/mpgoGTChGd5
fP4VO1vZMtsT7+Lq/0xZ/5WtMAOahBswRJBOd5YBS4v299aHN+p7UJqu0vTopFSV
fwOhTUHu1mvL2rbu0tA6h5B8YJ/ESNOHD0Ji4yAfs8MdywKep0AKrxxFcLXg9oGF
4mkGyx5GnJiwW8T8io6TJgdZd4OL5JyzeFTiESFebQn+EizNou8yfMLoGNdLulrD
N1NXxA6JJJIinOsPni3LL6ZHDUPQjYNl5nyYFSLqeKxpclKQ21M2rESq8vk0gUBQ
rCXbxxdFqFzk+JeEy5ofv2FCdbhaDnKjzvcgV29s6PtgGULWuVuBvqK3SrTGxUBi
IgYteitzGTFtWKQxscnhuJAZyqQKsiTUHlpj6YqyRiaw5NlgzM+5crvhNjtnYqwE
kQ6DB83BmPfgsrQ2OslyCuBDDtIlQKrYOAk/9oe2anfMvrc+8TJtBJ0kZ8JR6j6W
H3j033kpgSm/yCupESqWL+GBFX4NNO6ktuRiavR1/aw3Zu7pzQis0/KMWFRRVwMj
onMsfV7aojeZkwxmI4KWw04hLMqSa4PKXrmVDk77GfgsZYXWr60qtnQrm97K21g/
r+9TnbXKVvykG3tySAeQ70eU6cDHAGX09ZgwTcFU0panMQF89yYy7kAZnvtAqUbd
eWw9TfhTnooTRCPNRSBz53GFHStGi0e+NoYDFVjXa0gnFVs/CuwzBFaclvFUw5sk
DOwAUC8OqRkAj8ZD1dymKVwBTTKu7VOOd7i0UZCMhYynMr5+fI9qL2sWmKk39CcY
pnwLLA+YefjUW59bx5CBHoLEUhc6D4h9ReLvY1h8XPkx9xhfbFDBqsCWwEZxbEve
jx/u4kTWCiddi6sloYS+xtjuzfv1iw05Lq+CqwPpVXCiGpkKCwAIGs/aU66jwWpN
t5TVKixcYRy53XQVwvwbjCRdtSmnSKjvHIRJ4u+oWfXbn2s362EY7wPU0CkXUffh
DlKPeaT1oA+glIGegSS7cj2c0gh0OHCd7TtX46ww2Oee7Q5VrIDhUp4G2tD2je97
Ioi1c7FjTTTw19Me25s45fik5LiULlTokl2Tzvb4lCio2eyzQWOGNw8wk41yihnd
WQ8fWeRKSw+il2Cl/uon7DJzbD1LhqUMwIQePs9GfzKLHZ+jC6oi/eARK4xzQenk
NKHkKtiaAvETF1d5bTVH2gqLZXrDiWZf6SXQOFEWutTS5dD48xYx6Wt53tDZMTI7
JlSXtRbdfctjn+Pt/Xgle/vVa/MKwdeMprzBbUy+1epSuwPp8nOmTU74utHVNfWS
u3jQ/rLk1kq5KN8w7pGQ1qovq6U32eoO86sSk47RRPTjdU+eVe2efQCFZ0scd/8u
eS6jMtyzPrrY7P8nJ7FLFg9/szr44p/C1RCvuUW23mEjId9LJg8TywXMw2BpI+JG
lLoPshtuholny7qtSX35BhS9lccDYwEHPZGJviT10M5uzRbGk7VR/C93aBOamrMa
viX9qMXf9qzVXFdBuChnoBTxVqYmcPV6gDUeZLpTN5sT4JMMTbSL7RQBYUYegOHI
ZmaX2tcr7tTIqrSZGLyUThr8xHlA1cGiYBXsaMimaGQ/YV7YwQ2h7VguowQmKP2p
Jvtj3CIg7rLpinSpGpJcmHksrdIIspk6JCBYshhTqnjP5yQu+wZPqEQvXn5/m3z+
H3elzK4yCRdr5CHMVg8q+SCVvPoOHAb8lQLKXjF+5OyTRQ17oJWOaMksuX7sQij3
hPQkcjIZnX8bGhBeAeGBBDtm2RMo+U4uUMA/9jeHzER1GXBpbCcsGWOrzXguvFbl
l2o63DpcFijYRpqRMrOuZKpAB6w6ZP2wyOx+pQ8QYtxpORSxD7PPJsHA1uWoHb4X
oL/6XkJGUGB4QsaPYr4pIsCk5M0RrXqHwxlJK0f+Pvw92uM+1ZJnkQzHGMRC766j
a58to5+TRqdMqBlTFx8HDmnra3su98uMx8zo4W+7RvM9xlRjcZTL2MrA/+tf0DVG
J2InVIC+8Gl68g2me5/F4gqQwPgr6zIJE2KEoHIAcMq+teks96J/uIJMtrnv2+H5
Nb1GqX2qQgtPJT4LGM8gYcgMRjoOlgkqJZqoGK9M9yQvSeIDysb85FB++quoVuF/
Xl1RTjGQN89od8sMZ9F1LhR5NuVJZ28hJR2QJfFlFkV+QAPLzr+SQofLuuoEfzUS
f8ed/hLGIqU66u+FjS8WbN6YPPHIyHSrOweKHa7L1TUM3zHhDm1SvXNot6uQv+go
XtDeWkhZ0OuqcGZxVNgSIc8spchaUTjds+4Rdhvl5WiUu/RiTttBEi6EokUIG7/v
e6+Ju+3uGczu4MhUyLlULRdESBaTA9VEtWdkSeZUTRKzQTfoAQ4PUrj3faCnf5Hh
wYYFGaj7sbfh9TRrQhTg7gWo2SVkxsxx7dMdTumqt+7ZBLIEHKF2Wbg1Xshp8PVb
1XmLodnlTqTEfhOlPOtbuBtfTJPqergPy5Q7ZA/pzRpwVP9YLBU4Qz+eil7gVj6V
uKHRm3Sbl6l//LYzosI57bKheBIlTKwW6q28/jqYj+aeLUJbnPU5LoahuyrwMzRe
Uw6LNcNx4wj389f2MF2ErRdmYvRWI+pGg09F4xn6kXgVQOaJrGHwTlTiyrf0K05e
oxolMMhM3TWUZQEqiY8dhHqJwmPosWObqcYYjRMYWWWeaV8cJ70ppLqV4/ZyOAo7
9cuAI7SjeLrplNKKUUOIDhYsKP5XVJSstOxCh9QcxKg0oO+9evybRklEW10ipeqo
nx+u/G/gbM75JrRkc1g+j5aZoiaBSZm2eo5DKlCqNWXlphSHr3CrwlF/nj9hiTMo
fdx2EVu0LZEnxgqaXmrcFGWxDPnSsXLC+DssBenrboVFdY5SI4gBVWzGyuP5fems
NzpDAnHtiVGRf3Oau7fnWobm3P1Kbk9u2aCVC06hE+VFTBuy2CE56MZFUDSXsT69
OSA7ke3+4bpeeTc+pBKE7PRtzqUjOmixtJzpxyyS/whZcHWDsqBW2DrppV8RabqX
UnzZjCbZbzTLMiMsahrBbp42ebQHd9FUFAZSxLXDLIhrPdGoq5diUqtuYaTRK0CY
CrPMx3L5QweiP13rCWnYdj6nKFKtr/PGMtEX6SACBurQs/mLbixcy9pTi5Ia1Jn4
mx/t5BjHdOYxNHVGVZ71HkWcTkbs4dhUwiMK7iai2QP9xF1Yq1OBqEeGGVXU19Iv
xMk/eCORHEvo+9II+62gu+Krb01WPau8V1jI+HuHL6rVeCFMY+PqABHzmfosq8fb
W22UvjIWtCR9xylDLqDMSqhbGsUT9UgNQiiGIECt0By/0pPCCMJflcQox76MAcPY
i9QgmqWiVnDr9lrlJkYAs33nVhU3nlPD8SHYDE2edMrIk0Frx1jNtwSXWbYmGT5K
p+2ojPN8MG51NfP7TzvJmWqLXc0mKjnT1CZVHMinw8wga8KR7aqU3W+V5TG9p+eF
r5oNXPFvSOHawqLDbIBupiltfD/LMGbJCiZRAr0u50MVvsAmxLWYuNTPup7ot+zF
iwxbM89RP5qTAWh0JgpoqkrGBe6Wd4rPIG2gwwNDd2BRFDllWCbj2PWGToI0+81o
U8P1EyQmk0q5szD4qDh697FVyTKcSjWfDD4YtKYk+/asC0QittCV86B8wechLE3s
56ET+GmrhHlZht/An6ZSV+2q0OTZZp+SujIgwXCaUr5FZnDiC5HtL9fXhH24fwQL
lgftZ82Up6VYV2becr+OODYXyMlZJFShCisJ5hLBv7ODRCf31uPNppQL8foShxfU
1gB5OzRHop4zESE3ZrrGokTA4T/SNTWID9him8y/vIvUucP9sMY6vpwKjTFg13a+
tG7UaQAZgrbYcJ/sUDTSAl9sXdO9C/gYJhxQQ4VYMs7hiFK3DheFGPkgR344GV3L
abH9vSzDlw0E3HCEHJvStccmm2h9JZmW3IBxyo3kZYiWp2rXRnRlrDeIcClcUmOB
eJ1bIQ5BwIwpeB9W6AaPER9Kn6Gwfz4pGEycaotzde5MqY44TX7EWaxUM5rUR0bF
1doosEkSPq0L+UqMLXBWFhTZq66kZEVxEMRz+feovMZ8KgzIrnaO9r2n1orJH2PU
jxsaJIUe1hm3bEKLi2g0uTwFTwxXLRDhLEJ+eM3H2C+ehYG1sd/bfV+zUm8K2ybv
YfaZVa8nt+Md4GK9jTytm4kDrW2+OwgecgtN1qVtP6wjdWkgMDIygAO5XAcj/j2k
MnZmV50fYkS1Mm+HETHCrNYKH9b2F/Q79p5/eNxu74TaEDasUAM1xtPQ2NutSI5T
nNn+iHdcVOYGFW66g3pJFYpRbGmJhWKSS3ZkMd/X9QARE9LfJtdFHr1rkIa2K0sn
43FzIKtVqNZLIH6xsFwn3Ip7vvqofPWGicIHcqrklEAeO686P6mkYVEJB4orG9y6
MXYJLmEdyqP4tFp4iHrwMl4wpSAB6lKmimJj8ElYSHmEQU7iGD/6+Ki89P1SMD+X
nJTstyzpKQeioQUoyo7txmLCh0Qohll8eob0ck8SxEQPznZMw3/Fi2mafK8apNH7
T/VylL6UrtZQUYhIk1hfjuLrojup7CPlrNiUAwnnggSuGitwcps/EKpR4OpeDttm
a93Tu3HfBs4BOhqiPN8LYd/Xv1zqTHC7kMvX0GwgZ/o6RFQU9UB/8xjKQ+vGK+p4
c7DwxoZVtpNuTVBVJ0TDajs3C2i650Jo4cGtEgLdw/9teT7QLxvEuGfRDnSPr3aJ
1lfZnQMYwbXjTQ7J/VCoqsAUDijJLDqvENo+bhY0pxuPna6c4AEx/S9ci0mST+Ix
i5wYH+jlQKKJlnjo9vDyIkeaygiBD2ds395Ci38pI6N2teGzpASXeSCaD9740rvr
CCRYyIny145gjVTHr00sy5mlPA4xvGtEBGYMrVta0Vq/3FU7GzyYmHGjLsBD5pBD
IEKK9VpKF5ElkRthkdRgVlXe0s76d0uwKGesG8X1Q6yEmCxQY5HcOFKIR0p1Brsj
nwUP8DGE/9O4OyDi0hiiW9ZeEx4kEtmYbQa5JlrQYw2dH+kXCj6K/5pTcvbkaQFv
8eaYFgDGoxWUQaRsWGcc4zbrIz2UTfvidkrDftwCzdgvQjRjL4KZANK0Woiv/B93
q9fnkPcoAauRQWGPir2UrZlwOmxeny6jJdgn2D90zLJ9ZwdIYfDfM9mJ3iagL8Mg
IrSe7iu/Uy9BLJoIKmI5LRerE4isl28hw+3QVYISnI8rmh5r5X3wX+6ACe3280oo
kXtBVHsA6vPH00aT99UDTWwZ4CbYAwHUKlxX2qKbrEQ52/sG2eqnjCYl7f5pUBvS
z5+uDlwxkiRhR1/bfN1bWCuASrVHZezwF90o2Dr3cwT6Z0Y0DcIUQ1V0g/X6E2vE
aW8n6aDzmN+eN4SVCI/0O2DjBptwhKFxz/ZYTRhJ2+rG7t2OpNlyy7y/+/qSv7Ub
YnWim5Ov686+AnDGSdEgUIUN8EXoKwA7sbYggRMqEynwYP/2SjBBpsyCKRudsDzv
1qLoaj7/2tislZq+Gza+ikKpu4YdWeM5SkPHQxycRmYbU3Vtl27S6dL9nwzUNkGk
+UA5kV/R92AFuzJiVOY8ZNy96bhbiXZA19p13ax68UTnRICq3v6UtvIaa5zp2ooC
/lGAOeV9/wwEnpgqfqIPeS1eSKWrvEo2YlCBusmbjBQxpv4lO7M+LTvxj/R0rJOg
n0vIj0YUIeZ4ELDCPUsuAK1Ykzcxs9rzEN/+duMYzoqvSAN41rWQNCUFlGEfASp6
aiYN2gq2k9AS7XpfSn8jPJvdjLysikaEacmV+uw3NucoG7OpkusEtBaKc920GR7P
PtmrpeQZNQt5xV65UIRPWj3m95oIjo1EIKD4aGTn5VbVT+dxuHiRO84V7cuQps9H
JmtkLDAQYmYLQNSg4fY0JedgUVS9LDEoeD41vqc8j3ym1X7tpc3lkvRpe2p0unfa
saVVbfeukUNLDoEJwGfhDzbLHzgfjzwgHEDqlt4/TbQcXJZkkGudHJJ19OUFtqcv
7T8iF6KPvJjc6FPMyOQQp7z0DhUQF9xGzZeuVFOA+dKk6SubGMlFlUyb8JBlwvRP
I0QKiMZfv2QffLcPrJhLuZV1aYw09a3A8DCKl03LUKIVW5usEyeoQA+ZFlutkUo1
THtvZu9nKP03doio7E41LweAykVJTFIJpvXSBzCVsEf5/94k3ARHihZlqQc5Jagt
4ZGuvtGpBuSK8WHE2RO+ChCDnfRw0u+wPMmiiECSCFVbOL7A7LAxpp1QJvYgKOsS
dDn8QQetmGM4PoVMpapbPWmh3196krHskGzcXMgDyMOMozmaCWPmi7B9lldpb8Hx
cPjMK5UDXz06C796GYgtWm6R3xFipZtQcbRTjXr4r/9u7P3QFk0rJG0iKos4j1ND
MgpC3TZMWGoH0hDbizmZRFG1BUrGkJ+bwDzZQ8DiMx6AWMIkip9Sc88i/mXyJcKI
V+yzoAertI2lOutz7wmwuVUrDlOF5V2lzP4ts0kaGq3+RAfCiT1v4kCJlE1v8dTp
e5Dz29n9jbILyCLBh6pMB0fODjrGUAy5utExCsNUTkQYOtFG0knLagYuRyR0rAMF
rmRVvNJHAEbdv1UuZYBmzFC0D0b6K1IxaVCA1SDVC951BSi/Xb2CDM7yQwQ3mp5W
3i85ni9Z83p8dg66Yacd9a9ldvbed8LhCQeCnElX1OSyOF2pwVjlUEgzGRMZPFp8
sRM4rOOv8Nd70XDxQG83inWHNrd2zf7nMYZLHOD5MdWKOvrt1HYYrKmpJimL8clj
bP9UF1dp15tdoobMDXLIHOmXxq6XNz1It84zK/r24LYqBddIT4GDiGtOzTPkqO+j
JIx21Suo1WfuQpVxU/e0df6EGUj0k72c66SqAd1XsXz0KPENJFW3JAT2Hw6jVix0
+FRc0UH/9N2JmxoQG/E02mLvxjObl6oGCbO/v6YjXsReyetzfjU5trHKZ9IbgnIR
O7copDofMCxIk+w+RaSjpSV8b3dRqBOHLdTwV5eODgi/LELcPrjEeBGmpYp7mkYn
F4rIB3Xwbo+NYwdT9hqWJ4RyDalAsU+RxlQFIYU7EdZtf/SAsW+MDE8+tSw8pJsT
d9IMqnLHeoE6TNXJ998ia9By0gL45LfBe3i5YCnVCgEIT875A/UWw+RGFyHOtdhu
+TaROBTUY1bxCKZnuGI0HoTlcAUqTltFp4PDdD/aZR6MPxwoWWcp1cHIqceQwlUR
9jfzb06tGPhuHgJEq15LwDFBUuUopzt65hnCASWgTTPea3NWrFCzs3SAC6ahgXUF
bfWKKeAAHMFcWGV2qy2ad3BndowRiXOwqGhLWl154iSsk7EML64T+VC1DRFECGLF
UnNfd8NXZxu2/hY5AGm05LI9/rIvDfG9jJKGYpZCIiytqJ43kWxhPKgwGzqqbyQ0
TlP4lhc4RzxvrwXRNZd81PoWrSSi7PdxrrXf+UvmOZnKPR8Q8wRe0RPj3T5SqInj
pEkmTbNkriUrsJESRYTRsPFjTPgimejMrPvfctdEZNlttnIWkmMRiCi63pFobcPV
6qr1qUIS9IGNEOJv2LwK+3gYogZS9LqD20e3K4Mzy/nq8nFBcovt+c85eNEcU6ay
9WtFLkENThKhC9S+wCYl1teRJ4YnNSz2ydV/vhIqw5ez18VVc9GtEOlPNeOgnHX8
fD6pJZIL0dH2H0FpcY03gJuKu5AXrGjCJtv1wtG+u6DuJO4uiKqklcqkBf70aRUl
QL1WYAdU9d6TAh5dW/g5S1KIEcEromt/VtFX055aoAexWpmIuZUXRMzV/IhmdcBa
8v3rcJ1mEHC9bTHAhNeQJwptCcy+UtSjsXF3VYyIgcbbibwZPseCujrgwjNJDZQP
L67eObsvvR/QgtnRM/bMsFaOFvIDb7o98SVlCryL+J8De8RPWNAGnmpFDSkULmoJ
cEXM/164mDWVzI9D9t2t5KD+B4S33QJmLV2vykDXXQ11s3nqkrP+VnfdgAv8b4rJ
Ya/5ba1DWZU3/bcAE/80nIG83srwBZ/bUbRp1B0slusNM/wIwiYVBRjl2ks/fBUP
xVpZcCsJ6Pu+vMre3/ZAKrtmLrVHGL5LhMnTjfPjsO+YYsRrqWKAxZLzC0MjDqDO
/DlL7fLxCQjTZOnh7/Pb4ugBna2wlL5/6MYuZhNbOuE7ChIqpkP9+v1mKsuxGl55
Bw5H7c/HrcxQ/l+ZwlC4aJ5jyWBEA/B4xBjRbj4Z+nFRH42+eLhB8B4z3Ax7WxOs
2nUEENKX9PUMnPyXJdK7NIVorlj24hG/wIRqnX8hDCuDLTdF1JcfHCAQ3InyXAbA
WfubfaiZ6jYDUduh06iYsWS9DpvGVcRvK3tJ0NJ6P7r61anq/Tdj/8ovw3WKlmkb
a3F5iyMDxWJdnMsEMaNpWeNZVJzvB+KpdOhq5oNwXErQu6mEpoEpiYI3e9/rcgx3
zHGve+Bgv69/HwTLGD6HaNpIYKZ1+4i05UyEWD+LdoQpKv5CQUDbIMHOqfc+3zsF
tJmFc3jFJ5nCViF5q1Q2h5Y7CKFTH0nIvmmeCIhTRXLvI0fShXt3r7imSufhNpSr
v8AK3sgIk1hdu1GHPY1OZ8nZWFCZOnLQpwLfoKrvrOjqZ0HJeAThIaXoX+Rx2LAI
Zuuih2kkM/tLwO+qRBQi2h1Fjw7Dzb/j5kCjIHdRhfSCXlk2alr7W936vDEd5UuU
B5dV2BHsZcIh+pL7wjVVPtudJf7CL5rl3ElkRDtC456JWSepV6KzUh4vgB2AssW1
8hCsku6WpzwmJ35xguYWgasrI4IK0lSujkTIiOdsRSZnWylrKT+bd9/mIqIgt4fM
+rBKc23WAchPCAA8LuMyuViEWm53j22H7dewKfSNG3WhD3SyQmFdBbsPXR5yEPgH
DHp/WUm1tnFMVspj1VvqyQIkvLOvsCFXlD5DyWmN4dVLxRTiZ5w0lSOtMs/k/2pM
ctd6/0GLKQ6j9ya2mZ3BhjnJ4ZAX8S3drXqzuCBfeCfHddUG7BjNmWsOZLIZYKa+
gxGBmRsd9bIZuZM7MUwzyECNVKP0YF4U14N4b/6Pq5vsCs1OZmZN1iXLG2tKwbHp
Hqs3OrrH4JlOHIKMkwVozH34jptpONOo9XVx7XfC+hDYNIotVtoV7ijsfatVuhwd
X/8IwlyAlJFhrVKPLQHDnTDzQYTMCT1T6/b6c9XOolMUCPcaIJALeZHS22DfUKYq
3vNgKKMZOsGRLOyCZ1ldN32Wi1TcACjIsyEBs7sszZ6m4heYIfaK0Ro6NWwoWbeb
+Blux1Ylp5+ffWlhZBaHUG71dtMgdSKVKZjYagPerpQfzFpqVLpix07/knHzPnSe
9cdzZ0duxKPvOpHN7aKkTEGbRvzCTctx3DUjWFdJG8itj0IJHISqPLHAu/pUhK74
LTc3fQ5FXXiKWQ/EGgeqsABkbzpU85BXOtKPaPMGMWHSxm5s8oWm7+Y3L+ghaLEM
Onzre5URNsTSDRSNkru/2gUiFW3nL7X+3A6r0rj4xx7AMlAv8LAxcFfo7WO4QTQ8
KJcH0rz5IavvCwCDbgy0opnBraP8WxdYEb3HRdp1kGeYfRLMQheNFErp0xtD5wEz
U3hzJQ6gKpgNrUtNGfDAr5pQk28j18/uUyXuIfg6xC3A0SuRac2Qwh52SzVbIPhb
D392hhdw4B7EPr/dr1F41nZ4Bozh1kG+6WHZsuB7ORzM3frflOh+t6mxQqLK5zhN
oimNDofq6psMqASaCz0vSqPJ/wTETfgvpS+p1imSXlPhnQhuiY7SkvcgHTT67cyy
7tRrASL4KXisfLznlqeVS5TC0HE3nKEIJ8NBAASFVh1UZkcTQ5clj8wD7fGgBYjq
sfs72XXZeeoOlqDbeI5G3ypYLwG9FDxfPcPls+QmylSbuCht8B0Uqu0t1W50P/kf
bC6kFa2W1KwzdIR4KrR1n1NyntBWM+iDF7BEyrEspJq534DKPr0anUAF6Wa5G8Ml
gAMsdAiId+SimE0gtDSF+Qeq5wguYLaEdSX/Ojvda/DY7ja3QpP64elpWa/sBd+n
IkAiaD7VFs1JBVQFjGOnMVFxIZGEnzi49147N0iQOkj9cEDCoz7Ahmf1H+oiW+Lw
A/0gtcuV/favQLxZC4OqSTKHnp1FMRP351mXAmLB9JkuHAJg6Zn6cunNyccm2lcB
qD/nLsKQfF+66yPP9+2QzXP/gWjvASjeKDRXNcQ3ekqmN72ZEeDSaswnBBsM9vHP
EK80bX+L0gxGCqcNdVqy48+TqixGMUR82bKfnrRuEXgp3xnV1JvrucNroqF4z+rE
fQzj4jvJO4libPEzTsz1L0jo2+SBq1mhWoZQ0bY4dCmK/MnI/ElGsVv4U/ZzWRDS
jUJdKZme7hDavdb26g6Aj/Vjxp7LqxO9H7CKFrrV0ix9THBzu8Y5lrH2tjg3bvGI
GRVfsopPsupWEQrXOBg1FQGKKv0MVY3OhIw2bm+6sRL7WTVzNapFNZAqmqjS1j60
JXRgUmHmK3cSFNg7sCavx/liqSFGPwPtQ06uqfflZ6abhuvQ1qAmaRCz9/4yfIP6
lwPD9YsC/vXiDjx1kF5KhjFYS4FBd4g9VUd1Ry/A3fKj7HijvdU1c1ta2AtJO6dE
a6MjAWdHZtNjTwm0a/8apdGpgdwHS0w5YkCTvpgu1T7WrgNbIMHanGA7Ekb7AmyQ
Wuj84OS8ZpYN7DemyjtCrkjQ6qvMKGb1RC8oyU886sLcBPXI2FvlcXfqVrMmhEGa
qkTulUxKbVq2mCVVqeofTB8dB/EEEDxnUMJ0zBVk6jZJGyHRzR5WvKKCNRurDiEj
mbCq7tHqcv8TALFj0sIL2i0RbeWY5WL9f3xvytC/IgZwjiI1/sbMSuzGj8uA9B69
zkNdPel1ewqsVoZI8tfOZdQ9jWUevEoLsQAJemhTym2dxWMOpbe5rh76SO1qdsPV
sWWb2NpfT55q626+CJvjKT3UfZOg9Tcg2ym8tL5qZuk4fyimr4VCQiCsHajipC3m
b66GPjaKJjeFv5I+meEnzu5aX383a5pA76+5FmfoLFbPlrkIGekCX57lJ5Gwq4a3
3q2S//L4vOb0N2wq10o+5wLrNhbbhatuXF80JbAhizhipVphi+7zvCf9vk9919CO
YG454ITi2UAHEVqWnZGCT/vGTczj4zECzyXlk948JVZoXLzudrNlSzroWhdbU2J2
q0OfRsantIzUCDkZf/e+2k14jH4ptVfxopMms0WuQ2OJJoM8cn0N+6Zok80UOe5P
DEQWLT2TY/y3RC4dffHXH3BAoGl9SQYc1eF82yi/jPRQSuTI+/vjRGc87yiZlF4z
kYPwwSIepSp80WO/lYYXo6qbmghgNxXndaEHbdCjrr9J2twoxKvrei+09exGXZhh
Kz7kP1yqu5QpJYU6X3M787PPGq19L7sBq4CQwbllD7I7GSXF/EUgRrLBzjqNtC84
AWlQfhXffRZEJUB+d8cPnZs+7DzwXh1W5HzcSypIoiqL0fGcOeR5zt8KOHt0tPsI
eOyP4qFTJ1V2UnS4nbVjMMjm+BdH3aQHnK38CqZKkAY6vG4tm4iP+7Kv8NdKzk+y
TfCxQDmJn+rWd/3kaDyhtwIteJw0+y5wkXEdjfjeJLQudD0apKKTaVn0ALSQ5noD
5yiYbVjYOuJubdI+BeUoR7LQF9Px9y4AH94sFO16pm1zP5eQkAYNSEwl23RlUN10
pwu4DTF3zglIJwH1BvS6scET23sMfbL9QFgMSxnZVGX7xKDAv9HfDLvVrGAd+K+8
erX0Nbrsf85bTzQkpuumsPg4iOqPC4oD2SNk65wSJjabKPlZecrfXMiFe5p9rXLA
LTE7CDd9J7MvPKglb0Ln4S9RRtdeuFzak6OCD2aUi+uy9TlPd+oAFgl6/3ErDTao
7rMv2J4JkEwheCm2t+6RDS5dpb6Ow3lhy1eW7IUIIpi9bfgwCYGJH4ykVAjX6YN5
R3vIfV7dAL2iDmizAgcKcYCz8ImiST0034uaaa6DnggDqjWTetyC1EGlEV+ax7uu
mLZSNidcHMLjny5GHN0TW39Z5RGT521oq3ZRTOEDkE/cOTZP4Myd9gplsndplUPY
HnxKM9qJg8t/JR9ADmrATt97onoRCDhMjZHgYrLqR/NI3+ormrtqz+k/bD+S+bl4
VtiJqVF2gtmzDnDPKztW27hWyHllFckwRPrXi6p7/HSLMevycXJVpdLn2u+vrUK3
Y8EWKHCSSyw724hi+f1P1zdsdAK9hny8+LcH24Cn2JD1awE7TXqs+64puTg0x6SW
xj1ZI1cSIjChc/Y7+te/xMpOZa0lP6eg8B7U1AWy4bwdRFBhcySa7yWzQYr9bPJD
Jp0aYQXkQ+4QplFPXdMeRABoJhU+2NJ6emyVvMXWnjCvC/UC/KI27YV9/2EdqyFa
0gJqYuYcp0R1ajAAeN69nkHBU8gMxl45USf0hlbMcSeyVIuxq4HkIcnvl/PZ7yHl
XVanbUcvb/lLVD6yNTmCxf87CmGa1Llt4IWoaL/dvnq4DnjBjJbYI54nx6m3eD7S
J9Zqu3ydS18glxHwh21Z9PGxmNEDkj9dgiK2aR9BrlWfn7GGXmFBOK7BqwqKUr74
drkqGB+XGMDRnF3J2E5oMqonVCXBYVj3kxlQdUz0fzvVSvCm3GkB1VQiJa6aCkXP
qLkAyDZsmYuDVb6k/ymLUg0P5h4sXPBxHhAjSGn3HiTScWZPJBDw1A0kqr1pH8S/
Y8HGqmGXIa5JL0czBRsrbavrKfw3QEejsNsrgsa85/FH9c6vXd6wn13s4tFpWt0w
kDVCFGmv1xGBlUL1wNs0SxazS58q8HcTArYUJ1cHcGoRSXBcXrUmnxGJnRT4wfme
Eww4uwF0wOzXeX3S8z6/b5rtLQSfVdIcDdWt3eBPjjeh1x0Au3iX/1hvyYRM+WDO
snXTPZ34rNp1+exLbtM/SW1hirGBeidqV7tTe7NeBz+pE5+xNEFn2OlUisRSaO+J
Tyk8I5eWiR/dwr8iA9QwJqGjDTou0pCbTZIOHlNPx97FIqygge+oj5XPSM2IV2Ni
JPIugil/u+cq4d8GvCq5M+2+X4/6e/pWwcFLeJnHuudh4kY3+MFFyQs/iP1qhTYn
vmxfk5nQkLzHKhAadjOLSE6lphjJd/HizbZZk2piA2ROGxd+uH4id6RQ4+6Bt9Cl
AqUpqVyvmpNDddjm6YRIb1o/XMRXZCY4exTbIM/lnbmT8mqbFhZRqEBI2210jWcS
vU6NOvt6sK3eroH1AMKit0hVYvtrcvhdD/gGfR7eKBBrUxDaJDjjLkHXb+chbJUm
67vUTjib1tjFOHyICATBubxjXpFPQUbnr5XRd73IO3RzUKuemHBuKrJnOSnmGBdd
NBXYj1rxjlcTP9+0Yh5EH7gC7kMxnBywEdNODZBP2M3yVzdywH32hqVQhkbzns48
zJcNBvyrB9FSsTMaSrEYkwx4Q91eIKfIPwxseNrKGgvEgIOGC10GAN9EF/pA/p78
dK8o+Vow8Ozev4/D9pfwJeTeNgElliUV7yA4SFWPw/46Lq6u2UgJvN0ii89S71U6
ZaTmzQJO0ydeAIDUfX1NR7NYRQxuedAVqh2ODYLl/WqSshtv1xjsTDDnZp73tOHT
3OjCSXiCXtc4ye7miCVMO6se4LgprLmGiXsCBklY7u3jTja5gNLTGnATJOH/rCLp
1gnHLoZeunlKKqAQr/4yexNYE3CW73/LADUj5JvhSa9KUWSoIj7pszb+pq789i6m
+99n2ZBhwxl/KiBm83fs1AmIiDltuMPMjFnlI0JUzit/hH7eTrTU4PA/8/T+3051
hakDcF/+wum+bLKFMldBKoHEWqbYt0bOnBI1N5+zMAoGZAfPVcMx1YObsPFL/d1W
M8b9fgTX5jfpFfu2g5NTEViW7GYhkRzvDL08Wv96i3wnemuKMOFpDKUuKiRtmDQM
eWDEXckzcvdie8wT7wR54079fei3SYKHZP0URDU6U6/c2w78KfYWV7FCKJQWzRar
hcaUAq81nsEzJHqf90DZe6+V16M5UVgqTa9Z2VFKt54lcqWp8rafaxFPHg6ERaZY
gLHCdvkiZRwB1d+Xd47OgBfKaQHPiKiXOmCgq/TxUa6o+j0V/0zyaHHclNpZRK1/
NOMZTLzc9dSE479yt5bCNzJSL+JFGngCpUwpYG3fnw9O3qtS1Gox1p0LxUVm8qs2
8tQIRzhOUPGmVhDKSsVWaRtgaNv61s8OfC1gyRUG9n7e6iRU2BD27KAxvn4MYlvx
ShibZLufVPSl73xiJQ+nfdK4+4NqTg4x6RrFx3cl/8JsVke3v6Kz0JFfqvyZ2HYH
GtPOyJ6kqXgmlgRDx/p373mhET+7l4XjK17jEvyKorNu3MHdNt+xkGON4G596ShP
PdeRLVKl5AVGGZzhlFA64YjlCAdl6sHRJ3zdGtI76LBe60lBfuXwFd7PlnQd+Dfi
4Zh7L82Y1MGTA8Oh1Pe+5CA/6IBJVX3vJC59RPkOi9pom004M/lG8pIBRvxpElHx
EjdrgQOk3lAP0uQO1nkpXRD5sNgJeLB6UaTtfPYJHySEHxbuOpXJLkt3hnIZ5jGw
+A3Y0IlGlCthRa2SthyPIitefko8PK3zPT0CM4xcgyb68Cby4tYWw1rKpKcyk3Uv
Z+UOifl8ZieFhMCEkk7wMM+FXQhBklSUMDq5kINuAcxQJCghRkAM+3W+2ADD7pG/
xp2FtHM3aIC8vgG00yOaHFNzlFb581AOaxOFU93ryYtMX6qqyIl636zaFkOPUtg4
2se3gH79DzwGa7A+PfA7l1hDXgmP2jGgVZTRPzhG5ffH3wz0iTg0FSTL/Y2e/Ev9
tEmiDi2l2SLz6jY30r9lUZcG+T6j0ZUPbc06cUJVKMX5KERKhKG8zHX6h+kq/4GJ
M0ZOAFcgz3EvZi+x/lAX+4MvVO5xAfBLan7W+biCIIl3IgYYbby8exWPiL6gJYff
uk0wQS/7D1d5o2bat0sAqWf/vq/zg2VL6cvsx/NRyFZIQEJXPMTJUltoOqew0JPF
Cog1/EnvnU907oJvKvREl9HryHceLq3LNm9JeeWVtZ3tXKiHDrEF3gpPkcjItHeB
O/X5V6bktYCGfeWWFfvzmKehgLYwF3y/r5BTVum9iOaPsMeHpWrqeR0C0dWBfD+E
WUIn0hu6LqRUMy3wdWNxG2vSfTTQZpW1uC4VIFEEMqai4hPFXdPz1YZfwT0mzqsr
TD1ftiOrHlPH7x+yojlSK/gxaumODVLHjHCeHcchjRfqQzAlKGN4MzxLB7WR0XbJ
oGxDcib2/dyz7CrCq0jSdcZVmIvNToCoX9y+PYEhUwETuYxkdx40eP/td/0I78nn
msCIqrStGqe4O1LHhPqKOH0Srf3NpkHqZghwsws605u1rys31ZNUHW64XZf9wJvF
hBS+2iwF+Gon666fNQu/FQ5qFs5O4mo8VhSOrE3iYX0rvjwA3LMb2jWrsx5ggb+1
MAlgI9YlbYHhKm3wUSgqVIzA7cbvqLoG/KZXy4Zf0SgcqIDk82Oi4NdOqtPdahzh
Sg4ls3Nn0JRnKbo7EWf3UZvYI6i2PplG/Cro3JvGb1QPFXfClUN2Jo7+VQUMIuyZ
AMmvWYGN//+FURRIJ5lkWiGfRegLMtS3Ib8+6390DsJxLqOKczuKdDJI6LACuA+D
OIcOeeK7OIzc3jJHMlxXFUPzOfLklYCgRIDi2jm70IOyPyClO0mKBJ0A+l9eTquu
kqNrHpyvHo/NVIJigliIeTRv9l81bVxQ43N7GN1q/gVgRqg6F/yQXDDBVqrY5thU
3q169q1tgiUGtwLYf670pjb1CM79eBl6lma80RmrsQmPtyPIlxe+d1dYvbpoSfQd
1jLEgiMshmaCP5zt/dvV109X0H/0aDmBqfOAZGvDZ5QQ7+mK4OJrvXvBJfaCgL/9
8itiifOxiEne93GYwtXtogkft4lYYuxfpZHNy+aW/wD2y7dGP+xvSoPh1n8PjcPw
fwZmpVTvrSkY4g5e0bWgoDo5Z9vma4BDb4hfvKW0KYd6o2drSVf3GK4mODCi2b4d
U7oIKgnjrSuncKBnF/XFC2hyqcmamhjKAzfHp71WBeJe3K49qbGyHu2/pjarD96j
2KX0mdnezVl9Q5HoEtP0I4ch2LmUjiyF3xjPTyzrXSvfwPm6lJHeS6as+e8OFl6C
Pr3JxwZyBHVSihfFTb/rBWAKEsiKuI+P7Z1oc4pb0j3W2QW2YDYG0Lz5j8c66CFH
Tcl2iDAHHg3MqNvpz2JUoBcY6YliCoToSy80lS1ZvIH5IB+0g1ySysi4MSakSHcq
GhOmSZipzK2r9J06dnJ01v129LRnAhEaJ90hvM07deFbSPF3XVXp/hdPqtPPQOlC
B6MgXdO0p1LdrgL1akfyDmo3k/RlM8YiLN+d/JoV7isIQIgJApNuIDgGANgnOh11
HFm9EYMqz14fw3f9CyHfBIv9BS4s/9Oy6M3u8FXmz1HaNL69QiJ87TQBO5dIEtGr
U2m9rdLAB6hFQ96TALk2gJuPPK9zNsOMmAYVXyzsBTi/IdHF1uiMgfgNJflgamQE
TQTXRFY4ZbvqQrkYmXeXuepMxENEGeWQQo/ysUsq1YY1pHWYDo8dfvCDwTtjaAzm
Wjw7Pn9t1zBFgnqfK/QX66IioYuH2L4Ev9FWLxV1anOOacU02ataPYv1x7timJse
55ZEBpUlfiAsCDJ34c7S0w/VmCy8zy3+WqTENgEopoU8lRfefmI7Xp0Xakxw1/od
6NAmDQ2gaedxZIssGjf+6129eDQzBWat7ukcmBQfwoFV+MHzD/pTFMHp9fwbbLFL
QlTK/1AqwGs2/NME4Wf6sTDAzw2YTckvNomQQj96Dxp33WAVispid2A/r5ZYc9+x
vUgBzISeijJef8JLgMKZZ7Q5JFht7iMjbQBcRql6GRNe2TWT3qmAfeAcuWKXLgZ1
O80S2gb1DM58i0s0HYsFaD0CKA6wU2g3sw73cWzlC0qWLFQ+f49m6CaICdNUkLtA
ROkJFDklsKH7RmOlM3I349aTOJCvBuXGi1K48N/KDJ2jy8KYajb3xDRpQbc32CEz
x6WgfMecoe9J0eb5SeWSKhfTxDPiDqXbsXPTLW6hyznwmupCE9Kiq2TgBE273+GU
3MQaCJ+Q2QLfkK9oiv8G9sO6sOr9EKlkHs5FmVyUlkVuQnt9WfWbPxvYgl2eMehq
NxYibssu+V5Y67CFFv6i7N9an1BkPk8BkSWBBLi2NXbixBzdTBtoc5Grf2mLWP6G
1ezPBO//cKIE++RkBd/H+/N6FZD22P6NW8ZGmJqam95mU6SUnxnt4gJdStwUCnTB
0VZPz/XUAH4V4TxmK9PUeuN1RPcMEbCZQBAqd8ipA4Zx3aRT9HLeqkC/AN7ILPlv
+pxkEanOpj9m+nBJLhp/WznWG8RFdjNSgTb3F8CY9Cyjz2qm0OpcJVkLdqEkOSdg
TexImbENrFaG9mkPVsYL8Y/y1Ssr/4cjDHTLz/9SajBVejzDhArPYm5shKcFqo0L
Tja/VDT389qDMU+I+LWK+Nt16cbXHxn2nI0n+iMYVVLrVLnfMBjgamgiUDjazQjs
vS4jrQE56nGTx+jE2s5bi+zEqSpmEgZT3h2V61r+OtgQsf8OFqo09ho8mphZtCJo
Gt36LkBoiBqeGelW9x/b/RweoI17Cn8ozuYGfCFG2wH+fwN1TFbSJY4uDzWGy6ig
OmReQJR6htLMJAzN84r0pgOT2bIRCgvbQfV2GBd22wrZwuiAPBkECVuB394L44BN
vndb9gOtI3TDk1Cknoex/nC69JXPqUuQwnaub/7Sg3D8hWQLncfZ20XvsSkXFGs2
yhNAKzaxUmCiCkxO4vbIMNk8+9vUhNR4/2TLRwAG4tVe2A8NPoSqbExapwtOeFT1
hnp4a6gaZh7KA1G86mePhYDg/fAOfx6GzSvKnpbF0LgZrnIyZMbZHNTX0AdyAiV3
mBcnuGWNFnhlh8Rr/q+zodCqeEra0rD6Vlv2do4OqaW/xKvwpObAA3Fhp0ArPv9X
3J8tuqI9UFMxXxolqmTZolW2mG8vS3v/fa+DS8DnQgG/0ePybzV9NQXMCw5Qvyap
Yk4sgSu1ymgZrhzPEXAnOalHxbcSAp5R4qw3TAe+NMLvs0MnwAOD0kJCNgQ2cdOb
o/Jr4W6KB1xdAs/mkTf02Thiexe/SI2pfgPcw7XTjt7eHphkcoRf0nnLGC57sSWl
hUM/XJCs48H6jk3croABgab06FhpJCKFUSUrQj8RNcZOqvP0UTZdUBocgsTIO6ca
3IpNZT025razIb2y8pqn0og3W/Ew1kWwM7BqjnAeOWpgU86cN8lAXVoX702ORCMO
GV7Yjb4QMMt3u8QunujDQBhNbnx0ZbGLK5eB5N8GmzXiEZYyFgOT0WRqvOCMJydQ
r6FFvWCNY4ga4r7mbj9pEWL/l/zS1PoYzH+SQLKDUEML+sJwyZIz17hJ1F3h7sHp
ICTQ9jK0ugSvhw/e1X/InER5dPQv94B/sYImpdd03C+2JlybE0JMuwtxREhIpxnJ
H9sYRvuVdorfV3rrt90fTMJebydFBWxqOr2KhoiqoJ60uTCgTqadnZHIZWHvurxV
9GUnny1CLpW6+KO0xGvx77slrY80Fo7I7bSDnmHkJMwgzyNipmARAXUA6+YRoGLW
FCwATzSdYZZpZasfUCgE9a/GamKPatie7WEi8wtDDtR66hqdbzqyBc3q6+fZRTph
ZxvmvFMYKd1dFPUMBn2P5ij2/RpnmjNdtLAwXqSmEk08UXEniYa2dvqRQSpRa/b9
wNsj+oF4Y+/2tonBEKPHWK6Rk2w25l3hZ0nImcBrgXc7Fm8rmwWFtJ3AGXd4HUlI
kCxYzEl8ze8A+en4yrV+WxMGSxpxB05MsJI/nfnadoEF6cbg5N6miPag7h+D+Gwt
E7R+8/0bG7XCpdKResD0wBVtpGrF6rRkAbUVO0p5J0BUJk+xtVL3omSqJiSQ8DWk
g+Zd+4WmhiJ14Jdf8m7zQPR2M1DJPtckLz1PLja1Jvb8Jw/mKf9WxtX2Yb25Dl0y
G/Wz+asi1y3tmjdB8pzWoipuQOdySRsxcka9RUGU5Cdqx/zcKZKiO9ZQRk0VGofP
HKP7J3ZnNFnZlB9SxfLHorUKJ0qzMYoS3XKbIB6+CR+w7OFaYtKcTohS0SQTVeIN
w+PEsWePhImj10bfxkKmCm1Cnps/x0FiolBQE8Vf0DIJHe5Ske7GBC5rBF0LF3ox
D6gtdj4SDntR6nRXyX6zt87QPoojLTj7ZOAM4bvGAN/fqQtMGKmHuqXsPEEmCaZg
cy6uCUdVxRhbKiECdRgZus3gFAgXIL7916Eibrf161scKjm89ixNI/cZRS3bo2kY
HYMire5zlxLC+3MR+s0e6nDL5sEMUopIEkRvUd08fyLbFmqntGYiXwWrFPLnSz+l
0axVxF080sKMC+T7fdFSvJ+in+dLGIJ0qOBSxVZqxNGcKjTW6RAZ5Hi8//HrFiRu
Xrfi4humakTFK+SI8vGuTAY4fNPBq1/1CymaG3sA5qXjtGiCHcnUBBmweMP/kM/T
aA+yiVnMJXnvXejsF8dJ2pl2z4hQvSk5P/wX+LRnvhoyGpP5yb+ri0Ye1u9P0+Ef
Q1tscJl2nmM1E9l9uRjiB+iAfQjFkHsF5rDFi8jSkCy1o1rWKJ0SOf/YpeHozy+w
ejDn5RoaU5ht2YsPT3vFyUvaygzUmyYFHfAjWNw7EiDVtm4ISFaiKxt4ntNoV/1q
prjBgSuCWSxkyyB851oLZ6aHIpDQfWM7qwob7x1B3PABGmdcd6/eYwCMEMK84CJS
gYi/ai7VU/H/U+QuF101UwvyPP4XUyRZt8AenHObnt27RU414Vg+/4nvLYi44RhJ
qPUA4z1Gh/ukc6dfliLioHfxPRZDeHk0nKQUEEdc/0oOHvI/dZIOOwkew7vNoH4o
FbWRxfYA++CuaaUDneh5Wvj6A5AD7La9af0OZjQV1lBeO+w9AbeN2C0rKzHnEYwB
SBIDQXK7SRZ8ytubY4twjOiYVuq0DsjIMKWj1tdA5c+JWGwzSW033/bzEuawo1Gv
62fLc1O7v2FXQh8tl99+ptXvYBjg4MVIuxx9RLgckKpSRLCYBnrJZkBny6MX9Mnx
BxoLQRT7eQ9hfAcntNO/l55KfYM3RCaJjflndd8pA2zEkFs+9AaqRWW5NBjz1tJf
Q1CX8vCg4JMSpIi4+njD3QtJNgt08p4hUrJoJDqdvttoasf6Q5z4DT3bSvjNi8ZF
zSf0qG8cakPbYLvPp9Lh8ZZl4YSt42No3fH19GU0MFJYHVef+8aq8m2wYMuyRfnx
1tEeXkUjpbv/KHRrXcPXbAvKECrsP+uUM0cxAjb1s8djU28qDielDURKyBFxKcKl
9JK+iG8lC0HHOanF6xQZ6mGA2gZ9CIRuP3GpOb5JQZbvG6M+6g4zxND95kUHKDVk
WtORrSsSANsnrhJttpJvU3kQHzmlX171qWDDHhwNgECQqtSTcrETz/dbAUfQSGY0
t06UM6YhnWFA7pVDOO+alTrngnJKKWNoh0nSBV5N/paFhWQH84l0HPz6rR+E1CoP
hFEgZqc9mjS8xxUlekuCewjJidVcbeoEKSe/KmPRH+O+Tz/DymFLFsMJjkUUX0et
5YxqS4lH/beJsYCmHKo+wBSny+BUOvd58b3qlFTARFjgiNN90iMePsqY7SVyAvCN
x7NqGCqp/EctdrznohJy4+hQsk4zqJBdawvauydCL6G36Q86Km7dkVsTrvRJHQ48
V3kH4H5JV8xHxnkMFst9DcH51WbE6f52eJ06kUiSk0ihu6zzw/nZYtZICKJcqvFJ
vjMSASKtJqJaMCYBD8piehMOOV/krgkNZ/rmyBUvC3oP5PyQfznyZqP4VK7DRAIm
NaCqUd/v+hTYJZfy+XHGOkqvfSsKGoIeChL8OIpSqAWQBcaTYZ1CUcZ6gDJfgcgP
UfSEXaE3hSj5jR2ml0DyJKojMrpYtGrGf7jE058CykoNsyzcnJidmTCGD173jpqx
S3CJbAH/QZdiDyeOBsBAs5eePWLxiRb4RhxaTOa6LJfmBqRcwhqasf6xFa8CwlxL
zmNDEDGorxsXAwpeHKAThHs2ivxqih3l+BBAxMWIEfBTs6FqK95nVp5wUG2NhcPT
/tPLUckz41jmEye0Va8b9tWNiQmfqSo1ZSYiLFy6ssRZ98vN116gS1GHaDac2Akw
vFmMueU9CACmRWbPOyAnY7n/WWIVtLUH6AQD0LwTszBmb7wGNjUhskSfKn9LwRuv
TV3zfCmhYGF2fE00GEC/l5iazr1zOC3Qr0nF6vpfPE8Ur1f1AesX/r9xyNNK5pOy
nERDZ0az8/f1/3Hc92zzRZlYdkUdyj0Q6+D1vljMkVXC4LjJ7dKUpQpnDbMX4P1l
VXmrsmDnk39eFqGAsnNadpRvDi1hJ2iBB984c6JrpV5uKuat/C0/mDn5drgucJNs
lGU+3cG6Rvt1kK4aPAd369lK0lyhNkWh1Msys4aW3ybiOel0bkKYPupncvQ0dotB
s3nft3MF2cVMPA34TJNRnd+21S+B+ByuMr+ajfHOArdaQpVIQS9+vDEyBuQ5NEl6
cHVjdeaX7mTJeck2Dr5pdAGK142Fe4pqOwMYcYJaL9U3BAsaVOEUnYDgOuCgp1+f
fPdRcVOjbhr6qaL58cXUDBSQhO3IybLVWDRJPodZ6huadRK8ege/BA7PHz0offOQ
OIzEPJQouH3RKFU6pJgPbQyc9rhavUaG/XbXhZJCbY9Y6cA4wOiax0+ZGtZ6zHNY
RG4nDGplGKpIoPomBmCGx6sTzYBy0N/IKtc7A0b4sH1sQsgNTQcK/hQGjzmy7Zdt
XZMgDkE2f6ulcShB9RxJbMvtqC2RK48HfIb5KZqMM7ryznimDB6NALP4VBDTBUlR
uYewtBKcFXW0u3In0lb8rTToEBrOmc3XCxnk0jEtKfrmRAkhH6dB8nbjyHmFWCiI
WHfk6MhD2S/5cdKa158n6lObuGkyAaNPq1+T18jXVy7AOYgPQEsGRoCX29gdlhhS
U0trc7Q5t+YDReMJCZ0UaKrw5xHuLdUWqOUVp0ymjLSLMErQWIxbHTkEWVQfgm1R
Bm35feyivGlMIByZlZhD+upgbbM6or0u3kYMIeCTokYNH01FVyvTs6dViYfCHEcU
XhDXhnL6Xk7s2NEZydU3q4v9V9INMTcJG4HO4H9rBb8/BMHTSTt14odVtFNzGsAS
l8jSy6QedYpUKsY/9sjPwC8BABIB2YrcwX/Wz6eEyXrasyjVrwCKGzgtMhte99+6
dju5uQZhoWfwGI7E5dLtPwDHCD/mPfaXFun6MYJeu8bmp719NNGjqz86qDH9R+41
R/sZxYNEbZlKgnRTmZgSk6QCAoql5L/CluF0a8/1sIYWmB5K7MXUkh5JGsupU+cW
RF/kDgKaNBziRsLvOu+WK+PcDYPE3q3D3Kve5AYQUCWHm0AQY4/O67/q27n90j1B
23jKDPgdwVZ536b2k6OrAJpyir6Y5lr+Jm8EPH2bTXFkguklgCHCkL/+GiinQn7D
olEiDvNFtKKuTaeHiPDp49sJWJ896UIrEu7veKK8KZ0VUJxuKvPEMjFW8Cnmq7GX
MuoKU8dfBQq2kEfWnfU4R/G6Qp8UBgUcl9KR35dYBXoLuhbMORSBDUxR2/gwIt32
dZfLb5QDB6PS4EIbOh+CHj92JyehZXdOdDJuNCb8eQKxbGgYrsficD+jiYVr8qEx
HayLrOWZ19tjMzo/FbHEP0R/Gm6Ra0MSuFCs4dk4OQKZ3uFihlYza/BIBMdUvxEb
tsUj9CdLagGxAPEOyintF8rWz5bBUgAyxzri+gmeJ/EV2zTEGszO5pk/h52nKQw8
sL9wlQsAeKtx+MdqUvQyZV6IAHrnbo350Dg/Fgm9IHTWQRNwuOdgeOnzVjlnZb8o
56ji73NsJOXovhaOVjTn7yb2tOaRF1KuOk3FLJWbZwl21CIDATKgMBonpS8SkEjx
Oz9i30fIMjFzgBgp4zz6ZP9+24F667AyLj46IgYunn+gAqTjxqUCOU6PtgyePhBh
wunfcvk6cgbPh43so7ij8T5QFtF7EeGU7PSD6bYWTuI7OMejUkqrRlX4+Ug91ggL
NMIu3h2eoQsNQQaNq8Qd5Mr+4R26J6fpxRpNPuyboXeI+7oLTNbM5dGlxaj0AYU1
gFRkOj9dGZxbpCfr5b300vokvXhusPydsNArb9eO2trpgz3XvI2NcdsfNno2pqWB
Epm28xDzaC/LnC/8Exh5wNt0LK1fPOgrRiyrriKYv4KFYljyWjIe46YGhcpBwRzT
W8g3IQEDfnxAo3cxiZougpCdxNsCnClnd/bMiuKz/EUgIT6c7LI9Ud/g6zYmLO/j
W+c2cG/aPyViLHCjTIDqsyP4bSrFocw19paAJhzI+xrUHVI/G7BpN7tqMCrIPoyE
DguKJzzrK+fALUbYypgz5iHJNdDgPHOC7WJiUOd3QF2rqSy1RywPQFgV0bIkcJju
Ij0lpP6XRpa/nwpVJFt3Xz0w6yHWmXhtgmu2G/N2mE6J6S385YqPNSXXmd6qY+3b
7yo/DwCUHenpENZKgZBkTItmSKaiNjBKxb2s7y4f6y4iBf6jaaNzhz8Np2Xg5Qwa
EiFp3/TRKI8OhaR351/Iw90gdhP/TXDEMWFTZEPGR+sxGjiQk8DVKXLxMVxDXOlu
XvNGURjpDXzhGHAqovptCDeL7k+FtAYisCG0bIhugB9SoXT92J6HjVX0e9sdGjf+
7v4xhEUX+zBqkExEBuQIfZSdVZwq021sMBEW4gWLt2DFi3RmKw7fSWpzxDvu3FGA
KlGa4p+IA41HEm1C/Xh5Q+IO/jAv6minvN7lC2Ydq40aVu/iRBNcSBmordbKcx2X
358YRoBvp77gCLwhsOJ7ptaJEMzJ4PV/i28GKFBCvE1uQ2e7y2QdpbiLcYGyHjZL
khzgc5JK7bFr6DH7UGenjNXb7xs3P1iihbaBCsna5nump8ADYn5DuMv/XGGIJhBn
rVd5dYNJKpmLQdIkQ+LockfKBNjpWv1i0kB6O8tOtRbya/3uJ1RseHoqr2tFiwdC
DKUDc+ONVUFh8H+bfqbDZ+V2LeD6Z/vkvx7sFKear/K+DUK8vGgDs9ChNP+CStTL
V5iV1Q0z1t4/F9JUexg6VU1Iz/cz6kRkOblMnxgf8ccjmbwzK07109/lsNjn2JQ+
SK2LzD5AjnAIzE8bs/0QfpEehrjjjBtKzdSc1TnfyCYOQdJbsmGkzKO8BMg9vHC7
bOpwKaaFyh0+4qRNNmEPoL2wkwi8LavbbjN8kR1kc1cf9UlGy157GTxEA29066af
004nQXry+IuBzOvwJxfFUTamP6sQo73kVcaYHCSmT5M0VEjOs79VPq2iK0bs1Sju
2IATuV8bY4AjWWrRzLLSTwiUpQcxhOJ1gI9gvQSz5Codu0ObHNkJyTgZ26xRscgn
fkBQ6B7gh/UYFdgonkMuAZgq9IG3JsyZW4BpwzPn1G3jym60dKVbXQcUfDuk0yx/
DqxB3XVvH8wCUe56ZumRjoxf6dcpiBOpesEi1TeGHdZrfQD18vwMH2ol3+F/qKsc
rugrqseUjp6VnQw3ylQhSOmxWisFBlZ5M9UZyuU4dMO5WJTtHEbQ6ZovYRbBBmDD
QaC1DQporKt8RhqFIiIslVSnunQ/P0NUECCcpHE6EDWanBetMCVvQnVBepaX+Hh5
ASnZv6wwPwd5HSOV3mf66iFzURzrjSCYW+PHi/xTjKZZ9HJpPYCIjYogRS0m5c5z
dxktgK/M+bW93aI7DaIOAta5o8q7cPsoyJvDV2IgGvfIvefrDvCjcxlb3W5XE/6S
SiKCP/HXrbPg+WmIlQCmGzrNSwuGyGRZ4Hwl5XZV4Z7hg/M9BGCvmchOqoGNbx9i
cF8Z5fFB04NodYbKqP3YIS9w9GVX9lI4MP/2rMxmKHl9OF2Fs8TiJSCslcFHtlcr
ZP99cb1xZRA7v4QSobX9v91+j3MYix6Vhy4OPxU8kAU5RgKrXqRkCtM42RKTHEfp
74XBtJpKm8ILuQS0ZTPy2pVPf0nPLLpTnhkLjRLYGjK6wjUoKo5grs/sZeF8vw4g
n8rcfswqxarwaBEMOlWRpq1jTmALiyI2TEckhEz7FOy9hYpFI1ZeFAFABf6QFyr5
MA9MHs12Y2ES1hlWhuhB59SiAymowtb6GMy596Gpj28y2KThqQvfqBGKAJ0NBQZv
EQvzLyTQnic3KdnsTLQeWKNWitUuherRQ0yA4aIfCZOoIve3r+0Htyd/Km8YxRM5
tHRw3njZmSrkXzGQFAh5/GZFYdOakQhKbf84q8JBWkEIp39apAVyRz26UZT4ublz
maZH6JscgqBtWFRmm9wJRTNuM4GFtXOxV0LUff+x0gXVDPQ2yh9KGnA9C19RliaZ
a5n82v13RIDHP0LbTkgJ182T4W0yF1zroTTEU32cQAoMj2RxXVpXoHXxnZHpLFd3
t/wnUzc4FJS2zE8LJpzL/y3y7CkLocnbyF4nczp9K00J4aPJBwUJb/snOal3/Q1C
s7lDtJ5YejYMRC3ahsNSU6L0FbNOn4Va6iK0s1NFR9WmAuClpHdutNo6WPZ21pqb
gxUCrKqVJKsLpgJVfnSi3LZm0a7RsJeuxWtbqUjQLNZolwJXPDeYx0xAXjD6LxG/
krD+NKedh2ngIHPMCJXmh2NPAWTZMd6MPgDj6c+zftZTxiAfhKGg8yBhbwYtn9f1
B3oaQHmpfyo8WPmhxCKX4MlXPA0Cd05ucaw5ZuE43e82bvQDVP70UQCrS6/iZg/5
62SZjVgAEnAxout5xyYXg0xgO3Vaah5rpfyuV1REwHbisZSMtaU1YnUhvcf9G62o
nxnHErPGtm+e7miNA73K8YAog29tP5psoVh5CKTRYxg/FUuoKnvRO8VJkUD5BaZv
i0lEVcocf7Xi46tlEb+q2CHpt5O+qZt9MjVU0VrBvNdbZiqwE8hR5Pm7l8nRf3JA
ZqKmkS0VeGgwpsUT8igECYRcY6lFh0mOkhBxaZiTGxWnCfg0NI+lagDAgdJBdMS0
SDQdmo5SlK78lITZH/WfEX1KCyVvhRWTOnTBLlPqXGOtjB+invaz+fKSESjq6/Kr
W1x+FKt2Zo94HQJK5z3Vv/iJwfIbvEaQ8uGyinNyYuni4679Zgwv2+mzHOqzkeL0
2x8lN2y5NceHNj2sFV52Ihvo+gmcFBYoGFj3JEZXDeHt4JRhUcXVCnPITO3xRxmw
QJfBzaJiISqdvwhxtjJPYFrJA319QFHdoW/cLD32al9iliT+ngIYMPdaJWMCeWpg
Zq8lkAo3ZY2MxR9qmFeTGU2BrHBZmLhSDSV20NHqn47hAyzy3PAbzSf4Fpkicm0P
v1ml0I+B49vujXOEGHkMVOaYrM/Iu59M/WES8LZQnBkvslEQQGoNVQR9/ZhOHDED
Ieb13nzs3VTioPWT/BfZq4jrhUvFHjSgtFusxQyqYlHn2mbMGJjTYskDQyBnt5v8
0bJUbFNM4NK48PFljF7IjfR3aI7I6U8S5RL1My1WemOuUP/wskz3oOFPZjHby103
ge1n/ySGTk/eSaAv/iAvCtcGtuY5RHqrE3vvK6jrNM9udrJHvygwp8XjNPA4ZdlI
DnVsDTZIA56GO1x4TedVcyInRlzT2c3PF1rAfRBnXmzaS3uA2SrEX1vMDvZnc2RZ
YFCEFXwl3lbYNaB8495vCrjhmn4+Pz9UyI61/fPSMLDe9xQW5coJHOx/M+tTbrnx
6lW01k3y26OnO7WFg6p3ziyFb4ZVN+EpwbMpmCHWoFkKq5eL6mZTri9JstDWXNQd
msXzZsfFLdC6rc+/YTYzoo/5r74FBInrMAkPVfvRTpNuPYKhMAFE3fe6vAzPKGlB
pHPY6lfX9cUwcxmscjRat5lpLBkU8VuCXCUzLj+fKetAoZbZsNG4CcnXIITGjU8O
m6pa8qpL315tEoqZjWWU4b66WrP3yltM9kDBfV+yQwrBVT3eN3GQcC1k8R5Dee5D
kI+eF7GwjtIIV9y2Nqekjqg3m1d82xo0q8FnIlUjrSmeWNZUn3M0U9IIxfubhh8A
XuUeiSS1J0qXB0CqbJTN+Zb4QxVV/d5pzSDxikRHVYTPzAPi3tsvoSTmEPj2FG5v
1mrKevZlPflBtXlcm5E6rM/r8pe+uB/Y5o838zz7rjU664NpqBqZCF70ZpujQz/L
NY6xdk+PEsChdlMwTSaBdnpaklgQYHDIxjvCCKWXH9lL6IKrr/6depvQ8hQK50lF
2mezSunntj9+0ddumwmapqnVwnQAi8hzPdkIif9MUkbWXAkZYvM8xJi+wA+lOlkA
VbrR8AZPB4/uNG5UHyPfC17eDDvFASREbE0Ks7//3Fc42PgIks6k8zB22EbYFWrZ
zCG1MbhiqtIlTYsBXdCju8A3ppYPLb4COaOBcGN8rh3mFf59QjwUY3/aAu6iqSzT
KdmqUXIVH51+9XE7vuVMugYcYaIcwBwJ+FncvGdbmxlndGDuRTw/yw/nQWVynLpd
zKMSmKNRaA0kSJmnUZdg9K8SBE/4jJ7DYmAEi0+Ka47pANB1fjL7rh4Rv286YdSM
co/g6e72kCztYuJluFkwSbQ9Sj6cwboUSrBn1lbNNMjBo198heu6MFTnsIZRH6FZ
BJb0/pdYXHgZ/nZfHXvNACFnUCwrQO8/NnAOaYe+qc7RjmUooFMS3g0HlIHhx1dM
Zrkkiiolpf61hfxHv75PlJyojPF97EzWHR9VZHx2G45l0d1adVI6tfGNeVbSl56o
rwCYWLvnXbM8UaK/UBjzPKjLu0pcqCVsMMNCmRIGxqks1s2mU6yQKHAG5GgUlCnU
B7rOSSL+ZlxuA1Gm2tNYTFbRkkBZKOAjI5O36RejEF4GYwdQRwMQnPHTHRKtbGk4
sSa0KRjiHRfPdIVH1l7TVKD7rcza4HlF1ExF2hM8rEQaSS71JwH6jJ8me37k8oox
Ye3lKhlaBh922rzkeHpfKCysQTbH/Hz5ZIfmPkk4TyXJiQDjzfrXFzvsbEhDnlkT
gR5/jFpdEBWBF6PqHwcn0ul5aVR9KMJ2Jt2xFBzJFiA/Hb+Q0MttEQ0nB3jmAemJ
yf6BisFK/o5Z6Syi0HDAeTeb0D/MOLhW7+gdfTlZpNZjKSO12Ifzk2eZIQXO519g
wy7o3XG4mnl6WNzI0ZiXawws4DZ1Maw2vmuD/GVyYNKYGvhEtHBQd4dfxvT5Rhjv
fu4sPcHK62xYp2MQWqi80kNxbycSVkS5Vmgd+X1xRoQdch8t3Br7B5F+fFfXzItG
e3DMps2A+b3ZGfPs66v7c6axomZQ0cWZpVz1VTnyIlPtX8R0O0TRMotYJ2QVx7tg
F2LFmp3beL7PiVE8AEzRq3B5oCCSDS6wwK54aQ1cD0EkfyOr52VGaFxT0po136Tf
xmHLhTd7K9a7xDgrnBaVwDSIAlt9WhaeOfKfrvlD1iXbTg3qKX33nu3BHIDx+9tH
utmQMrctwsPec5WgEdd1uxg5t/lFErcpArWV+YCrFzvT1Evnfslhzml7ETg1fgv3
vm+83lTrAh10kADOtP5eeKKaDB9sSOYwE1VprFBVnUDnhw8NC0qCIYbWBstRX+ZW
J2laDnfq4RjxLtVXQ2WtmV1r+QEvIWGRKBpODFxLcAe8Ql6FDpMRB419gNefrHIU
an+aVgOcr6QGLDigoW/1xqxEJRlrcBuVlwXnMPCGJG4Tab0pcO8HwqKjjupgTwQt
hWb0+KFl5oOGLfEvo1r5c0JdSYgOJQ3w223bKM6tGRZP6dUvCVD42q/Z9OzuG4yY
Lh9Slk6LShOWNBi4wBjpcF2KAj3gMthykYuTmc+35043jCI4jZ5TfXW4jK0pXJZu
OvO250jzrbxKBeWDU79ztSbOkjXwdl239M5WQdWYoQPu0G6jAQ58l+eJOtxutsxC
yzT90UQx4ttfv5FtOWJAWt/jlUutjWlHEr5YtFf083s2TIMg+jC0Mcd/zQM/V0wv
dyCWl5L7/T8vV2pav2YeOnSVvCoRQ8MJwXC3xh8XlPhAejkAXXhH1oA3hTuJtW8/
DGA1mnCGCiBxZrQsvzgaFOKBiYyBY+tOCGsnBi2ufqUb5pMmvixoDRg8x6r0wphR
ooAIitvdO0RwEzvavRhuzSJJOeL/j2gxImCEVX+9zlyBw6YY/qOTlN8HDYblgvaq
gayfw352imQo7lS7WicwbhlRFwwMVJgD6Ql1j6WNBrmGjZIU+drIWhyF+kw80bvW
FkxWAEVNJ/DUsNCLFfvGb1lFQWB52pzDeDruv18GVReer1IfgICa0t1gH/q52/1E
8nyQ+ZnIYLu80KwDsKfTvZiiH2SFXEJYXwRr8gIyJnJ4j7U0QrVicwj/9VGqksax
I2VU71/uJ+HqHeQFo2NTLDRbc39l8xaGolRKeqB4B19SyxxGYSl04SoShq4VmDcn
OgeYInA+4FtPBu99e14JLHS8ZclQnwiaf3E0JAEIk1Z7c3CxhCYbPkG26w3rlXGW
ViiaOQrRUB2a3zOtiYit0mtv2qVVgrXqN1R5O9+JaGf4ZFRBkhdhhDOln8MMr4yU
R5+/0t7Vw9YwzJD5wU+gmd5L1vMUS8+OPGE9qYPQpKbzJSOqoBnxIFJmyV0A3YJJ
WadYU0F6q8GCC7XAh4sKliiMosFHpDKgzGJqrMrCoCvkpCy6xJyLy95AKpMNjpQr
yDiwCLQ7oM/u4iLKHE6J1oG5+SN21TAB6MYN+/NiiLn81IQUbTzuIG0Ti8HwryX2
rhFmdvGdpy3PkLs0bMawf/gxnCSnPmopxkty/vsJqy/NI2coj1P8O2yzNnAw1iit
JBnOFB8CU5T6h47V3aMFjSk+O4WCDag3tw/yjSp+eNIk1KXRkx5NN0oyenLoxRPR
qwe6n/jMJqiO0wJU4h38FX2RRZ8YHgXdnVNcADH08Q79SLcSyvf6HElPFtP0ffHB
4quckRKCWWlLPsh+NV9zrAi0ebl3OYlkF3/Lv6J4H6RHhGSc/N4bs5PrpQhhvgiE
O6x5qYtEz9C8Szb2Z0Jp1a++wyFsyu2VPNvfP3FpZKPD/+kxN/erEGRF8mZ8bkfV
KSJ6aj+fY4Ozfj4n8TOoe4BEId7lSC7A2UH5vOlST15Z5h5mUtqZtSRGMLOdQ/zz
dKNpQ7oslMrzpwRiAXmWScaoV9hrwz59R5PeLA+f93A+lpnyZ+KM7gHqA7pTiJK5
KkTWqFKuTnhLO8pfyqF403kVD+fUtrkljR6Cj/qOli58kCAGeIH1+LY2upxPR1W2
cAyRvu7Qn7AkNCBF6uzfz7YdWXX1Pl7vCuzvUPATkO15VgyIO8b6BVi6AJjuaFgC
Ik+WJUjGZSZwlkyfcL6d/RiBoUvF1/CHtcpX2Ri794WIO3uuRbBvy0fBwhezlwew
0B2kJkCFrGFDcr5z6cwrBE1S+o9c8OZVRal7GGNx2pWxpjXv40aeyjYnTZ2aklCZ
dHnf3yC+dsSMvW6mK8uAxBV8kzoWv3ZFeSGCzu7nbAJd5XNGZs769PwpPt+oFn2P
EG8p4Zxqr3/eMrQtnIlQCrwBiU89R0mlmBzSk8+r34gf1lwFID2TXbkY/EnQA5GS
mdedWnSkmE9fOaWEF4kTXdfolKew5YF+GVxRNQeLmXenq7FFfQcKNIA/ojM2asql
k0GwfqXaW61DCJVMaVlYTnwpoUpVB7EG+ved+zCtNSQmIylE2bVPpZao/yEDWoJy
dv/ZsKNymHsf9NIfEwpQk07Il+j+FBgqGbxlKIKNGJcW6I0N5u6eNtIcTzEWTFlG
maeBsmGftp5z5MbjWrUAzqT6VyhWl4xa+XbqWSl4q8TvX/U21WJ2feA56OD2b1y6
TYCn328ZhhGsbEqBbwoizRZvyUxs2mWzyL88COePb/FoCI2hplGBgIaZVkpJLwAK
eWWJ4nmvedvRIU0TpG9BJieiDjDzdaE/OyumgSuPYwfF7mzp/0P8iHkF4RYGBjg/
WCu9Oj70+/8kN9Q31CIPl47HdVpIXn6tfXf5QdIPgEU3zpcLwRP/lb6IWOkG1MTx
yfk9/H7Bpw78ORnieW7IeuEkMQQiTIckAN9rT6E1vOg7m5cAe1vHf722ymC3PxCm
eX7Yb0FHc8yRDpf2yCeB9oo54mf3DJ2qc2WhLnlWRZCoa6ekSomYtKEjFxI3WRiV
ApP5NdxV6J989pvrUKfqDPIDgek9+beN7lMbKPZPJw2QyPFuMMmaEW/ZV7eOr7fA
MqeldtSnjcrisjOdGRlQmZ3zzuMj4WMHM3rjQMPZXcWd5CTsT5NTRIRFrCkyO6xM
3qSuZXQrrT2WKvkSex7DTNc+YpEH1sjN9+AAd4n/I+HIdhhgVwgJN3DmKZnyWw5A
6AZKQjMbqGyfqzquFZfzUqH9KjO+jCG3iON3ud39DSxZt1pxV4Qow/mYoUaV7YcL
gImJmhao2kENeV5iHbyXKBYn28AllsQZIVc+/FfZqCYyfHaBGadPkfYKfJArGV/V
pJ85wfc1DmQ5oqap39XlrDDSE9SQUe/zpMFGsz41N8FPX9Sj6VFBGel+5yYC1ex3
2TdRg90ELBnLwe4ZgtcA4p3xlo4PhZjaLZD+tnHtbxCpMZ4+6RJTXJieZCr1IPTi
91pbrZ0IfuXmM+rR5uSZ3N4Pv4FRhCjSc7GEvzmq+eNynHZSQpQR10jt9CJ9Ywt0
+I3SfwyjdQTLYSrglZ0YLRybRwlYArbygu9uO3/ZhS27oapFF7dKVIqnyqxBNwCf
pYucNOmR6xKEnZ0SMuDM/0KIaFfmKp+ezwQp8Umr7T4FKW5abYMHGHmRSCKsXhS6
rCWxve1IpQstAbwpObdA/Iap98OqhLxxXM7y4/vkvDPMnQt3ROUvKmi08ko2BSKe
dXwmRtb5wy8yGwtHwi6RCvodtb1y9DZktLvKv4r1ktJFiqYw3xFTvyw/FaodM6IP
7b8SkoJ2sDZhdOaC2I0H4LaNPh3u7/7Qg4j3xKa8Mh2sd8zxpUchjwgpf5oWmFPc
q9FsS1eTRyIAjWNiaqLxFiOhZn5ZOQs59gZQqzTBMYGILHm0nhxM7vCQz/V0hTW7
JMIpcfA/rpFyYPlLO7amoYFqdMY3XMYpG/Wg1yG6ZGLxNROa4+UwrWLlZXBL/YpI
WuKKa34kXogYLKVUCgq1TJci8G697e91q+QeD8PTtykKbcRcMdRK7G5pz8wCE7c/
7bw2ikq6V/lTEBUOkWoal4OIMtHfZLmfEzxeo+IgWc+vbaF7XllO3wZPxIbixC16
oFEhF3XgNyRPO+y+h2x2GZdFQ3S+Rc5qZB4GOlo1k2D85SxOqWi0dcHyOGk8riW0
bbCm8PK66RuTa1No/kpgnJgQkXrtG3snAeZixa+pOy4OWXZ+POrqCXKaoK9fym9q
67ou4Es+Ksw+wpSrYLJqhQUDX/QI969HnmISVoJX8FfxvN+vH/KIUy4lYdduQHwA
wiRQPHliaVaX3g4g+VWjHcvP56/eFc7hdJw/tz0tdSPxzENGUcDSWGs2ORS/U+vD
WD459+2YQV0sWnN1J1EounH4C2i07rxzEDJLnwuTI+e0R0Hr9mPXTHMZyCEx2LTG
4XhH25HFJiyWnNHqXEpl3OWBPCXGVhz5Ht55T4pqdUKhGyyGE3eR7wWpD5NtghTB
2Mv/WAdYWvVAuoKI9fam4G+BcR8GAokeTMT5W67HKeO2JgzOT3hsRehlKvY+eqM9
miPB/QI7quU8rrFwQkkEgBXihezsP7V6r18NQFLMDnDmLIRbpS5F/XGCSj7njB7Y
o8X9wD0CIHGMug+dUxzOvfrXJHDZxfP4GFMrU9FlMjyXwkebZYFK3GCB8AnMvcPJ
tJHfBjYFF8zrAMG25VkMRbY/XG5dy4fuWp9J6XIxprfVIoo80ttI3Olz+pQw3fZu
tVZwVjit+bRS1agJ3f0CxDcGJIltlh2QLT5yqRVHAZpsFnHjK6+Rr0f900twYalK
wNcwqx5iuuvZYOkgGtCDYHFBRFxCQTz1g8t6A/lqP3u6puMiSXbIyZpERISGR+LT
hw/c8jnS6a3mlyGFcWfLw4zCLuGKxFo6iLZVXw+Qb1WUJiR2F5ZnRjdCpVVsFnOm
z3tX64R2DSF9XRWLH4NqPfLtUTB3tYhZNBMk/W2lWcQQZUrbuCjXDM9dImv7cO4j
OhrrU3zmKB/tcjWxmA/SBO/DWBYgiZAt7MUnD/g/EzV8Qd6EzqXfpJgRVdiNKcx9
vnZfJwOfJmLeKm/N7xXhAl9zwSgQT0SRmoHr73GaOnZr6HxLvcd1oZ9KAhqywaGa
z8ZisP8BCCkpfx7rxyy486no3oCy6qhHMkuZWLjPWKQar3I3htpwGg9DC5zK8d84
gy8dSW4EQLJ0krvSTfuq1qk97Kz/bRwdnJfTaR/q6uRSSD9TsciOXXDaGG5HWvnT
M5CA7lAhhzD+nRsMgLqAX2Yduyh+7k4UOqiF48EGpW15Cmpb/TAZk4NFYpNsoC47
bTugWYKw2XDt5UqXe9kUPUkBxF1oOty3XNpcGlmdd2x/wtuiT3+vvAjPqQkSFBuh
fAHvEZTlqSu4r3X3JtS8e0h3CzQNcKawCIUJvCyejX5yxiW5ukRCuEmohK60J32Q
ywd+2xAlhQnENH5zYzpG9nOt8ekHGOB8s7KyZshO4fy9zGygH63cWO+dz05KHrmB
lgy2yyd+nHUdbbQESPMaDIbCftJGZfDsaXscnLbv5Dp/uF96GirrBvg1l7eOKlP3
U6VQ/w7JfWox4khJCxum+Yeb57L0bapkHlwPhh2hSIrMyem87uT0Tk6MEQLtvf4L
qQgc/9XrlGx5NSw14QgOQf6sa2XQ3KZKbncFWqGu8PJrvxz6ouppl5Wcm1xs5DBq
jWIvnao2K5Blh2vbd4ZFJe6a2b8PgHaJ2uM+EBENX4+4CUUHyyKJtwMyjxtbmKBs
2R/MD65z+uYKu55DIb/2Tb1BgNc8mj/WwtoZ0Oz3QGy5nxSKPMVEZ4ZkTBSApqMk
pV3z4ZP65VtHLnLTvQ0HsMzr2ofWSvgiA3urvMHNfbAWv8kqxxcWqIYGjYEpgWU/
eoxzHavQuRRayiND+LIaN6M3xFWfnOjTkupYahasmb3NVtppxAwWHGNqA5+XsHio
ykjqf1D6uu4d9BcPPxa9nzLrT2PftESc4X+ofKQsDVjvzeorinc7uEkxH46R7MRq
Ks+nA8kcvF0CvZ+JsZ2lTfXelbMbwex3BFPYf4QcvYuZDDtkt55h0toOs5UYSX60
ka5BJ/NMmspiMh6CQDMZimyQpb/gYpVPFPD5vEbjI/QTrnMUFukr3r7zNJHsI37G
/o1pfjq/ylsK4jN/icxZtv8Nv38Jq44ERragDOMchZAC5f5qzpS2MXVUGVO8LLFK
ZsEhKhbvirwXzBHtfgJ3bySqeyOwtgMK5ILETLwu9aYRAM3ZwSRlC4P8QYJmuM4Q
J3W7bXbVd8lUfklGB77d/VzJCj1eZKJJtZ0/a910lKad8xnUJ0UhzncwNtYzH8ks
iz+JtNFwKG08rcAg+7r6LztXUBdRuT0ElwjfvJea+TovJn7cRPvrDmWjU+wQWF7G
OhsJ3fjFAuQSLJXvN/deV0V/nlgX0FKV7AtUR0fsgNWVAKWeo8i3xVv7pRWPaPAP
osblkePsUDrc/mZ4qaxUyM0oxqIsJJjcOLXtYLhCq+g+RpBaRWoF6hMK4zH7ViLD
BF6972RIrz3Q6RSckDXaDjcyCnWKm+4/iMgBNfUhKrsSLEyLkyfc/YaQZ9Gie2OJ
dEs8hDO0oCRL9r9pbUdVIDaKRxO10Zk1jLARty49LcYGmZSoWwW3TfoCANgFLlM7
3nBXOWzIA+4KfJCvftHcALUfxMyjcIPopDSTxrNew0Jl8V3ZFWlplbfwT9VD/vqn
hLFH+Pkz5u5fxHT2UvLGOJP77TowVLmk9IZ/7y2OuVhRuoMzBPkBbs+N4bX7m8lt
U7fy7LUzX1w2NE0qtvkeIbo8lgDxl4dhmlWWG4s0fxwuMLvw3Aqo6GYYcd+Yu74I
2nBJmqhz0S9ExTMBb61BbuL8sBwKobt6yRVxn4U83SJTBP3D3ndaWujBrE7QZ9/Q
3V5hucfNaLdLasqHDbC1JCcvqLJKra4PmWMti91BysgZbSOKevdQumUZMWvXX7E7
DO3v6h8q07VoDuu7bSn2gR/qbx0V7UClb6CP8pZsz/50zBjq5UE2VuO5iS9bJj5b
MpS/SZRMa9UQ78NfRMKhHViramltT4Z1ZIxeFgUuzATV1r0L7ysBKDIEo520W0/V
LgtGxRI2A6xyXo8dda8M/EMdrbEDTwgEUsX/HVdBhxK/Jl8o1mEVRCEqsCe4xVSK
uJL4VBoBg6UVcoIkujmyigvmG59Z0RGcssMgAglx2PoJvKmF96B95c+fS9eLH/Mx
h2YiFkvrF2AYbHMl1p0BXESDJUlVmv1FpB45xKgMrV3GrKU3dIMt/MehKqhjVorm
j8ZAhAj7AaBodmLVsVrGV/cumiItvifK/Dw7vkCpi2GnKavaRUdGpbCS2St04e2W
Qdi75HzYaeQ+ThpPXWeFfMQs7LWnDkERpyRt8yhs4iPPMSAO4x+/kmjnKWRUMRkT
HBkikeWPkP4a/cEh08npe+ARFk9l8r4jLUZ2MfRjNPVJszt+RJIe+wD3/JC3CKxB
iNQ6OW4tLyXiwP0h6yXm03v3aSSY/jEaO4t488zrVVVqxFl7XX7hTcFMtMfK4LZc
Fhqc54qjsXIUS8JS9+VXCFt7vUqfuagilzi5riyYEhfhqaqY77hQfkC5yn4HvZo1
KAZoyNHzm5e4Ir1d2EXCqzn+OmQVD+JY2504KZeK37kovBd0oICBJdRgeP8BIIpn
OhzRh58FYBdbzrzcz+Tx6XUHHjpFgYh+PCJIEpiyWqpZIuU3TK68aIBd6iSmafXl
refIOKdto/MZ6+7pYgXsvE3xsnmq6P94GmywV50+I1Y6JbZS5QX5ZUX4y6SugBVr
fXr8NxNx9MB0Xh2/TFtFOZzw+6JztRjAsk44XYE0gbQ+BV1UXVdUsT84yDK+Iy93
UE3lKBI52A+ZOGwkJeGVlKz/9tIdR5I9Bg5oHDqMKQQshAm0ubt+Y510fpyTlevX
d4DYBPaDx4YszRNunIeQJE1YTo+4UUCpg2tsADiQZlgBpyplPHjBSn51aiXTr3WC
oOsad4yv/nsnwCMbU2fzeYIu7iIKO06vj4VX5m42xtNs9/VqC1nNmN9JmGFgtQ0a
/9aS3Yz9SAMp6wo3vsMF7kuE7V60cVmSjEoG3cKUzgCZgM7YdhQvkDuObV3/gysZ
MdYCf94PgvnzrjOJ9zLECvkhej4EcBaOhB05E3D8XKxbmaKjoJ/gJ69MOzZ7dJwp
cWy19qtPUNBOcSmzWo3tXUvfxnmzXSkrfQJ1tTOEvRo7eUw+c8UXKaoPoHxMlSa/
Ai1r2juon/ODYl86Og3yAXto3gjMaDcjTMsRoj2pmeDhXqzscBb3tP7vsG0WYLIE
YO/zz6/DMFAyA+j/CuhuWhW4XuGec2jvJ8k5iM8KRRJ2PUFAMNwSsoMvS25ZqgsL
eR1HxNDXpiHHDcTL9KEXb2q182b2zECRhQpS17hEI/yPrXsvwvn73yM5Fbb7/n2y
e4Q+wlyhDtB4XVuW7/EFRGjMsfoifpqwPhgIZ6zt7db/JX9DhJ17h9wTtmLzxG5X
7vRtBD+Fxd5wGB4tnJREZ/vZ7Dsa7fnrpHx/Cm9m95ZDHeU5wj10+yREwi4cHJ7+
DYQW9OXvmkTl8CysF3Dr6OoSnZsWpzc/CwFMVo0XXlZiuy8RiPZXtuIWkT5k0Zza
XtONt40U6+ME0F5RX9VEYX13yE/qlKDASIr7k3oM/6Yf0RAulI2aLzuAFLXkuHU+
qClgbFtH4Y149pZ9nTRv1zNYWi+WInKuXM+7fDw+PWc0iAGAGYAmnlxsmBl9pbYd
Z6qMSG39mNdE/6wFmRZ872QFqXUyEDaFA2YoAsgnAIWVp/AhJi9Vh7G451sEhh7a
a4XlT9JT9mFReejKiJ9maY0nk8lps+xns6vT2oX9dzvWg7pf1GCARJ06hv807gf9
rftWzAGBXAPWKnA6plR21vmPfA4RrROZUzD9j8fe6XFDV2SNd91U1w4cz+06BEbE
4VOiADBhQ3igdFVvdZD2YBysQlY+118bsKv5jvItBUGQmVPH5gqceZPpIjuwxE5g
d0GSQUUiz8GkO/6wmkuBBIeuutsvB3pD0AgdBaYZPp3tnpORcexd/A0M8cxmktTb
icy7UEQw+HGbv+JG0HXZYtTaF0JAun15KCQkmwGWNMiICPQBMkXZXHobdcheWp5L
WtvU3snZckiUX47JYKvbhY0UL5/gDwbHpeNekxN9rJUu1aLVNV8c5GmCDDVcRf7L
89wZ+LQ//Agqk+8k7VhJVwjpYfmbjrWnHztLJn8VwVLaUO3BJ1ZDvNXN3RqvJvcx
BsnNKowr6Miqn4A+P+8YJaq6ClJKVWkELk7xOQ0O1OUsQW87YCfn4oUS/eqJY5cM
3OMxNG4uLwsKkEIL9Wp77P3E4g7hJaxpoPjeWO9t6XkgJoDwpMdx5n6Cc02Manys
PF/cHoZLWwEvO1KoQn6OWgEwcIDrzn2I8tasjgCb08x0u5eZvN7LAeojFJ7NFu5J
GaafMlzfaMlFntA94JcWn3UN1JRX8OGkQJHKIFuEr7KRNOSxREJ1OlJy8mWFaaeb
ErRUwNWuyCyGmwnRjkcG6xMGOP6Hzj1TBKXV0MYvGp8uqhFRDBUZb+S/IaTdZXky
Ry6rVjERsuL3aZ4McoSa0NI4MKiknur0wMzCPaztNv0QZwEP6geGhm9T19AtQ8OW
I8LtO4/aLM34oQgjBpU9rsPMoi0+KFKeYAzl9KoFFCn/nI3ikK2L29oKpGCKzt1+
gh8bifvZBO/EMu0XRZgcXskQtxzg/+VS5paeywn5mjQNCIDKx6UaBDYDgKrOwd3a
Jtnu1bQ98JKCSL4r5fkgXAFav30T4YV/u6fpWaDQTrhUF/g7PlFGQ6pmJm6tBtzb
XMXVeFdMpQ6+pLyqivBair4i6UKn8IgRuu+MdOUVV3I2kuX3zAUIrdouI/42xLKS
WCgwnHYc3js9c+5d61LcQaDKuek0xOMoInBHEQdlYKHwpjTx2Q7sSJXIWoAwpX9g
Y5nKtTlACnRmzOK+hBYEVasyZA8YWe+82LS/Ap4vfxcUiy6vZPRzjy+14xeIjj6V
s1xGZpwy7HTRNSvjGWiEa1iLzr7pOcF+c7sGJtakVP/0Iv2Z5CHOxf+yKLsyKYAA
LByuwfv+ofi/ZhhHHBxD7CMoCAhYr3PXV0FWm4nqpozm7moVb+QHixBqehIhHnd8
X1egbta8l/0OP+R2H12JtEf9wQrC2QphHON59j1rra0BIyLsBKUj5Z2Odw1rPbKC
uj1n5U9OOuvs2RgrJ1GibWcvxfV/OQCNSiddNNtUUxin3gu1t1kNX6EOCtKV3SWQ
9rgAHCPGV3oW7Uv5IFt5P20xr2+ldNSJ0/rWpOgBVPXAWMyMtz+piwmXyPMTJ4P3
3J+VKXIJcbHxxadeD+hXIn8T95IvWs5mgPWD7tLhoSPEY5tI1/Z6JpHtTLvBeJdy
YBAXpSNpgQFh1DewrwdgRMBNqC3GwtBNu3Tp8/JfZtudDoq30MfryxOE6ms3eP+j
omlEM369xU2Gg7D/72cXiU2tpQECwvJngzOPSjY9zYnVkpfVtLQoLm/ZZo6ciO3l
8SZrrNbxYUxbGA8Tu8XHsNnk7wp7FA/KMuqFjDsKYcqk6udRo4NnTbHm8FaWvJ6A
RqbFhtipUD+FzEgn2fRdWidcXTN0gUdItcJn0qLpCSNezkHQJqRZbWXZ3+RLEu4v
mX/BSzbcAKM3AblPvM9HCkTPFdNPsrWLmXhJv122SzuzcxpxwP+BUd35s3zmXif9
vQqRf8NYrJT0HVG5+fqeAs/P4x04dwmORlYjxMseq6U2cbNQHJ7Q8TZ7jyblcZgP
2rs2gR3ZQsSDobcUUPbT0sa5JjVeeeNgAKtOYZb5WqqFlUijfCFowMyU50C5PnaL
4Akuk/Is/sWsXBqQJOthqC+kQ9HkXDi4vFI2Hw0pMZb0GrETlFXf52b1/deskGHJ
5TsIqPGtfDEfbJYXUMd0IQVvbYNyX2q9ZcihHGRalHW4tRQYYKWZhJ3A9YSIT+4J
5JHhtfugF7V3ReHopNyfYCJmdK9IFRa8SptlG2L3ezXAsoriEpxUjCDz64hxl2Mx
nYLqbMqilyr3r2OjKumfAp0J+mIy/Ul6uMYwL63WSEUj+uORAKybL4BeVf3llDS2
71js786opWdihKbLeWVPTgBC5MZyj3HFQI+9Cwa2lDMPli/eyOWe8sjWL6V8FP7y
8Py+UngPY8QJrYr5ikjlib+xHlTKtJj04Xc9MU0FR5FQZF9v8rQw3SqfwO6KXw/p
ewFgx9P5kzY53P9/C13Cgc/sTvSyzBqM/CszG0yyEsdCWURLfeyu56eJO4LdLBaj
qvoqhJh7E+ftN3vPdg7Q+we4xKxmGksob2EOpDAdPrw6tq7/OQ5tP/LkWgj5tvWJ
9doiu9sdklTgzcPSzX3M57EMPf2TwkQ8UCXeqx5d6i+MD0A2NDRr2ZUHCEXClUzh
Fs9eKcse/oc10U2K9OYtfV2Ka441iVaYv2Izj0q9ZqayseP8hoJyLXu2oDquvVe1
cpAa18+ktMMULsB1eeNnbRClPUN4VccnHapYevNJKdKPggpum/Hsk+5b96m43G+7
yiWai+6NmrUNt8io7Zm9HuJNuCWJXP4srW7xx9Rqn+VfYSN6g+wUqY+9wKtbkzCV
R6kaDBg6JR/j2e+YY1qVU2BUGJGwQw7tlWgh7tGNm58pJkngpo3z8dTYyxoh8QGn
U3Dr03knPUXNml8cs/s66iLF/9UoAZcTi2PsrS8VbwoF/5v5TVO6c88Hc0WClyHK
N+/tFxCoLU79Lr0M88OpQq2/JHYXax4Q1V4d3tvbdEMZTvB184bucidJnONOZ5R5
27G40P4uw2tA190Hiy9mQ0BCPbhyWA2xAwRsSXndaej6mePdPRzUyLfkM8foQuPt
t4RbitPSQ9v/oK3p58hR1zuyr2gh3Z9/rEW7JP8IMfAw2DYNY6nChs7Ax3of0TUc
ais2HhAuannehvmYzfHGy8+BkG9LeCgd7J9qt+Y3RG9HexI7mii3gxTYR57G6rvH
/1bJ70dpyHLLqYaF4lLA3OEWW5+z1ZnT45+JV6BcQqov/mrMGO4Ip7Np2j8SSlcw
QxDYaieywWeIGL2cjA/CbJFCfsc7GbeFkKFortRQiDJ+J5sDd+FJ0m2DINbC+4CS
LVLE3z/6Ru3Ov4y7Cb0Y1RMRDjjiursIHu9vwt46MN6+e/YgvwyZNqWWQgRP3U68
az3etzsXw16BzgczqeTpD27Ut8o5dVdKSP4CDR17bIYkYpTem88rTtpn9zzaOtFv
R16+2wP6CNKwfOi5+W/0XH2JWavgDlxMdiZC4yN6bijTAa/YvfO1YKjTT/r/NY+A
CpJW8d4opxi9m1qU6HNJAvHsWp9lggSSaosmhQ2U0+vksnYjj2OJ5da+wF4f10zh
HZk81zgDZQE8oTk+CG5fflh4tdbz7T8KQEC+CxVU6Jp1DBdmZZRaxVnrHJn71wEp
ec2+0cLFlmtiOR8ayN4kMLru+mWtiaDFCBAfNTGwFZx5DCqnZoay4b5A97lFi4Wa
g/T7GgwpE62OnnOC4ER+3xL5V70xkb+fp2ATkY2LAsrqf05yyyAvb1lLt65WK3nm
wko+kl/V7O7iGFlkDtOy7Q2cnCKbN4qWewfHoeva+t2yXGVP5QRfbOQW6AlPUTy4
zztfejOD3t/fyMn5vSyOEzqhNcxUs+TB/FVtUl+J/vioR+raF2N95K1jfdG0ekWo
Y9qBLpvPC0WDshXo5qyqRdoOW/ScraNRKRGbXJX4SnxMdLPbLbziTG1d7tUKrtPj
wO41z7OJ7CXmKZ+//i1JGS7yGuFFN8bcYMmXdbhbM77ip0MXMkbLFEMZkvIcQqUN
I+c6GFkZNXFK1giL8634JX0B+9TzAAqc4IA5y9yEy041oMQsRjSmlaPag7P0yWYN
JsoMZtn41shUIMjNY1I/WFpveltrHPlnFYNZ3OUrLD+3C8g0CdzVjGpiMFu/aJtu
JC3d7ZnUYjG43v8DfnYu2nWn0St7SSoa508Nd+VXzdt+S+2elZMKmI0JmYsayxGN
hDU8MZIPqZkWRhpxYn0ZodNzVB0sYmDaM88kIjSq+kEFS2Ex5HWSOP1pdDEAq1JF
jdU5EuB/wW8jcTEbHLHRiFn8HJP5l6jwut7XHWaB3WmEhLDRZUMRCS7w4cYcCEvB
HEdkpRpRroMfkIFaq5KHNFjEWUBNdb96hYrED4OyMRjUFLTzEGXFlbrUNmejDS8M
Jqm+cDBLxVbg+mQFfPYvm0Pq8EzVrFlhbdABFq1f9zG+HDkp/ppRA06yzbHCDN4n
ogV52MIat6MgC/c9zdLv2U2NIN5BsiUSfXGOk26tPDvWAisSt24b7eAkYz75fmiQ
ZU/sQVy5pr5E19TXzlHafXRnDH88A1ieZRD43U7AouQsuwjhcvLsVpmJDRYl6Mza
KC3yjRUgfxg0OCyhbg3katTa05cQWSolIU9JIPfeNOBbPcdz5ZZFi7DbjdK2v8hP
IooO5PzGyDS2jWQRxlPAgE2QNXPjEqLe0P1P0eTKtIPPrJ8wxrv+oGWY3Ul/1ODN
MAcGF7oft/R9XybLs8FgLbcuBth7Wb8gPic3cKwH811a5RnbTT8GSyHnb8e99yFu
1zhIjc4QRt4FPfAD+4wNyiImKQCwgCNHRPR8VpPAlx8jT7uQ2YRMZHHDiIku69fv
zOTOyfI4kgYMiG39+a4iYKJa+q8e8ncw2G0k+YXhT4VEqEE/MaGiT3r33HOtTOvo
H5c6sWh3vlAHGyPoQOHSV4aIFFiuvqc5yB+fEBkjs3qzsy4TqdFuuimshb5AYnAI
eXv2cntG85S8rHNXnBcEGttePCiDrqUlnGMZ5eHHWAGAU55KiQc6KSNWo7KK2JQk
EKLazayA9Z4cEtAuCP3M8p5BqKIYGAu/UIX61EJid71fkficoNw7v41fKRjNjBvm
Oz0AkYlUYF0AQZn1n8lEGSW/6S+EA6XA9veXNf1tm99vFrz3gsx4XqGr6Pp/Ffp2
zNGRR6POUClcdVcZBgUBpPY5Hn/wX5LAca6P0JS6e1Wfgwg1/7Jz6EmETVd1HRoB
jFKL7ctODp35XOC+g+2aRml/gWW7t9til6jzwtQ0DH7JhZkdxUuMQ/LVeRVLoG5Z
JBcFhJBW+l4WwadOFgp9HaKN4u3mOm5ang5xpIMAsS6st6SoSjACDtcllENCDxFP
xL+hTNPf7/0yMNNwpylG+QSI5BUp0yPg6YNf1qEmKexUCbotqIG84Ou0O3ZZIukZ
Np62xdk5cxrnnh6iamJbxPCEMCm2lVM/6mkasKcAjiRBqGl7isjxH5sUIR9TQu6G
rQTIX2YXsw0+mjk+p6Hy4NRHNDVp5UBTIDCPliv0ttS8OrENT0x9jkme2zS0EIBp
d2zycxiL1JdVSApPP4+/Qi14Vx7OwMSyFb6Ho7Jw0vaP7ZXwZDsMPSGVh6ZihXjw
FEIBq3Dss9N2bOxyJeZtvYadK3vUOH5EDjVrExWB6bRpr/RuHyvxhzlwNlXxUDoK
mWmnQ5KSW47rfIsHiTyuRSUDChsGsOc/l3txnNyqAMSr29UTOywz1QE7wXxBukdA
Pd4Vjwv7scyOzSJREC3REBJPswd68J3iz+L2du1jLNkh4yZi9LbXrBgvO93GezmB
sx13/HocEhbzA4bLi2dxAFpoaWeByMXZZZmjYLweETzPigJ3OYY/b/XGN6+kaRWG
eueKTo5qTDhp7U9QtLhPHwsNlg4B/CZ7TTEr1qcGJR38GRmv7Doq6HsNREAUQoLm
n7FBAuXgAvv2S92y9YxRm1jjF4nn45+1ZgcTPkjNt+7cos6cjDFEnM3Io41uNwTO
gNyu7q3r2aB5wg87aWf1YHNeMf/IqEIVUnrs5O/U1uNE72cmmb3MuSlR+QqRHHPH
xO/YZPvMljicGHAxRZyRoi09nCY9p8ieWKtKygFuGcZ6pK/Kh4IexejlJBe01ICC
zhN3Yw/8CTjKHQwxOcxZhF+02jKVF9j8vAGBovZ64yrRoVZx4xW2yfoZGixoTvVK
I/6/fs8QREfrCkK0XYTjtBrbWWRdP6FV9CA7HLyN4BEoXFjdpGgVmOSoE4Wf4O2z
TQCVttVdgk2GMzRaNjUR2Vg4RkWNGWaFS/bU8Ln3M+dgELKMUzi/U/9FWWVcYZgc
iJteiEabFuPytd8Z93UQdbG00bK4BqpZ7qC1nKRvTv3SoQ+urs58xDkBkS/TRoPJ
gM0Tliuuq70P3iuSSmty2hbat+GSHGgcYtyMbNDdM8Z2sVnwFaBFQteKkVYl71fL
UXrx7+zRfODDXkzj4itF60Ir38PIz7KkOY3V3W2AObFYyLw6NSf0b+6EfdRtMUOH
+S3goaWoA70AWasF8xOvjqS5njJ+uIsBYfEsmzmBkqVAoAjoRAMvSxnZ2F0BlVvU
vDQN47JhRTzgjsA7r8uEJKRdGNwIOU4IoHKXwWd56ek67T+oFE+gNiwc9YMwBi+o
FjMXt+AAps5sZgfC5wMLDVnMk1b79P1rVi061RGVTVbGCCtMQQb6CqeqJgMHDq6q
o9JcTEfkHv3SEoEKpFgkir2IFZQIjUSimfbvRxQsk8i2B7RWpEHI1rbsavtNH1XI
fa+AGuenVvSApxkfRedYqM9KSvNCFFA5ryDwdWRdzLNq49flDuc6jGIE6kP7RtJU
Vx6uBumbeR4cdot6AB+LtJ/R/b1otSUHJw2nyDy68sbNlbDw49crANtYG98RfQra
kCySXf+SLagmqYb9F62YpNPAexzwHAm55mmAzfAmsxcjPfXAJ0yB8MRsriiSwgFw
ytwJF0MvV7083aE0WQ9YBUOOrYBNDn0/CFv0/nsxRdfhu58SMqo3YqGC0LbHsE1U
jMoGCI2cyHPEKQh5B9hO2+PGwgQcd3Ti5vxYcZ/XtSpC4AVaoQ/hBMfmhWN/ySPz
eXBy6YEC1ajd2LLPtYKrW9HaaiyVNjf2O2KX8q3xuJ/L02thXCC8QGpak/90pNiG
jlMtWsK/NUzmgOXlYZM1/usGNeGNLKTA809QhG6oi2WgTJfeHaPSd31i3zck8oVr
u4d4IJvIESXbXXAyCM6+B/NnV52Rmh7BWA18Ir8JWFa+O9M6qhLduAGmfPXs3RiV
rmhRa5Y+jk5+ujB4E7LhwX/qIHC1La6EBN7etwQvHXP2J4/a44c14mGCIcm9YEb+
6OpMyJ92+Uq4siSkOG5pEG+ZLnsaAg+G87KHKN1wO0uNbRH99ueTVZj4H6GsgRuj
4Qjk23NkFkTJNlQ0HpUEceQl3BcgzMu0fi8Ww/gFjWbw+qJ3j4cQp6b/DJHu0oMh
nJ+LAsT8zednulELqo03KKM4sCXtjXow96BdYiHsct5pkT7zK64DRPBR5J2pDF+q
abE0kF7uSwosc2jLeMoyCob4+5OlFIYVOT/ucg8Ds022IFTgVC6cnkzCOD0f2ZXt
fH8rYHcbcDfrCDGVX8y/t2/6g4CxkudF5X5A6i/mHpo3TANz/bmMbAkwgQpl0jSf
NMhd4dpNj88+2Z4HXUoZdoHxVp8tCgOXEII5usw1Eu2AKdDNhTK5sG0Q33txAZiJ
RQeag2vLzFu8BtXQa8Z6qbmp99iF2QGbBMFGJAsGMgL9LjKVVi7vVllb+qq3hfiI
4Ac4y8gkdqYMuxZX71tI2iM9qa04ufTiaHN21PpQFNaVfSWqDs0itc2tQG+reXqa
wW9upWLVlHc9BLIsm9pM6G+ecm29w3N77P9pGpS19VUV5s+VFuiM45U+7tKsFc6Y
VRHWWkJYEqqDd7lyOiF4EJjhvrTAWR/wp5pyDzUOXMgtxQmpEASuaMoixP0uPZ5y
RA1HIPUs9Sx60iTywLeprflU2Qd4Xea7nD0zTkqxqnRh5WFslw1PqgSkIqNZl4eV
Gf1XU4bxIb44nKI8GZpiqzv4BI9ecJNdpq+A+o/asao6LkwsWiAEZgiZcqWoEk+J
7LQUTgaKOyDERulAbKjoEgCngGsrJNUrLquzhC+OxRxCgFIkChofyFvq+/I5GMiP
N6XtQFhl1BEEQPYuQaYi9XHCJxWkiLiL+f7QrlzeFREAX86v5HUpDzNro44prISW
3Lu3orXKTOnW2CCxZC7D2FbuXIZGZAVLahEmKsE76OOZtlp1rfW/nY1cp3xshKwv
IESJzBfVoYjp4vnqOEmMzVnFlYvsrNpi7zfXHpGE7cU8n9w7xKnZVTGMgr15S7Hy
++y4folVxdvcQcFnHMUBP/mB+ijM9m/K7s/gZGZKcRXWbgPwTgs2ZmVebFA5atAP
HEFHh/1JTPP4C90iYzZ5OtAxnA7uidLxC1eXewuzK9kErlicurViounVYTMKMdsJ
zmGE3cqY6XPKIpRPyQrQhZcsF8hmkZ6LJek39RYAAUTBycy3/+pK9gOUAglwoGS8
lvg61LiApyjL88SdhGtAcjR+9xh7NbJmxZjZs65oS5LQkQS0Ro+II5mD90JUwOKl
lQsoKNQaWQfiBQzuViCKPUDwXWMvfP5puzfTxprG1DXGish45dUY8C2ui0vs8ax1
dwl+IpLGZcJ99XQq0YyUipQScv/hJ91ynj+loNckrZheYCKx48v5JIum2ytv64ZL
KaxvFx5gwwh1vj2Am7P5itMVuyJr4NIdsWZEwPfFO3OT6q+xb/hzExF9miFDLact
F+iV5vIEpo+u05CbJdHI/ecCDu376LLEpFo3iTqLDIDE3Vf37IT8M1yK71Pmih5Y
M7DH8v9OCVQZRkUHXHKaRNEqhaRLsg2q4BZXosBDPANOnsMyjDzmJFwFPQ9WoNj8
bPDJJ4wpqGXyu1MzLmtvlsnD1K8fFtMVCSr4hLOLjNXq2toW2m98OPbEEeExo+WB
xcfGufawppSNgwN0U93ENG7xGb7uxeT3hC+yh9PT7XfbexDhpEbfub1r4gV1IdHS
Av/IL+MNOK8HX1gy7C3jD4WJlruXkjQUnDjMOqqSyaVIgwld3S/Pa2L6gglup2Ab
AvHPuSIc0+oMSFH3i22Hz4QmWPo4KNDaRDRYkgFAuApj33kE/FOJb8XWKXYGEMjJ
eiXJedS1y+pTG0n71sJp7Hy3sHKxxgx+gyCfsELjj11uNfbaCg+3jquBZoWVJKFX
doUxyJE/mE4r1EzSpJaoDOcp/9FZQXqBS+hrQqUX6fvCGdFN3kxv8hctVFqwCAbo
eyddhr0MOESVvdug/q42MC9KS6BJcGgfMHJC2IIXwR0quODCN3eDRrRWo9LJobcj
H/06+05/3BazpKPfjB7OKWFGDDyoLOp2aDxXos/9PNDRBt+OoPlQJHtzRSHrsh+M
xnlu8Rkcdhi4nJLY8YvQpc+Cuk57VyGjyqORuFY0R+P2mC1CcdaLsidyjQic/lmI
dbHFMqT/U7Ep7gFvywtGTuz78foxS/IVai3YjqQYMcWMZViLj1hW4eUobS6jO4pJ
P3z2OsXAfw52uVgsbZJ8cl0C/076r2as2v6rZLDbFDYmdkf0h1egt1RgQKYgk0Qa
WgPMpTHN5thY6vNhGekMzRhxL83eALueEqPAt7kkouLeGCQUN1WY4mgGSGkEabB+
PPtmjCSl9ckLN3tj4wk1p9D/UhH/OnZl4KcMQiPwJHFTfR+Ln5diohON0sGwX1GA
chq2KDHL2fibZ6vYFG67hrXi4HkxjCjZ8FUmn3p5npvsE9AXZiXmMNk/fCLVaN2I
9Gh7k3IICfmc9BtZ119SiBCKFpnpMT9TE3jLzHk+J2VJ5a57vuKTUVdCK4NS0NFH
+/JgPsnudzbmbnnVux2uHqzcaikS/pTa6MRm0FZpFbKu9qHvMDIDua5mKbIHoYHI
A8sXcTz/yVMdXJm2XtvXEsMu6SemBYe568Ko8cZv0R9rXeMOepAs8Q1KNqGFDFPq
JdX4aq1MU9UrReJQ+RRGq8X4nrSENwnXL9VggT+mQINJ0hv6lM4hrrlYcYvKTZOG
XSyUxPbXOoFhkuAzApGvnvSVGJt+RSkUzbG2TomLdoPx4xOKp1l1QhriVMxm1XaX
MiWebtBSFERUXff3W4Obisb7OBWfMRwk5mExxnzk8HqqxvS+RBk7sfJJdms3Zs0R
dozbpXpopjUK+9p141Ktykn6yEiOpeNTlb2vMO5/it2Qo/IZnuYODCN/vPI1QX9j
UhORkIG1Gu6BlHqw5TpcyzZRfsluvRGrkL6ufw0PYgXkdvNnk7uqxSDGzo3LhcuC
Dprbq9b9YM4G2WISmXgg5hSyLJ1jmUe42sgJNvukcUs9+mB2qUFOZpBvA8Yv+1rE
nBZd4u1BEvA9t58VFyDytfbHv2uxfx3/X4hdPJpOkg1w7MJrdB2TkEYRs6rnXLjb
nZQamRinBXVsn/sNMJ6oiix5fY8f5s4D3Zfgfl7wQnkVA8DYqxViHYpd5dszLSbo
CTLsks0AvWQO2on/GnymAmZH9/v+uMB2qFUDhfGfxhrpMxxUip9HQfo9BTQw/Jcx
lYBsRqe0t/rMrcq3GihkrRxhZ2pmMBZkYHe1DORZO2OPWU0zK0gsAuugRoAl4Iup
FKaPZaHMSzGQTsYsKGUM0CAMXMeO6l2n3gVvxYpfhnCLwAkry0hG/U+AE2eUBAgv
/dxHxTifFRYEghc0SWrfdD/I/qEyJJw/ReM6TLbcgdyLOdKGLk7ddscIKjVlVa1j
CQNvQU/4l0UCWNeD5KxJ4t83OWvEowdVxJ7BqU8EoBgFBqswdL5x1thedg294ALl
lxxnr2hQkjn+Q9qeTHZarO8XHCpH2KpnraY1MSbr/Y3UcmbMrDdbuN8lhnMI9223
pbkS9IU6FTUcEevi86NGbrvLPDrZGqSIfiu78BnkfKUKdreutfe72azht63v9fMZ
8vgTwwduRVsyTc3tkzQAUO/j6hb2eYi9hHYYXJWkd5K+j0AK/TUpQZRnMmXs991W
TmfEQPTWIafiDADosJBrTnRuWgB+3grF0sYxQGM15Zi9lwwjUE3DOkUOQBPgsxw2
rmO+9LCkoomIulWJfwG0ckRyWko8QvZeoH6HBMbKiMSic9QKOQGl1IzniR1zttO2
XmYenY4RaoGwXoD8zHyDHwW6/ovcQhW9H9APu1tyaYg6GvHHtsd4acvepskDxeP7
F7ppYkjhGxHpaFt+mTUT65IcdcUBcixXJ13rs8f0qRffkn3LO20TfZf5xtuOVxXV
4v0khsuN+UDrPUPwTreTpmHtFOu6l8pGBM5TRNhbp/DOVd+PHHaU7oTENA7owJ0+
12LSJnrSy9z8GWto9Jfp5rSrPx5P4rQ3aenLhUEhRYICswxLjtnM0kSMnhAZZItk
e5wcXnc+LbH36Z8L7R1sIsL40Ctff9UQcIR/RGw09sm6kp4gCSa/bKms2AQN+fW5
l+l5oBrPocz4qIMxeThNohx6j1oMePl5A5n73mK+Owxh47aGN5sE9zlsp28OZvEn
tBUTOykmR/nLYZOjaQ6gGF0BA19i22JtzUrt3jAoSd9y6BuxuUQy3rt3iqWCqPR5
LspxvFiEQmqhfYFq+6V09i1ZWlM/gGd8HYSA3rJh1yzGA5S5pmhuIDc0r3qmOYrq
FnbbXtpiQpN6AY2dlK7oZj9jkffSbmch3zLzgsSf6COyV33U2YAKDyjZvb9Pr7vH
eo2rCewYXtXS1couolJuHdpH16Hw7GpGB2ACdFZdbJ9ca5YS1zGtzR1k4T2YaQzl
Ddw2LiZmfojYzfq5iC44Rdo0p1Ond92cU/n2j9MvSBFgVQkDZyon619xzAnsdpK5
8zk1f5rVC4ZJY0vFME+uh3MxYQXXnHa5zK9j9ZNpXjtXHAFX+q/5Nw4NZxW76+oH
rTTW8beprdaH3+7cLmk/3dLaludKF0eTy/6xHtqFeBrNjmFJ+LujZHknkcvdJDE7
vlzDKGzuFthCrO+oW+oL23kLlAUbFwj2q8aaLdxtf+k2kdccCKvbKJcaFbc4BuuA
Emxa89W/NXqLr5Uuotest8v77OxA3/nTb6yb9g9Tbba2f/rq2o57nGOKp01H5TPZ
ZfJ9Fi6lfkQgYTuSNAiEEYI6Fknw0r2jKLJt6rhYT2yQd65pbshfC7Ygq0zKg39o
NI8PTW09Ts4u3BwmKcf/m78N+AgmINtP9N79M1ME0/R7qamLorS0wu1x5+/TqKN3
Cq4pOv2E4X7ujea07mMTixmt6fyTwqd1rhS7iBpSTQDeuy+dmmPXQQ/kbMjjWy9C
p8aa1T1a/Kg7eugTiyrRrRVjSunetIesOZCUOH+yu1Zk/Blx/A7WmWbIEnYmzBx0
nRdFxMEbbc4fXzdrie+w4VreEa4/sUpproi2IuH73fXhL96UURv0NjbrVPFTSM8e
cQOT3dykevXhFxZC7aCr4KYtg+Sl85koWo5LrKKGdQd76aluIFztVPVHRP89+ebd
x+tCYQieCxxcsHAurIysBYBLamX+aus070dTacEKucUxX9CpYUsghMZVcsdVLgIj
krD+xZgJCKcm9iFY7divnUnRsUh/mUyCAE9rZT8T9ciBTdS/4eWizmdVPR3PGAr6
LQanbW3p9XGzugNOW/+lCGBkNyCn4gGAzXJ7RwnNXCmB7SOlY0DsEEuFVrOz+VzQ
swYVgWoJ0AebVfrOKVwc8TzoX2KP1WKHv60thZ7oNI9d53WkdkjJBq3376CywTu7
mO97DDdf+GQxqy7ZTKRNuYw1oPf6DY+cn5rwH479joOAegLqVLcnTEob4ou5TRpD
aR+wYIQ8km0OfojewAQ0HFMwmSNUHmWCVdYRUheRk+J2N5D9vEgFhhVMDco5MPKA
eysG3/tKjAj0mcO6GRwnYH6TpWeXclECZ8LVszPOQMtpym5Qs2hsPNqVP9T3/Bfj
gMz1hs9G4ik0JBuRYfmzdo/99WerQBHNtJzDA4CUW4VA7nCFNXKt+ynZRPoj28SC
+70bKvn/EJNkT5JNnhDU513c6J9q7mzZTb/eaqC6ESbXiS2UcAD2UO+RbvdL5h9G
MugiCAVO1eZXscKUtpJpd5ZJiOqXOwTJTulD+JRz72Tdd48h/BH3/Ggfphua5iRC
AzZs8yHnbFB4l+tyZTyDbvwPDhDNRjs7XnGTiJxkdR8M8wmkJYwiUjfbS0hWOAXC
Oq8b9Qs32Ah0V0bRhOmAggyCZQjdkhp17YmIO7+mRSlDU7WJEfe01+1VUhRhUL//
ReZDU6Ic7LMB7ZwR9ZLoawmAdApMVmAMLZgVYUAkMKGgSGgQVXBvsiBk+v/yaChT
3vMIjf2j7I6pBVuqFOBwKwkAtnPoWeUPpS4SOP6ZGDCUN2Aym3qna2g/IBjmZLkh
OlHZj+oSDr5f7GTbmIc5AQuUlAmwkr8HoOnFk/xtl4rxt0Hub2Xdn7WlXjWbKJ9h
LJS77FBKZYWURLbIaYnvJ55zrzlCrS23dZo1FD41bTt0SMTYJZUKokguIfRWKiEv
phng5CJiyWySVHA0go05sRzeh79Uv8Z9JOHrnFjey98S3D4dW514tjq+54QmeAWQ
CjD2lbVd/ERa5XHSvyHAMNhjzi7znPNx59K1mO9iN+ErcBcZRfdjOz+uuGpDNgiz
SLooyDF5yEE6XioW9ArsdDSiqvO94dOCyXSwj8jprNNScx5TiDnvBj+7sFqCPs1X
d0RbajsbtRdnOOGIWg8LplxLJVdqPvRqpqM+8j7u0sJWPwP/bkSSiwCVHcKrkfSI
KZmsRu+Wu4o9GhHE8M0ajud7o2r/OeePJTtYPa8BNrntpfZcujIgbO0/smD+P6p/
yvGNwK/ciFoqIRR3A03I9qhJWPq55g+ExZLWGAIwlNJI/nOENhHxN+3WmnGIesln
7pqatPfaBCpM8SkDtdeVQX+3IbChqjGPe85OxObfuysx3VFmDoP/EB0MfUyCS1Ae
T3b6fCMwwq+d7Q0jT2nrvoOtqpHDyR/ps9i2HNsm+wf3LFogDD641s2xcVV4ef6b
DzZcLUsA4qbwRsVF0ss3F7erBGRbIX+L4p8xk7hhuIWbBXMUBmIitvD5V0krRorg
UI2mblb+m67BAO+vQEdHpr+cF41x6TI3hu5YsSaGdb38h/sRSrLZOe/fXdnGVFqC
4z2Dy9+yas44JR9iacvrmbvUSZ7PGA+4B+K6z2xnurhOhhYUS7OGB9/S6nqPrDN3
L3J9nyv+wcpR/9UKSFWVM5S2ipkgxVx/o9DRuJkAW78tAto6Aa8FQ7+deNVpbnDg
X5Eddk+q24Ti00NehAeZVSksBORZb4OryMppKVjnLPo4BIj9WkNBo8F+9U/hHw+Z
tRhQhNV4BtkK+p+dUMZyCY2E6xNrlZhqnCZ4nnj5aLk9B521xWy8XX2ghPBmPI5A
NnoTzohhE+ZQO+L3oPuJ3exi5/aZzqHk78KiOxCj2GP7dVoe6EB7ast3Zv6cPQVt
JxKERJaAJlZujzkD9jNnD20jxLHAtiqSlDPkGr+cr6nPXb4QBEM29kADrDZXC7Ig
7TRtDTK2aYFeyf5kh1XwbaFVVbFr6RW8h5ynE9o8on8apGuVq1HFs5ihvmxzvayg
V5NuY/RYH3oZ+6xyOXxFfoC5eS8Ooy+6/vjZamL+PRoM4NJVPTTIX70wUNGl1x0u
iBheFTEIo4fw2obLc0UzYl2qiW6kCFiASopRx9ZFfbC6L7oH5uqUTinoiE0VdZNr
lqgXiHvykuSB1ATr9i3rfIXwdGDCH0oAgVrsLQjHG3Us9PIdF+3yKGxFlvgBu20f
INOVhDloWy9a0tB7AXc7G0XdwbWHVuyGO62VEQ9WcAxLeRQ7ADML4Rf1nJD/ji8Q
Tek8yuCrhHQmsorTYgQF6pihSyvju6eD2vBwvMAyArQHAPRI4FfOE8hFsAeYDZMv
eGlXeorWrx3T4eBvsTlICQDBdWRtXqgCMUKlTrTlDdm+A4HmKR+gSfJlag7ugUtM
X20mRym/Dtw5zmNj5d5yQ5OpbiSVyC41xt+3bCLkVLPSRIzMCzNocaA+htierlzN
x59mNIsHemQ/p4IHGA+JkumlDHKrwukWwVfdkT/15AnlB2M6+cRYkfR+QAF20+uc
a7n3dA0RU8I0forUgW+3IwGJ2uK6AUqe1rat33jf8JOzS75RZueM/xvGla4+JzSp
nRBOsGru6OX76BRkc2qS0krUsxX/z6By0agJWfI/F3wjkm72GxzOAZj6aO1wmPzY
2fEJs4uwUXj2OCEcVOV5taT3lhXyXztVHJB0/qZ4jNf5+VQvRdQXHbvCUO4FwIYA
frU5MLjutlyD6iTdu8IKDqFJu4lqejfB5T5Y1yAL+ylUwTh1avJqyJiDyhDXS4vh
bCs6rXFdvHO2Q6Ccvzlgveohi3PoYrl5GiX3Kd1quACBphCRiVEPIhrFzuNfV9dg
QtLZztQ9sE3bhsEAzcw8FzfaIJHxGWjo0jhCkxhJWxVRRAzWc/jMo6LzHtZ8UgMW
FEGjTR8mApkiRWhdfsr34ZVyDJqxrQG4cB67C5hb7OSjeqkx9IZhN1zeCxttnSOO
DsxAL+X0834idlepBS7/PaRowNJiwmVKXzWBfdqhAIq9QVgSoKcWOmnoPy9ogwsS
CFaHWdM+2yAJsGD9KbXTQ0DIP7rRIIzyGQNBo39anXSZ8tv26jWsBCU0t5MelCAA
2O3Z/7boqmUT9l5nIL/qOA7CQaktLsW8Zf9Q479plbEuIicYns7+WWr3xiEL4Aq1
2roiNopEVCyyEguRr+g2yiSBFTUmeS5aYY/D88FbYUAJ/d/qlrscK8hZghYiw7/K
jHUnCakjD6nr2pBh/ZsWBvkQqRkY6WX5scgKiTp33OKG16Wp/HFB6MxB9OeaLatO
SMTrbXhJb5TOSKOjJSx6wV0rz698e0bNE6Sn0NzvsYmJ+AJI+Mnu93UGcAmO0Pte
t+6UhcKGIYAz52otRow6g/lvCO5yurlk6sWG7mydtngfZZStG0LQ9LjF9MhDkt+u
xTDmN7ROK9ISxJDwev4yzgEi5DaOyqMyjWlRajzSCOH8o8JY7u0wmOfdsYFAcIvZ
1j32232KVzsInaJ299/A0Cw6AEMwnkL5jPVny1jppTBbRBvpaGellX7ZZ+lYUW1z
sO5no9lZ/jjwuEn4fiYvNbscNRh+5br+LxawQgK1ltnougilpg8KDhA85BoVHLwQ
Pq0yqs2KXMfdP5pfGraJmoG/VwNbjUSuKpsacKHYZ7/OV1gHu1XB8miyxHybc3HT
Z7MyYOsfuwmURP3OscCRHP+mSUViby90WjTopzdjQdVecxGXRQZ+xUL0kNg0NmLV
VMFfbn/JT2gp+O3rHtMTt0bvOC/r+LWu0VIRoa7hJT+6B0D+h+BX/fj3cLWygRJL
FWvnzo60nBZQezV9LERiY/C1tAo3b59bSIJzdiHvK0WUKTWWI5iFj995XHxSwul9
3btomY8a8MRxSeiqu0mcKHlbpzoaJRC70BlLulCsBy0U5UTZaaejxG7ps4nQRSvh
EE+t9lMFUHpnSyrUmrKH218tVdfiGvHvPjxO1xJx+bWzwx3k51KwBD7C/B8FIueK
j/AWjz5SVOTN86l5Q8SpTRHMASjPAqdOSYu0UosxGUx56lNDy5rjeV/7RVnYkxwJ
w5UfkIRKuhr6Xg8ZHBdDvLkZ66XlTD6AZyKO6GjAJJVj+2jfZJOwfnQllh6qLpOC
ywywoKJS7TvnhZtHrYphkXEXPoo17TSRUihhidn42S0yNK4F+U2Y5YeaG1Ehg2Ps
nbbvMESOiXIiOmyhvpgsXjBntKNnwEYY9On+I40HtWcAjZpSE8BBu7EQR9LjD9R2
tHPc9TvzA2hSlz3FRbt8Kt4Elb0dHysvukGCfZGwfBOEvV/f880GIX7AdWyLyyNV
zMUCkpJ9Rr9KJ83XRtmZDxpwuPBguDpBYSw5jNNshrWgVL8myMZj/6XX+V4I31k0
FdRUFp9s864zISexl3GrqSYcb56DMj8UBfWc4rH52BrP78Ox6JXKV77vXJF7HYW+
D72Pg+flh89c9lTh1/AUzHVuNRt3sOxzKdNwDMDQl6fRaOTlVuPhfhZi6UjqD8nY
1Rn3s6U25iuEAX/PkwcuGjSsUPRhg2i1C37N27bUR/8jJ1g58y4bsCw+gw5bBWmf
0BsjmXkAx31/s7oP96KDgaUvy/lo+EV+nES27Y+2IGwT8LETD1gVlWy8Pr73ntoZ
S9n1JQYQ6U/QbGQUp51l0Nqlx3udI8DbpvFqi7IicxgMRcjgYcws3MoIAalOLv7a
CNqoS4gg4dM72otIbsTQ7JM805q9zoar1TqFWjiU5/oIhph1xOSLxRu1SxfI6d4q
ot+HKfrOroDy72Jf40En+b2LG8Hb5lHQCTMaGBdinJHiFZ4vOuJ6QXpy7dLMPyvn
sGLEGhuCS9FWRtqt6QnuZDawgVVOHy3MhPMvfnNEHMgPHB5TTG/Xx/ZYwxlDOiJu
BC+vGYJ7wJmKj+zBxjfkj0bk2A9anK9tkALJhKjZlV33JiwCoSSGVHAP15HbrRU9
XERs2bfVoLHQEgfo9iJHC1bTpokQjXZ1apBjUZiuKKb99anpTv29L9b4b5udLpmN
OENrhxjfe6tz35WF/fbV5E0hipM/ABiuFCEi0qBF5OKuSKhms5eTA01D2dMRldcN
aF59CtK3ceou6Ygot8TCmguqdUfSnudTE+Rbu08c+zsv5Dwjq+26JZngSsg7y/Vi
sZt6TExMzWIYg6eZzoUzQ7l0WkEzBSEGFJDC11zX2PbMn5o3kOV9Pd82h3NVfBcJ
YllDdYLHBw5EWvCnAV9ThTumeIPl1MC9sg0RqyUXfge3ytA0PLkuqghGD86q4+yb
VVCfgDvG3W64/s46U+hIvYvnFgyiyEt+4x7DNRZVhiVeWspIuub5lPjyMyBIvhjO
H0arBam+lmI29dA+kSk4qmQDdqdCUppzs5pTxNrPcd9Oj58UoHsgySIg4O1JyXDu
oMZPK/bAWXh5MUSoB0vxs1Xdt65S4UtjRe09WuRF6n4RnRHr3PGhYQkC7lcF2EXO
ry51M79GP+NsBdLp2kmHSJWx/iyWCOgnTY02dZXFOFsCeQmtppxTpEDfG0nSYmae
Fz4twqY/C7zY9mlltvaNa9PW97reaoTxtleodjZnr3rBARqnipK3RAjWxzhq7zkL
01GQzVj3cfLgCo7G3sRBTfWS7RTNACXM68y0eOKJZ79hB8sMi9uY76BwNPoawa5W
FlqWHaYJQUITI6pzmwyVGdKI1QonSiYbp9pup5iNTs12WONkbP+Lwg5+GhY5s8PU
JCD1l7V7O8v/2YqBnkFptNednAfKrs6SKQQD8I9KHjf/QMWBr89gjxwYvUy3ETtx
En+TbpCd1ZIfJQ/VdaRUWAsgGR2YzqAUntL6J5o9ssu4iCd3bPXV2Tlw7CXode6q
DwTF3NaiXRd69Rz5wPkp4L2swOHoiOYtFx4Bv5J59UORo8wkdvCDB7L4ux+DoLht
jrZS9XGVZ/T2VJ0gGDKDd9v+4gN215TSImx8WJ5YRGtAzGGKa7OdUpmmiBpOWh01
DR551KornKM39JFg2WAg8d2ln78XTZhxoeZIzRRhbIXZpjq9nehUWdGRWdeZsLLg
h2xwSBQ9Bu8ehmQ+FnabJLfhvMAnngOi5rNbGIw/lDojA6oiiWiOt44qtMj3puNm
AZOrRIwfTS1o3k99kXubkGzoN8LZ2rEUEvSS9nV5xiAsBHmKpfgjBbA15CgOwBC9
r+X6L7y0/VrKbTRfT1dW/dlUiuobPOsXzrZMNGh3l7xlDxNaKKL3bvz16CitpIKx
8Uq6byHKZF0QQgh2vPrKpDu2PirVhz0nIlTD5yDNBzrDv5y1L/kEHSp56w2d9hda
Yxqp8BFG6rfTGFeVtYRRW9SldEckOselcAQOeVUT/UEuRE7pWfToRWu0C9JaYbCj
nAj/l8J8TzEZcPNyAj4XsJX04Bm/d09GHZX2Vd26eqhnksNYmm7aMWLR2huypc4A
oJXUr9a1DffGI6Wj0N+EtgkeJHIgYA4olU6a3Q1EZi9YknV1jZ0HoKm8Pd9gXQd+
kpM7wwJFyvDj0o+qNYf3u98p60WHMH0eu3Mjct/nMfncqCiFZYe5mbZkd9vETmuM
cBk21AJXUL6qlGNyMeYHlcrY4Rf4ANymmmEKlQIalggmOj1qHxmYawYBjXNeVILr
LzsupEtJ+boNCfSvu7vJBTSTvnQs9hC0HG1jNzJfCYwYPnSnpQ2g7BqEm5uelMnY
r5UG8N1ol+b0Pnli1xAKfFc2pkOIteMxXBC4lKowkiqWMuSjKFQT26QYkplnXoMI
0KZCkdkukrM5R70MrbPIDo+KIIBXohcH2aAyI6eCGcYf3BQ/P9ovqX7f7kALCkvZ
pHFxJZh+czpvkMQBTLdemhaM7eAXP5igWMRaYCL9vE+O/QGYzyBoTmB8DIq8Nc3P
v7G1c5FC88KjHExa0ubROrLGrPk2y6D8gKv2rOAUg332wbd2hQxfOGUerHUenHlw
3vJNOPPvIHXZSilxJJJYfgej+Yxk6M3pN3dmnc6x9SKwrEwG0W/akP4Qqy4FdcXX
G5QfP5VKeWG2AEBTgNzx0BXc+N98Q8lBchuS2kV9dGawtkyQ9S/DgBefJ7eVtez1
CbXCSCUEnx12EvOEziQ9ULoX8UJa0CcSQkuUYLkbqMZ/+H3emyehQZ1q4J9GHAp1
noppic4+ainEnT4sk8M5foToj1Lo+8sFqWkptUbCmZ6NOMOoeyradufnfvKEG2VG
sLrfpRa0dhjPPPgkMRUMd+3IjL9rhSs1N3B915rLqDx0QabXXvMESD6jWf18SkXw
Zz+Vd7VIDw+ZLFA8kdFpz1xITlkk/n20zp/+4+Bsvppw5JbuV/TkURbu+Dl5VOvd
omTXfRckhVmVvDSSKVeU8bMIg45hXD7kd2mIHiKStlcC2qUHPFpQ5D2nhynQZ8S4
C2MwI9RAjNdF1+1zpT6JM9qd8pyU9LAOl2ZUf6OyjkN7D7+Xc1ZxprTj02GLenuu
KTFbJr8SbNACOvRya7mjjCC7d+dJybKdW16Q0xyhFIQL7b1KncZZYC4EMS3wl5ec
uI+/e28ImRORAfSwBQJq6LjkG1lrHhoNhdL3KXxyGV0IE3eXKBCAxhO6c6J0FUyg
h0HILK1XRoPEEHAVLFQhq+2avCcMZgeyDoqmrNFSPVcR/w+vPP1z3Y9NUsbjdoOb
zEPTMv/lirkh+dI/1oCO+DoQ20eVzE1lA0ErLFqgUoA3WKeD8WioorPOL0xNudLR
vKfrPDJ69cDHeSlQr+LlRGA+dIyKUQK3mBUw75y1SOkFnn4AozcQlNTuoFapurcc
+VM0crkjudw9cioKkcm64WGBk6ysmWgCwfvxRRYp3X9DSOCsg0VEin3SYXVtx467
axGZzF0UY4Jl3QUixk/+26sNFxfl/kRov1NHHova8hRLsSlKLtHX0RYSus1/y1nS
Nj8ICo08sSFczwAT36K6zp/pEHKZkm4U8jZpsyw0oJhc6OmaHHAPB/5A/2hqxw3o
s1b0bgA3ofpBvTGSO7nltIVvEcdDezzNCwG3Fcq7R7yuaBzRSnNCeE3sjiGChMVZ
i2KTr0pA11cACcGjStZ9MfdYdCN6iKgsjaPkStUOKh9DVcBtgfFxZlWSra7aVvn2
7g6qM1/IxJLaOEs6mLCmDzJJywrjmgQgcN7skVk9CA5pIQEZbaAZhPuMI1atvLhu
sZJU12Eij41sddwKEeRztOo9u4U1VuXG7gSVqry6PW2rPGKZgegITwcYvXaVwg6Y
RO31XyqJowlq5SkkkUx8dy0Lg8hFOcuQiTi7s7BDIYqYetyzcdgVbb79HUvd1z7+
fMqHN5gbsGj3/dyxIPQKvnFxYaNZVB1nb2kTrKO2/5VRwmCa5gR/9XRpaQEzU0ck
3qomYCosmMa3qzoPVyycDTpxaIh6Gb9UM2M+DgXSh+lsOyusRSkJXu3r7rWerUoI
NgZ3+GJUKcqeOaH2IpUUxG3+f4lxCxkF3uJZFpkpeG2D2l4TYG3jJn5LrEWhu62u
KyxAzzjJyx7d9vvtePzATjhJx0Hp/Ngbv/d1l4xVSJrKtOdIMfYevAHmjusBHmMH
mIWmhoQjeCFRdBAg38x4bwdyXgBNUXx/NiRIvH/ZtaaN6ub8mPDtgKqZOTqtqEdz
W8fSvZLcxYQcNIOy7LtFWTeRBg9Kcf3/dnzfTNhvg9Ylnm4rggoNSkmSo9MSpjD8
5fqvqJzOcoxRueBoRkubam3bF29IUXJw4H8r4dAuEAYxC/fyfB/qyRF8dJgGo3xa
UyjFqLYy2xm+J76bozdsUhdeBTD6iTc0U2gWEj1rjHnca0zUauQcxqTqiGQPkydX
ooRNNNZWr65zB3tOzoU2unO/40tzCKdsw3sS4+Wd1/EhscnFA45Uv7xJkMbWo4lG
SzM/WGMcAvBq4dJgFY4AGPIJQ+UIQKmQSAX0cPna3NJpYsjsnWsd+sK8X7TnDSP0
2AfptcvdivDdmU8ZRU58PK0/GIkUcR8IEaFpBzG6po3bOQg8ANr/K1tpSXrpG/8g
1vVAYMAU6alW3rIvielaXDDrxg24UUI1HildHdyvFd/5mUyrUoClgfhMKZHhITD1
kIZVKCDy9PKQJ56zba46ykSzIbJjs02FKWmXcMK13G3ZZGMzE3/yx5BXT2fjqlLD
kMKDzzAN7QxtyWtPS8gUo+JGno3+wkC+6sgnnTkzUsLhcMbeNwxaok/GJXEKfQvU
DFTI1qGm0PjEG0z2hYKDZ8WW/qZqWteHSBicy4BfN9DIR311h5DjrS6LcY9t3tMT
av6LOkIV6IMITept90GRKUxfmbh66Sn0VMDAWCYTIo5/LZ2DRgOUOtzHvoMvRAVF
DPUzIMWHqYITQwePYLEHLkTtv/NXTDYQPXPqC8auCpsXZp4htzBCs48G/1wqB2sX
JALgGePhkZgpxy0dB/ostn8U6PfUCvJPS/oFJ+2PVF+a2yj/Zdx8GHkLvaB4jy/o
5rfvSYWWy/gWx25asPyK1fafHxiQWBhPa6GVbnAcLGWcWu6W3DZ3PgsPWlU/06+p
YNQcgFHLsK1lruylreW9yVUG2VXJbudWSMnbLVLHcSwy3TtrWE6bByoIQqSnoGaG
xtnxeZRAVA5/W0smkXXRZ7fgujF23ue8++HMhQVwumoqr42Jw7017ppYnTw5mge2
0bLW6S8HGx2VKUjC0iEpB6KyarGUKBXWQmYN0mw4kqiSIeuNZJhP4uExKwElg1Es
1OX4BF8DoH5rdoK7WS+V7h7TUP0TS2d8Et455I+KOJjMraDeT2TR51KunVbnSUoX
AbKxnaHzesVnlUIIgufIQQT3kSJOc9WyptyNoJNFeNlK2OZJAoKiv4rruAnkfmqz
yCqCZFpjFklahY04McFiIkP7X+DjkwiRQ1/110/KmmCZzLoa+aYM2+FTvA5G4HIh
tcJaxfpZJEj+Y/+VmHMaumUmZbMXOnJFdlKVFvK4jhUpAQFa/ntLeI6GDlmQp6EC
3+nbbSylE5pvEaRwbJhhKGyKnnkbmnghLkDNIHmgDY3VkK4MdYFK/m91VsYrHFd/
bRnIpyZjxIWqtcQduprWm+f9MvFWH7+xbTlt7O1iRl5q+nz+o8wKGIff2FvBC+U9
CKZDuS33Ze6nNoRwJiJujbgLq5C7dhK1dchTGV5uVLSf0Y2rukLiCbyUsFqwocOA
qJGCebVeN9o5rOhDC3WTWfygVOIcRqVQEwpim8NxR1sIcIlWm86hBBZUnAqtfwcN
Bh6PEtF4Gu4fKwsXxYnZLs1R4URf7xD+aYOsrMkPHCJomtwMgG+6N2cGPUZz2ecT
Nd/f60pLs8ORP5Ir3frtVNaUSL6zpKZz8Z6V7Vp38+2LPRdcWM3N4TKyJ8P2JPMc
OdlY5YnHvXKpfbhidkedbHveB2AyNX/ZDl2CzdRWyp4T0ClXxtr1MCpFmPBh+xbD
iyMS03Hi0kd4Q7PH6MjLQWOSaA1FTolY5iLsz106LQEdTRiCDYyhOVymwYt/Vmax
FLD7UW9mYGTDyjFZaoZuuWZkc0RQszkcjbqTN2gG7tS/8J2jlGOuMITIrE6ZAldK
zb5A5Wb37GtbRmIzWdIQUtBh6jHobZQa3W1JNZCG5KUfKY7abrXgNubNz/FcHeO+
wMFT7Hw9QlmcRtYVnQQhVJzZ9RVhpSNtxIGXGAXD5xTn8qT+m0znBXTIWQbfeeBJ
+we34idah+qsZyD+ZdfqR04WRLwGRrLuaj5VeU8e9kcTV86tLd5CXhsCtsCJLhiK
j8t0h6sUjY5qYbWy2c+YNrMrrf3kUSq+lgKDb/xF0o9NXLd99+Q4sr7cgoMbpaW3
CFuJDlRF5AqaMLl5fRBC+DUKZ1n9fAYPnhOOy1Jop2y1Z5EaOr9l+jkskDtzHNNr
cp4hdmxhNSioFeUkuCdGOMEZvjt7xnC/Ad02lkJ3TqGYVgZyEeOqj8uSx+czZDOo
Nz1G/lZL0EREKQ5wxzpg1IVbYhPcsCKQx8MyKS6XBzhN6Bh8pVP84Xu7eDAYct5k
9ZzZAIpvQvlRW1ltVOhKNIRs6InteVTYmhvbZQG/pw8=
`protect END_PROTECTED
