`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/n887EJbjMqAt0iHm1MujJb5997Fz6FJhckT8Ngbj7reNJpgDYuX1I3NDrq4UG3O
GcYcccUceUJTNMt5vIgqw4n+LtZ8kR4zIPaPjb4j4OBsTQmKeEgaCXLtomGFZbom
yLxgOGLLkTI1Ivi734gKih+S4q0BMB+ViGcnCLYh9vNj2JKefJD7DtTDe9vhFu79
a6SzNy0ojMirGqSPSPmvHc55aOye8LHSib0FU6BUeDTXsDDQSLuvjWAz75O5TXfm
GeSbCGUZE9WloqvokQ0XfIaweGs/5Ee8xJDrzeveZhSHtDdpqmxXY0oahZyYmRTM
RKNHl7PjKBUdG1TnaNufJo6sCZuhGqcNE+I6y9tHv82SSXd2OyZpCjRaqIHkrYsA
fkexA2vr/XwFYc4fAMFxAr8ZDnvJgRFyCrG7IB5lOKaX1MQg9oaPbSjCuSWp5i6V
FskZ502HGMPdG91ljygHMgJnDLrJBHqEx3bk2QAoZhxC035Lbn9QoBsvUeNj0jBn
xVojtpBtw2HJu1QC174w3Bua3WIOPXLv7AwXpa/RuZi6dg2O74t03GLkae+3QpVL
aszmpjwNiDSukmS8I7u2DElyUdKIlaB2HRv8vG7iwSk=
`protect END_PROTECTED
