`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V/yhLYp8EBLdl8LLS8BWM8/OqgbpDcIgh33YEKPsh7hcX+aN2C7JMu+MZOkKdn4T
y9KC+GR9hmrFFzpF/owx0u3tT+Oz58wt5RH2lhickteemdje31T9Ov2/JrK2jWMg
5tLeUxnRujvkC7OjP+xovpiK0k/ZmPQeeDPpnOnFJ7yZjTOEhDSdSBXQxd9DaYWq
4yCIMin4sPwlAmLHjbX86gPUIcCULP6jK6os/eqZIFfg5dnMKvF13C9jw2aW/76A
KOwSS7sTnuTOK72LKMzHqB1rWg7SbN9Tm7Xvl4KhGsZMQgmmzdAoQVMZNGg5ftFy
ZycEh6EwWodfVWT1Cwx7sCMhswZi2x+jg2a9r3sSXbhALUqd1jlTIVYRTV7QmDZ2
8SNy8ZvqJccqwGVmhXCUsCCBM9ht5MDoGyLmB+l0fvk/upHNNccG0YxPrm7JIqkH
FzQ+1zMd1JJiWzvBHaZqsmbTCZ2sZwGLaynsnVKYb7t+WE1WfVgsDS+I/iOayBYZ
nlkSZMiNp7ay70kdPe0DMvjamvbJlYArvY+88JIhR1+dfaNk6LmrSdCH9Uhkqr9P
jqkwYmxLHEdM0LKQ7JTcWTonNfYrW/gzGGpup/yQ7b3HxDNSoxDoiR9u/OIaiPlA
LK2tTFKn7faHAKinVPA276RoiXvSxOzk+brvzFTu2Axk8stDmdArtcf+2gPUXsVR
t9j2czjpEqbfDNv5+qNMKG8XyFi6FFamwzmGoKgUvVl0xHPgxvbOdv+/ZK6ekMnj
GgvNEzFKMfhg/vdDya0Km3haZGIbIa7gM25J0DaWhCx0DGoS837/lLdU1EFhYkir
3gpr8qOWMthd6jHbYvNviJpTDbMbeGxhe1mqtj0mlQqifJzq861qZA74UYvmIZmS
GPVhgCXCAtZH2tRBUJjveZAkeRKLkzndXLgkoNiTQxOdBC2wHIsY/Igio27JPfXY
FDLvCM1UP2I7TFp9gvLWzBtMuYuUfE1Pufu/ltv8hoy1t0owbg7S8bq6mS2Vkxa8
VjisSIY2AiUmkSTsnM+aoaqaMtgahIab39TOsqJCB6XHuZl7NcQr03SxCFuamScM
F+39DpzBCBNTyegW/JYBdo4VJhiJh+K8XmD1u+b4x+lprhoV3ybLygLBmDEVvCWv
mBBYDdtgDk8dOwii3Iy8FGM46PFvH+NHn0tUGs7eMp8M/vRnpkVrm5r5k95pH2AO
yEFa8k/KgyHhid1uGAZVJgywMVPvPAUrZqpJwCQiWRP6UZdXiWyJLJQwPP+SYuID
OHfQXWyg6DHecYfQU1tJEuAoidUn0hEL6JNJl7c4CKrGemTVTw+8O091pssoh0W/
L0Fz+W5MrXwrRcNQIawFeqbOtsjyBb3ZytB9yeWvX81Y0xWGFPGaR3n/TidDporW
P6g1OOtvZLpXBhHK7dEZLpL67bUqHt2Y4SLPBae47bTIciL8ZuJArQHQj7u4Biy+
SYqcyKWf5HZUmcdnrGmJgPwXSVqnt7LcdyiBGW1Y+jjcCKcqIcG9L/AhbnT7Umnt
nGta4zgpOWQQLDf4o1ILEle1fQwagMeyqCgLMRoj2V9v2C3AfXjNm8py5tSCyHqq
wC1L2XqCMmho19ilmso2hfSbIx5Z7kPjVS09pNuqB6fpl+hkbdQmrjWH5EkWHh21
ftVfLwFWXMFnqdx7xc8W3tafK8lZ6ifpf+YqLqf4EaPWW7fJEbaNqvq0p2RTNVpe
Ukqi/2cSBKIKiP58H2m89n5pFcAJZTc6sky6PVbLJk+Df06J+5+4v4bQYwK6QQsn
TYm01pdVG61qjKyGPBCoo8HEguo82KOr8Xn8raowUYMycECZJTvfcl2QYm4CHXXZ
ieZgNEXr/91eOKPozAi2BMaR9XI2vZcVAFNbIKV6uuFVi6keK2VlUtUwaxjFx4iy
O34a2VjByzPMa5fNalBGdmyUnfmCAqW1oPRu/2IoWNYYOUnLX0dBr8ZiHiTzg8YA
aI/rLXk110htF6sSPDGbUvvzJdyvA55dX89CGfPJ9oioZdp4UD0R5q8FiIpIxezl
oKN7qqH6cSLdt91yOFC5S7hIchpGOrdgm669OKEUn4V8DQmJA0FSSK+18N7qPquH
dFMFAFiwlHf0Y59FhNw6mm+EvccoMaeh+yG36Kfr/VA769FhbRDkE6ellU75OYZK
teSR/Dh+XsyH2IGmRJd1V186MDA+n7JbZ/ziX6EZlw6EIax4xvqWd9S51BGm+ROT
EgKvAk1LQopTUxiKlDqbGuOXtd+DM8sK6D7W9orQM8/JlNS/SttXbatKXynpHKDF
b4pmsumU3v2y0GQRmnCRUitTt6rngS0lWVBZDc4iK+e3WDPrd6fzWFTGVCEgGo15
vhEgbtA/uOr9w3Ofcq6SGQRRh27lelrQux+sCH464taQ20T2JKfK9GxNy82O0Q7h
duEhlBMD6f/cIyhNZ8Qp2e0IWD9NK/VqViw1j0cz05WljIvLj3sf53SkJL8bfwFt
Z8fZeBaxHeDCoXduW7IMbxBEND+YN+y37KGJJ+G88yL+BJIf71e9WJxrMdIgLoXu
VIYtkTVvzTUnXFc6qS3SCuIeW+i1q6v2zEOACpzjks7Be3pZgrrz7I/ukv0AK47i
JN8Dynto88Xqzhu5uy9gvPtWAPSgAO1hu2bAYVKRFqqPoUaSGMfyDuVvfmGUZNG6
iJPEN5BBTverL67MxhQBTUvdx2JGKF/pGtkU/xjHMIA+5cJjW3+FiAb51mJKyzdX
PuuaQuQS7JoCKllqemK6pxs4OsrOnZPXflNFAYDg9ZvcgMYfb6iw8xqugLPsOlg1
KRvJxk8B4tb97wIQHAkgMS/YxnKcDKRKYR4iaRLRW09kFQDZtTawb/A8Qjk74EIJ
IpHQ34ZIUuR8wxyWfj/MrfBlNtB8BlB/1J82V6EwCJJy+d09TJDX3Fn1IqZNBEcq
OkbWzF/+U8i92cN2NavjO/fbWwatKFigx74DOOfweIwevzN/c+gQaL1LSDfJYFAa
TNt5mA9n1QHajc9AGmq6rya5qzdwDgL9ah/Q87fiSc+AOa41RnDEaq4Moi8hH/Kq
zWE1IbtpG+pj/S1TOQMydtkpIync4/PjKj+X8cvgkpiSgZ+ZJYFSY8MwRYaUlwYh
xoeWlB2OzPiB3xi6pDQzdDrztkVypSJaDAfKAiAHJcmGduw77blFeg3j1VQUKesP
oARMwmaInJZZ9zkoBf6jbcAJhODQH8iMPf065qpg8GU+p2aKorB7CxQf0UyoFmMI
rBnnwtHJXHIxRfeQ/0iA88Bok1dpnvPXwWWKDT2f7pcg0dlTEW4ozQ3SUy7D0zjz
ftgclBsN9lgXQHjD6WWtRkiNdcnCNWWHanmIDqfHIVLdDS4ZBXd9eokNZf3oyqLz
xWZDPtXOqmtBWoKyi3/Tr9oVdCL6TVLR/DXAXiDgSSZqIB+BlPBq8ZGM0FRsvf4i
kmgxrIWDqS4plu/aD/n8BblVMqRtsYpGGOIdrMPkqeNvKwUOSG1zT5BylEao/HyK
YwWlrJxIcfXSrd0ULcM9rfELxd0iOf1V0SZaOFlMvW2ePxjwJTQopx5PhDgRLwyt
N0rlCdfZYOoqDObGoUfzbGjse9dJQqC4rOjpVSmG8DC8EYxLNfqXS7VNxamQsFaf
LOOng3QaKtttMAPUSxkTAwlw9UpvmArDehts/2miQvhVhitzbCMVfY2ru6BvzW98
sVKtSUmwpluRqhX3X2vaNm6KBqCi6MagbrqGw5cUiMVCv0lvTzP5DCq39Fwqm0lu
Rpiwg0e1KMs7vwlbRi7lPx6CF15Q95ZniXQbpXxpcbg9G01fEsTvnOIzIdFbLqMN
eBaBdaCsNUQCWmDYdwOrsmXyZ+3fkefGDrvkxUOVaYL0+pxP84z33Bx4UXHqqNdE
w6ttwbaDl8f+rqOws0hh/jwLMjBFo090LQZAHkZhQbhrWx/fgGv0usVb3KaF3lE/
mONP4olyK2FwzMIpWBkJ3SNis4k1qUdO44qKdn+a5dO0Lh77p6NLSA6Gf5vG8/eR
TzZQIZEiQU9hYUdngDO7mag1Z+CsBO/WcFGSohBLuXjhM2rjQyzSH0C+ttlzvGbl
1fzKql23fcQBrFAxfNU30AlV5telfAmjO+Qb2jP5ZCAs1GXzkRWAHuo0zollkMXL
Y+7CSCrBVwFgy3DeL8ULhQ0BJugxC75ZHhYFhu3ujD9iLei7iRx5kN4NBQ5yDYKT
GzTXL9Eqe0DL0kfRS/09Gd/feleES33BHNjUoeoCIHHdvttCQYU3MdvJQU6Cy3gc
kUSOoKQRG5o8kwpHemFUncHPFDxh2FL0uYS7BJaSnrJtzVNpe3tOwlbKocqGNVMc
x2l+PJ2CyGvuVjz2Ns3urtvhYr5n/IuzNK2fMA4Fb7jEnCeiFl0OGfj1cPPRx0HV
NQ3sFb58TkqutrS9n0M5n5wMrmicF+iSc/6ToVEI6eaaO0EDf5DKwlijYD4/rJlY
CqUF2ZFXpvLtPeCvHlIcivMrGYrfsnOxqvpCBbGkR1I3YYgmXWrAylA+Cskz2V43
/sUDxTUQEaRju9FMPFtaBnnEGm6PbblWISkElvrBpxGkGjhGUUNea3kf6tT8M8g1
Co0oJCNirq/g/T4NbN/5zdG18rk0Wb8vSjSaww9zISF38cPxc3V5oDN/XrNiDqPu
+M7IXK47bfnCWg9tNHUEQP8wyLQTrNHDVk1yfVVg2ATIP08LF16Ejpr3w3qBbcBs
DsGIdADqG7/sg4e9abxlv98tv+J5iG+vsQheA/O6SUxg11Qo9nhUq6Vuzfit8kcV
cc8EPMgfG+elAakHPH3Jp3jHl4t+fYAHVHxGsZZbbsWz48QZ68//m/t8PpjdCirm
R2a4+bqVrgXze8bpKffIUT4vZpQTisR3pvmpx6zG1gl0WiaTZYVxazsFvYAyy4Pw
NfuZ40cktGD2Hj6RKmpWqvrd5tl4h1hQQs31kt3xSZ6kyGr0xD0ROVmdWOyhMx1m
9+ut1/fha58Oa5c78py5zhUChCa3wviRkZ30KkYORPwhzjim3WhUm2caIhbcQ+jr
y2Hm6kwUp5xvmQoth+WWUIzexCWxvEMYLC5ADrYquPYYFwhrBCjw+F962P9Y6MRD
rlpWEM9nHue8HKn8ItXpS+qEAjoVaSdNgusgGjbOu1QCHdXNBr0ASQrBbZa54Mba
Z1uV5ElLR5OVKADBVVoKxThd4Xmkb1WIa4MPd6PiaFKeZH/Nw7DzqwJyLoLvue6s
O0ov9ELYGCK7WyCKFlhBqyRTzVtkdMV4I4u7gP5nlyBzRiZE8aA+ORtzJiLDdB+B
1Z2sjZFMayjXeIj7fCPh62bSfb9qg0ogTPIzkVepL3NZYg6rPtogaDvrBB1X8hv3
b2eWvMgh+0d36DioZUuSTe3eKf5j5QwNTw0jJs30Zdpqsud4hsikxiEoA2BCSOPI
hnbDYHXTVpiHQIIYTD/OgvokGzruW2d5mZ+u58e96oLS85CKG+IXJu8A012YWBVz
/TvjsB0hp/eSBfnw+3tSHZWBBzJwjvbA424QBxPgye2fOogtMz4sQyN4L0MmuqQS
7OkdwpWcyw88UaQtPZ4MoOPHeNNhRkkSZQpy1OxSCjQ0q4+me0c9uQj6I5GtqzBW
xwg8ub/Rr5xNFBmlhdcoze2lW4rkdXQqIjXMgzzF5oOxHJX/GS8ZpC/1vOm+1AeK
8VzZNxRCxFkLvXTxUbllUsg7tv0h8WRopJyAYZekI6CE/sL5C7M/zx0jEekO8Xsn
zK5oyAXuTp1agvW/lTLiqk49gmEqP7QNWJucl28z7PjzeyFboWa0QfTdv/13Ob+c
oJkJ2bjmnu+4yC+NT8sCPxTAOccIlaSxtqA4YVF575R4Z56O78Z/RdYEnSGssZmM
nvycCZmiJE39mrz2lzxeU/JXfIFiqKPMbK01qdjy3sqBYgEf5uqcKQtyY2ZN4s99
5OFXC2LXSLUbhCAhWeGWD4pPl5XuFQk01F/pjPibu66Sgh0Jqn5GDi8FuUu64nbS
8LGP42r72ED2OLS51s1I0lLfk/WEpxzr0PtZ+Uv1ne8ozAJRmbNBsevRNSJHBPIj
wjrVM0UZnCduHZ+GHEnL73dVCmsH+/euXlGTxbfPDZT2/Fv4z7Sbp1wqrMrcZrWM
6CEf9lBT6REYTucLk61B9IO8n+S0Fk/aFE3wgo46n9Xr6CqFzht4ZBqOlPHTr/yp
HpyUtth26nsfI97qEhMnLRkcwsxrKQb9pXWjSulkYXijYTxO+o9PqKYG7jH5yvIg
ZcSGAkR4iIiMMiQVC0hDFo6b7JyVT7Cr5uK5btR/VY9Otq9TJK8qWSv2WxlyyCmX
dwQtdWCVPzTVsp9R37EN9rrgegeghmS8D2Unw0DjUHQ94qSlm/sZf3kIZQLYmiro
00ujJERT9fNeA5rPx32rYI9WhhUdg77oPL070mqm+dyp3zuZwACBl2rplmDCcPME
2LcmM/Uj82IGfylBGm4JNaqjfr/dUzN2cUFWdzQ+dOcvrPL8IMRM/FKCy855Qmfb
yWGy/oSQCfDqrnBep3WxaNpKjge2DMLNNkmdtUcwOLIKkcA6K3N6/bMsfD4nTlCF
o3uC4JDNTwgKnC9o54wMJ5T6GeU9Qz4RmBrojAxXmByngs74gsYiKAx+LZwpBSIx
DuvtaiUi6xg/Y9mZXi7xZzYErkAzi8x2BtFQcIDa6bXKuiTep8ry1irybK0CkXtW
oHkfn1g8Oj3Q76QubDaeuZQL9w5BLo9lsvFn2Xgvwlqw8Ur8xq6pKv36MbfnqPUI
hj0OPmFDJjH8/Njdw28rCY9+bOxpZwAffn2Nly34SLEIaZNLpX1bMAC8tBInSpqq
glj6KG3arFQ8vKrfWkoeZ5UnL1nTIQrKcLfBvyNXleZQLrxxx58kGotFbwA85g+G
bteWQd+UWpmE1v+TIanozVmfO23/JJ+XbMk7fIMxzDcFl+dNDrPfbYaniNlEXs+R
W9SSk3yhcqo5yZ4WFpIBYXQnvxp+1PZxDNCg6MrD92cHpgtJxqrgLaguImcR0Bu8
0b5nSdmJFkB4D8CsBogRi6fTaTksB6QtyhGII5hhDUtaXkdp9XrstV508Azc27jQ
xuhVC2IRrdzkz1t15rqkgnj6kG7aYhpiV0ECf91zkMO66M8+SkZuiFDCt1mWDNFY
Pfwu3Y8cP6y/DIvllJFBDZYzH2mbB0uKBFabfkzPex5pRTA+7a4ZPdnrZkumFlAK
tnJbcFjKWJW+fzkEBLnQVDNdO+muRLiVArKrlinldvu7Ra2v9DT7Wl8KVH2DNioz
kF/zxRP6C7Txu5D7+76Mpr5sREqEJYj7lZijlNRv7ijv6GiyLko5vpS1Zx5qMGk0
9z3XpiKabgHRD/WPHF8u3bClPg45k8HGT3eZtyIEhLl+3U3RY1bToOxmGER524ru
3vDYYiexexlKu4c6eeXM4HiAYNo+EBliqrbikCCTl06ReU8ISIBH5mz7T7IH6Qgg
oeR/s2ROmrFMkTWBv0FXV35p7q2M88TnHsEMw689BcRr52aIOyet6B70qN69tb5I
/7N2Iawf2capLg08asz7LBOXgTZjn2G9d42G1e8n76ylUIapO02Sz+pNqUIODJRY
szASGe/3fMR83kltnDHziPDp5WQYaJWfwFfstPJUUrOdC4knyvQJ0QJOr+JyiPa9
YgEMpsmxP+FUmwEXNGfcMaL0DAVlaNTY9b2nraAimcy7nL6h1H+QJwe925YpbjG6
AMRG058Pc4eomm8f7/erP3sw6KDsN6RuruL/zZYjV9hexQ6RkAgqldMI+ESKJVwC
qRc8Y/HHDNUcYFgztearLCHTJaA5+IePoWzEyacRp9TDAMOiycr7CVpH9QRzkvlD
PwY0QuZi8Z05rztFE5jDVJxywC2gJ6KY2Os5SZpqvyqQAKmww2laEMUb5BQhPAU2
AvNPoakhdlqc31V72x5HmMvQgOUfPWF8wI6673ApJYH7CUNwrdYKj/8rhlPwsJAr
IjBM0msnSY5yza/LZY69IXMlJwDZF8m2pGAOD5Pk/k2famVlkKJKCBTdyntvnCNH
cPBe3ehoBzomJw2UxPIi4simwkwStGgLhgExKx2goChd8RGit17v7GLdfgBsoWZc
T+bouAHoms2ezW4u99swngEqZ+VuDIuWjxU3SM1Tms/wrTMpl0Ta4Ch5n5ofCL0m
mZOrYsjKNDCsC/xcrjqsC0bwyhXIRMlHxALQghNo0SwUwFdhpj9WZmz2fSdKhwjR
Z28LOynXDEMQZpkvOUX/szM/47S9zghndw9Nor+W8tQe/6cjb4f2iKGogYS6zLpb
UaJq5BE5w51pjewB+EMM+bmzB3Wv79oLEkeG2WUFbYQ4ckcLxIdL0MQVCq9uTYkP
BidXdoFujHQOJTnAuR9jrbVFdvpwbu6c5PAKzSIhJSVgcGWTZZ+u6gsWCqqxK0Vx
O9fPqQ1UnL3zbWqzSmiOqt7ow4CCk1Bfm4aP5wSsk8MUpLEgH+9D2hWi20kwbW/h
l4e1z8y+hti5kfq5fxrkqQO1oRTeFv6rBPZn826zbj2cbuvR03Uryfc/CEKQLhTq
OmWCwTZCYqStZwtXxsws/nnmDqzBJuZUo0vD6uBXYv6fIMOfjsbT5hmsaqBeb7zw
dKLUe0FLvfdu5CI2NXi+k9RnVyBNkvQlwxTUqEPBXNJg91MUo4BxfYR/FPDCptbF
YwG1CRwmu0kHvXdP3gXkr0LLYsHCErBuC2cBSSydb3FO8kpaTXyuoJhyPt+WwCO3
Hl4Tic3GfkS4JkKEEtlzh9aGH2MIN3XraKhEnXIxIwq1hwkoOHm71GLNUUaoeHt1
Nv8icZ8PlmHHtidcr7Vf+59ZPrU+tL6Bczqyh3YzybMKTTnOzp4I0xybhSS/sUxY
FFoFDdKFZmIJbddMiqDHYwZpRHDpe4whlSus0W2rIH0zZGrnf4cGLkcXvdWbKoDe
NeyvJgPpOBqlWmiVDDza7ytjgDQP+Ek7++IkK4KnxV95z33baJNSkH/dIzsjn78n
80UbMkW5PT3etM9gNfs71Z7z5jO339jdt3uZHmeiUwP927Ag+3RQTCbRJ9Z8VaVR
ZfYRpbpbje3BUo7/uaxkU0IIFQfRcpgeWIaBfcncCFIBViCKoazImz4CFKOhfPi/
lQnJwy/QdTLDQlngnxDa31N752EsK9RSaTwP6dHPhmadX82LZyx0olz8iE/1uL2D
MOdUyAVV8vz7wR5xgveaP2j+On8+f+QAzMq4vmGpcOct+UAAkTGTY0YJt1Bmkf2z
FVKVJCpN9RZrOnGyHod/dKbvpRcUqZ5RhaC9RApvqZtEpyGJZ1k9oGXnO9NgMv3M
yicgYDqv9H3+rYb/AcwLUEfxOOaO+OOsNEyAGC13WA5v91SjBIprQo9ohgYUmbba
deXpNrOJSpowVM35k1hF2uiU6n2A756Sd0LC6ptSM7sZUTngs3W6WhxV8n0iG8by
nAruvUsyP1FB3kGee12fvUiz2OvbZP2moAjwf/UUuxej9Pkmvmh7CMCG72lTxoMK
Qwn9cIvtPj0ZTGrpbPAO8iYUjYBoVUYI9I4DA/Gs7ZSpFpwPhgPRfDtVuvpyYaSQ
MkoJwqdvIN4R+SJA3Dp8YL+7B1imA0B36LCdNQ6I1S/Q1+bJjeQ9z6rbbvnhhmjJ
OtNySwBpcjUFL52wBJXz4MOAorYnPuRsVRtw72Aj0zlzCqLOKqKnAJM/23qMmYoS
+A+iMYESOE2q9IuXk9N45akhpZ/bwamYW2BawN7uB7CoxU4v8vyg4/TZfEM1T2jW
+raobS2cOW7XgM5DEC7z6PykWX9ndy2UM6h+gLii+mxmsds+2rNUovh/Gr2Foi5V
SN+JL8WMNBrL/uQK/VNOiuyfkLr9jeROjpCT7lr9cOtxlBnO6YnW+faKXO+BEikY
TLMlsdmaHHZDFO2f+nCjpcIVIY7Mz2h8tQ8F85YB+3s/Ou52wsnlkW6adliZt7Az
wWAiXyMUnW5roYhvpddi0WqM2s19WKsAQZzViCwekn9DViYSQky748qilplw0sYu
ce6VGpXzSOPZNM3QcW3jBuIX5nd8KO53OLCmWL1phfhzw1ucRiTCZItxo1iT/xga
wNgBKIkYk+qFrwgM8HlI+Z1jLsD6hsYKWMsjMSwARalkVOBv68S1E+tZGi7cvEd7
fMQpqcdZEqixPATpeTHiLOjRrnCoFBmI2aRVvyw7ADaKDx3ZlDNRy2w7vaJJZqgu
xx/fNq6hMdC4af4+OnmkwiQIFPFwmszZqiouEzPeBilGw1ZSqFuToRYjHI3c4xb3
pfMVQ7CPjJAkK7NV5OvHJr3pBXgmRB7Wehv/IybwtM9Z7CHTPVnPzNa9Lcq/9uaC
kHrTRvc6kXnHjiFlNNv7IXwzvKYtY+G/d9LOWP3UjzQf2xFhdJm+BP2YvoQbyYNB
5IeLDOq/TCSt70e+wZkmsQmPeezLb6jYUG8urHgFMDtF/iteWF34v6wIZfJP46Uy
+fYJdz7Rd2OCc1XJ1jshcey7/KWXU1Bv4zJBxg78EwVlxXrS3+2DbMTncgyBBd4X
FjTdJpj41ZS0XIGFWPy6TLeJwBqGSHiK6Y5osF2ur2w01pKE9vSPzMi2hIRWEGU6
zAj3PzFOBFVJy0FLoh/x0iHxEde/3XrDnRhk+CchTXv4OwD35KW9W5J4k7GD2JIy
iXgPnqzKzUBHf6TsUAwwwyK35TYMJg0qRDSqMBbe8Y+gd/zKDqIbkqi0x9ib8Yda
weqgS8lgzKqsIwRY0LBLzI4I3nl9YrmbxLNF3SvTYKyZsrkhr/wUBz6rZt2MpJc7
mJAMxOQs3HXL07tnn91/l3u9BlzUShvfuKT2bycG3zhFLi5JXlwyKsjvq0AH3L7f
/Sex6NsqELr3AjBLfujnV23O5aHIW/V23uu8Y972cpAU5e9zuQfJCrAN9SB7LZK8
xg3SBgypGjK8NU6wxo8QsUD/AhXFvfnvw9Is22TK462KqJ5B79aRv2+fDNZfMDyC
dFaj/lhJFMHRJWARPvDMrhbM66ImnGUmOhvYRaE5CwWs0uGE2Mx/21h6XvMNLbRL
gScmwcy0Zai4oigENuH6s+NQ2e6Hd1ECsT/jYuEXvNWtqDz8AsOXGGztB5MRn7O5
o3KkKcYoealnwzvkFZxcChBYQfCpSss82o20PQWV+M/e45LNO5A9xqgjqTvO1ngC
wcmy2iZ0w6MWc7pySIICezR+U+dGrpuPB/I85DBfgfXUOFpShpYFl3SaPyPlYSyx
+Oq0nlJOAuX/d9FSXV+aZQetaE40h37/9PU21himSL3vYlFjjk3f75TTMjkWhRxt
TZ7MjTw5GEkmRgxV/g9dF2Aopd3qBzrJcCOe1ryH1QwgHLy/EhlcyxeJ3p30f5p+
kYQtwf4NMkOGBSr1FRToT5okMko8ED1m12d1vda5zHtCHgDFgvHYsC9CDr8xZ5wV
9bN/LLz9278P5ZH4GmH5c5vOCstdcHi059S5PQvTEHc1ScomK/cqLqRYfHW6Hkir
bAtg0tLY5nGRIfcPieYkU8+ZkKjULYqkcrWSTgh2PpxzSB4l9g3EsyCu2z+D/TWn
7t02at+tiB0ixHRVsFsOQ5xPCx4NCwmmw/dGgREQDXl+tc72XgioFNDQtxiccnfZ
/CDSYn2/L4qakO09tdGL+uxLqZeOtleG75bgNB+xtFkz069Jsde5bD2wBXj9kqxJ
pD9haThewZIE+Y8a2Ix4q+rizwTKfoax0qYE0uBkODwjRsL/dQPFJDGdG7rRNDBq
h8ObhMP3/sCZi0UDAG5Pdg6R1iQmmQdSG1Y2ER3IBIR0NNacr9RCeFmNHODmQ+Z8
0iqoHLfZJrahvjrpvjPUafhFEweB+qSjeSit4X5ACWM4EfYm6hA6yYSxDgqV52AN
R7xoNYFpPaXAO5wFpAiNpWM8H67PWjml1FCzKoehc2CqwcPsUOztQNCDqB/StSNf
ns1thmI4ijyYKodfms5GQvvT7InzXz1pQIA8Jh/n9BpnY40L0LpBIQMjh6TtswOC
JS0NrLCAz2/Xa6UlIaTCIRNMh07Tja28XQcO+QBv5dnLYfutGXMvcvCQZSpTRYzI
F4yLl3YEsjIf489ApvnBE0WGNGvywka5Vd2irX7plmQv6BxVT/2MRm2wBeMrKtBf
s3pF5ZjmKakoH8wIAVvwzlp0+iOZ3lXRWpVi5KUKiP+mboUALtKGsKllkgteQcjD
DVepH0kyykS9nbcRssEagaq1UpwdiUAPb1Oqe9e8/mVyjhwDVl6UGpT1evvE+yY5
IsGiqMuSqM84ipZCK6E2PZCcLcdnsxCgji+CS6gytfmVl43N96ed6c55exES3fHk
kyX09/DVBiU0MjcdrnKVHiGBTzKS/1Zj4e+wwKAxnDdtXv2/v20Due8aG3PqJ3Gw
WMpL2HNmBKB4FVhLfFD0nM1zN8q5pN24IvDPjc7AI0kTal8ZrY4GSOPqfy2aRs9f
5e9XErJn5nwyF9J42V5DD8kfcznrFKlcPbqSOYJg3wGgk+S4KAAxkE2DcjKDJsPM
E+R6DosSIJYx0s3Vud5xYSQbMiEqdFflGg90wh7DrPAF2PoBbs5no7HX+S1gd9kz
R4tMh73/BPHpbER2hSyJOGmRSZqxnzGopoZCKL2SBIC+OrPMvMKrRP+yOz9+JSDc
C2qySOirPJ3NQ22UNYnD//uE1Hx2Tn09SAZ9HpXSHvY1vlJNfSE8ALCtEjkalR/s
hcM7gPm2sE1fSUwCqLB8N0aFcaWmZ9RQ6HxUfgwzJ6r6N4k3gEmxQMUbikQIeYn5
hf+FAJGfUCxDSV11jbh9cSYA6bbMCz2CZdSQGJW0xg87LJsdcd8jSh0gw0BTazwo
ZlzZLvvoeMT7JMc4LxOmIBOm0M2RVjOWdBq4sj/EDoVFOMrgGwAsXiWWzmWB93Pw
RDsvrsS8/6pZ/xSLpJvTIRQnJB6pVOJlodF/CvZ95enbgaBdvCZk1tK1N3xrfXQI
niWnOi/iZwD8Wj+gKIDAs5h3zdKrHLrXb6JoPpXooeabcRQY60QYtIWkWDcH73GF
JcthynJKktNZSlJsRQMuZxyvwZ1924iOnWz2Ago9rW4Umxb5oEX0yXEIBA4HDl98
kE6ZELhg4UszGSh60/+2c9DAP67K8YCJopee1S6OVUQ3UrP6Ll+pX8DjrIyZRYy7
PYTWFdVLQgXViS1eiuNh23Ndf0LFU/KwSIYkSwO2hKFaeO53lus9/juouYmamo18
kkvNnBEgyAuV4t7emwz8jEjMp7mIfQZNATnpZIvKQYtHGGeA02yaMj5ex+MEMUFc
djtsWuIEXDh1Y6dS7KSVmpcasN1i55x0y/ONLIu2mTc1zN9NngdBF51G4BxuRIvR
jqP9Ad8s0MW7qTK5oqiPrT+D/biMM+D/w/9JPCueP1VsWTLfHuSw3gOFdQ0LC4rG
sxDGn6qzT/BbXydYhZscIkxjNVzsn3SE8UlEQ3VKhLudRpdkndxQSfVgM148/VyD
NG38cjZyAoJWs9p5174jjGG0g3TgO7WEzH+T+w0FNkdGBW1F8KaSRBBxn9d1ym64
jbvWTCwqFG33Cjua/pH4yXKJBL7gDVTj7nlJIpykX+O6ufD5DD8TUjxXSsNPy3L5
i0pm8VdIaXYUCj1+bwBNLJpQz4GbMNUyWSLCrkEtd+53vQYiL6vnRedqVW9UlVtw
qZS3XLXhr6TXHEF46H9gpO7EXifA8mCjdNhZjfZfjxGY6G5f93jD9nWxKTU512We
dE/l71zN/TF1tUAe/Uz5MTfjK7vfWmK1EGY123r0iaG6mNqdepgdZiN3noCjdZQy
Iw+Il0pEH0yqlaWeHL8V+dNC5qJYVByVqrewK3/GLJ8OlPkCJ/gXnvdEd9zaYosf
yfsjmNY4gWuXdPJiYf+YAD8oq+AVHMl2cDyqIYZcY4+406Dgxq3HJpBvH+0iPdBH
o88AKqn3MnrGz5kTvK3NH136os39SwiYElk8M7Fu9CMgscRvHVpBePmKxg3aeMai
TQ5JcenieTQ7nIsnJLj1PD78G+uhZAbr8YBy0JfEY1rOe8dEoe+8FKMN5IU1snL7
h4vgqMLuCofJd5SG/hbefQHxWeSJKHAxvt+cHUDiDETM51r76wLj89wDK2tddYVZ
lL4hRU7pa/Vy2Ll/wjRa43MA+OAgZuqE36j1qkto0s980Kkmjdhc0bQblO+SF4Om
Jlo7mRLc0I1nWLPFhnZKOW+Gfd6aLCDnzmKD0BPwyn5DdAmIfdG2oqkfM9ZhkEVc
PwhMUBSMER8o2A9HVPJGl+TGd4bo0EyFPAFtGq33Z5lpaSV89rSd3P6Iu1pcIFO3
IM1V7v3634tisWd2eUvcS0huEfHEFoqb9+d6Xh4TfhlYCwxY6/ltyeWtYkFx+2AG
1/udx4pQYD4UrzfeaAFyDgvAmjdc2/W1s7QTSYewvSwEPuJBpIdobANP3aVHrWIk
jYDGcLv5lwRfzAaRTsdkwTcvQ947+sWKTCBvldzH3W1GStBPkpYGQU+qUXN3x2+m
/2dbRU2IKD3TB8ICeHDDZrYDFSv/e/1nz52OZ9tsBdpm0DgIwhnLNQpqoVjYB4XV
VbsOwwc7pPztc//GLIt5YkaVBfwCKm02QUE5aTdcPn6TBgpMSJC/MVEsNfQjz1EI
1ymRs2RmchxxP7EiLvFrsoHTe9xHnHLyyOeJ/MLw3uiWJ1OxyALrB+R4FAp7uxcX
+Z3QmvYqurEZ3QvIbxxAEh5G/M0Wz2crGQXmOtB06lWjP0v8nLmicXcXv3b7BH1c
KY84gTkeEKtmnIBgwVEZMkinXFWs9lYBcRv7NycCSOb0u9sA54dLl6UfIV+d72Yk
vZsGANehwF89rY15WXdWepuf3CypfMTf5jdbxMoSXtfD36KeUXdwosPk5sMyVn1c
16CPmwCO7a80zXgOgfhigNwv2Nf/GxIci9C8NEZ0eM5Q8lh1V27BtDjrfJHZeIBi
M8m9thzZcEZGL6JNwCuwAIc4E5RfzjBYXyc1PMHfFEucDM92/Ru8802bIR3w4/2G
+PjN5ECgcaYNy0RJqTknyy842KDm4U3vwBZ5VoeGxOLbGQOoKQGPsVUi5geFb4Kl
yEXrUiKyRCHjUm9mR/fqHMSmhcUrDQgxg3x39gieWSw9BrPFc+3+8exftWgd+Fp4
Zgm2x4bZAds0smCxbiObbIHU4rAw3S5qQTLZe+ZTsWXhkssI9ApuSbycwY4a/lRp
pK+NGPtXWtmdnvfrR48oU0XOghZMxMebi33Nq/1d2kDrl1qAo0ZGVmZODgMk2pxQ
cy3zW43oP3nA02c88+eG1p5bNFrf++caw2qyI2ac7NV5D8ORH6oossLQnjIxO7f1
W3wcVzAlaJmYNeVX4sD6NN88SfVO8ej3Km1pakl8GyImdcrxJ7IBdwfSa/8AvrJr
oXpKZDZIbWzjLxoMMdOT4aFGNnnmrzwACIUgLUWmAeMrgrwkP0WIVjlF9H5K4u0L
jw7CLb3Xi5eWJ61IIB9zhsA9DWkrO1nrj0Z/J2SNDR7L139GJlDtJQOMGVGrsD/Z
C1zm0Mhx0dEb9t2olmGMTLoTKu7DpcZpsua2Jrno7IX/QjkBHU0S8dqsOptybx7a
dZP+3z0bLrJwd4RIxIiewlC3A2vh+0dgOox4GWUZGK33E/3v+UezMBlLE8SGdFqj
v+1IC1tozgWsUNz882MTGvZ8KOhckx7jVe9JoDEcLvM=
`protect END_PROTECTED
