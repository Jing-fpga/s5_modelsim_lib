`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jUwMfND5+zppFRCFOKM2HULruu4xUST75IKTlz5axeUD5IgwE3CcBPJ5x2E4F2xz
1scEy7IBmImIYpw68YEBcq7PdQMzjAWUGb1pUrD/ReBio5dVot9O8eA6Y+jKynSw
vi+IW3row40Vs+2O13HjuKlMwAMQRzctbukWO3XXwhFxFMtAfLjfdi0LpCPJ8rPl
H6k7xTJZ7hI9wO2CGYZ1xgvguUiPCenjlGpmPSA62MZmYdrr8CShv7B2UvYyMsr+
JlXVOMAF2BRWVZBKE4wHZ+ro4s4i6tb3fE0eVFlvFxNiMRhvT7iDIp8bqYk/7Yin
DGp3WxwGMZwG0UyDWPHL86fuYZfTr2xmGgfEJrh150mwKaGtNI3VnBagSue3FeGz
J7+AMdJb+76ButudaE/he0HFylNjXXDyjvPL64HF96ikIQN1teN7NOrqw9zZrBfr
mpSos6V5MrJp4/RLSv9RXY1ZJENk05G2UPE/Ja/aiJFflcdGknf8Pw+sAq03+EEq
vkLvr5L5/NckXDgDJetZLnEaYKELTqaHhGKMpqF5YS97oHfjK97TIRwKbxu6Mdkk
j8Qo0412wQsJew1jGlIgOUEtllXvscMA0P2Dp20bCgLfqbK9CqAAYNozCTrgr5rr
9an1q+b4ZUz8+vQTarbcPJW5gVC4A1qwkanVuKjCEjX1HmIK4MsGMVymBIPCXwSU
`protect END_PROTECTED
