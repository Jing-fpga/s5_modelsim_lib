`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wag1KVNxYnnSohiiKpF0fALTb2XBGRMoin9LsUGP0fyz/BM/ZBk0c/9nTbDndob6
UID5ONrc9kRB3uKhUmijGV7dOE1XS5VJxYYzct/TLD/DSLCytZfwQ5julR/PQfY4
7w0kbzYbF67uTHtVaXor/oIHaE2P+3zaPxHQNF6ST6T9sVyQhUA94WOwPlg7/j+G
fMEZCqyOgfnp5i6P1AIMUWwnKPTX6crhnWHAmHEx/L1hSXR1JxdwH42cYA96k19M
HP6kH/KzYsgDq/w56yFmOmI8MomY5k8+bGlg0izKNCI0C/4oI/OjfbsDKyF8i5Gn
FtM5AxgbjHdp/n1tklTaVXT94urNOdez48MCKKz8xa/eIYagvIlN1JBi6jvFtSqA
dLknP+8rtJtFFlLSyzgBQSyUECXN3t0XBB6zV6yCRvYLyEYka4+MYznGNZcNnRwG
YAqkwi05e+vgYnEMr4sdk3LREqCNEorjHU+xohttORPMh5HnBdixdS7yMEAkjjJj
rEpXHF3AisM9gnImv9jPVBIB87St2I81gacgRsIq+oclSxXi3KldjuCqbhemd2mw
dDDjzk4b24anqVhhi0r5iztTa3IC4pHL1aFGzsG7ZH3qCet2Z3u0exKPBXlhsIbj
6bp9LJhVsEEXCKjSzxhoyL/s0ZDUNFPBeCqPOgnNUnyyCXhUzZ0LITtmvKzenMZh
W8ji7b5326114p0bzSBl8ANvEyOvykM+GfwLEyTwMhk=
`protect END_PROTECTED
