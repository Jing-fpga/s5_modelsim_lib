`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EJPOml9vugBBfXpiulYEsQO7JOK8hfZDLfee7n+6VxjMs3WGzcDnAld+U54S4CXZ
rfeGn7Fi/F/cF8VO0tndUxX4UXtqSo+9czzYsjb2ngoPn1cLnGtPUrbS8gglc9T9
5V7xriTvvuSVTK9mUHJFEsPDAWOH+BRYaJiz5vBO8otZzTlfMBlBfXGEjfzSaPL4
7FMt7grkJCfrmAtIsLE3vzaMM3X9EF04SAHcIQl2bcwLrd4wZVlcNqzZR6I+ux0l
mkV7AfJJEJB+S2f3SEJtK7WBQ4Mh06bbgqUBTAAQZhwYytnNS79vV8maQb083gg+
l4Fu4aoUhP0awNAj5xgnyQ3RyXbLmgbQK6Dsh7ODCXvJdqt4ZjdNiMo4XcuOEzx5
qA6/twpfNnyc4xIwSD1T2TdAbJtKpeNLhbLAsaboda53IODcMY2nmLymntcbi9Fn
PaUpRMMEOY6Qk31mTpgrm2IveeI9ALmPA4h2LzwvFSIJBBxtozzwmKLzrQZQ07Va
L/rTUEb61oUowYlU6POp9cWSPb3heGRBw4jj3C516Uz4D8WYLwJrwxfP4l8zCimY
PVQGxdc+GtNJqk4mKctZux3kD3ifn3ShPKMuy5PTRTBCvxBApT3z69I3XnPo0hl7
3OL9PW+BCGhg2LZhdUmi0KEYHO8LQzxvgjh/MtJg19ZdjQQeRktTJ99skUDxQwEM
Jv4dt5MYtb2YqgzXh37wloR1C49jD+3Nk7jr+LpXAgVoT2772bGnhxcNvTA3M+ci
f22KMYEwZO0QTA2T4dDtAyjzh17oa3feRbjkpXG12Pm8lXIhnlm1ryZ720oFjyUT
HGhZ2NZJP2r5gBVSfX/6vjiiqq8a0rmSUjqjuHwEczuYRXOWDPuDCRqXz2NalQ/+
TUEpVWsM2XjQw3Be2W18DlZpj7AEHWlGIXYMq2dDTJvS2L3d8f+EnZYstwx17cPX
bVDe9Ah0s0zTwmM6rUa2VrcPOoc1H/S/q0LZhsxPnuOgSq7TxsXu2R4DM4aJAjtm
K5CijMY1NWjZSZScdSBl4OZKuveSv2JD6jtopKQFTo2+FAZLRoPzxnYSBCT140bb
05wNm6JXaF22cRV/dECCb13iZ7M23fRikze2xHEle7fPvAkAgGL9OcmDG3Dzb0fb
bu4I80lRGyx3lIBKbNJZ0eH7hCuQP3SUv8tFsSKH0jbjOmA1HeZJsSx3Lcnkm8/H
dUxndTjzudyRq4vue8q4UlZkTYDGaLTOpQO3F+uKZjWJkBxOYzipY/ztN51nMpoA
Ti33inuU2oXGa0xyI70RwKM0AYYaeUVaiUDnyZ7ulJq+LWsyaVCdNXho0A/wBodp
laFfBTr3Cm1fvlHIAZPWXIH82Uxj/xIoDLxywwii5NC+7cmfbcz29dBD1bLAr6da
B4g/szaDyxCxJu6DPIxe0Kg4HiIBmwiAHzSKz/QYF6fv7lrCIrRxI4+DFQdD4hSi
w3FTFY2nE7EbN67Ixc5X0MmU1kxp5ZHw5sYVPgjF9d5rbQE/Ss6u5bxLkZJq714g
+HGqHMjaMTDNs54sg2T6/YF/UxGoUCAE2SXw1k8ognsV3HF6sFf9zS4DpPHK3WeM
EmG+SLOLoR2PWfUY1yL1N8jqewxfvSWa5hez7ikFYtJqcaaAkzhBmXvRcfT36p5M
5WO+qBfQCfjL2K2AEAumtLBxbuOFrchnn5Ew+e7y2X4eOQwckM4uFVyd+ZmeqetJ
4ZN8Lbw5F+80ytuP/UORNDfjL3iifAjOwKxrTAKUP/lB/AcSzCWoy4aIPmBvC/UW
G/hWPHSIVNnUrKiwxkvFmYW7WqM6Hx5YlUJni65cFy1+Ceh9BhS/bcoWpv3wGx60
bkozs49PnszrDeF6v0WiNYdyFgX40UByQNwryco07vQEMHWPvuzctHIYnxNb8Z9L
60TizsqRRYZQNjaGvtTaCXboKHCvNHDpcgmfcZAnE2gxMBnxpvIoYs0KeJFaQg2q
TuMw8yFMdcxyB/NB6BwLJyuvsdyFHUiIqga0POBzneXz4yOyc9pVPHmCZZ7u76Bf
0OurM0dUuN4jCUxijGm4/qdoLjN/ZJBaOtTihsJP+QEHkqzJOzI/c6udLE7BOsJt
`protect END_PROTECTED
