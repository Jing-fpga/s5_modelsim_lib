`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TEr6kPKCCiffHOqUTTx/1xOk5VBFEErcr60xT+gAL7GIuKKiTV7mPVlvN6WxafTC
nTjcVIs/rgVOABW0mHcXjaxkrutf1nsW+d8tBH3bTEzMki2G9NIx1theS4Lp0h4b
Sb5JWN3RWOwPZHhrnKT8ymmyNU7VK1ZtSzbjEzSvwKqXhxmibrPk+0sYUAShu4PF
Xe8zzqg4Au7/IgwexyuqqOLd5rHbzb14Vj14rKrIMFeelhG7C3vytg7bvOKkUI4F
XMyi1ZsSqGazGgj2HZx+rYHvkMkO0JVzvYCb8u2pIDaJ2sMROu+1yn6StefKaD18
5Wdf6hB4BUnDi831TCFnpuY3ddof8H/iKk7p0poQZWQiLt2GaYbKEw4WmAkv8K7P
63HSpb92H2b91WyeinhzOsDoJ2MM81xapn6uUUY2YMRsA1cL2Y7DtCADBD7t8jrq
027ZX4QQWXeNMIf+7RwHlcb24DRXi9rR/IEISVt5uSQ=
`protect END_PROTECTED
