`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I9mekX03KcfisSDCOFXV3+NB6GQfeKWYOny9E1hJRbXzGjhg1Dj3cctjkzpRRuHU
L/aqhoaiWIDGUdqgb7Yj/betFOVZe+d+og4pqOJxfK/vQmN7P/oDn+PFMObElJAy
mAigsgMJH68WgKv4YDiqChV3v3lF4QPz94Tff4+xGHHT+uf08npQJGW2vdFy6GYO
jin2NhfPZTGenor6p/lkYBB9Ks3QZe93z2oAuGc2JKrKUW2kdmINXYKj68HE8Xkm
JJwJdjoDmp4J1iH3QRi3JnJQN2OGySULjKBLW0xjHfDweoiBZmMma0JOgFI+cuD6
TJFaTdDaMPdQbfecc0MOuIXn8J/RBWvU4VZ70ipYtQ7coD9k6wDBoM0yXgFDQmbU
+DOPofyzNdSkSjE22Cek1ifyubmtc4UwsdbH3RuBzN//QfZEbfSVMMFBhxGDuBAD
xiXuAvi8/4VsSnNEWAjYTM2JE3Ogm4uarNcnVFRSew7eCTartg8jvieFQ1fbJTKZ
`protect END_PROTECTED
