`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
84+zKpdY0laCMl9zh3NJ7OL1UgAuXh/8GH615/9hzFFdI14yGTqy/PUOZDOkRyF4
3dElDM6qsm6TS+gPitI2ByVnUw/vYySSjPIdxuEjsjqBnkZiKt7zO5JDb7mQ3KKm
4nr2ENhsbApVPaxuuFIIiFFwdrBMZMs3MWWsOiyZUuHrSGE6zU7RD+Ij3JfAyDmG
BNgLxdpBaNyqNmEgUwb/FiwhVmmPgN8hymsRqG0YN/Jt4CjvqW6fFDERjXtfTUSW
3VgY+G7rO1mDI4eFqOF08WJoEoFIuRHKPqFujHvyekmNiA7rFDqvfc82mukB4fgK
TNIzwVNWu05yiYv7WVwiWw3Yzd34ntfy5jGyp1TbIRUeZg48iFlrBQoWQPFCL9oy
EAJ0D12x9UUCVfYDCuaoVs/iBG3L4zf6VzYbgI2sXoi5aJw9IpLcBNWtwtyX/+V/
mmCVXsh3lExjSID+WEmLWen6cysyEFngdpHbprOUli3bCRydnPnP/SlE25rO6j04
o3DeYbfcnLq07Fqwm7NCHqLFs7aN/rx8fxKYXXcM/vnXF+5u7iUW3PrdPQchYrx2
/ecOfBev2dxfeeNNR0jKrbtTOzt/NXx7qsc9XGqdGJFpgDcA/OJHM/LojlEkWsJy
OQfx7V0VVkWlwpx330aE6BmE/QlkMf4n5vh5zHEXBuMOPhhtI8c867P41u89WDWT
gXjggxmnt6n+ax1Cp7Z2BUXrhD94CuoeTwH+EFsf+axPUvUB13yRXlxxWkEQpjqE
tMmvisF45c4AdTmGutIOOwiIhdjDLn75pOYzo7SrEo69RzK7d/A11FuXMT7xW9eC
rZuRfPujI0wmxKWH4gpeNGkuQNx4G4yi5zFwjaMZL5qd2jSdcUc4AkiQugrAMpy0
hKDtJ0eKeKL9Cjx7CnlaXYXglrRdxY/4gjTO8quYWMKHIA89AejXzRKXW8KQQSKz
TIFuG2xzuiuyG5vWWJE4cGEWIoz1NPmVZHnxfwke2YYvLU5pWA8xOqlz6+r7NI86
bPKMyiHV0tNRmB+iMganQh7L8gfpZfbAP6rQN5g4JfkTQc9OfwtmUu6WqFOdQoZ7
UXI+EOgu3IdHx4sLfE5vSq+H2gs0nb5OXdGQ8cKzQ3XjOxaH+fLZX3z6hL6IdbED
cv5iTd80hdSNAXBRj7rvk9nJNNIcxbezz+fxCvvmPqbYI5K6o1IDM9AtLESdOwvn
bK1I1CukMkM6T5F2PjMf94duUQp/gJmgOgradMVakYp4Y2lQaSkqWnJhkBAIdCCx
JrXwyy6smQ8IA5f6LuFXQg+qaprhai5iRwJyfvJ6nOftoS/6ZPn6wsAT/xUK4QC+
yMNvvAgITuKPO4FXtq4RVASTznKYJMWgsDZ4vUDJRNDQoF1Xkd0V6Z61j44SflNz
LPvptE7zcSj7C7wGwA65gDewGNUs26L1M2Qv/D10+OswMz/jZQbX1hKdwU7yN5Y0
wScChmRowtVIlvlkpZxvoH3Z+pfsz6au6YDO9yZNKLMLoNua3bX7zggSwqsPzeyy
u+sms3QcTt+N3wPVMRGzgZJKiB0QtMd98135BQ5+GOhmb99GomP3SmNgZTeCOorT
Q56Yg1O9kmDvV9F+5miwihnid84Cju/N5CHB6B96M9lNVUmlyx1huG8T/dFRR5NK
BxQDZzm+ENN3LSUuMBp/9l5O1ToBABsyDb8V9ltJzhMlVLU7YF2cDJ32FlxdqW9Q
92BrV8i2H8MNn3qgJ1lbPC40qXaU+9+F3iTKABKV7kTYceFs0wsf+md2QGKWAhlp
dHjD0XNB0mkmT3oeSpuL3cz3M+tFOQg4LOlrkvRTyxQfd/j1t4YokJAH3ct7m+lf
QKt9kRpPbpYfec0NP/HbZoVMgOQ7d+hw4JGxo5Gaap5LA6KUrrFOca9pyblgMikH
Mt7s/B9sr1nDnMPuoBiYErr3NTBWyPemU33rz2LWEavUo4EQSD9HPx7O8oJW44dQ
YyhTT1KdhVE2/tSXNDMSSsHedN62IRBWF1AJ07M9XoctO8SRHG6YR6xsmMecvMyK
1wflf9DSHxRpHsuw26m5cu0M+UJIDMdihzhC2vNo3AFqYPhULJe1Q8iNfKrVwD4k
3ZBLjZ7y/NrjIzdl61T+9wc4KptAUh5EPPbsbDPzQrLcCBCU5YGJH28BC4EgSzzJ
KNBM/Eb/z5PxK9IyXGTmug==
`protect END_PROTECTED
