`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I2i01SaEKNmQ0YvsUKxgFElzazQw/GcNMHehmiQoLb2IcIVwDU/aZQ38ublsi6k7
SHr7ugIDud0FIQdBlgTlebVBV3xoc06AnunumGHTUgNiFC0Wz1xEBokAD1csCn/h
2rL4QxQt+WTE62+bU9eRY+LDYjb7cc+HIVrmyZDvzZTCPFumMk7dYasFEa3S5WPC
bL1G753509aQEJDaXEPOyjGQAJHBDlb1r55eHqQg9XwlV0Hn7iagM71ScvK/l0I2
ugdXuukPuY3pxBWaiLBBDYuxuQT6SD/9fxgBngDYFz4u50dIaA7n1VaFVPS1cqVR
Iq146OEAaVdqPZopkEE3IiGMV4zNjhZ8INt09SCcsJm6fGKoN5DAU9LQxadRUTGe
5lUVRElgLVq3f4B7hW8y8ryWUpvMWAeCdnGGmPuS4nAVAQbyFiH0cLpSZaQCozEW
8HkaEUpkGPzxVkUO0GOeaoA8GuH0c6cQeDT97DUj0BVT7s7R9QSNv69CsrHhAdJc
/bIfARhScZvj6c7OGnAkp60hJftJiEeCzp498PJ6W08t2xokQq0Lw9rBKm5j67X/
GzmfvtESftzzYXSj+bI1Vcgns4yvVNFEEA5q3e6ksGfrTtfC7kAWbjWvDoEGuNMv
`protect END_PROTECTED
