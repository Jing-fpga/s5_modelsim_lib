`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RkO43y2o6xY6lcgNXQcy9d5TM6xnLC8ZvMvWzFRjJ1YyLiGdZwTirwJ58f9d/7cF
Da3KwWk3jWzHEC/botmBM3xAceJzQZkSPQOTHkbBABE8EUqFsiEtlXDY2q+DQXG8
rBDK0AJW+detkiEUIraTlr7O48nmLnplkshGbdJTMwJPmSBjvVz/8ajVfhA5rNQ/
VwCoGhMVoYG8wV5X6ZQUhiv//xUe7elv1M8xhmmx5VG6zToTyTxEbH1+SFg0KWuK
4rwMWEstv45+UuU7o/6LDJpYNxo4eV1+iRbc3kVN41o5HslLHi0EntlsjwQLNhoW
2Pe7iYpPgprEWjpSCxB2r0IRWaRhFD6zR3DzkW5/NwY6vS+/p/mXCnmDOJQ1tOAf
OI0JnVoiopLGyPrweUJQbfJw607vB5YgPkF1VDDkS0ZaSzdG3P97pycz1LbFifLf
5+Cyi+aedwqm42zxGmP6QaP4SOhjL3vAxDWGLYdQ7MbIMC1ce1DcoGjnFbbJquvl
SquY4JJ8E6/QvicTE7ifJJB3Y52fN3oAQBcVmtoIpdzpXjmXoFi7QmKfru9dURKL
6dxjXvehpUpQP7Otdvfloq9n44joUrZC3a7FxRPzior6FBxOWRCpc2kYDc5JwPhQ
X3J9l1SNsFSqoUlN0pCgspOGoXp+Czo4fmTbFOrpJer7EiX8/Tmyl5PHxy39wCd0
GZu7Xk/jhFRu+Ad9TBBAJld85ncR2qpzaC8RqMN9ZuOdj8nClyL3NEp4zPBQ1ZTz
LArYUnePnh8pkW3c5lWbsI1ffpzvAYj59zCYA53O51zld1HXwQtQ1RdVI7UefiM+
0JMKsNeFaDZBFGZqhBKFxwi76T35jhSTF7LrK9CxHyn64Ll+JE9ldRVYGNEq1obb
IgZjVhAXTUKADnqE2Km0CqB5JV5qK3MD18vMe8bQ8VbSX0iXC9SlnMq5viiZmZNu
tUxonXhWhBYaoTu06NsJi1sQAFa9sVXhd9S1WCQ4Al9IbsAQnROmop3R2ES4RAez
Xy+wCpzfcOEm19m5dJfOYVPKL/LLna9TlTSNuDiaDAKxC6idv9NVI3192+ECYGzy
hLEhX7jSpU1GcLogkIvfzVq6wf26sxfXG5zuHheVhZKw0ulaG+GlHASsJSAnwZ8p
5xRKGZLZYQQJWyc6W3w+A9Fo+3Ta+4hTp0R+ER46UO1lRvSQVN70WUF3xpna7636
73KnH9B5n0Y6f/V7Kw1WofYH8tJzznCjUTwhyF22e9WVHE5rJr0qGHX3xOWfPzqn
Rl60BHs46yU+HDt8L4rEPMlcw9Icwi6nLCoI66GJek7NqnZ5YtUFehgHS2UCKzAp
trNdV36ChA5TYLgdJRX5OEiQzgBPtv1eLO7wEEfSkL5r0cVLQmhiOMEUiVjFMXjS
G64k9oV2FInFg+pyJKCFMiBltAbHB5j4Jjg4Ze0btI8AARr0+N59jRLp7h6sqP4A
clqDZ9nWyYsBERM0x0cOuGKu/QNBtNXmpq4lRL5Nf4YxfyhXI1M7/5ighrwO+2Rr
uCyfclRxY3eh2I5/uj5dfNIQeYDXOtaber9Z61bAUPC1YbY5elZeWKuo3fqQtWXv
KgCbZO6ucKoS4InhbkCvpY6C9GTdbmOQn4q87OTVvUS1YwzkYRP4L+13n8nxExfx
GebT/CM+Xb0cJtcIlfCcfNWzZHJQ0WDfsCfgyuDrRWsb7FXTV14xFYsVdSyznvui
6XI47mgG2AWqkUjKKhLNe4VUn7HLVI0lA7oW+8DsWWsJKXJRWjyOWP5A4aVa4wdj
6Oz1vCBZx76F8R9vJ1yLuF/NvsoFmDtjBRl7d+7yRoxap7g7px87kkNeFsl9oySV
WgB+Ddn6oIO+mQRlFjPzxIWGhO0xT4IVAjSrI4dm6+hK8aQulERw2hLdrOLHYMpO
rQPUXLkSIRInogTYw665Kg2LGRyG86+Z+TraAzZQei2hBk/eWrtyMu6byixmIlQP
NG3/v1hECiq3zs5Pg97FRv7SVzc8creAv7GXKPJUagf2TCHinnwP+sruaJU28eqO
JvyyOamjeLX0JYmLcpLUeYFjXUgYlZhiybrH9kDmanXox6/K/qTLesPDJKvf/p5F
c4taoTQinQD18aWk8FeEG98EpCkR07mhMMFs5TmEyhBVLfHB0wyl93f/q8h1w+rm
f4BexecKtX15dfwRrwYPFYmDGNUjcjtiR7cscC77zE1KMhycwdmTeI2B3rbBREMt
Zhit1rpl9Ln4GADwc9Z4oSerWk9rR2VbhUgErv38DQtLUMAAIJfGywkTbMIZKQ9s
gtN4JTw/3siPRHlHAiOCl7sPUNUjc3/EhKHPPRzvLq2SgJpEeWod8dHOpnLSCjSc
6nZPxnP4w/mNUlOO6I15hMwHI9ZSL5ZHuBd/ZZaLx6Pyq9OT8HOKnWNvMt1zwjjU
82VeQ60Awdu9aNZQQWPGFNnSo0fBJN10BRyH7XENu8ts2mCaTmCIon/pjfN1XZgK
YGO4GLRWCXwrIxuV9Zer8sItPB+NUXp8eJ9PjfEgAeXLh20goDNjEQQFxdfP1w/u
Ix4zGRcr1l0UEUutdj2ALnRsa2I+n5+lusCsPOsEryhDuGnxxBXwsL5/tYgnWvC5
`protect END_PROTECTED
