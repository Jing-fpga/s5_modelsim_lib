`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j9xBTSiU1LBdQ0gVwqqLWuSNcOmb1dRcshMxyUEclrI1e/rKGVd2ouhaaGhXnPql
oy9rme3W8cm+id72w3uSvwbpl+9Aa1V+DSNqgMfJLq1RKn8NmP2NFZ4Gu5DrwJ7N
IO0ywjAO8qpg/XhoIGRJWQgOGfGs3UPHpPSyU/gs1YMqhGB3G+Gdw+u6xESqvnxt
4HZ1ymrIaZRQF28hobv9yF06oqWlq+sEXlgrT8QfrUp9H+9OG8Oxw625o/uOAFc6
mn896wXeUbAHBW7BSm+LLRZEB8TbA/uCpm+wBE6w9/J+6B7y65k8Dqbftq0hbbNM
zofGBv5CxJIb6iah2cmeEyvz4KBZ+tBcsldM70c6fGZbpEeSBfyvdeHA0N7TDpE5
nCZFfEuN3WiBhQomsMDneM90xZlesXq6GwVWpkbp4ZWbWqfp12TCZVtYfsvF3aPu
TBvSgcXHiaSoUWeWXR1SEy2yFseibWcyzU9XS/ydB0PBtRjdReZTFMpIWG0loJpR
XeRQysyQS3+2aAaD5HOpAu57rVkafab236Tuuui9+Nz5ploOlDzBhmUwEA9ctQVL
7zU57bHZ9huWaB5z+aOIecBBvQXmMTGhM8J/OSSyO9MFPOloclsIXebF3wetgDp2
ulCBmh2p9roD0HtONET3prV1H0WkCuEylzLLH7pi4KRKm46h9OR2kc3B2L6sv4GU
wa68YWZWkoifi0LnS59jgwxRcuy7SCH3rDA3ThlsRg9EX/TTVJCtK7oFh+K224kh
kR9dzMJcWr/CqX1r4o5oYLU6AN3coM+lIIBJlupneAEuaS4H5JSYBNfR2e981k0K
p5FEzeE3CcFS0om/tsnh2MdGQ2JPWzWZu9FPLoPn8PBMtgMRUNI0I5uLYuG0+4gD
efNPKWAPKvUNIQrr/z0sstLwcYkr29G6VBTl7YjzukKJo6WksTgUzD35knbYE5pr
xt8sVJ8BSoew09wPJ32ttYQfn8lo2Txzyz7jWhTXdRiYffm4Hgh+nTo1mZR1Xcaw
R9awZ7AZ4qOeOvefs+0Ez3WNQds33FWoTCP4OIxcb739BJCWWZX2nzOuwZy6q1xK
hD+xgtwxPNbuY2w2SE0p674ZDv3mMzJMd+Vxhlr+lyAvJLQRdOn+VBFrt4oVou6d
+o6w4CY72KRuOW3AVNrHgiQryyrHSuKyHpi+Uon4lvih1+1qQwEVjXF/ZbclL6gv
Fu9GC+qffMD9yv/kRGwmCrvwP4R7FE9QT+RrEI7y+bPaCqWib8lb9zuyJto6ganH
4bSjb0W7X+/uzxu4zCHKuCqPsvDKx4FocOpRDTgrXlqmuxPGN+6GQIJgX+7lMAem
dBeWm23ZLFFY88IThoVit0IQq2PRX8sctAucy5R3NeF9psBE6xiGfw7O7qAamejf
0y/psIQUCsU13UcD1m4NgZRJungfJmJ8wUe+bG2+zuOm8CDdIyozDY+0fAfQMayV
B/n+lwX+8u1lIB9PQY1V5w==
`protect END_PROTECTED
