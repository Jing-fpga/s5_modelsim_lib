`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b5pmOXrh2FdaSLRyJ+DcImuuLLg7LOS/JiZfXoKMwwHSghOXXozccaosN6n9lZ4A
mk6375EjL4hZ2Ez1Z4/6pnJGSc7F42RKzw+7TbFp5G7vobGiDOXOqoM7JrV4WShK
5nPuw4gzROt6njv7ePjj6EMDV3eOJv+Txk9Ebsy+jqvDXy75QkcDCTMU+W9CSY/z
Q/Qve40Hgn2mxHzjW4BCLjrsM7XunUXb/M1O96KPCim73hwrtwE1pGsZMftuSMi/
JuRen8hLPdszR0ODUw5yl9KxSg7d5KtNwl4DPrnjbUQ1j59cHmByZnhpotExUlyU
xtNWZB2tWhU4vG8uB1l8HHqJSaPSshRUyY2qwnXFrKG19v0zJ3YXKFfk5I46W90s
2HDmrNX3iqZgUVqMHVHNmnUuJElniKbx/6hBy2jeW3fGtcn4fOLbFAkFnL1XE/E9
lcwlOY9Nr0eYaQzS1Wwlk6K9fkeoMRxnafsby2Hss/+xe+6mcPDwoHxqkThSaDuE
5DRWSR0EjP5us2Jc86fd3nnfmVKGRToAm2R7PNg1GoYzPTW8ot4vneNI2VGufWf4
NwoE/g106MMi6S7yrGravxDcDNRI0iDYgTGbMlZX9mE9WTSKEdc/aXxEkMogwQQT
av0n3uIlf/lR72xL+cRusivB/Z/Hi2l1iVLrVO34FG+PtVzWut3xr0K9S0p7WSv5
WqxOLa80nEh+k6aOx7HKH6FeLmJ6oNp5O+/q2lieqbeUYKjVsih/R6rAFykz3/pB
ScdBqUTNJ3z//yPBmOOXStCRHrK4DULXRE5tltvP1MdWbLFnM7c4yhgWui0gvmop
ZApFpyFGtZoiOICJIDHTDsoJTT91UkjqMejdUdmN/rSJoaz+a54fs3z27WdfS+sg
GJexfXwGq3P+mWlfm1BgcFpWX/tuYEBOZ8fSQeOzWYQGEdQAij1bPyPe6QbtcHk0
7Eq64m57R/Z6Y4l3R8tcVsgWJTbder22i5GnzcgqyuDdQXwz7jXiPhE508SiPC6P
yHQv5J+UNvnGF+aL63x3QFcvJPtkavF6NHzw6oe7Xx0PyBJ3+6uBofTRqiXMD8C1
F7ha2SV9elytaCQ5yKz+sqMPHf11DN7gHVC8fYyv/CT4OEPdIbBz/ipsrS84ru4S
5UVuJ/VJn1nijuybWOqPew3JWUbza/fJmOHGFEzsw7E2w+VjjNK3X4WFGQNN3BY7
q3NBvcdI/Rm+3WhRAc4+AQeU77Do0Rv+27v6HHoGDSELQzeA04MLxpjPWIlyetoF
axpkDvio0917Yd6F3vKtQBH+PLmPRDZ2nOulSi43loET3VpQH/MNKrbelKIkakVm
wZcpv7E1BDTs1t2WLh0XgbhTK0NGPyHKz2wvRwhPfb9L2T93BPiuZuEf7vLR1R2W
v/4j1VUjARZEMRlCg/HNzYpod/h7p0qo6ogArOfNiqakkH/bnJWljtBkF+AxyjwH
FT3uIS/tJF+UOaZvj58m/x4RwrXZ3RpeoF4xZ3ECyjHlwXbov0rsol/zfwHyPOtn
OHMi2oA1uph05O0AmT7VuGlVwfT6rzkpFbNkdsmNtD6pjXRKOgUC49R5VtKs3ZpW
3SewsBnpLn/7rvR8h5Zt8L6z7bvFz9zib71eWrt/T1YjOUfwkUiGkt5N+geCSznR
ibxaOqNxTtArlghWPEjmHcetta7G2rGiRQLAxh0aCbD06j4Y8bCIKuglrYOL0wsi
0ox2vTXWS14z7XXylxxJLHtQs8fBsL4WT4lFErmmEhcpWXumVwWoyO3ps+dwL/sK
MDrlLEftSuYG4Q/waeamsj0RBF5wUqj1M+3nhqEUw39h+KCCu41pFDX9A2OPq220
QZPPoX1bl4rNLa23o28Hx5HN07d/xfeIvQb5oUfXDWiJgdUGVg28d9lwAhblgQaW
ndPyzSdnzlB8UGPn7fOBgcZy+KkN8CARghR5SR1+SOSInCNiIy0hYQfNVojj2zLo
6kaBD7Yjr/7wr7G/E1/FBcBsPgKmZJ/BBl3LQR3/aw3+U4UYvLLiqYwHH047adH2
xEji8jGwUM2iUvhbckcH9aeWeLjBL8gUd2f6VIUGU49BuFtvNiR+t9U1EFDK5YGC
YOiqgn0PbZmLrgkA4XLlutJmMjsLvI1HN4kI5zWYfQAB1j7x3IIXnQmOMpv1NXfT
mP96jJjw7hWArL3Y43RanaplFhpUzbs8ydpsKRomzpp1HDZUTpvPXLfZkqoH15bg
CbVdjNp4srZ+LzVhVj6JWU7EQ/iUKW8XCLCTKczhBglch8trudZuOL/j59yvC1Jm
/VW1RAqo1d/zIQjfWjd5hEHaXI7TBdw3iDX0gEyXok+aXyLBm+uEwopstGFpGQEl
reaFYSyQU5nIZiFPyeGUnGvoRdBSs06FfG+Bjp0xGiMwdEGw2yc+2qzJrst30VoE
S4QQK13xtIQ7K+fNofVNVLKY9rzkvnnJjr9gDsJ+Egk=
`protect END_PROTECTED
