`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mdL89JMUGVDZnGYrIwOsNdgQVUXxCB1Kq0Acjisx/QRiUrx6042+mXtZ9GMqsKTD
pzH4BKLitfeE89pWCDmUkbHUEJByKNvb/wN1aVl2Q1beKtjF/cpBcBIEOtTeSmcX
5g/R+icRGLepBxKF4Eiz0UN2C/5qhAbRTkLWfCUyDWDV6qHMsof/93tQkGZ6mtgX
WCnwWJoyvs4+fVZ/MKb0VDk8H26j5SVa7c6nWLyjOgAPBoxBLdOZzeMU7j5LpJRr
sECwzUVOc/vIGvsBpH5GNiMVY8nmpK2f2RFF8jnnBpoPXlfvCSOynq+zrGKXrcnT
Wm1P4fybVnruK65h0YA3mhHXQjx7BdGjMu7XU2DsAhuyY8RYYl9gDiVV0Oh0p50V
onIrL7HNWOjohSnSRaNFPRhEb52InpMtwmGXZBD9sIW3+h3tJEPK5I8xHy0QrhY+
RUiB96/EL44luG48gmaeUgXNAFsJmXmjQjMOzUh9eSpJyy4zPU9P/a3VJzndUw8w
GNF2nF7obTZy0PTW7S57gBOVvh1lCNcHTsJ/skY+QJxn74NeT8aPgmLf98m3t/LA
NP2Q6LMxBvFKVv2xA9hyCPedvuNs6fsGzVSbM3cMJhkD9TGIMIeDYoSpG3WHBnI0
0JViFCVkZo+h++Uic5AFXJmxSiq1spisifhxn8/oH8nHU515xVOjEC+0iGm9exWe
Teb6xMN6k80JRKUe/Yp9mqBE/IzOklwoq3Jz6EJFWIDqncl40Iw0zNgiJCH8l4VI
3sYrccQ7ZzCMY5oMvJK9fauDXb/EvRfU4Oots6/BE9+eva53w60COdvzVf5HTs3L
RPwxMy8HEohQQo78FmcjBGi4FsKlP/a/T85LYuffsHo9RXhkFZQA2VP870tUYLvn
GZ9jvvncjbiA600kHZ3t2Jj0vXp1fROZBWhnoYs+o+vGMPYc1wgYAHomyOqTu5Ov
LL8EczxD6rPmKqBe1opE/3CNi6n95WRz2rOt+vrpZZDcngtZOJwqe+iAHQYJk3Wn
B0JJQ34JOcWxov04cWj+1//vmxeskyr4kSYcvkNLw1v5GR1eiZg2uFfiu9lhtL2P
Gt+JCyN7ST11A7aVtc+WxlQXF9IgVA8b45kwYQct/iK0FI28f+Yk5jzxruA9wYqi
1BL8+2nVl3sA7laEatSyeXfDAg5g7DxAZKQ9KPLU5TCa4gAb9M/PoT4fJPpW+LLg
cNZQ/F9uYHMNIjC6uCULyxOosAb4k5xsX00WdYlI7MAO8fJTLyR52QoNMSpWMDOa
g4KQkqSv/LRqfbYFLpT+Qo/20FK0Fq0XPy+5KNl/aqAl52aGJn1l3e03cYWWh6uK
7It/4/TnM//SyDZxDFxLHhRTI9mQzuJik2mtl9W9XnLFF32F/na4id+CnVn/0sxZ
xNg7gjo0PTarqsJoFfgmsR9fCIC9xxc0/d3Zay9ZVQ3+C3PnjMy+na/CKhtT0j0Q
iC1WdVkAeQDkfPxOPRpPKmqhg1zcOasvWMAmEIMJewtr6oy8NLJ3RZvhcTkRO5SE
nb0r58BzrXsfieEqghwPQV8v97kKB/GcqsWwEH5FuHzYWgOErx7xXtdUHJn2y373
yqBzCL1HS2o5FiV0QhwgMiDSw1uLl/HBCT1Ru01sZO0Ruzt1cadCi4XLsZ7SWzdE
I6udeiIh8iT8rH2S9kaAVWHvCrjGlNFwKv9RXNwCS1V5dyVcYa0duPSbQkvHw3oP
cnNB0vpUp158M+PU2IvJSvxYHF/SQNMuOakyI6MUp5ZHy9OGf3r+U+YGpGySR5VX
w/UMca8YpfYJWS8RsqN2TNM7AohogNCc5oY2oS6JQNKOo38dYJCcUkUqyJLGiRsD
bHECTKLoG42oQo8UKZCzKW0+6LxUVC+WmU7aZ+eC71xjT5NSnYCq4rIvDVaEOU6u
QXwIeTmbsBHQZ1ydHrY75fNHDbf3LxdfT6iYDh061g6vCCz3DyNFBuFXw+APhjuA
WIbxNiuMlVqWSoirRCtL8OUUXb2f1KYlo5EIgKG7DLfiy19ZaedYVZmUw7sQkfyR
0Ddt2MVhXT6nC7qpLRohXHCTqxlbWrfBgZIK3Ntf+IaV2BxaATA4NfplZCBBwbqB
Rsbc82LINV9d0v9rghhL9mZozpRw3JXHswLOgaQfWjEfjA75+0bdBwNODb1iO7JI
AhoBENYPOudYmuou+Vks4jBnY9mqSdPcDoj/f2TLpuNjvdCWjcFFRU9g3tsnIhWp
KrkKjNybaQv8u2FejJIvZ5fQy3j0eyPM8+PBn1G8LH6cC4fbCw5Fm9emL8RjvA2F
cOlnkEBH7G/Eawtu5NoPWbq7OpX3Sr+HClQYrk6yhZ+3dem5hmoj9rADpWI/NuPL
W4zjHQqmzVKTHWdr6zT7j2g3bJx3fIRCxV1kV9YBph2LqYFgHm42F8BJsZAAKcAm
22mngxjTSIiwpELl4nQiM1GO0VogmAhkcRpAwrWiNNKi2gfDty3dO2jj07faHAJN
zt+HBXQa3pfVzkt5vv8cA8+IIENDp/s3gaKHFDljU+eTiGI5brwsqGZN7yf+6V0I
qBSj+Dj088xGmYvE4ummqg9b3i2iIf/HqA1omkezdSABIxnvWBhgJiKPZdk0kBO6
s+6FeooHoY7mYUkiAPkfEgilS1uwttnXHhcL7SqO/FOF8VIjJgB8HpMg4yUUEMsA
0Yt63A6Fr/jSqlLTPfeHL1og91KN0rL7zbIg5w/3Fk7ug2USZiLI4PCNHgen1LR+
zb0gAQkQVL+baVGTJmPnp1Ov1dbGwdFUUJLM09Qcw/smQr/vVciYQapyIq0T91V7
Ha15xJwZkHxPaaRfmX0eZ/pn8I0PJqFnUabOYbPGwS3CM+39Eo13W4d8j42LytDZ
9k3gCZMYSdNOkCCq7LXX3jNDEy2KyNmScPyyp8IQ+HzYfqhvm/g6ls19k1cZQ+Xk
BZ0g4yEQg8X4PEN8G3SMRLSZX8LPn9r4NM6wZjrbOI4e3wPcLc49tLTGkHK5Coot
BHQSgfqjr5WjD1+7vdCHtGyTkRjiyleI6ErznN8rph+dtyipI0nScvPCKDXJXwkC
0vU5O0RVFQBrLlsWqeuWJBDlNSnOOlI9kaR48MRXZomgArf6D5jSPogjoSRoBmmN
k/ZvYS4vmNh/HZUQwfwcbu2dEXbdX+5yIF9KCZp0eC9sgPE5qSM5pxRYkjsp45gO
dxJLLr7Y+/xOhIKpsX7f+RjEfhh5vSzsH0z/WirVyoOTfHMR26N5lrP8pNg4J6TY
b3MhSvwRo3drA8pPZZy0AKPdcxAqNmpLW5TDJTTl1qrwjdFK4wohWUER/zeDBPtB
cSypkIQB6CyFbn8+q+zNb2vJc7xd0C7SFfYHEjFMeC94UbTkw1a+NhVO6A6PHtSa
cjtOnYKp7Sm8/mnemozJUI5wD7pq7KLFzN3IZLddZAQZh4ezyZD+qrdNdn54tfyB
eBv7EdftXzppg6O04F+N2i8o3SDvb3Zu+5NZ9ghUNlmAp9s+377UW2EB2o9UkbNs
dXQZqY+nDngwGdUqx4NysprsTresUPX/1x9huXs65Doj9NHDySiSqm74Dhj+iNqn
t6UtoWMJ+uE+uMWbXLFKe+ARYxG++IURRd5hJ3gAS6uFdo40/jFuT0XFofauz+f/
hqli5QOhXQujgZiw0cyEDijrnSeE0sLZCmDhWE718UexzZtp53pJzxr7HsWZjsLJ
TL9i/NEQMejw8pltWzhX9ovliXWgD7Q9pvQsuOgLwtBD+YRIRZlk7F//WGcgH55Y
cVl7LX6bze1PN2IVZtm+YdHasYeI7Zqz6dPNGfMAmd6ZqhpmFA2oVUMgGguN09FA
2LTukHNYATDWlGRe7oart4qJyxGd/y1Y02lON8EiA9l1uLmeJBysAILh8icYEhmE
Ic9xqv5Z1eZ/GOeblgYNbfDDuSWLGs1D0WucLQLLcorniYiPSJURqV2qMgcZV99W
hPL5vdlbj1a6kpCsCJHLnQJYAg91pc7wdwf6lIJDCd3YzCUzIdFz7rugq5xMj7bM
JGpMLBYfKZZ1lwjSdG0hTT7yOjyFJcep0Vup9p75iqJwZMI0DBHrWkAyhxmua08v
sP86IC28PH8EpFv1TweZrR0i9kNfnoFbd/wM94NaUzDOGjy4WoiO4Fm9En8xTpfy
juzg3N0LBN9mo+2bQYwvdg==
`protect END_PROTECTED
