`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9m2MGsoFVhBENBOEziPH6hM8VSHqw/0jfNWU0WtV2bnDQ19zWxlOasOfow7hdYVP
PVICONbPHQZwVqy9K9AEKLVpjRvxC7tFeLHMRH+NMcxX+ytpkIuQUT9PwkcAk+IZ
wXpOmBU+r9t8L5qBLg3eSSU5bKNrFfi54OvwU8q1khynwGWaS8lgKQD2gH/ktoYv
kSOYDCns7PuTx/pE4T/cwYV+rN4cLzZ98KWWmf4toKmfQ0RA4dNBaJB8C7VfO6nZ
4Pc/XG8TD4VYoaORDt/cHIFfPQPIvHuIGUV7bYOH707+XLhEPXGRJHfTpx4uPnvo
MlQeeZk+7PuICr97bLOS+yLuwYf+LMsJEr4+oEYujhzaTWRwvCvQCwglc6uRFM9S
uFNKN8LkdLQ5QKjXR4Og0xuEWiqX3TvG8cYPxeEktZrDdhaZlXbwz3Y67PKvnqWy
iIxjoDFY2U5CPraL/sjMw+/Qi8Z/Xqon85qNuakD3Qz53dKCybVc6UH81IouddQZ
V4ioE2W5YgFy/vHV1vczqpB5ORefqVaQ1KtPka5cUo+0yEqSeWqJIAb/I3Or/2wG
5XGUB2lvg1taRZ8j3YS82sy1iDulHYGwGHXpQz8fD11ZLYkfXkIwcJ9huXmJQPrV
X3NFsbpmXmH7d/DurV+kwV5/Eh31Cnn7nzjUGkz1FT7A+xiflHg46yojlflETuVa
Pl+pG1H8CjTcB0yj+CQzyP8ZlbrQWQ7rGVF6PMBs2v5AbgKpAH5ut1uQ5WtOnubo
t/j8QPiosKfoZtRPlhYF6znFEQmYg8qc/BhXGvV2dNaexEktk+QSAqlZTOy2+90g
3eZQRj6vR5ui7mFbjBtk5BR3FGwRuLamBEOkdn2fMQU=
`protect END_PROTECTED
