`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DnjP16Gt2aqbdvARGIuyYLp4+GwC44FeuOQjnJEWz3FZLZlHNnEFSHnE4fTOGkvf
p5WeUgoJGxFMKKh/oSuvb/F1uslcXI39k6hmYr1JCj5ujEPCAMqQfEbpuun4xjht
zGFfMqsGQQAuh/UDHhBHY0Qc6EvifYw5GkqOHS9kJTP9THeg3L4D8Z76WyH1qkxk
TGBZEhrqIV+9WNJ/B/cu2PtCXOiKA4QEDFKd9dRTPCvoHVcGoL1kObCCNxRinTGV
keABBqCXhrJXoz/oQahaFOCt5pqqAXAjpWoBn+M2tiE996A7faWXx5mHmj7aBI0J
VBFMcfv05JIb9Hqyt0yOg82IGGphEZ+ExRWu7FvbWVCdp+allkz1Q/W6OC31aCzb
aIBgqpyt9SMWRwco9a+bk6moY06cIt9NRlWlT19BJs2QU3xHPi43sYW5hYQsfg3A
bYppVabCh4vwrIYtGAMRfAjaD1mkrOCq8IpyYCaVYTTeEb9/BYThaaoBPtfEqtZn
Zet6nOkvbwBLigeYJ6WbuwxYXkuAM6OyIygdNTuEq2hs+C89+LhBElQtdgy5IBBU
IGn/RVB1B0gB8xKzU6P+PpwE+cBwhH87S7Md4pcl1cU1Opcodpr0d32J7xTVbRPl
6csWPkmbSOMjviH4OkIzCXygnGdfWCGYYPk4RMO/D44Qce3F7IUnZ9sqO72PlR0y
LLpnF6P7HXk/31FDtD5Dyaxxj4xSNr6oCE4MvVib8GOhsO5GiXPz8ZQzJStbtoTF
3CB/211R7FzyuO+w63rb5eaOT7Rq6gofJuDfbYfljd8Vkq3TjwQfyx/pDxPwOzOb
m2HjMToW2aHx/ulmrfEb8/N6n1sJaZvb7QJb5TqL3lyzGm99627w2ggmt9vDsY2x
sxyXu+e2UC+m6w7OqPR17t5exSVNF6bHkGHN07A9nSL+qFnPD/u34bBIoYRvmG0G
HSa07PR7nKy/2UPVf2vBmvWB6BBHpnnKZzoycn8CsTFnaSsG45o/1z0FalV5Y639
3V5odAUxsTdyVRiujD/brJCzUZhoL55x/BGmfGwqPmmynCFcjXzcvRUhVSfCk7Xn
L4YGBAWd7Vs3QH3DLhr33crfpM5dw9u57rOq5jxKj007S/L0RHaFo9jxnvrtWy19
WyxKBp0fvs0dyCYtTXx4Jw3kf1LhhTpxEVDwBJGxCQ5S8B1DljEds5an824hDJxP
9l7ORPhR7llW8y/YCjL8YLbYm55fwAgim/sojsGS585ejt+39Qfj+77yhIO02hEK
Axb/P4be1dF2/HbW5qzTF3xyQoIE84MZCh8refuzaE2q6lU9OFqVeWsNUZxbUKEg
PfRkQI/2nAT2Pnr2yMKZkkmguTnXyixK56KimfXuSAJNxdShAQg+S4vyrnGa0/np
XZ37ZIzITB0YiQXOzClkgl6i/UoOujst7Ie3wPJxRa6DImBk15jkuOzSnonMOIT3
1VFl0Mg5HY+lEbtIozr/OdDwWq+TLaaoh+HAXfa1pE8lq2bE02D/HjlDGlVtPu3q
sPf4ouQcuXzNPtgBHbha7piHVKRDBjek3LjW1GO7ENeVWpFyjOhaS3a5NFDgsfBl
jnJ85aTQ/u1upVVsI42pkx4PyhdR2L73VAEuFIqZIqsra0xFKrwdvKYRDkF15D9k
HoumLm3ppzTzOEjqTiSHjOFiXJCjE9zz+nqd47gvOLiPv3bpU/f6WeRlVaotmVrV
lCBa7h0N4axzHXKmNcaJhytvyux8WNCpKtclEq8VrptP5lMl6DZdb6OLnEgm7+oR
pA/qoG15DL1ftpIT5rbGsN+kA26L68XbXAsXBW7oIB1pNzGMlkgnhbFdV1O+uzyd
MeGT00bxfP35EB1kPzJ89D9CNkB2e2w8hvbVr+1c/w7dkPWzUjhrQGoWjubBj8fd
akvhTa1nsqpftf+XcJi9BCIJO35IiKz2sxdzPKMpcqrBarp+oxO9qDfa+GoQJinR
+3ULPmnE+QcfPL0/Se9/ud46ilGIoUQ4Pzcc/ZWLJA/th/4OpzoC1CC8DRvtIlNx
CQGSG2T6joJwxtemhNSZhqJUpP9yEn/3nlgwXETJRHqC6nwJzf0hR4fWbHhwMz7Q
SEPdFm56s/iMg3BAlv1BwKoQsuCuPZuOCtFASicGVc62/CC27Jl+fnfTPXiu2mtk
1UWDcVfaGu62bzGVNHLf+5EQLpUS9bJAKrDCC77qDZ1y1fIvMF7UQfMArP3t9/8s
jMsPTB5vMOtp6jRIV5mnHOijel9w9nJ+NtVykoY0MpslUKoIldcL3zbvxq7ln5EF
gTbzBix2EtrYgqgxRJZj6p9FTwgsqm93bfw9H7PizUp4le+/HPc8hdy4iXoCyfrb
8nktMkXi5TJljUEUPLfh5QWAs9GhzxtGBjjodv40JyyVl5YwKUy8hRPAJqrBD8HZ
2VUZxgvWnTZz4pkzm+IrT2CX7/Y/VSy7XokTAPmNcU0TmT6g/SiGzC6Rrzx4OGUU
AOd9tgbkZpUCgOpGfLAySsW5ncGn9DzwzJea9UL19XdcmJaumcxzPSHS9axGvA3U
Pt/L00rpyAkk1nGVdoNCPsDkmXmJztFZ1JDtLLVOOd1KdAvJ7isBl9yDBu45s917
SAeo2B92jqkNzS3hX5Rck7mec6cBdiww2fM0C8X6XLTsg89VRji8ZL3LdXs48nuu
3OLGlbPlqqpK9i16tBoYG9REclrKU5WdOUR/4+Ppfq5YGs83ZnMXv8kKfhcTxqPk
joBuGGxKp+LRVsKONB8sAq40FuU288DH0RofgtLVZlfw8mQT3vuJvcWvhpqoEWVi
yh/vV0OF/y3+PEy/SzCy3eHjcY/+z3p/BH9Wjc0lDQNGF6Hw0Srd9ptCFgOxPfVP
7LyLzBe44oj02ePqeuWdpwaLgaRhstWqYTXwwGAaNlpgOfqoyl2l4N8BdPbyLWfY
CG00q1jUyKB6BEC8cV1Rz6GhOWc5Vyx43BdAAl1Q6o8ga8HA5GApXKKxn5BpPt5Z
X9opga1jLFWbPUfQrrP20Nh8Rk5zotVvZCtr3JdKm5CX8EXIuuSX7E9ftnbWSqFx
S5XnA+ejyjA40LKvLV2IEP7eEBCYMP6T3RcnwKeSdrcjgEbRPn3xLtH6xruY46OR
ZPXwbEW/+yBeP1SeTB94A82llCB4W676Yp4ysMJtI/9hBUncN0g6vww1StWIToVk
YbEU3XAuNeBciIcEiQGeJsmOXAIFmTXZS/KUt+gItIu5RA+xM2onnF+RKfoD/g2d
qEG3iTPxAU1VA/xJr8OLJY/tJyvUdBWSocwMwkat7yv/WFZjbDqY9iwF7bQ4QVWD
59eYdGXqjJkbT/N4ap/J/n7DQCkaa74QxbDga/sV7A5pc62FAwkn6ZcK8t36ewNU
oYqq8nWoxS9M4VDnjJPX8xwz5Y/mJSGrcLxVS20xhyP7zHYiKMWG8mOxYguM4F+f
y2kd1v3e9OzlzW7Z5nxLLvtXTMccIwxXzZpuZK6opFYAt8Rx/Zt8lx4Wtq1HxSAp
U9ioRea7JPZ3A61dZS6j1y0dJDBVZnNu2YsSkPUzk3SkN56nFLd+JDBgmBODsDq6
IFKUopH7KwDgcQ15YT5HiGmh/kKdynU7kCY7GKd5G9HIGhlOOk/KaDM88r0EV2vV
YlQ23lMBDb01P75YXlTDBur9546PtteKzrhCFgmjz1nRJ9VD1mp0O/sk9kWEhI6r
PiR8ItuhMW8fv3/eWPzdQF1cBr7llIaauO+Ql3AClDd14sfaS4cFe74eIbI07pAO
GULWTt6r62zuuZVetbUKykuLJmK+71/loV3F+RQGqlcnRUmU4UfMpNHuIwjPbJj1
wIrVH/pR2PjbXcF6Y83Y4IRX4a97K63XSeLYXxYNirbsx7NmVsof0PduZoFKUmKd
jJOjCKpO3ZyGrqEhbJ1PX5hqj0luT0krWPI2CjPZlC0P6smuVoSfZek668l45Y6f
nNDEE0xUtqbUvBKgNicyor2SawI/ig5iCB9x0/KUlbCFA9jL9dl92SSGD+AOd0SW
+vnrFg1Jps2laO/drdTOe17CtkWDAU0gEw9DcGZAYfKeqHgwch6p0ICQN8ZVstRc
dbUAX0XY/ZnV21IcUcn39hINIHBN4QtdCZkQLQ1skO74gGuPsSEX3xl3OSi0kfQH
bFPVJ6uyixY9195Z0ZAF/NUDcB5eCaPQ4zZIC5jp6AFJpjHqqwD2HnHuhJZa4CyF
/6as5dvYeaNdfggxtrpIif51Blw8NceLDIA5vdPVsWSX5wbQrMkbqT2WxWQA/pKJ
leZKDi6tew/7QEeifwY+Z8VUQLfd7nCnM9jPWoYjsGyz/plwYdRMIYTCXUyQZf4O
Z3N8NxiikfeR6MGYv1OBLP2N0NgEm6BD5LJK2mWgaHSAF/9X0tpoPvnE2qbkSFXA
GFk1OuSRDjwQw7K0DTzGhOOfQUi5U+CzmZxAaITomy14oYfRLWBtaZ/XK9xU9qa4
yl9BrIH4KGX06wnWGjoN8iTYeQHU8eFzLZ4Ibcm8LPubJqZpHLLOGGHQ0NG84gNy
D0aOb8cxkhH3xjKm9zrhRFWIPIXi8ZLP4m6pzYdMOozDoD2mrsAQh5uOvvE4XrMG
UMK+hUiR3YnikhzDGPxHe+03/y0v5odALAsCdZdhRlH4r8PqLrOHjChEv8L4MKV1
Zg55O9I1ww/QiD81r8da8rffk1DSyQPMMzB+rJpGuhkgUYu14dcGlPsBQ06Avbft
QKvTwR7BZK706ltvrvtPXI2u9cuSkpDltWwslu0pqHVKC33W177fApBak2883Fml
bXTNsehbU+vXGhQNG7U6qRQgkR2nEhYQRzUCrRg6mMeu3CY3CMJD1qxt42wadjqd
CPTlIW/BlviIBbfLj1dPRfGpQsZJebjtVrgVHjw2Q+8S109zgDMLZe8UxY2QXFVx
OExiaoqvbQEjYuBVmIkLeKnDEvvD6LfRTebyIagoDtTbE9WRm9D3+WQLVCTPzhHv
rfWHrtcNsCSMUBoVY81/kYG2HKM1eWhL46F8sozEQHms0LtPka0uD8xNVUzj2EmD
uiVpYBtZGKFYOL76LxoEKhXgAguhGaKoP/3p7GjOQhIL+uZVbZNabZmVyxfqpykK
0jmJ49U8K9Q55ykPEX2LNkCZcxCj76RMNOyQSKcL9X9akLZ2DpPD4M1wUcEwEfkY
kLtJObwIPVYeLrJ+9BwgRc8bgVay/nQPlD+vd8OtdGdLTZB48bXJAMVtCLFNuClk
4opdzAWU9LHB+CByVQxbp8VWxDiVt20YEWUAxpfmkKS7cavsmEHcrZjUCrUzsXh9
N+haFOdKVteghBbS7esw3j5xzsyk4O1HfOQJn3uqLWCRXaD/ZnqY6pkRXfL2ZZbf
ehgq/avHNme+12h1QTWLbo8jxBfYLCvbJUsUhah6JDQoxjHAgMltG90VXks09WJf
kF1LCN1TAyd7BF1g94L+Sl67mprLxVnDdOLrzyciR8VltWCxRAykDd1dvsH5BqWY
RSwc90+g+qWcI4jW/irgzaKECvXQ9iPEj7XqQnOtDBijvXkdzNfXnsMKi1djcbB3
/RL4lZPKSYsqQFXGkpwL7A1bPY1EEQZ1Dtf51/n5ZRcSXba1KRPxZ+slC86l+kGB
W4Je2fixf6WC3ael+P1hSjmokLi7e5CAnOA+lK9dhOHWX/Weg3SDcXCPWCntBX/P
5VJJXMyZzy7IYpuJ300ggkX6vu2MOffY2QSEdX4jMvgu+qi6+6jn5wZLeM9FV52w
QSqcRGmLj3Z0Es+wATqfXqpUZ1yD8EziZX1QepLvi29grjgutCD6+iA+EHAZJQh+
gCkDSBGaal1PLd+J2xY/cSe3bEu65k+bTo70WNA1qO4rks5TfM3v5pk6gOG4fnlu
AYaHWHLSlAczD6nzegvC6ipX78P2Qw4cRkjR7kXBANwvTbZylAtKBqYJE28OBF1z
DjEqZnJydnfMdjKxrwLAZLrbWu/KjTGz3hnzivoIN0YlNUHLVRvqCiP8dO1/9Hkj
fh/HoyQZXTGX2AUaKhT7SJWU4GC7ux1X01T50aLMLc6n0Lj6I89c5N3ULOg0W+QM
TBqJTAN3SGerA8XciXa+lc2x6Aw93U3iS5qYqh/7y43MiQPIXzDENQpouIFrWg5Q
XUen0BNehptXl6880rr6alUlyW0brS3ycTLTkmqGUTFh3j/NVTQ2kyl1j7K8FgcC
L/9708AzNvDnN7Cyc7zo25jW2HJN5NtAyavqz5L4DkfDMPpRn3RenJOlB6SVT6dA
H/CixiIdGXQRBdm1uzQL86o6A/qb0bTnQVmDhYjIG1V8C4JciiibJSgQdN59D0iF
2r+OfSpfSV2Wui4gBPAacQcnLYMlvCOhNgadRq6L3mvqA+8Lb5JHgPAwnKkFOZJd
85k+s53Oa1YQYZ31t33nFDpX/QWO+YO3QZ7Q84lEhbGqAP3qMainerQBEVexumNV
4x+nWyOMn2XheweVTo2nRufkRFhxQ7FJK2Xhrs4tg/55OLaedF1fJtYVIywVkXNO
YNnp0YyLToRyVhEvbhJNDGWYOE27LvQ6byDNCykX093IQ5ySEiScAC8KQWwZqR2x
foit/5dH5WLQg3SlTBKfjPLPu77PvfrYFGWoBf95gHjuZSCT5ffP24limfyRaVZo
rXiWhMLQVc4jzlVwciBCo4w0mf5D11ckkLg2L02GPsLRKuGkL2lYauNWNzqA0u6O
3E+bMGrS7zSwfe4iPm3SChLStq2yCkBRsqNjP/U2XthEhfVCCUxI42F9bfQuDvsl
QJMY4s/IlIwll5ozQi03FsTRf4rdyXm+G1/sasM/qCnPJJagVLT/QeFjKZEGm/lv
vT/DwLU/VMcffcf6PKEr39+LkB7PP+mdueTMO2R48EDqCBA9Os6RfU7YrNh5EI/N
pt7uhFaNK+gbps9NO1DZV8ZMdIqdieiyYBhj0sO+kY1vIA9MC9klmOaNRHpNZPHu
NN1FqNnxUui6w3YRLHaGUPeShxy8UGmdjoTKBMcB7uu0UIbPUdHyYAMkAAhG0zjZ
f3TKMVKjRlF2UCEcmNNNBY+BsPnJxj70cSywRthKijA+NHmyaYFUNEmcPUl9qSWZ
xss/zs6g+Kh66zC1V2EtYib6fcJkUY3/TkUOas171cZCfRyEstCabjwqgtotAPp2
FfLVsHxzwPIdIMaG4sq0YCoOAFI2ZL9ZAUv12iietAsut3S+4usrfsj8lHuctNQM
7qPkOUcaD2oYFRoBAmRO8skhJ0C9bDg29Roq3xY6NvPwS6lwOO0AKgetw72vSQN3
niWLfD1Q5opm6iZVrDqqA/p/2N4HfVUML59cxUaaZSERDqYqUZUpk1V1NsPAe/Ki
BXb5H/taeSoAgdE5lbnYOrNAP9HWTITvCiQcWqFS8Lbj/yaxm+iuCObqc3wU9GEQ
OOxuOAoTk1q3tSlWaCvyX9Pqf9O3coyu2xL2XkkZXDC20kn0n2v4OleIZ/0w5Uaj
Xl1vvt7uXLUtXSFNE074PmJQCh20wM6q9adhEZ09uDwBJOwl8KfJHPWxUIQQFA/i
Ipq/64TjpAngBohIx++jBeV5laVgJ2s+NKf0nVMzKx9xju+Eb4uCivTmG10KssMJ
pxmafJItXJTGndMbMAHkbkxPNnQDz63vB2ssksuMizTm70OK4QNncdmgMS6n6fdA
NxtMWcX2V7UNrpXS1QJPbyslu3x8e4WgdYUHumzQn0L/SMsFsbF5YNcRVX5GgnxV
DXxQJm2VK3mmDPO2wTELtdOoQDpXI/8h0yKcz4kn/lCE/4fpDdfcCkfgHaXF7+nE
2lqorw6v5UCf/ZdNjvOrk1/vHkZPbOg3ZGCm3zM3SMJlJioloUEUjPz2hz3D+KyT
rvpaB5ARgQaaXak+zldgaCdx+hNe/LwjWRXXy/+G2+TcH/Iuimwo/I+rJ1gafLWc
z3W1H2oi/0HQ45iDYVc9hQi31GwWPpDSfjLm6fNqvFlU9Xu8jsDrckZyKQUnWrSm
RD6rc2uyDhKYXzzedLYOJJD5/sqYGn8X+ZdT+wDcmIVcCjqfm3OfGa64KJhtuZLL
gOm4L+GWkOjd24iq12nqgb0kjb8/JFHVKmWkCtb4oGhTxRoupDPvwS/QWvQNR2rD
YHtT6enf0N0zs6Q7WD2KGgEIUkETMrxcgemQIQfMJkCcvUAyX3t7vrozrvXeHxt+
X/nIwPnK7UQVIXrtMKz0tFDHBV+R1X9t8cc2oarhBUUmFZPw8+G1FjiLjNTgU5hF
R4HPvazRWbGuiJdorbm3CMYyTXOh5Arpdrk7pcJkS6JiNkfYtFQNJBB65CBxpS1g
5X8yY1aC2A4z1/lGKy0rH5syZV/uYaDyqiczG212Ej2ZRbULtdN3fKGrvxbIa6C8
jiNRdWiVJGQ5uPHC7se/UnbIHm/KhHFUcdgVKXGco7MEEw7228uLASw/s3HVfPpU
uFGcMJRM8u9ec6CvNHfYbwOb9At0Y75e8RxMTR2xjBuL0CAngSp04qsMZkgUP678
GoYMHT8ZPOgPmazMTYJeivFPmrNAvzY6wrr5qUMHhI0pKCE+DDuRPTKCiN46Uf6G
1WqG+2PFsK5JRdC/yhi7dOZ1F3suWKQt7Bv7ytJh6tPlflDk397KRzsHKf5C8BGH
CcmFbq+SiNV3lftXkZBXx8DOhxCovZd+BNunI2zwA2ZzAVYZGqKMfETDh1kbnmSv
AgD9AUCDYnCffPQ7ASosT9GrfmDGmg1kHh8Y797WRrjeCig0byNNv6o7makj1l5B
Q+gJi1dlfCVs01dQeFGX8fZZ3R6W/5BphoOSXBp/ADR+k6BgkZ3gMssSfm2jDtXF
LSqXB5pkk8obVAJmqyIJXVRnBZNkqUsGoWmbrUDMTBM+VxIGYZEJ4LMCivua6phS
HvBjpFC30t+okxh8r2QeRnd6XDOBDu12BNdEZv3nB4xGpbUzGa3pZ0eE98jMtMHX
sffVDyiIgANJbxkx5KAaUq0LEahePlDvwnCOeAKycegUhf3FwUQTaHATD+FBn/y2
mKSPcnriqgMZATM7C9oW5RKhTGWShRf8SM18Hn8u8pOyqGplpnPrLwEDSqfL0qa8
NH4ONTmt+ipIQsFfItOP42Rbk7HvsP0EjtVdf407ytvUng+/2ve8OW440xSFOgwe
WzIYubk7/d4vVOdUYBhzkCH8S155FaZVlQlSRV7bemgG7h2xBW1g7XbtjXygFuU5
g/MZjTmUgfPJjItJNq+iIxFos3a3cjGEzrs2hifknuc4a/+yxyygqRvsKeRiuHtF
3YbyyMf7IRYYFHYXN4fQwo+YBenJtgb/aKSmCgp8ncMgL35YBEEQSU4KvN6c5aN0
uBSwFkbCtzFWP16G03e61KAvDWAIOpyNxKD462OhxwYxWBb/Sheumv9cyteoUvua
CZ03EboDNO7vCaLNRvRVk5b8CVSfCQlHlptZqnMUY+edW7UGBHj54Uhp3pyKBjFd
`protect END_PROTECTED
