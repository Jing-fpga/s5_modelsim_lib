`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bdSHZVypifJtBnbIFT20SJTZgtykJONjpj4GUC+kTWG7wVBPQNDF5jEg+dTYPt3I
F9GyLZKrNVG4cRL5dIyJllC4Cpi2h3+rwg/eC2cNQ8BTEJ81awapsti7E5z2gl9o
X4ZjGKQNpjHJGC5OjkEPhWN7NJbmRDV5f+tGUfpnvLPtspBMkAYfY7nHXidAXng+
GYnio0TbhIFQgJOdRptI4RVrYURXM5Lx5f0vAvYiJ3wWYxcAFIlQCpQfwaLWb/ZI
EesvTDj1v5ya0XTR3rHTJgKb5jv/fLuXCDGjJYQ05XCfushhImMVm725MP4FhiFU
673VvROXonLYidbrGOGYjGGUqj7DpySqlUWHcO/zmjuaZfF6fQIvR4OsEtdwurq5
ULr9pUez6rEZABvtdkRT7lKJEPVuBQFLhonVHIKarQoqKb7YuiDkKhOuzA2bxwnm
++W7NhmBllYhg4TUHl5EafOGS6aeD77MfQJsU1a8Q9BFcZLCz2F9yCMERPKDf5Wu
b6Fj+eHo1JDU0fuhthQypgteVf+VI8ZZBQRAJuRQorMTPCK/vZAGzekp0VYiaCnI
n8B4fJS/j1SbtXf+PyV/WJMKLYpj0CWbi68y3diINAx7VusbnDZqcjMW6rdSjWiv
Eodguw4Wbnwe0HZ6pwIcYbAj5CCLywxb7I6uIyoOS/1LfIOa+VCfeSVoxM4goAZe
6rNOcffU5mCsvlxtunOkHSTcaZlfCVvyQbPY8+6r1voAdukyCGfAiK9be0Y8XZRS
WNaS3Z/NCGCST799K6WtDugxICpyRCNlQUFR7fSlNKQZY3gs7T++NfhbSYDasgd+
1glIUs7YJa4BR2y512XqOPECaNd+PZTkfRq3AVGoxmF9PRSsgDL4wedZlhgRwkkP
3JZOxesDBrnQXlYwTbw+E9W2GsAFMRHE+a7JB9Del6ysS+3r874cgwwZrMWwziPT
`protect END_PROTECTED
