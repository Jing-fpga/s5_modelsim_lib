`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OBBo6MpzTOStXSsQcaD5zSL4i39Jwy24BcUv+OaTYneoOjMavJjZFIvA0VepmaGX
ySfzKYKkQwIT9/QRQYGfpJenbVwHi5+eIRKwe9s+tFZ7SSalPM46GSRH9UAzFXyu
t5zCkDq7enlSyaOMMZjWWRRyeDLcw0WeYjDl8aed2JId75SklANc11cdJ0441S2N
rMRtZ6xy7XuN5+czzun+yYVLxHnX0e45Ia2ulpPQqPjqLXBEAHdP8bDVaGdaX1RI
db7vGybWuBQCOtHivxQEJVqou54kMc0BbVQAvDHwFNEWZZou/6jQe57oYhjAh5tD
4H8fYARWSkCEZG5qySIgxTPiJ+yFsFJtMyGDWG9ZgFpxHnpq45W2PmUM3cZc+dE+
uxTAVWAInV76grh/LQUjMAG5Qeb59W0X16ntFvPiT+bxBr9v0MPbjKlmD2CQZNZ6
7mW5h6rEJHzMvjzx7U8qMAkRjplq/o3moVfYg+GRiI5bkoBDTen7JACUq44JkHi+
N1gHzlI3u8rvvZZesgU01FvcK6x0/dszl12FyEca8PyH0wq3O0JjaFMnZXpkIS5z
GuMHM5JFV7vYrggmz1ZUUsCYftCnqXGDtXG8WXOhaYKzTWJRJ5UXu9kQcD2Q7xyR
EYVtP4Xrh/nxPmiNPBfMpUaAXJd2fs2YR/9LitfLaIc1bZEV0QF7OYIjRSjg5PaJ
8cRStyUB6mri5QIrghVsWjgg/hwoC0LldLIHfLqDBXM=
`protect END_PROTECTED
