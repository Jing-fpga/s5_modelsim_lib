`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
44CwH9hSaUs7aVQ7r51Us0nkz23Ku7rH3t4Z1p4t/qQB14K4INHT2KLSSEK4A10m
pn9dukNZI6NkcTzaiOgw1sOYk3SrqKJOyopZ8bkUA+DZVOVcEV13uOBctOG5w0xD
6EocI91ab3S/wxL16BHfqTIx3CwSOYLUlqKwpfY81Mf0Omw8nfphrPzoArSeM6/C
u1ORn1BD9+qFBXVecUvdIsY1lr7OmIlDRmtMLHqYb/bybSPcwkIucK8mgB6aPV6T
JYdZj9Fvg6NxtGASylkYGleedV5aWP8FL3et+c1Chf4rT1GaQFJ+h4JhuK+iLoR2
BXYOJRKJ6nfIfcfRDgS1RWZznmEHfz60OZOR2itEwzRL4zmtP2/1zBongWZQbe5g
GCzNyP34XXPhgkEUuinbtg==
`protect END_PROTECTED
