`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lmOFdobXB/0svEUNsGJrGQLhXc69GLNnTGYB+g2mollbxyZQw02fgEfKIwyf59hy
aaI7JF1HxJoriA9CE+uLnecDShTzVHJGlaBrNvdxIniPHVNPaYSFsntaHKHzHv7z
Blk+WkBhkEZNcOwvyx+ocaYWE8LMLpmX1/NWHImYCAindjRMt6vdA+6ZtoPluTla
xSgyWSce2WxFnuI7PLz2XDLyR2RvxnoZnN8pqTUYVAhyFh0ICxAhUh6Xs6tTL91p
2e3LWW3Gpo6Deyxclia+39KV5PUEPLi83Kw9yMXGlU9KRDH93+HturmBdbhopwkm
SUL32ESyl/V5D21ZiPXluJvZ2Lf/6mdcaBaTD3lMiA6nq+crvKJpvUxbZ4+O21B3
tJPOCSRId4/L/YHajSus455NYH3lfvkYTB3YVh08eDSDZtQHY5V0KdSKwq+gjMVR
mEgHnp23HWB2027ghn0v5B14Q1m3p5W8Bkv2TjlVat4b7Wwaew/kcKhIOYJaiB49
BB2Wi6qmocu152abvPVFi4ft/sUM3yBp8Zt26od4VsOZxY8jWIn5iuDYUGnflhJa
1pOwMZn6w4ES5aV3I/ZQng==
`protect END_PROTECTED
