`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rU6LOUttDtQwti8apkUobFnMzy3Xel7m0GCdbymjW5WMqlHP8HdSTWF9CIA5t9jr
dXou7KfBdz2QM0WX5xAgDkDzB1RYC/R0FCon2IdSloM6KqlPnES0Ys50aMdOxeSy
DL5Q0+/jaBCrx2BGHbRjUvL7jWYAOOSeTcj5I/fu23Jz+qZwzyPq03nzhiozixQ4
yJ6k212MfBVStmsO9ZOiExYKCRcRrZXP3rj3n7ugoO7jVwsn83aL1dWZLpfg33lW
ubni1qgejzXlxlQcVBdp2wslUrcHUkrHEExQznThG83Ykis4julWTVgx1rt820Mw
V+LpQvSxiEcjEzqBTkYRHrz7O6MLnoNTToNbwwJcEbB8Qu9f7rsF3CMHVzBv8Rho
TR8NNs/RnX/7uz5zYLAaf84i7IRSObOxvLchysPITw2x/0Ze2pnLrpak388aXYZt
fIkDeltqqkc78W5u3dHjIQlFhj30zwLqCe0veXCcacEocCmv6dUCkwOEDu+8DblS
Iu7NcCgJRKvwP7XvlDlEMx8uwJ/AY63xxUy26JLXMqWWHazbehEiAbDd7mQq1lYA
NCSo4opldpowdLkKu1fjIyUnCSKNP5T1rHwq3tTudiD1HyuZhvOyAbxN0PH/t4Jr
rcfMSoRA9Qcj/jGgnB6iLefJuCcVgHZ/JPl8JSp8akV7oIah6RSi3j2F13umwfw0
fHSZxuxoYsDlNYmIH0pNNbxXl7j4aVD1Ite9T9+WhSL3Mljt1lZzRAQORMxpR1ci
hEn+rQUlCMBCOrMcZUtn5BujAI5bi2QmZlJCAX4u75AHdgCQJgKD9Yyt44oSM9iv
5UM++pzpE6XfWu8928ociMdQokAg0oee1v/Fp+pffdY2Xsem3tfaUt4ySwqG8Ov6
FwErGFPiQxNBD5YrPvVQGDj+o0csQkzIKLSgw/6KPI22nWpsOcp6NJEK8ZZurutY
xbOWCvFsNFpsJsbtY5Xd6qRWAC/SfN5VogCyLd5z3e/UaH9lHtTFZRe4ydtlfOau
6hf8KCWfZ001SlHFvsihTQFjJHNWityyB0onNYBWLrEExQATJNkMmB2Lyb6xPXxO
549XpSJ6UwSMuE+7KLDQhTeD2Ir1MnanUYk+2lpayJ5/jgUp9gcfUUQ0WFb9rPwl
GOaqzF6u7Kfs6hzCjNmaeVlIRF39zUaMW8yBcW2ApPDtPFDVpM+Inq3sWWBtQTBE
ZqpsOjNZj9Cka3ZkJWDCFA8NwYITs/PGcXlYcFgIibvuJg1rnZI6HjlezB48fa2/
UQ8RsqXfXi6VHVTUv4v1betHrRxe4aWVNkKYVBKiVmU8H7hRIuEMm30PQqnBmdWR
YxhoPhGtDnj6sTtq1Q4uYTfQLGkFnr1ZDJ4bHOMG6eaWlHGkq3awMPQr8tkJpP+q
kEbErFqpmvWbiApMSKOr1O0wxB5YiOXPp+IdfW7nY0kJHwy0w28oBqfp4wmAgDXo
5U+5yGvbjQQS+KNteZcXzFqWZu3sryhTBxve/CITK9SFGT9OgAQBFVK9kSk16isP
RvJL435cn524ICLinIZ7u8TVySzK5/7K2wstO+Rs0QMLOp3ji5RpuBQ9Rrqpkbyw
QrN9zrinhKxvMuaOOeOMU38VKpzSAoEKTQIUogOIsF63zjBn1eyI25bCmrWsI9XN
JL2jfsUo3MmxdYPq/UurD/QdhfbAdxoc7n15Vi6Wj9oS/ik7loRdDRtszngp1lAi
SfMJcowbVdouv3DqOm+d8iGFzK+XdWf4QSBBWLuap7P6CJ9x7qymHVjFBbBs9BaH
ErxMbB/dI4/dCbhfjE6hnZ3Q0qiFCGMZN9Td26dDrB6tDmUqsyztPDp+vscwp3/k
x6BKMzTsCiJM71UsvyYTWL2gjKaD7X4OcUkPQyu+AFxmPLhrUoveT5Cl9uV0Mhjy
Xe5r3P+QJgaRRgH5Wz4Zf7QSf9YZM+KY7V9YqDQ8chdDJs4tYG8mSLc2k9VeV+20
MBbHQL12/P94nC7qOSLgrSKNA4Y/1FhKsroh8UdGRZchGg8NMzkZTyuh0GFyX9QV
IWZsmGK2h9J0NXUEUlSGiNZsivT0CF1PM3/rUnnXU/LnmnL9RST2D8LXhg/TOtaS
VyOsogxQwMgpoX9bApJjRONazD/qIKJ46Rs8GiiFpU/KcO6hGqT1X73GqZ8ggB7O
Fea21ADIgnxqFwUS4kd62ftozwAMe3GpnnG/hRpE55BbmOcStoXLDryEhQARddki
FlFIKQtkGyHyQLOwve3thfRFQo7GPCDvXdZh9tG1j+SQ76+gG3VbTaY+MErjxcOS
pYqtzwGtrlUWKx2kV9pBATukyJPC9KzPoKNrlYJosZ9ENKhLMiV1LnjjFaVjVmhU
HtnaIQ3VXYaNv0nIzsPA0vDw5iKCEkuHh91wyj3pcPMoUsaD8/nJR+VolnSolF5Q
q/ytmJIJgTWCkbsD8a0OmGsSJGZRsuZlkJQoIi7pDGyw9Edq99CQiYpfoVF14fjI
4LSSqaGgdsdCMflCK2AeJZQT7ZvqHEPPhBwHoDQSG7WINCBtAImu6g9hUpJVpYBB
azF86pzpXod044luaVHTm2OiUmDYSUDikchocP2DejhsXf7MstY0dLHKnEcDvyxa
CBkfGz0UPY2piahTdwkxaaRsz7rhInX0aHG/W3HYep60ZbB+GZCdxZjGw7mXxuDN
MuI/PRKT4m4TMg63v+wLoUq6wFcqwojNYGhyVhNHEpM5zEhB9TW3h73xz0xTCKpX
poQ/juqmb5yeC4aAsZvk78y1JCmKDSaLyU3T8SrAigoYOjZm0KYHJICXJL2tSndZ
Nh18eIS/RyA0QzTDaxchtxt8C+Rm++5qogQpEpyoxs9uuTOQ46S3kt81PGlQ9FgH
/RfJW2NMlqCkoB4i2NUMzuac27Fax7XuU9q9Lt8RyRsICJ7CL1hXZM0gpurDvO5G
yGXIQipPR0BgKZCdjaR/cPyDPUalQuYbbDRwKskU52IUFNNFBhjOSYC5SwvruDxA
KcTEl4DMNvmp+dyyJ23PDyumKuZh2detdmNjol2OGpMZKP0KgqITI861ObLzqagz
ywcOQaKTyGaoloaN/RQUTN5PBWMEK99YehIYogN1VryTpRFyro5UoX8Nk6xmrP9t
AoX0q2WLT8guZHJ5rPpir0/WxRszHGe+ohVfX9gTUgsSwNLt4jX3eE/fO8DKTEzd
lQnPXeX3lTxXZ16saIOKTXl3/dyNMK3URwuE6ujd6P9XWbjABsS4D7bEP1I4RmPC
lXDiEjgh9pbNgRGFiQEAupZwbOcvB38VP8VRwc0vgUAuo21yhmFDn7Dns8MwCPtn
cOfQ2zrUboVwG64Kr/fkNvKjcC0F+1GM7zsp7+CBmDZ+kPg/MHEixuvCqVjHuaZz
LMRfrQ79UFhEYHjrQ9uiymK+rmMBaoO4rssG39SsGbMq7aaGlMHlDEoElIveAHEb
UOwk4ieISZ+YK3ZJinyr917HUyGzzC1pBWmPYhdIQzIjJ9r5vSNv4gsG6jdq09p4
Fbmqrjpa1QeLi1wWiMrX+ZVS4nxGmHqTduGIH8K5YRLv8LdUOgzigzHak46Tcdor
AEwsM/oTZORpmF6kFwFSoYZ9H1OjIhCtwMNpf7GsMNr5+6f97kggHhsEN4nCm7YJ
sMIma2HsFqkmXNKIouYRcX5AuuYR0m0tPQj5mQto/zV2yQs8mxbk5eO6iDRg3Hfb
GLtwXLLlc4aEdffxBPAVVaD5LPkJXtwINRI+E36MEbFRN6XUGp02FFAjLB5m7WrL
PfRDixCuCb2lz8V8oH+6Br6o24u+B0GrwzISRYziOlypRG6k/rWa/Lvw3XsEIz1d
50A/KU+U8uZEwjf7gG7K99Jmnx+BshsfmkaOQ/9BK6mz2GYvleRFNR5/38310pLE
S8DhBTsNwUFKLoJmXJVZJD3axaJHCj6sXNFPOGK/r8ZKjOU2PQYMPLJJSytCaJ8N
3QGsYB5ofjHh6TRRUfaRKpciBHsgv9qrjGwhNGGAFicDWkn6X3mWqrtwXX6/pKv4
8k2Ugbb96fTJRxg6eWrLO7z63ajrv3OnRf4zUBYQ0OrvADtMTi8y5p+rVZS00iPi
P5dqcwRdmwRelJTXJyy7D8DRJzH+mWFRYzPNcn/hvgKrrMxlMtWJKa9ocyGCzvBH
FBGRXYT36ziPKmLBGfcEqLAzSILYSXWvNMP7u90tcIKDFFVz8zYyYArWKGTi2Nx2
n7/5Bj94fVAaQnsqJnGNVsoog77xU9YfKewsfPyuNv8cfVIZZ2TBKgaNA8O7vI4z
e/uJFtfGjpsyU4ClIGyNMxxTVAXI03kBOIhlLzfcNkWRCZD11SpGBE85nHZcQCpn
ytVgt0wrERpcugzpFzO+lZGVbc6MQ7ldvgrEVdywyT2IUblXA5TyLhkPjgvSzcZu
+qO0epN4mRNFUqp4AN3TUBAP2UA2QjwPwde2mBJVneOyGpEH1uyx9WqIW6sDJUTs
jBSceIkkrSpof4su51Eg1CTGa1iE0EoexUyxgN2ECXI=
`protect END_PROTECTED
