`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yK7/bLTnsTPrOsMiCj2CQu9I4x+DHAFnJtiaxQVMU1kwAiANQ+7zqf8gR3u7+l36
e5fR43420U5Dx9pVwlfmXmkIzKFjEXvUAm4FtOKVwj8EVDvUTMdLuHu+xl0GfB6a
yau10o0AQ0ntiXhNoZP7wfGhPffm5xdUvIfM0OcsSzP7egC3T58royKrtiA91ceX
s7t4iDaNH7I5aEWbl4ZDPtzIoumVv9HPBS2xl3zW1ZYnwEtgNpAGVUhes9mOaVVz
FTpixlCwOu2lrc491d15Sbwog8sNqd/xGGkMgdn3VlQV0Wk3n6TjIuXGDyJQpyUC
37Y1fJtOOet3EjXyA9vpXvY3ZehJ6hUgOEFcuJ5ECIypBL/HhR/lCrqS5eguPRgC
8GWuuh/dHa3QyaKYdx9/ee01o6YGJCqk6w1IBg6BhXEdgyS9L4u3SuZNGj48WnkF
BGFSCZs74rInelF7hbNaKvTdiOFJtUcz1FyMIWBYK/6TYXnIGqAIVGdAO6mC5jfS
sg0eERHkz/m0zsYn11wQ5iJaEsyRqo/Vi5jyZszufx4pd4O/x3zgr+iwl0Qg9Esa
awJ3ihR4oAO9fy3xfBqyVnN2osw9hAu1cGlxDZTvWh57J8Y/G/GshyzLGi0iaK9F
C27kN4G9DWrC6DZmnlT1EDRVb8YKq1gKkhSkkEQh4QWWThVqGyOeYOQ+LDun0B1R
2QS8hxeDBiKWRJ4jilqyjzcd7UytuPcgC7R/COqm8FIvyA8sXnu7peDIX9yqzXxk
aL9zx6J51BcFhDW6XS08n++ciK1IY8L1EOxbQpoowXZP9Z0LGJ1Qn7Hmhl1c5i1C
O7ki7lZIb1X55bPwNq6Nmos+upIq7/KmTiCiNeMF1dUQaaKEZYVohv8oyJIy/xIT
E2vgQIE0u/WQb9/4Yy5O50LjvlUQv//CSoamgaZbzqdKjCHjthzAOR9Zqxm9+idn
IcVxedO55Xa+jHthkiJkgnGAZPwghjRjijGTc3n/+l/O5/58WCcKGAuJxUqJCAmm
zxV4X1e8qRMT/NK49+5N/lSlVAwjc3M31rLCtuoDzbg8Siepgc7idFLfzm8bUlcY
JR3dKy6g2qgMmmD+zTzJ7Jcv5p2TwX40+b2LlRcyHFEkAS/n66RbfsKYiCREiagZ
oZJJmyholHGUT6IR9QB4ElqJrb8CHos1/0Yx32JbFA1gv4cHDZFXbyQQ/1R9jYnC
blAG8LMIfSYxmGvhqoLnr82s25WScAJcVGxT0ycGGuvjJAIVskJqlDTBlkIHxEYG
hEZuyO15YUQsc3g13NDthXR8Ih1SaSL5DDX5rt3J0bKSR8BjoundUYUeduXLD+iX
YxedpnEIcQizFj5Ro4gMzBfYfv3P3z7wWHqlYUwkxbZMrdHeuo71ZN5ZZMlVk1el
NJBIfMM98XGe54U/rDDcGEG9QWKR6UZUigR7465ieExyAApoSnHw0PS7kSivOh4P
uHVqJZuFiMJ+4L/ADc/r+0KNppuYDWdYOsXQX+IKPl0=
`protect END_PROTECTED
