`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mSZ+k9klDRSCxB3xjznFWA/gq2+sh03tOcLtErrbVDhZJsV0n7hmMSCGqHbGlzpG
PePLicNYxYJtklm12nd7VK8kVhez/eReNFtstOCoi6FQtCCQaCyVimGg1qeKGmEx
yqsqsKlHlDQcNvyozm2bcKPEi+dVnBlImKeG0Ym2oWllwOIweMqop4sCcF6PrBNV
sSv6c6RV7DIv6udpvgSblkQ6QOqCcDQZ1lRxRtAMyoV6Af70zxK5UUrNWJBQYaUW
SNfP8fFoPzaMGjMTgsiKX9IQlphFcbmIra8Rfl6xVeSpLrjdPZMbN3fQ/yY59UNw
+5obK8rMe7pO4IZU6VSgVE4FHOqg4Ro5PIYl2/kt6l5u6IbcsWQg3iMnw97495m0
STBizcNoyC9D4pmBkEcmWFHzTkUealwBDMX4AcdwzPmLq1iRSLCYeNP3PqQOzXlq
KCUDJHQt3PhZW++1r9BiMIVwOkINWXiO7FaXcVDl3bBdXhK4web2N6mQ5YI+dX9H
z3kpETrXIrlGv0Gm8PivJVGP4HXWPBdmWZApOEQbZ205P0yKQTSjPPqGMi9dA9bN
`protect END_PROTECTED
