`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OaGxdDYkq5bTE34NRR/P6XI5y6UKT1UBMyl2L92SrlsscQixVWreGAhTr+XwdcxR
DY5pRQ6CJ0Cy7Q1gSKkIuOIggeeIiBNhYpAgYPAroA6DPrDTkAeiuNwerrcHXnUT
X1pL9dX+i0ai9ZFhWhoyOc7VkAAEFvcKCE4ezFVT8dsTTuJhkKLd6CK3BgmDip4v
xaiinvt+yCIlN+Bpptq43l/LbJbxtneifZ5esuT3flWCPSqnk5MFJ9u6YEc1DWhH
t/wSB+3SvHFCLCakLe4V63/miLmVD1AVf+4k+Ak8GE+ZEPlQto8zJFiy/1AQK+A6
psoYllwzGerNS/SJxMLatR2JjsrRfzNuYwhnZHYqTQLqbrY9OA2ApRuywbV+NuNN
me7hP4NSr/5JD1l9Nu4MIO903qUfFa1ViNp5TbpwKTjNCHbHMT2m2MCt1WKBnOxr
GKL2SIi1lQMA6OUrEyGJ+BtTznNzv1R7j4Rrf3jOGr2jQchaXaPE2L1iLKNhS2Ep
vYILNx4yKRuTV6I190AKFBD93wELvIht9pcoE+bTXM8KygXknaK1egFMjeFiqnWF
W0WR/pl5XTxusvux/uYbNOLT9tsMWxMl8T6araoY00syohGcW8FyVhBY92evjbla
siIHI9fi3Z1m5/M2Fyx28W4VIgMKjg6T5Ki+fApSOyCHm0xfWPk7LdsNhYz+VDV2
0T+i5VKQNZpzVK8XTZws2KPuiKz39g7LvaK6EJWBnKhy3m/Z9bKv+sqEGZ/mDyCH
/zHbP3l/pWvwfc2VcAUYlaHjfLi8cB6RVylIonkC7xN6aopequz11ze66UwoppW3
VI6iESC2a4n2Yx+xbDF8vlCvPaabT2MIC1u7ZF6uGGcXWY0C0H4C4Kyt/VTnWM6M
B7ZQvJ0gbadz7pSU2yP+qu7mWUKxitnmmTyZQTt6Cw0V+oIjz+uTtlzXHgnLK3Qg
OyFj1AoLjQuKmJhvxnGku/GO5WvFEcDhQMK4pBkQn8wsB2vP4SIkvD9N1iHpleLZ
PEpstx10cTgAyb75s9HZrrH/YzSsaxHlGJo0yVIm98svKCmi7esDcitu+7tg+bOZ
5wcE/bKll8XhctW1Qyf36HlFoB2d92z56fJ5dr20ezG1aK+3HjdyjXj5omsRJCox
CqDTYrwhNC7jBv7uKlxTe7Emws9J2MXMQwXimKt2TKpyEHARIfkKQf8XKNYsLnGd
Zh9k9cWv590dQuRZwkBUyNWnr045oY7+zvV7j2H/bmSt7Lv32u4JkGyY5Woby1JL
Nc4TBOT4+xVPZvOfd5mmoaIAj5oLsl1FGXmivzFtmZzo609ZvhSL/a3l1G6tQC0T
jkkj6S6esM+wLytZF01hbZU3ghriANhgLJ+bI1/gWoawZvTOTdDEFNY7baw2nm3K
ftGByknfXGDmzOusoB4vhSyq2UAohDmQTlEU8nBYCK2ZVtY84r1qec6UnX6N0Ykn
nAPEeCxzUDrZHPYTGBQkqt31IN0RjU7vCW1HvhivCLXEIU4lf4BaXrMqjYlKdruK
M+Hfa3zDeOOYUcHdHZgqzWUbb8M6FjZoy5secoMZ/oFgONVX0aTdg3cAo053EtSW
RkWUMrYo76cekVRN20wH1s/tvYMai64l5RVEdyLjLc/bk3AbkPgvwG2N9v+g46Nt
grvouvdDKRd7vTWPNizVH0WeIMLXXQ8O8yBWWL40vfhr3gLFUHpZFBcLqttTAmWS
IsY8PgzOXc/CnbxwJvQQG6eFiUbEGMW3WeIMF/3rCxtVOh7WnyriBHGIJKG2L8Jk
PXbWLO+T8qPsO5EfJEDSz+2Wu0I1Gxx5j/s08VOBTeO0iUTjVC8zZviyU3TBGTQS
qN4a+pfrdrYkxl8NcVmVsDZo1NLLoWbFcA/JYl1I2heejXXuXT/kPXOQfYsjuOmv
gLVR/NMhALp6Bg1aR0E0bdhjMrm9Cf1u91hvBGLKeH+YK83w9UxPOkkrYUTLa1b5
uzW5YzxlPrNqt/l2715uofz2+yjx4FaB3zVDpva9D0zYSwBt5t5F4yYvljbHxtqk
SWcgyqHe3o8rYjyPI7iuGVohJrtbCOZiUGqLDgVV4+xpqjXJ6E71hmToSlvjdFsM
4f5i/WUXPl6F/5EIImCCN99rpiAhunycwEHPbwpSc/qKuMLzDwKoyNAley1t/l/8
l3w3WNm2L1iTQZMBQqr34maf4pqhc3d3iOpMO/dN/8ydsLFKgaBwLJwvlveJ18ow
m6bg27y4Fuj3GafuC2K/44Y8frKodW0cPCchaTwmbaHTS+aU1vYaJKQrU9se1i1c
502TK6LQIz7irhJ61C8DwrIjjN8wt0GF8sEGkcCF63ctOrXkMod2FAR5zOnTBJUK
Rdxtmd/2LEyt5n0qI/KN6Qsuw48jEv1BO3F99Ybr6fsXUEibEHZrDE62Ht/d2gQR
H3fgg2u7zrpndus2kvjsD3uabUAIW1oJhuAKbtkw7TJ9LAl1IkqguUyiGK0P4ltY
`protect END_PROTECTED
