`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wgBd25kFxdmU2gQH4B9W0rqOh1MC3uZ1DdS9t4nDROxGaYv9mVDWnWnIhR5VCq2O
WKV2T8MKo2Rk4x6tpKqDJNiHYJX3J5acxOLkxFTEK4JxtSkh0unslT1Jo5C/bVHh
LVGt2n2UewCFGVW1YtJSx3kpANuAMlJ0Chw5dmSBFxlG1V9FfCpwaZvJevNtrhH5
faXnqV4GU5QcqMDTTOzRdYtFi9ccJrPSiU33b7GX1oDSmr8vTPh250JPA08WWmF4
5saWyj7XZ4Hg2xQx77rtGC6iHylp6hUv1LpZQvJ0UGvbON1vRq6k7AzMO/zGtCe9
yWGJmqAt2Bt02+fDW3J06a+cAX4sb9BUtyZhVnLjlFViJOJu23YKTdhhiicE4T4V
Qpp+ZExKz5/4061K8Th8byblSQu/9GVL35in6kvdGwfr6nhEliVC5AjY6PueeUc6
yC/U1ssVo5PlpHWr5fQghU/xtTK6lLQilwx9CFfpclrGdiURYaP+KoKSBcsgZJaR
iH2u3TQFWrjKhJNAqjjGlkIr7FI5sb1kVfgYFbyQJy6XdSVuNyFzXz6ML1twxEXg
KG94vQYPfveE1xchNJ2wg8pIpVmMzweCzSgAOyeMZE0ieD5F7psc10WEJTv7xMAF
BIJqXnS+fqM5V76T13eIJPE5WNFxE34ppDm9t3NRzn8ri4nhvI8QqFcEkmFgMFfU
Ys8jXpZlu9hKBAfdd/JfVXt+yqCo5mIGe8hrVA8LuBe2QjJ8YIUIv7ie99uZxzWy
qbRpLHX4en8WL3O444lLxDMPsSknLohzPdeOUY1doYg=
`protect END_PROTECTED
