`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qqGvcB/Rn+fBJuD/e54QitYytSNrp0xz3j9ll1hlxrR0sAVphlVZkRChIb+Zsxm6
F0Wc6FeksXi3r1/cCceGQ8jLmBRk9iwdxwH9Sijf1A8ByB/yvUQiNXLb0KAC5auQ
q6laKtGwSm5Y9mL08qFT8Wf8tv+xlzY0EkvT+Dj7LAuKjW6eLfUh49DumQnd4oFp
nZKz/BdEARCIkKutYKZn7TaTuvqZUBx+z8scPRPreh+PgGaQyZ4x1tdTWgQamgOm
5LS0tWvSFwxy56M1jhzaFhgD1fzr0B39nI7hlc3nn6IJTUFP600PDKb74+eWDH2S
8ffOhyAVmR0fddrDziNukw2bDYNUNpq6+fzsI/E5WOtoDo7kSvjd0oj0246Tr3xI
kRrJBime6507oQGBrFVNKujOMzy7Fq/JWrTTAcBIrCmDQmZlO367BxdTxznJqR5a
vjj76GiuekTHAWGVENtGDun0waJS2bFz4bBL+p8TZ9h+AHjucmcaZypGS91C7WRh
k92hPeRwpgRT54szpr+cLGt42wcgjcBgr5ArsUOFGDubm0jeQKPH/qyJ17NN7mR5
UelnHdWLD2ym/ilg5EzAiRljqQj5UpW06dTb/70ZcWkey0JnElOOiONVgBws49mU
rPzT8D1UWtCVzGRKOoG4tjLgIOskaOKtPawT1IZIcwM5+qwKmG9AIBTT/SLkMq1T
LS7G1rLo/kc2sOhNsP/tuDtOe1FAgmScSKIrEZBuIa7m1XG6nepOoFtPiq1jrCsv
7keGrsB+Ldm+qRj4l1fGWJm2+SmecyZugER3SV3SlYbNt5bgC43t3HgrIc1NMhoJ
HtykMsser3qUZpQgFDjkLv4jt+5jG0XsbOwaYmADxEOKs1nRcjpB13MeVzW9g7Ug
kxJYB/jNjtPD7Fdp3cxVEK6WwUDi9S4L80hTD/O5CppPt/GLfs13vi71QOYvLJR3
nb19RfqMdY2m7GMzv3f6qDKl+Fte4Ohmu9C0nA5yP/d0B7TGN2yC9Z/QTUWXbDQu
8Vo2sBzUbJGYteY5VjrP/ftfhFec404wkeoR6+e2989zqKOIq/Ok1FQEAIitvkM1
XUa8rKMFbDN3tqMZBftmu5XYXGZUacVcVMjWMCXp4MnJV/RdkFgs48cXCYfGsIBV
45EmLpP1ovWUoDKHNLop+HM9t1vpeWc3rtz+IKc7UxjBksPTgaecYyBWOtJMQ5iH
sNMwxgPHiBRKJv0r/NgzjDfABqCrH9LL4DfOE6KgyvwTKiSWMs91rDv5IxDuzpAS
C3IvdftF8GdqHYkuQtLa6J+XXVjK0/jfzfULPMf4tzqltZLm9VhhQHgGcZX5j2qa
Dg4Gvmnc5fiPzFbqoqQMVasPKk3QWKZH1h6oeFWc2SSKyzIowQl686tvBCSFhG/U
o+PXSf5s6RM1z4ZiADf6R3PkFSARir+IVxGTgtbMFuTvJ7hu/nNEgkwmZ59PGGnU
qGAHOlSScpehLQqZLw67xGoZ6VuMsB6qJCVbVm/T7JQtOeDBFf6Jcz/bL9M2ZMBU
WejLPZdLMOrYcCHYh3tQ9uAvpkD1N+fB6SYi2yLPqA1R9uFkoaqG7jVrlsdb+kHL
f4pV8Qpm8X6tZDb6XmoDL4/HsOCvHAC2ye1LD/PQUemExT/3YuJPBtsFQ1pZlFyh
n0JGzsq4k6D3NMkDXBVvuFmFTFDLs/Qu3r1Bm6BubLmwPIu3lKdwmuk5YH5I0pfa
VVTGP8ApwhrmVYWYffp6ZilobT/gBbzOsEyUtGow1AWHjYR+jvfsNeAMhcqlc29e
1rr3I3WxNfz8PxCMcAFxrJUIn5+tGVSWnqlWjncEFGkrvRRRtWPttIlLRCmQGGeO
ySzJ8NgLngMQPQVqRpa1p/0W3yPOv1ZwCy5ALJo5QbFqfCFgz0mhLqkXsGeaMqnx
rNsOkHLnubXWG1f2TjyWfkQ/Bkc021cipIyerZdaSCkThFuyGf2XAGtaC+dtpais
vqVkOtsF+C97IxXjbTtyNu+LQXRgf+VaYkrhfwLoq0/L5PsOT/KsDstDSCP0moGH
XdtQc8Yv0OMc7qIjWF9ojwvIHCrepS1fyaELXH7+LnLiFUZhAQCWjj2oA7IDIbjl
hWXVYLKvoM9aLsSUbeND5VIxeTJZfK7amyWvHhekuw/Q1GYLFtwJXL283PRp0unX
0uRzebtHQL7EMCjNRlihvx2H2d78Ata5dtvs8wn8bpga+CNB9lY3ntPHXDxcT3Sk
il3Vq+gEhwrJqOCxNeN2U6t39XMPhA80bp9rn3cc4MeM7PB051tyt485YhUXrFEu
jkCgHfewIq6T3DlKgux+vs2VW7dnfFlBFImsnbT7qr2hUbYmkk8C3QI4AZGvGuHQ
ua2Z5fLbmR05bSetBwWV4SefeZ0j4zFFvIcPr5WPyf+TbjB75qYTuNaxxvlC1FC6
mA2nAujsev7Q96PdiTw9X80avsOAmIXgFcPpUBZDzoUYxnIojrdr3PbYIuaKwH0o
HQW+Wij511E6nGMg9/LJEsn9cSX2qmRWJoEspqLR3vsw0IEXQlydO9JbOWcamfuj
zRRygkC3dvZcs7VD/toC8lKTjaP1q11Wpf3qfRNq1R7GjDiQ2BSor6Q6HlmHuL3Z
Nnex72zrRbVMQBdWKwjW+GhD8+qmVeq9sm9IQ6NDNQ22AI9wG024ZAZGhBwBHXB3
fUmYRNmjJqCpZ3G0wWZhIh8HGk4DLYN9RYwqAx7Joat/jTwIpZDGVLwvKNYrfuiC
nC0ISDGjJNHpUkR6kc96g6btiBc2KdY2k3SQxTQ70DsXLSMP8isYFeDc5cuy1IcF
IWU6iP59gllX86P5+AuftnH9luLxYegulN3zX+vRszolg19aEY/vTPWzQC/CocRa
7Ajo83WI8SGI+TRxwqIHZLmBzeZvoLvWPEjhfIWpzuvXdyxOlNarhAyFJ08DSQ8I
/en3yGrXJVbxTQ65bGE4tBsNXAB2sWhLcPO8NT91Y7o1WTceczmpchYsQRQ6h5QA
VldyK/QnSKwUAneXGm1rtohA0c0jDVx7WAsvng4WybknvaJmofXk6k6YKqDIeBgj
vUIMJr/1C5x04o7WBKBjl0Hegcim+9CLTuF7FEi9kmGFv0/r48gyOwOF5F2Nrujk
yhMySRAxWrEm0/ucL3nFhlfnTYyh9SUJoq5caGjzcCK5iH8+M9cRk4cuSGYvUeSP
5pVFkH1X2PNbtSwU1e0Yx6gyctlz7ugjRjHB7lwF+PLolTaw8EHgoHVThcJfAaE0
5dKw9P8l9afcbUgQXwG5hB+H4e+iqW9/f/3ERqerSO349NcIdL0DNI8/wZgeYE77
ace8QYdSD4S3ogTf2+Qofzs3BfHh1G5DJb3oOh0FAE6yrirNPM17X26xDoJI3jF/
z1XoYAO0/tbTQrl0g75dF/ZiUof5yPPbatr5Hu5xzwYc64A3BEq+Sxsg1ekdYTiO
E8KCRPqNBo9kYNdTbW9KpfjeEtzoR+93+TQ3m8ioflMK2jNYiLZwMq4UK2UEkcW7
yx6200N7YYmni7vHVgOsS5/M1vO2QbEarHvMdTdtI9rtfSUTz9wmxNA2pkFCycpY
7Es/juDG/kSBDm36quWrIvYBwvec3zAGQRmMeXZ0SAaEXJz1ZGRbC4VYYykPQXHO
i8H0AOKbCaMWL/cguNjU0i5CaPf5OS/+nmMepHqbnJn/Klx8WFFyQ6UR7wllNZSD
xzQjyyiIZg0rQjxeLkVALbjLr+1pttlmwX419mjKcYwwUj10CzPp0UWRUwoTod88
rSGpMESBZ0jsV1hkmwVYzmQzBDaTW/L0XRwLET7jpWKvsYBfkcYdFXPZFbgVBAgF
jhbLq21EMkfb90swuQInpBQGJ/Q9lFo/wYeUQMYo4xMJNuHIUiAvIaPtIxnwc3tE
8oJEsdbNcE52NdyF1f8uV8snSlknDltZMDerAp9XrRVxmLA7J1pjzNWzKZ6LC6iB
HTbhLazIKAvW5AAll7nLDbXp2OdYOjPrSnAmyedOcAnlMT6I4gSFFUhuuFLeXJLw
lBcO1rQQ7L1XvB+uVqxvjLNTzHb3FxpaRKRub1kOqXkU0zhTfLwsVdE4aC3ggatj
jyaJ65WrPklL4r2WZpwEqIh9XsM7tiPBtZVyNa7VhFU=
`protect END_PROTECTED
