`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D4MUOCPVcN9/rH0u86ZgG1eNLkDpxuEYEOpKzwPMxoJ7GHiFTgvZnFw2azkMPwXd
E4GJ2T+XeuHjNOJjm6CdskgppavDaA6h5eoSzde9lqVicQqzYfbGLglcxMw/nP+p
zQaBYF8aSGr2HGSxmnR9ZMSVmvDaDcJvq9KMfAbkinzyJc+K8FsV66vGmcapslOV
aIEhT7EMpu9yCCCEaZSAizigg4XVLvcd5N8croIf3oZAH0410FpfnGY5Zhh4kOKe
DJ1ffC36rhIjmpvC91gPeaXCKG16ZrV8yR0m4NLrEehC3aVvj1duwdupUb3rRKZl
NKFgIB0j2NELcIDCt6/tPc+4EN/wiTGzZsfB27A03LvCk6ZiYOprC/foWsCZl8Jo
62JhYY5Ac//bLSf+ZCZ6cC7tmcpMkLjef19i+MlW+QdP9Q5/NJ8hAQsk2FsT9Q+y
waj3qyE1EFgCyHR6qaZaGgEs7UoReukMjnZMuK5uFo1dx5sKCsbTT0sab9QvM78x
RbM2TyP1KlmPRYQDzWUilVX2ZU4Cl2yIAdfjQH83a7HxnnRM/9ZceCF6e6yh7IUB
btCZKbyjJ9Gt1nAANCk4ukfPiCF1Pl8BEWLQ01EK7Jg=
`protect END_PROTECTED
