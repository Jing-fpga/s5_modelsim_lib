`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l+YFbb3F89LtFuGgv/SDayHMAHexx41fwPM/DlQJoMGY79+Aw6cE+aN2zQ9a1xKk
7xxl21eh9VQsVo5uZUP8314OWJJHRO3RLV91laEe6L6damiJfBdps5z6Yibgjj5v
Y7wDuV/dSm/VYyUmps/c8iHcacHnltSXlN0lcrBJ9w/iBbVcvhijPdxjp2U/J/WE
7JPxdsBT3DQNTsVuyrpUTqJI9fAC6jyp6Fxvg0LJS325sE03CSYWnEJxwXxxHTl0
y0MsGpBjdxaUCto+8ZA88Y0GIGrSLfxgFJdEaF6rnJnBAxhyTSql8+UXVOgzOAnk
FrGNMHO29ImZ3hB1bv16ioiV8FtlbHs1r8gI76GH3liszU8k6YnvSwrVXZV+DUzQ
8Sdh1N5ip25Dw8ou85yl+x6QzlYN7yjr5YuHFEaWC6ln5rtTwHRJU9jIDLrgGwNz
75ckz0dCKnf39Bas4sfsbxVuvC5Z6nA2SsP5ykKfV7paAQAH+lw4xkj/W3O/MxJL
jWgOK3ERP1mjwDr3QsU3p5fmXQ0EkeetVATRJ2C5bfXMMwbsZoz9rXuvmdWbBgh4
DwkQ1G1+I5cvMp/brj9zR3qMUk/SeiGIFM9lVhtOl7tNuZmrWIwSQk/zA7E9109f
1VbUHWvNFLe6CQ7WOMZMPmhowhMfGJhdUclS3ILRotQ=
`protect END_PROTECTED
