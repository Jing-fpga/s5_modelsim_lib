`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dkv8yHIN9rl1RzS8rS4Nse6qeRlTltpNZeIiHCG51JwnnlK20JT/hMSt20hVuwzP
8fw8fLk5y36/5ojeUpYHbbv7yWV//44OFclFuxug3PMkqTwEnC7OKUE3pKnPhVCm
EvnbcJHDIowG/WfcxI/toIfiZu/hCRmh7JQGXm+ZxWkT5zZTeOdgyscW8Gnhs9/W
wWb31jMO6W9xrRQ7ByrBZgWgplJ1SXceK03BlwleoGrmGPT+BEuuKU27cRDTfm5+
nzF3fvjSTrQHamlbK8v9Pb7OeC1dvJgiKiB6fa1aWkcoPQCxCrmSfUjtjVL0teRE
sKaBB/YGgmElCGjFRS7DcmdMevacryovdunAYGXD8AWycp1ukc7XCzXm0TW5GrEk
Tw457EFpIfIwuMegEbBhIyu+vJDjvlG0ZttcdBmjVkVHDCUzSxuSJRoq/RCLuG4U
XsL06P139Hfku1tu27xiaQbC0duylLIvFhw1OmKIolERcbJrAKULIlwXi/4jew1M
IfdDomUU+aR92ex9L7wl1zndbogIf3sPptHNBPVJ7I6AVWELpTCzJHIgHhUoXEwp
Q4v7mj0hbevhD4GNicExYvdeg60ArhwMWH3AdMCdJEfIcC9Y33eQvOurfKIcnm5L
q697S/51w7gXglN5Uq+mo6+BTkZECuhrJ5AgOKOtISwp2I8EAoHsp+Z1Yfpac94J
5zWbpL3Ezh5GhP6j9mUerrXCgX749wQqznRRX4x0AYgfRjr76mfMAWOooCUXZUZ3
HaNQUY/f2UncYEAIZjvhFwmYoRFepMOM0K1u3S69zS65MXIj27ubwqdmBk/sX13I
eyCZyWWrq/dRJn6cMLmPEyVmTb/CNNmUnt3rJzu8TCoO3Lmv08N5bIH8P9uCtwdn
NkBWvyFwEalAcd/7l07ahawn1jYN4jepTfycUL/vlvsmzLq2I6SE8dRjxIkeymf7
PLg+cKBz55lFw5VmEfG5qqrhqa+tPFCh1SYu2WRbIOb578vJZiWG0pTpjZYTvK+c
SFQnkcV+5ZzflkrqJxaHDlGhmvkOYICAW4fKj+yZdnDBznF7hPE4kRTvfNsWWxOm
B11Wv0MFFBB3LJRNJL7G2wRckgYX5k84PGgsyCa9mUDiHi6VjmWY3g6KlhsEE9ay
PhSo4of12asr5qe+rGZjK67s1+Qpd31c7M2IPA+YH5ydX7FU0oImqPuxHtL9+Uav
gcZu9tATgS4fU/gvC/6KvQJA3wxupt7+7EVeoALGNFvR+wTlYUnJWQHbN29mquZT
MwHG141LwI/d2+TT2/jG6kqv2Zig/7lbabrrChca2IZXqUB1GgxJDEQPKk63ZaJd
KVdmJFEAkvaoZyQkLyb8rbIeilmtlwdAv8MAw5otOnJiXlw/u3Vbx3Kpbt+GfEi5
0EzYmBDCyUJg33d2XA78Z8ea4UM6aPD7oETojEnYchYDglEh50UKgv6fsvK7MZZN
8DYZGSgdnAEXIoSgsVFK/HOHsx6Jnu/YgCfO43quKLWgstQ5yyoDw99RwD+myP6e
clLQx73uogLOZOGNZcjYWfo7swO2+L+B0o21bSbhJufAe5OKtQUYpVhtaR/0uk6j
o52x4H4WbF90TXmOHog8/41CdrJ0oFlZyOgnyPv455gYHdrldeE948S5M9/7/q64
AUCcCIO5ch7Um5PXi/fTYISSOPrEtZ1EN0pfknmw2qJvD5autnxaIw+0fTNL3/4r
`protect END_PROTECTED
