`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iuJTksm8TSBAD3rjqQqYm6UMXMvwVQ3VsADJcl3U2oRqIfMZbJKhaeVsVbTE7JXO
JuDs9ZEgl6L8fR7CuLrTmSA/Plp9Ef5WTya0lJywxpHpIQIHOrXWjKsLJm7Ho0O3
Sx4caNDQ2JUfo9O8EE1iTLgLPjtNpCV/Np+ykkK34LP9TQmnIKx1eBJwjdgQWau4
rgXagWpNa8jvLEz27JhOUp9cWQUUoCSqF6/uKXDjSb6sGGyjpqHRAv+vTuuHauYM
ytUjN1RA58c7BP9mapououyygDVTfprcGG4ON+a5jfIE1c/ddWldgwp/IXZu72jy
VFWjeI3P0nBeIpRFO63QFWf2MzNF9B8BON0c6qjRoD3ocngkk1cohktuMd0UNixQ
C1+qdXqoQ3pj+Q6jzhGTe6R5W0xWobWsR2B4X61cjFpHfZwnNNaV6hSUT2pKmcYd
bdfGx/9Ks4Hz2PqzA4tamJxMj1FIE+i1k5EfLWs5WVS1SfVVRf8OYZ3De0P8PEBn
qSSmMcmRoO5z+JbFq2UmgzQvBobfQ/NgygZAcIJELbzdVcjT7qY0WbPavoPe7vRi
XCiKdEjvl9CFR+f+zwlLrM4TJLc08kFlviBFwwFySC2GAfmznHqgSf7IGm59+Kho
JQ8GtJYZYDbBeKDcIC0V3Vv/iihbP2Api3h76B+3rMAR25RMAfW9K8zvfVdQVdC/
kjUgFHESddqPS/ZSMaD9u07gQXy+PWUkp652jmhFFCc=
`protect END_PROTECTED
