`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VE1vdquk1idMWyIfyQwdMf7XJBsLkKgiIxJrO6nrZ4kTes9HbeK3e5Xn6kmYEo0j
ADkESqzjPsYZ7hP9eskm0cFeYHj5NMate1NLmmoSOR/UlsSTXAHQCCNEyee9BLTO
HMFxU5uPXc49UqLJuDXnXhTDaywLyMXwvNGmQuv8+aNkQ9dfUYpWG0eH6+ulEU2B
ZuImJ0BzhzbqtV+oPHaRs+sW91MRLHUeaTeh77KZcKL4717L05yi8cDiRxFwv24K
8rniJfaIVCMGEMOnOz9n3NrNHwlhwjlJ3nUTsZOy00HOZGLf6vjYXjxSViG43sp0
EXy200ZnR0p4h+sG5Pgjazkc8O8jtxBNCLbCzY2W8KCYHZaB8ACRLKq8g1zR2WhF
VK+3nzZO28V9qG+QuBMyHzruu554cp5rw44KP8E20BERH+O8Yhr5eBzxENRccrPj
/j/ZUfs0fZT8xqMfHs7lHVfUj8MlDR5fsAYwqT/ORO9A5Ja+zFDa+F5KcsgoT+RY
sSGlX++E7CeGZSPLVi2Vg/t9Yawl2ClfyabOvZESO2c=
`protect END_PROTECTED
