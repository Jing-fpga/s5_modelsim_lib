`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JGdafmUlhU1/zyMZSy3rszcrK+rhWTynEpy1wG3UNIWZsSI4QOoSJZ1NpWkH2OTM
QxDx+00gIatRu1wYSG7eCPcL/5KKPFGr9uUf/dWqrf/jPaifOhKJtDsrD4lrAIF1
XxeH+Q4jdlGyscilih0nLFM6BD3Gc43U66bUghsCK1I+MaXD6ge/PZlb7iZEWaOm
t1vlnzWmoPpXo/1XAa6lEVNL42xn4oNuVxNs3S+2bV+lomX3uiRc+WONlXG96M7A
RYMNCWRc3S4WMTIEBNChA6G0uv1diEIVZvrsXhYSZgsspzQ6qvF3kxQeNd5Qb8qh
WhPkfdJtYvmOJHFpexP55ewkA36LSZGdOJnMluiYnD5mwa5H5sm0KBDU14uDPdSQ
7YecEmuo33udDE/OTxhMJa2m1ppmTRdYX1LFH1hUKWL1Mc0S7WKuOChibcEcYb8b
Ym2seSfOuIq8mond2GWCactRVZ4rxCP9a7wYiW5K2R/u2EfhpLYU4moKOclFP92e
lFg1vzrdYJBD/gvc534sc7qhfGB0n9I95dToynZAdYZuKxFRR9WI0h/5eTfPo+k1
fSK8xA//vOVEYUUrSajKe4mdqKXsovSryAAGShEGkQn6jOrvCclcbo+5GpNbVXIs
K7PSoD7Km3/E0OgZT12bL4Ee9usNd7NWkZT8CjBkuNnq5q7/7tEzHqN5WJFWH5hf
I917T0G3A9NBZg1uTFy0uHDK66YrvZ9OXMssPiwkJ8tCVw7R+AYU4epWPxSNpf/p
P4tRrlXjM0w79gohwq0E/t3hSP04+D/jNXKlgKtKrA71Jt6M9pxF2SCzLo8eeKZE
EE1J5SwEgfJ0vN7wbjEQ+ZD+8/zD1CMJSejFIM8ut6NdcKqFngKH56lGNUH1kvsg
GLS7jO2KUxoVEwMLaLrilzgvyoAayI+dc9g3IxJFBuvZCjcHukdTee096wnjJIKy
Y4D+PLNhb46yLoaHk/uBPVeG7cvVaTTacD5P47rVLSex9xFzrHFDV3kT1oG6TEnn
jUWgi9wu0yAdm4qKLh8eYs/J10aLFZhhcQYaZwcYNLj+VIDEXM72qnz5x6sPCkUm
n7srpyJiSxE/MnfbI0gD9A==
`protect END_PROTECTED
