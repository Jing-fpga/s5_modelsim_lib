`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bjH6N8ZA2Jnq6Z14p1V4U8B0elKkOfiJJ3d1yGFMzjB5DXHEVHckZAPInGjZr57C
lVy+M9z2hcK8qYJ+fiiUeg93j6wi7DHb5PtpRy926+L4844eWaKUXqVQkrmblVny
+pr/I3IUuAY4kIglKjttGCVknA0HSCvrbUuy3Tbz3Q+yZjwAmgINiy3nBd9mWtFe
B99Gx1GGeWllWAfE468kw2lRL7g3ZbBFZBQ6JViUSYE4p7chIkJDkNHK31RuPBIb
nTGXklHsT1XLGHuU48E1HDU5CBeoa/hXJgpgYeGXBI6baZ1XPB6cim7rF3pgDrTQ
JxaMZVcWouc9CNiNKFTyh1HICg/TQt85reKcGcCAbhMb+WlARdrUG7y7MSQnQ/pW
mInlEVs/DaWv9qVUJb+qeTgVev6wDTafFB8nYLH+ImB/hMl3o9tiFCrMpOWltPgo
9H0FL9n3rmYjddaeTjne0DbOEpi3eKlZLazHyJDiCRzlM5eU2C/T7N2CEhzD5x4o
qOCK8tqi/NnDnTEjFBTMhYSD7PQwGdZ1xFEiofW0FCc8q9RbUv55+M3MfpxKOUOm
QLqvYAeXoF860EV1ctSqqfAH5AyHmzoNz8OAyX3TkXGFK5HOwy9knHHk4PuzIIxu
m9UwHdfYRZQd+5nbmFEna0nE6Yhs1JoVnwnAsfXW7lixyqOkZYCStsUIqKqz+w0z
ddR7GU3nzlIqoa3ZofrdrCwnAeqbsLhxyU8gyv2uaIR71WDxyNIvyDy+IfXpjGsB
iM+nxu0/Kgiiu14PvsyJKXabT2uvXepAS9ztIRLUdNTnq9dDj7RvLTmsYnCW8AK1
jzKnh+hV/B+2bgR728824QJxKA/r2qlJGZsRlrAdpQI8C9firM0uuhYyU/nZDDbp
6ThDJ8/O5eQ2kes0apZXXE3DaqPUMZEHFvLhoCoaow82cx+t55CxggvoxRCp2JSC
BpDKhFSfxt1nE1/xFnUhwtGaOxUvU6K2cITMGIU9CJtt50rFpSTQ4tWvFW5sCxQC
OR3qHhyDV3/4R2C4bm8g2pkOB7BY3QhpMNdawfFbGeJkXLUWrYL8cQm1UPvEA7q/
GLz5J7TSP/tKo1I2l0nMPpKBWytxp1FD22mShxdeoxl0L9t3DlEhokZJqfo6l3FV
C969c9sJOStGAJHofYLEPA029e0i8RVm8+M1PQogDxYKX4q1g4R+aCLf/KwLbo9H
tW/LdX0aCPKrVbeY8q4Y0JmvTzy5eLkbV3HLvupbBZSHrHBIavxJXOaZGPrbtPUP
LJRp6WIHCcAFDytbbamg5/qjxhfT/eBdHh3M5d+Oc7jyHlFDvLeOp80yAjqPsM1d
pkksityVE1XAl0lFA5PuaEYuI4nj28Q+mH6gmqyxcSo0fTiXsN0OhIJn6Gb1YjEP
w0gLLiI67KFrpLGnR2GKEgxWRJv12ziqroKIU8tluc2p5Ip63blk5pNQIai7/YR/
3+xL/JaPeZlBd81VkIAm8d4Xd9iPHgzThU66vxzBH6hWkI3qxRdCjGDPMDK0YeaG
FrhpHkwIOs0YqfM67Mi0qEUXOtnzzZ+VSj7tHNXlosAgIRXqaY1AxUhq3jCCnR9z
ynZvq+tPEatVNawUzdy91fBWgv/fzlMFrLDRLSxLUZI63TWYPuWnXHZ9O7G9s37r
l5pAUhNf/EbzVR+mh/aMEbBjjV4jjvLH850Sea7Q0mMb5cvQCUmtHHMd5QF3Nwpc
lsg6csXvoSbfJoBRGSDArhfXajGieCWUghK6PwqMOG3Mnu03e3quWfZPgLpHjmkz
J/srmq9X5ARLfsiOTi5bYE7fM/UtZparQ3ZOPahznYySCyOkdXG4C7mFpY/US6eL
aaJmsjs2MZn+etzCBulGOo7adohT3UKx3SZZ5C9Tc0m3LOwZWFA8cQD1ZXV2bmCy
fB8H/8KDplWmjznlJpmshAXQOJDWR66meewjPtYwEHCfAUaqSXJwmeftJ00kOrFH
2HjQzvzLFDejXwM3fiuWLDS6VHO3LQQbAhMOCEBjsxGJOtqDl7jTFEFqsecnD/SM
pKtKz6tezb1COKVmEpCaGE4aD59WmUJOTTlkF3LHNaK6E/j7FrljKb/i6hKnEuDw
qpGaftwbehrOJ9NhI48tI27JdhljyoAdUN0c+noXrfQjCxXGXeg/HvWyRioYG0ue
jq9A85C0YRDo8cjRytu5jDkdTMu+bkpDVqYfb9S96a9dE/nQrRcjBgMteO4gdOpA
3+ICOq956ZjZZKn7b+CtjGUzNZpzeZl1UU1aE/xg26y/BKvaedpgqfkemzInZR8X
WMqqdqim9Owc3ce/hIRqSjjHkiaKLHsmC5k0jBk2AcG0Gie0C2An560fIxMcnf6T
TeDHQ9VbwtfVhqoRAmb4QJ3pdQ0oeQTNF1Ra5iRo8MejZcKx/BxpU+hyd8hOPpW3
tH/Q/NGRw5fwUkU5jJM3X18JB7dD+2eTUuLS8ckuJ4tVCqhtSIIrZK1H4CT0mCpy
dImOURfig0KTfsPluItGnKNjmplogzZnNQwoSlFu8WWJWDK3YzDP2xBPhMMKSSX1
T9tILJBZ0H3ra6D6NIW3pBfm22WlzruzBdOQ92Tgo9yQw3igqvlPMcEpoOPawfuv
nwkeGG44T7QblPAI5nzyTNN8zq+jd1tSeEiKWPGpd0jNsbhLMFNn1gfzH5ZQKrdh
yqev/pTYh/D+Lt03/kRuBe9IhYf6R/+sxNaTN43tL3OETEyCaRV3FGL7UIUAz1pX
KIUV0WR+H+sxQrhQgFHMAeEBn2GluOkfSE624r70gLH70g48y3XlHwFy1/Ufqgd1
Ba+a3k8bKl4qQb237fNEkGejPICGIojZoxI8ynBn65I=
`protect END_PROTECTED
