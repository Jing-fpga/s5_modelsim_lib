`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D5u9c4MUMqjQUpxmCNvkfkpuwxVBew/RWnbd/j4sCC3f4Efil7cu8RndXmPXTfgd
JXsh25Que7/wuCTOPFfoc0/WMSgM5AwbcgWadm4PTFGMb/m1W1kqO0flPgtNy2Np
kVX+39z+nvZtuuEsr0gdCWj2ZLwItdexsB1vTJJ96jxiHFMc19ir1uNKA1DtfCjn
jlrzz8GgPV/flQif0vr5PAZd6jOy038XsnVrTlNeN6BHh2FTtdyM/LnJJL1+vocu
2+Vn8Fy1Mp08A9WxxOfe7y/Ij4y7VMR8lKf8i6YEnERzMMl0J18AXMBwrCx3Sta1
jONs4Bp7i2TdLfKUa0NWrl6F6433zsTmMn7n1Gxg45H1mtJ63L0ZiBRMANU82QW0
mKrsTtpwE07dNKHkLbHz+3ozOTwk3IOdXxeOxftbJsOQzbNdqSmGxDB4JKn1GGje
hxrHEDhV9NTd9OCx218htbviK7NQ1UYzhS+ojnpKmBhxZBfv9qKkoqI6K3NgoWft
EhqZVhb+80B8yNebLYQNSpP5b4dMBvYwyHZyrkof6L44ONNmsQ6KZ2B1ublNVyUV
IGHgIUWM1fNoJQd0uIAAuaYGnV2NreHvS3DfbtmOEOB1aQnxiUOdQGUuHtvNko4G
DR/oybPRb0FY5HNzJaUdITGmBALI+Gb/Pvmeo9fMWT0p8b/z4eHGSA6J1h6Cppcu
eiKQmKOsYhNfsuyufq6xTRQdpjIRRc6CJTuelIAi7eVwgfWnyhcK/7gkKU20BIqg
ak/BkhRErUcvJnyPgcai4QGF526I6M7x078jQq5J9RDGE5WdX6RPYFo5MEs7Ey3j
zRzM3jMuETn5T8EgQO7ieIJ/dPZQpneOlFD4nF5LQwhvG47iQn76YOsajgVd1PYi
DBKXkItbw7c7q/udpQRfal46NP8ecTBCG9Uf/ptolWo+XOEbdm0xCFNN3ou0XxIP
kSSh+1S63q1Ju7INChLDnsAKS92fg9s5t9k/4//nbgnG171VZN1dLUGbWHtUUjy3
TCQQbiSDr6sUgTUTCCFg9K7lHrbz5hJvyzBG1HDDdAZ6rDQm31ToV8GQN2iq26gS
dlB8eFss0zUf5sWLTHjtxe3RNyvkJ9FRRlkGk7dUmbyrJZ4sIebMAVYc+SiNSO43
DUsEN4aliaAe6WUy57CCzUhGtYtx6QOwl/h8I2nwdoj518V5aTL/PbvwQle63iQD
wyuK7BPXRfwJjaqjn33iZDaqxytLoFJXVTGUj5iF/Msn2lvk1Uf85eXeWJRnLVYW
`protect END_PROTECTED
