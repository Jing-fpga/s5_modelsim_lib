`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MugIHNWb9WyAlvZjMR73R/TzQfLMzTQIoe2nnia4HzJonEZBjymP/str0mxngfBh
N4B0A1PNWtGfL02rW98aSVS1ciOGT0oCbFRUer9sV/l0883xA5Qehch/j6u5FwSQ
PgKiqzoUf13VQr6rjceCRpberep2gvUL+a8o0Wwup3LmR1MowlK2Ps3X7h+TIYf8
QxwyL8bUP8JdfLOErTqoE/CwzFKTzAZGOkuiTLb5hmY8Z+K4w9TqyE0RdI49brnB
3D0zRRGWDMlV9srvtFSVgH1fjL1fr3F6nt5Pr3JpNv55NKoc6Dc7Jkn/cNFPqbXW
8b72bHvTNWv4xCx58d0oz+H065iSAOLEfAMzz5b2MJwWC3idJx/5CFYPCiuXse4V
kycVtUSuMmi+q04fBLsvg4xW2my5SZPx1easTjA7Tk57R+JP3ON77oMIkaJ2kich
rsH2qNNCmJ+hTcf7wOO5+JdGOVFpyAJo4XFGlhETgFGtBplk8nhK7fMknF9QUwuF
LUVCYTCbcykiVbH64Pz7M8Ov2TdrIurPMZflWYR5jzGROwu0y0LLHIk8geKXy93a
Z5e7h9z7dtGUKsRr2zEcbg3e96KNvmIwHqf11UNpL7XYWrsCmJSae5Tc0YuU/AkY
V/ct3dN1QgHWrJGOTKAfyQXWzOTVy6rRITd1OS1z5jEWe0nIP8YUFeGL0vdx5V57
SCmgcfSR0yNO9IGUdlUpITWdwW3hPcUpMEizZKLQnFsmK3N4lVSroMbOyZ8FaHgA
tV9lkMC2VIaoypIaZThnTuE651JOsPnPRp0HqwzCrtKsbzWfTCStmPtqcKLI9Te7
FwZkM8EfqHXXw8vqzUfpIByP7YGffb1Nh4yBglHhdwY5s1o5ROQa+a+BbMtbqpKe
ozq98dvFvGns2aIJqUwOAr6OsDsyReCswRrSbCEaegXs6659de7dOzfkwlaOk8f7
gzQdanyjnXTMYzy3wm6cD0hsUiQayIzjvqXpEW1UUqzUUuxztoE7INYMmZSZ9tDX
01jONHIjibSfaudkp3cHfdaRUtCSbHLwKLZBCyF6uEHCP7EJedJB4H6EnP9f6jzh
Urs0WRrj3kW336kXrSKmXg==
`protect END_PROTECTED
