`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
56gFwCUc4KwpaZZ0NDq+vLa2cVuQyozqm16k4I3IcJ+yvNpRWESuBhNgPMDPLfxb
XxVQsQCzl0OWExOLSx1WNldRzhLupHBTzeYN0vPkjMQUIXWikz/2mJH1ydrUqr2Y
EbDvWpflYvWibnRV7XFm5wTehL9NQi6D1ViiBxD4tUXOX0kS5N/N8QGWVOxij6Tj
+6m6bSeTOB/M9xGMSMV4ugTtTslh++BW5iRQ/F0EHpuY5nal9JvEw96vjaQyRma1
ZNq4KeQ83EsK4l7tVRVpI4Ou5Zy65PAlJYjepThX1RhihV88z9j81NEpPj6dYf/f
WCG3wW90rTdcIei6QwCcZnMnpj1mQ2GYWCenDBWPEj4wuNovWpkgyNz0xg3oJaM2
KKb6TeRHyqWs0YaSSiG7GuMZAHtNI9FqgOYpgD5vFEJRZJQD1hM4iNuGN9oWLllS
ZZpLm/kkfg8DeWz5Qx1kl/oJ/lhI54zCkBcibIU7RSzGvPBKu2nnscLbx9PgJ7Ri
VKOgTXcpqShzvR5nCT21iWAS9vtOCEd0DSKKFF1XQ+3lfBE1alZDpov88aMf+iI+
YJJCDq/WD/929tLhtUM8Ov20Qp1eEnObh645fnIG6JSNRK0owwoIwOCH+O/Cd8gQ
EHoWcsZoDbGdxiNvnfD7TdDUXSqH49CrExtzxM4W0sCvnpd/nKE3rhhmqUsVj/Fu
NxntJLkz756E3WsN+lIQ3tRa6WF5Bj5cwShGCp8fKzb1N7/ZBMuEOUBOjtIQZ1Sq
iZZwosgU9qMFy8Wq/Lkfb20+eVzchH8qwfq7md6Cj4qtsA1FYhW/Lgt8d4YqPrco
j5/ymg91JEvlxKZGweVPKU/M4Ez4AnsPXwnimOaooDqFFJqinpE7Ue+uIzHyeHLH
buax9BYQKd3i5/eFyixVXe0i8IU4yG8b2MjRT4SKeCVWGNE+Rb7P6bO27q2FaeiP
YT/OeVq4F1/o1JKWMIoFt+UK4Ij7KzdvflGUJh94fRhS+G7ruPWfo2OQKJzEdqFp
e1EfAAYEJQM4eSaPFo9SOB7fCX8B2wh/xWaGzMCCG1zfDZfZxt94IC/JReGlxjpF
PoTVZLxJfGZSn7N5Q34OHCjvIvnWbk0y1y5ZBuglp9E=
`protect END_PROTECTED
