`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
odBw1CekVX5oRqjOZSITgm996g+/7Dwuew0EhSgTu5RIDFqRu/iynSAEOk88C6dc
X8bz2D/AyTVg0iKKLMati74Fq2N0lzDJFN49WeHxZdTx9bERyabYAg+V1WcMBaI1
E6G1BQvpShCeIN/6deSCq2jUU8NyTLlAFOIsP5gPS417m9J3H9Y7MIuBx4SNm0bT
n40QMipitw5iI9Ta4B6L8aR82AJbRZ9NQU//bbuRpKjQRwqEmEbsPnrFWmDahY/f
U+I9TVByx8RAU8d3n8FavAGPlEmdF3jdMlYPUZPKqEVEzr7pb6AjCCrOFBPGNcBx
KVKzF0/TFicKltbwRS5yRA+hg0NTKexieAV42zXH4sx8sX9LXsDjz7etCSfKCCvP
Ubdlm6XrEMdPV6TiXOl3MKRJp58E/Q+GsFcneKHxTHQ7M545GZtlC6poL+wDiKJk
JFgqhwzoDdG1F7rsu573aYs6Nr43mF22UylYH/O7OA2rfQgoSv2IeaUIixCct8w8
cW4b9nSE+j3W7GB1KYhK6ZH/CPM3tEiuPDHqwa8BbPdvETh5xxllLePyjK/lFfzi
VLR/3QnapZ3yhVJTFME2yDsL1/Z/FORf97E8GH/DvrjHGW9ebDRIl24FCuvulN1y
ACi7sdo0egx2H1zT4KbDcT+i371fxLnXmQVZHMAut1JnmpERzYR2qdrkIiUmCOZe
pQ7W7KNSHLghJ0lJaXPijqh7H17ns06QVaLBJzQDb58UD+S4ZKr6or/oK+KOPI6U
SxFf1UH2MtbQXOMAghfDaNLDgTjpwKlL9XkGxzeMYXDr/yGqoVplaubwfvtqSKtq
zZa7g/b3R5SwYkmUOcNXU4L2AD6ZW1RGL4KQ21GeaPbjOF+ajl58YKeBSA3JRB/q
14K0LNnIjXZup8gUxnaHmcRJnVxZxS4ZTBSleZ+ZljVPq5U5d8Dv7KTRoJJgCJcX
hDyh/3JIueNySb0nPMIsEPwto6CQHBEcVUYk+B+OJUcC2FL6novkPpzBt2ic/EMo
BoDuB0+6xy8nORooonWpfibnRZhAc/a1ypRX+klpLsqUlDecTq9hP1C3EzRWMuL4
DfLO6r0BLtEKNIOQjiY+ND9ua8+mYtGdtmxY3M5kfgX4XQQ7F3qvUa70YsRRk1/J
YNX1klrHDATvsQ1BuezvrbetH7Ss9KTuykOFIioiehDjCeVhu1n3TOe604GTJMoa
iYPxFP+AHpVWs4/ETD/t+Dbo34d6Qszpn9dihSXA9CjLm/7V20tsG7BzK9LzRWTe
aLZncAsOvNkUOyVULBlQiR6pEKD51j65CUzD0kAtVQNVAPh8WSUa8BMLPUFbZ+TD
IJyFQ07fjyhF2189VMuTmjMZU3sAqm1vAnkyaZTQOglY3Qnswv0m+FBV7En7g+mi
kxoz5fRozNqqjHfSabQxx0T7jKfe7smCE08mKw+s3h7P3KWbo01ee0dxbvoZotcV
XCUPmXt7t7ceiKfF0NykqRvcjfdr+3oAzCq5wXjYP1gUMXhv+d92DnsZaglgRgdZ
KkUoeTmPG14Ovfketj6HEaArpn++s909CH2IzZiME8IbVSqgfrmWreSpxUHT5e7i
2+zjbsqGamdtJT4eFFIDipm8WrH+Ua/3x1hog+rO63cndUzr/9retMk809n2q8k5
Yw0ZMqr8N1xjQf4627Y5eOnpGBaGdnsEWMz4NuGVzF2PFTY7bRGinBU3xxScmWrw
CDFIE73ieJB4RuQqpE3G4zfdu7A4JkSz0njhytqGcqudaxl7DJFhAkh+fShi0wvP
as7qDzMDtJHL6NAx/nMWgayp8igJa4HfzeSG/ujnJ/+FnD8KE5E1LMh3qNzVfVLf
yyDN/PMPvIFxr9GY0Wx2mGjo8BjbzhBLrhB1xAp+vwTYUD+DmA/Vf7tSUa5GaCL4
9C8DqtzqWMssPI3BaIWEkV35s8Z+xzVabv3bZ64zJX4vi6bkDgPy5LMsXpfGUisu
zMuo3y/f5dSGbPh47Is+7tVjQxH9ftSXFKOB9JYMAMzSHbmHeiTOPg6D1V6gc2Od
MSrN4RKJeVFmjDHbpYqSxDGVZzpwN6J5X2FOESCxC8QfHBy0tk5FDDEjD+xsogU1
AZn3JYFvqCNvQJn/DDInVyxs01JIuwTipKgkXUoRGIxbJQBY0vcNPBrjFzF3C5uK
a1VqjzEcWNusVoOayYh4uzdpz8yc8e1eeZyjr/6PG2v72Kv3iLs/n1wVLkv7HW+i
Opagre5veOHm6UcZXuNxD3UcihhPuIpXgsPOABgF6a4bYlzUgGHPDACuUnYT+Ur3
YulGpke8nFZOpmYZAmhe/Q==
`protect END_PROTECTED
