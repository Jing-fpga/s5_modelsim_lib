`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n0h2+aAx3l/CKx5RnCw+g8tkhg2vZlrE2RtjDimyvh2fMnXRv9n1OY7YQ7hfYhcx
Lgi7/vBsoXbArY5vSyHkiupMCQhuwg/CzduzdWf77zRJ6XwgaBsjBVemIg/NSgmT
gD2Wu/lU4jGz9hC2E74DgIvX4vQtabdRtNtqeZuLtjkoMnciq0r+ctwF+hPKUFo2
0Mb1MeFT/d9ZeIX53BzNY/gLWN/ltCOlKLsNhRe927+UDKBejmpmEaaovI06SDmh
5nJzc5K26QdloN6J+k8y16Dv/RgyqakU55YSFGT6oL8ISOpPgbE9IxCoak9STHlL
O3QRF1txc6SyJVxb+WjesJrcRJrBEyFrNkI1FNZEzPCLZlLPQavXlTEtQtR15P0x
SEE9Q1WOe7R6X/kD+kNZqXuJghUg5tSOfUEezChdHXy/jhUG+kpO2FgEpmNYSafM
L3yBS7lPTP6OoivShBUk5fpawEMy10uSwKPPachkow7c735gBnyhSWJQIPCTG8G6
Q/fcs6TPBBDQlMPjEAdxjRe+KiVXcl6aIKpHdclIECrb/ED9iGFuTDyD2S1z7/NQ
YU5MIuCqW/AY2hCjHpE8U2M3YbPGIjYkdPmdAPZO/h8npYQKTQU7WNdJSgmNrk8y
AGOivb6ZE8WfLzpuJa0Rl50SLw4UXQfcJCZkPr5wVct7PWJILFWUFQJ86KpH6O0l
4hEg6Km+i7Vi7WjjUodMpynAmPbRPA2fVKd9xG26qSsPVspgkT/kEVyptDHfgVGT
RQC1+R5dxAzOgg4qQHIHseOJ9ODzsKCgoT8z+BwnEnouEYgVTTgXZBZxPcYGHw3o
uWGhlaDCCU+qCtRk7YW48u8BPubbIZtyz6iJ3bWSJ3MZcSwLWsNKqebnUkxb3oqN
DTM7dM+WZUg26FIey/C6fvXTJkdknCSbj7mLPj7kG/r7J5Igc2PB+gaXxe10YLCe
z9/bnNLiJJ2bKI7xduZyqPKqKOJbpRmnuS1VlsEp3SyrWkb1myQx7uEhMl0O12vv
Urg4i6Im+hZxAzzNNJIEcfcXCn4OYTalOkchs8crlifZDLxz/ljPwFID5cPiTWK5
I/NU5/DMWl6IUYwIkxmnOGIagiNmp7ugspZDOLo1GEGikvJNYvR0Vk0wBY4fjjCf
i9tFY0RRYbKc/n4ofSsMnCsA1PzlUf1mPofqxXhBfLORKntrM96tjn3CnmaZvfd7
tJYdXSvQUpQ03KHClCjxCXm3tLSe2qLH5ZxzUa+fHT/BZadppaLOzXELqnDIrF+P
Dlzd2zG2YbGQP8SXrnWBKg==
`protect END_PROTECTED
