`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oLrEpJ5RgWns9K6zh4Yhkk3H9yPTo+W7WeYX5ONpRBp71BCBActqM60liReOZ4cC
2jDod5atr/CPbJGf7xWKQ+l/jSo8+3iLIv2aOok3KSfSGcmy4w2eRCm6Gb4K5I5x
MoYq5dNq89KSYifgyEUfTKsP85fkwDWspdpau3aXpbKZtLIDFK+Rpln0aulQeQKJ
gEzMoTQQCapPkWvUtX5/P3jgCMYrD9DV87rC5kqFQEF2Ekur0RA1z8RBPebnxSFR
EMKmavap7N98e420BVv02Yt/m9cT/7aZpTWhAHfSY6Hlm4Rb5s9SMcVHovIo1yoG
Um2tR/kskS0DuwMnDT5GvzzQthBo1J5MtQxfQa327yoWznt3TdHjzuMyI3cglS5u
v/QD9TVApH7dwuXlTW48Oy95wxjo8G95GBXXOhS2/NFozwOKusH6CrC6EDXDU7Na
gWNssIDz1y/8MOtX48QDdDAP73DYgWNHTmxNSNu22R15fDAhrNYwAqy1Maerurw4
+iRZqlqFnLjZ7TTo1Wfv6aZOFRKfWh+qdwQwqNYl918kqvQrAdkoZWJ0P+K0eZ+p
gI9zIO5MHHpzzWaIS6QFIDW34QTcfc8ymsrEfiVLyjzODEBqML3z/tNxI4L6rdVh
Ipx3FBx3ojFTw6Pz1gj0kztXsWwGHCenVLHz8GSLDCZYvWBVCDBZO9m3tQwkW+M/
Bptn/C3mnf9WSSQermlxo57FkOlIDf1L6D//bWvN3MvVWucMNcQat5LzQxJG61VF
HbDDCDmwRH1sQ5A2gHehpwMiru0HfvC8lCEc05CdW4u+2LQ25f9JDWQSqgYnhX8F
Q7s/zipqWZgtuNl5h6kN2Q==
`protect END_PROTECTED
