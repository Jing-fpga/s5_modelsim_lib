`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d50ao1eCCzDS4PorX3KyxM9ERDO49mxs0P17TWmSvOLw3G6i/IxYtruYD9xtwjeW
Pb96PdmYKlJ/9Le2N8YkX/UEuys1TXngwpfaLcPNj3FELaf4aJC/DbEICdkh0H9G
/V/bag20YNFB00MqE+KjT3NIkPmiH1a4FoamZBNk6stq63dJMar+Hz1aUUOs7+VO
68LgdigkZlngyF5ZnEPv6+X3G3JnUVkiKdJUtUEV68w2ZcmrSvWWGKKwG5zn2a7x
qOfBrtZnJ6lkke3Gl8GBQCnrz4lT8UWyPenJDrk6HZ/qgCxqkwi26bV5hKjpwzt6
i9q9SDD9uozcQ5PdXScKXZ7e64ZQgQ3mQzWHP/aP5u5UqLU+6lJMNVyikoFMw715
ZP80duyLDd6lAkxmbFSyCw==
`protect END_PROTECTED
