`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FCkzroQOSJ8jPpWN8bHBDq6m4mHj5FG2cd5z+nVH1m763tBA0uxw1p4/tpOuQVOP
xrYXMSv0OB+P8CbT8y0E3OhjKrdOT3uwzzsUprk737QqtHzTfYCn01r31ESf+Xpj
JTpWJhn7og8TAtMmLIFcW5dUXCBhTCHlc/PGVrB+wGDjKv0jbXzRxTbJ85bU51oy
ojcDaAH51mKOnVA3ZgO4hDL10k29mv47h711fIJcetP2DVS6VATdbQFMYiYLPDCD
/QpWaVPRpCMQamKzddhl71Ejc1QaQmV98qei5v+u1B0apVXf15oQwUsYpBGPMwTX
6qWgGYpArvawbome5YKvV0JdooGPgXUYLdLOThxTF8J6NUah2BabO8hy1Ve4y8RR
MzLe52C9WfAErn0479YVyLwLKgTuGjYlJllyAzkYAceQvbh4m+HkCFH9JZDARu8V
LHpvsFYnqPbLeUvzaYF7MQz103veiLkRnPNWkEW9Km01AlWHS4wNw9Gyqqi3W13r
UffpOHBLENp6OkHHsS7vFfphPIc8Zfg1J7wyCSPhoy5kN6VTj5tTEYBs6m653x7E
u7s2/Kb3n5Q9Cp/WC/Ldp2dEIKRz2Ne2vGrcZoXFILXAZMyR89jGFaCSDNYcGZFG
QhUuCaCr1hun/HXCh743/y3HN1RtNavMhGtiTbIgOwz7/Pd/9/vmturcCqN/BGLn
HuDzH4vukxkgFjy44XBX762xDd/Musl/9LYXL+OolKovS6CBtmL6WJUhNEuYTJlj
xpmoOZ3091dpxzV1uCgHDFsBG4zZ8G1W0xX0pUX5qgntr9EbIRuOa7xwdWBK8mdP
WQPYXTQwpJLgVOZ9JbvXvH32GdnVGnR9yuxQdAmF0JUZ8oPRAddjgC8nTesUqzGq
uJVsOI+4uzJ6htX/nFAKTUs0lUB5klW6JY/f4ViPYsHCzkszQGF3chYw/HEHxeDx
BB+P7XjULbQ72ojWexHe72KGHvWYnyBqWbmWqhuYh7fLU3e8vZkAi75grfTtQnXG
YamWyZIVAkjw5W/pztiHRfzSgImMOsieNcd4Sr8FZq4c/xcjJSeJgUEfdFj1bgJS
zceD8RBdC0/l+qrCvuYbCZT5MqfrfQv2/Jvmz6juhUcEiEL/KuzS5F0RX3eehVLP
u+v7zLB0Y4ycB2zLSh6L4UYBcdgJni8wnBx6Z+yacLDkHRq/y1qspXeQSiD1gCPk
uyBI5UlE9cdEAVwnImQnimArULVQY63qsMORnvBH+HoaIsUiUErrL2YRe+8gwOw6
`protect END_PROTECTED
