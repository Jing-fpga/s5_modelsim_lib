`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3E2NSgIPhJ4zY62sSeR9iRCbRryf6dqhWTouzLGC602nJTl28EyI60VDJP51Eihl
9LgDZfFY4yXYVGSKl1j6OtxiZfu0NPeqc16nD3tvoCO+EHDOnMVQfosbktsjK67z
nMI2do8kQr3CZhVIK8jdh/9QBI1IV8pv1vO+X2nnl20efLW+6BjNhM0RjaOzzyc8
vX/yfob6UhBpLksvmcsvV8CMNFD7INFBZXxQuAsEb/1p4pA1opwxAJY+k1k6b3SI
n02D5z0e7+MnZw01jtzfshP8fDkue1d5h9uTMFRvpb0b4JbOA2hcz2troaPebdY4
e/MxAm3rww5F5/md8PMh9ay+kpbZqQCTLqxCGTCw+EKk2oY+y+LP41Lo8Js+N5+q
ILdheGYp/KuIMMmXaNE2R+ps3txxOinbnwAXjVAmn/vxNKbCGDfdXkszOjapY9SO
JYmoDXHvKKGjtQlhf43C0UeXzbNvq/j3B+pRxzvu1LyjKqVCBf62ThF72m7ZRv7z
Oa4+iK8tIBPfyF0cpfcMig8FFycybVQUYs0aLwrRfsk40gPQEDyyzbeqqYwQJ8Dh
wN5leUtCZXzQYRvgTV8M7uvbAGXPa8UL5G6TKiQ8dggSIn+svFgVNDh4Q6VZiVTd
8L9zcq4W/5sRUjPE7uC/kZaCVEQwZDbNlBLswuqcgpKcH80OMWe0MlvnwzCdyl8S
NSpULMb3ayuRYF3eZeUBvl89COiSVvXw2rklQlWu39WoCDFj9jTPgjHE49UjbEku
KkA8b4g4sg+OJwgjEcdvAqP9czQ9fVmrCSVpOZCCqj2wk5JSWR+/uCKWIS8ZspAJ
Q1aNz4HCWDAImlsTGcrQtgGViwq+R6jyKPL36InikqRex54qjOxTyfgq/OAy8umx
I0X4Qt6QmLSsE/+hGFHAEJA4zoRUQCF+E3YKdoYsvrROQY3lQDg3H+ovnVDD/2P4
alS/c52VMIPqkGN3JdO7blwA58w2oxiXxoyfGcbNLPewISvkKUIycQNsEPbuR7Y9
hN/dJBjcHaX9tkIoTA4hBVMFl5Weaz7vFNb0gyYFlK6L77gSdiCVwwc7hTQjEB2X
R6WqZmT6AVB9HWkuzUvcr2Ga/7BEXjV8YP8XLPz2I6jqDZaDi8MxUW6Esx31cfT4
7udJo5IYVTAzORh8p1ff8scvF9ZQKk2YC/8mjMf8wYyD7n97UhfH3ufmeRzZ5vyi
ypc2uTTQl1oP5R8bKn1XEdMEeb4GGrTfkLcXym+T+jd3eHsUm4hOOTnfwjI7rWEl
chmAv+F6sSHrXpTIMhUfRkNuY3AmRh4a7W2V6ld8sWU=
`protect END_PROTECTED
