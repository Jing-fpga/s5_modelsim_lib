`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wuB/TnNEC/ML+DkI3y9O/7wjzk0hP5xcEXkM3jelHybq6+9RCLlFUy8BgwZ60xXd
gRHXq2j5DD15FOlzSDiGZHa+iqGUZPN8o2Bz0MNwxai4q9AU87thbAyVI0oTuZmi
CDzuAoDEIQZrgKa0awgCjqh7EA4Gv7VNr/oWTC71cK5wHa+u0eQws9bw/Mo3zK66
u50smkOliIXMKt+JjG4k/aWXr7d0SWtdsEyw2r23FADYNCxVRwIbZedRY7Y5JLKQ
/C92a24NZ82ujWVO1t/Zx3xGGs3MoM1RAGKX3fM7qzu0S9OHYhVd32ERxqeu3yW5
j9lKRTwh2QrnU7DVAt5bfUbdlJ2tvTqaHYU6J383z6fixeKNtZjV1ZiJ5ba7/bGB
fOBhuT8sbPrdsMbgGr+U5fES5Z6xuCmuJaGdla60eIjqa8Dj0Wk0njQWcpAe+1fI
4I9nWsOSgMiMzGSS0HW6PhbGKCCMmQcTEdRZIlteYCg3ZDjfwCmjaey+M4VGPzGB
0gpKTjbpnc20AewWsT8jgPYkeIn7ppB5/FxKyshMSq2B+bO+ngb8cyjSR3phpDKb
URTQ8tmj7j2v1sdMsb41wzGx3bDRqPCMpIykBScjOQ/hCkBowkeEPRpFUSyeUtG6
gdi4dnTV5C8XAuc3ZAFondkyjoUV4jdokp10A6KS7je8LFpG8XPMHx4B0eNEtFfb
PSdyPGb30+T0PL2jMkL3FiLULyIO0jhJhG6/6qWm7GEPw8WQljdMKii8KTb04BxZ
+fOCcRGga4DqXnSy18m8q5Aq2LpZhTqIBTnhs+oHmgG3QmqZlElPoVG+nos4cJZF
rNVXbRG75O4J5lpBYi7XO37v02EhwHvWH1RBEM7SA165VX5DI7Hjul2Osm13py3e
yEeJOw+n1s4bww7c2iuahnswcoQQgvlcGPWfRf/AIadp0VBELb+OIB/zxbcrbk/j
Phz71q8wQ1HT1OoN6RfDtiZT+tn6xOinEN20+2QJbDzNTXmptMIbbOivNTAkTNlC
66nipQAjOtmuVOR0v7Bsc775iUqrjJxUGdWANqq4GRyeOR0rqvx83c7tqnnd9eDE
m+k5TVFJcWbIw6rY/x4nd13MCG9X4KBNMXFonv3ToaADPUJ0gZj7MO2IDO+8r3xE
ENHvv3vFf2AAxqWVM2RGaGdv+RCDi6pL1nvEJxsCd+K1rSzEfCZIuc0YPKp9bN8v
4ZH48NKa3CuUpghzrf3/TDAwFRvBb2YTMz9E5p4OZGUMcOTavkqWqpxAGzQltDgq
qcYV1fEFcbU8Lxh+qU1kCf+C5tp1vne3qQjvkCKCnERxxaIVe24TO5GmXSPeefAK
1aRt6NzKiPuQkygRoSrt/EgYtsTpUDyjwxp8G/EP4huD//CLWt/7ebfDhnZAn8RT
MnCQ9Kgc/4s/gJrmyj01U37G28Yj41kf2HomnBctEOUpa0Fb+PVCOUaQjJC8XdRE
swvwrSdGlj2ac13/FSYeiVBaxU761na4NtPRlaa+UQoSYDXuUvoUTJDL1It5b/PL
NVpkQzdaFeIMe4q1UmX+YEVY59o8y2/sYI/SazlJEHxT2gVUzFXgmONplBI4Gjii
8ZY2vKQXEPuPf931ZlMzYG162vu5ColiCv2lmzjR4kjDJDC3cmRohy1+UZf3a+Vx
ee8OpYPZy0Fx9wo1oP2JJ4Tfl+mwrGGFVzO3/G10P9+rZG7pi3P+YFOAWacFerxV
kT+ToMPhprEbD4zL5asrj95G4hCVfMvy6BUu9OCRmpXkdV8UZjXsyka38rWGDo+b
93qSHam19zcS1yXm87OwQ04kLpQvb++PgQ3uxwfEZfCVYvM62f9js2F48fGP43aO
GnyOVbTW6H5DU77uYR0jRMJ00Z2M45CxVq7u38p+iJH25ldD9dWUh6+1xotHqmgh
Ek+NOMPopTr/LQOeB994yZ2VzdoF811Nnr9cjsUjLs3cQ917dSUfXxCUN3VM/lMc
lHO1Ytl8r/cfU2Ye8toC4Sr6cJ+BC7Uwus1E3zbxBOim3DqqzhO8egE2xiInIDop
yBoXSsW1MIr2u7PlMiB8NNW32DqKQX9Px2NB0KxMmdtVUyFBGL5FVuypnLqVjT0X
h9D4ImhNoz7NCJhz/E2szqxyuSdnNmxtI15F9tOMPMH+/992SGkEs2hl7sgr4fON
G8BmonZEkgOYkzX2BT9ZqCwN4t78TSBR3N674t3341UaG4m1i8kLMHyH5IDEtLWM
tIMIuKmW2ma/I++mZbT5Pjc7f2RtFltJjPcKBRud96CT8CP7+X1ln54M2uF2xZen
7A+1qb3g17AsH2g6nt/K/5HJZtcrzIwuQtjdquu2n5OhfHBMM4vCIRAY9DuNFAGy
vjnpQvNqjyRjLE56ndJJnjq9ULkfleoENvu23WuUbqt9+POAVrZuGamiMjbjGpkE
2yGdjhMIhfMPoKBDVrDLQfXyknq2dnamAgu6ERszNVEw/bG/qkmulKaQvNbPWDAL
E6+hj3TLMxWC8jWVlwgiJpVo85KMONuCUzHCdW4V80KJ7RHGcNQAOqU67Q6PvSJp
0ewuHL+3DjOXUKahWXC7JhV9+I45T9yP7j11+6KcvSRTEvahVaR4bFz8gS8grt2e
u8MesIBw9rL4H0aFyCqGCQQtQw8bVYe2pLsM6yW8RqQVS0EpJ2mgY2vMK9y3NEAi
0oZ/FyM3yl83Ua+Gl9Fohw==
`protect END_PROTECTED
