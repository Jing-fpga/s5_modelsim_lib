`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pIoOdM1Dx+mPjwnsmiJLII2UkOsvwNcTK6h8EUvli1gj8XIueccMi5FRd6NKS/lK
uDA0wxF3EizbTVumGYa32YtV9OtF+gkpeqUd57gxFQIN8BUDPIPKcKMKr27w/6mw
dK7ZXmpaGUJ+wz6G+xWK96dp/To55fTt6eIPw7VetOtHvMGJ/CCnc+n513jquDa6
eOxc6NhsUYLdRb6ceozW4yPERRgpsw2T/GkWSQJz/FqBRVHhwZxNf/33rXSW0bJN
hHSSqEPxGnN2257J+UMnsL5bbb4eBA/9ZI7p6fzN/8j9xfIt0XVXdGw1Ile9PkcS
a0baDpu0HBvfaokg/4/TUgaMSKJ2BwLCCnx0nq0VFcJgcwi8LJNKBSPrs9R8Se0a
Mq4ASID/8VoQh/lpMh7xjAHqjDGM4JioK0/dvoKhULWFKQMUuBRNv57xv/wYV3+i
cdBiZ8HlgRFdoUnyhpYuTVojSaIQgRrFasp74mNmtvHG8CAANefTxkCimIp62ffh
s722dU9gsCBg3/lwMPSHnL4P4FcsD9xhCAhz3t5MMVVBNk1hpaIxBz2UbBkJAorR
EdMNTLj1XcYeG2BAfeFqfWnKyeg4yjGM4Ntk50SV9IxFfsArcCWb1VCKvZPI+qTr
CL+0/xiI30J8aL28N5a7O56sKtFUiRR0HkijBDzMf8nL1ar5E1nYHc5cIbX3Mrx/
An8E1EoFlUwea2v6AdYiyQLXPU9akNNUU1HYuY3IJnSeh5jYoXTbWWkf7XZ1q43S
FVvwQp76ITTQJLaZ1prKfJUvgC/8/rAs9m71zcPlnJKY99Vbmnk8L8/U5LRo8uJd
Ed9EVyPqnbQH+dJUrq1+dLKpydUJ++wmcxxPcL6bqfMdHgrPbl6Pwao0RPspwAxq
kirpCJ5qeepOry7GTqHo7wQ3U9BNiVB6/APkUv0Uu1HTzQhlzWj+07zBfPjSzxt0
Xj3Nvoee1WEVoJzltiydDu07hj5PeFDsQ2wltY8H8jB0Q9WYfuQH1k62g4Yqn2ip
+KZDE/Fm227yj3CA1635VkzZG0o9BL8OEgtJ+XXHHnqu3JdYcb4eLCc0ImPTBkL1
62Il8eSUZXCskPjjYx4yCv5NO8MVMYLlK6NuftgPcytJHqv1rGVGmv9I+bFxTQzh
b1iXY47UpacQldilewuCri9RThdbaxLTWrYwXQ3Gaxh3iVvO9E+4XPXbkSld/iPq
ViAbV9ap2y7VYGdKLE1PVl1RPJn5ydDqqxvsRJaZR5o=
`protect END_PROTECTED
