`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
txvqQfvQai0CYYmvAo0lC8J4kjEwXva/ndwSLC3BaRZds2tE7iBsBtBNw5cW9nso
fvDwIck46sXDFJHv1yJIlmpKMAwCpYnEo9nhV9JdMJz/KrywZsIO3qSjvg7uJpEu
/1iz6uP9EIEIN+YAR/TM9GKsb4LzrQAHFBsxa3WIVKEzaD8qc69kCZc2/H5Ythrj
4cFqNBJv7Ne7eiCmeS9ymeG7tB1Dql3NIrx+lVgHh7SZ7wLCUGt7F/3Mz791UdVi
SwfqcLNPE1zpS1duLnfltzB+DuRMO+0v9IPGa7F/OjiYTaTpM0mzCu+nN3nfWav+
nrZRyHZjCZxN8kU/MQvd7TjOtyWPIK/4NJKLGbI0AXDFwaaKKa7/XM8RURIfg0Jg
tDGs45un+TS3rk3yo17lYX/dCuZhIqdJuQCukVcsq9y/79baP2ZMykD2bVwkK6dm
Ip1DUN5Ak5O6OoNYMbPqQq1Rpwy8itYyrsA6QythO9jLLla1qXTpvRSg3UcMxTem
GEo9qtO6rp10jLpz8E+WRiNNdWsuio6IIDc6Mv/zgTKURsJOcLkf7eNNIssPHyfI
EYzorl2B0blNE77MdBfwaasPWHsVSyKzoPMS8cDVxOyvug5zvjmKPKBsCpSZKVdJ
zMnQV6LXhse/UEyJHOKAMFcmwPEVRGURKNMBc8Sy5LtmEDQX9tpq8JtyPgzXbse+
/UT1oH/GsbGuVJBpHHXI9NV/0NRrZMFltAq3pdT/bsYGwwhGtCx+bN/znRxiGeHI
m4m9Tsie1n78jkZftOnGqZs7JORIgtnxQLkFbyVFznbZQN+1GSecrVrEutPx3X0l
1Tacp5+jA+VTcp1eos+kqhCkgivmwEjwIXZmUfe3vMj3BWOGqG5PwQL1JdD8geFF
jbw9NDbj6VEzMvgP1i7iynDiqmTJiRT12dYjnIuk2tDXsSsHxcnjw6kPGrhn0w34
+Zjn+ov6p2HZ0wiBRciC0miDQKy4+jjXouonZIYD945pDG05vQuvZ2HLL/DFQ8Qx
YF8nOBU8oHelmOuFiP+94HI3uPk6Nt6A81HP57zpOHB7sHv6G+jifM+BNfoBaIOD
`protect END_PROTECTED
