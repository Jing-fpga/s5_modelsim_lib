`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZrTdiNa1KLwEBm2c7UJYdYNUt3A/F2Q/4lQ8EobHuYMfxB8SK5wwIDKZP/Rb84gI
40arXGESXqiqnxTC235RKgRRnWqE9TmeXagcXKAPIwKGqM37R0E9Qx0ttI3WSD5v
scPHcv7Q+nYda+8nMR9kuGqp8urshWQXc0VH3SqEy/gTXfZdZIYKEYykut/rUk8g
TlFSAfBC0AyoxgZojgz2qkRRWxwfSy9iydh4VAc2TshKlJokOUZECmvcBRmPBzez
OwrK6OUNhfpkPs4HfRkeUrngXnG4w2NG8YUxZGF11JBGxLIjXcK+u62xMZJDGQVd
0OLlXh+kiONsjtODseqLnD3yrIIvxxnHU3iDwaqR7JCb4PxyJP/pVrd5Jf72BUcQ
MVudYsZ7F9bau6eiC/CKyxFUmKf5nUAtXFqjgNB38TX3CGz6jFtIxc+FRSVESDvm
iIIaqvQvWnS+UY8cDiic2HP9lOHoDJ2sl3KSJBdpC0JQS1X9888oulvaxfd8QbnQ
mGO5ST91QzxyiIfRWGRpyxUsiyyyFoOHpSXmYpMMb7thdWwyKirgjv55nGXfWpDr
+5wAAgF0xdUPpXDRLWo9DWZLPS8xVjHRagP2t/EFHz/PVRLhSjBuMtBlIU9LgzXq
sRdBGbjZ+cYrnnmndwoVGlSp9anBlE5rXJnrzOxcEBtvvlPUa/Qnzrku84UE/VsX
2Zv5itwPmztVv0DBRuX5it/sdaScAIUVW+daQ/Y1TXU7PpTypBbWEwNYPyXQ7SUV
SVc4cf4CdOvhbwVT0+5zQgdWwV+jOV9jJcZGokPOYGSTzrNungLurbC96GXQ4GdJ
5Vco4Sc088xc18XUHJX9xN1rgmMfEivy6KGzthiUPSKVJmRBjyQTQkIWBKpC7ugq
DGKciY+RA96hxCg3c5Jv4qRy35LGEtygYS4vRPZVtpvg/67nZUBDjt2xGIb+g49k
YKKzViBwD2B82uCskHGwAcPM35Mxmry2vuosM/f3Uavv+eX3+Yx555sFzxQ9mi7r
GFiIBi7JwvgGvPyZZ/XL5n5TwRA5yw5WQp1M62We56y2pe1o6cYIjxoBx/dg3/+z
OiwkIc7767+s6rpQScHIXuGbd782R1NacTD52ULjVNHonvJgqg1SRCiz8/VjfdpL
3fn04ZvqZrom/aRjZum3VJLA7jxWKafPJc0dOMNjGPDajz+Hdb6WQSHDYjZn6MXh
4P1G75cwjLvPW2CgQzWwLex4G5zWnoDhjOw7iCdNNe8=
`protect END_PROTECTED
