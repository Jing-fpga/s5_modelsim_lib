`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3SZ+VPQ4dpoEmXmKp6fz9tuFku0B0cioLgotP74A0IWMqgi4asSoVlOKyJTCu7Xa
n63lCalpMQIK447crNrXQuIM2pOvbvsvUs6724dGdSd04/zetw96l6HPd6BPTEP6
G93Ucj3xsU+b68Os6sGOf6cm7szt8I6e7P9/U4PPPt71YmnE69Zr89EDVs370T/I
VV936hnr2/0eTI5squgqQK5gCIrvXGeX1D4gsqURVLUxrSBQ/nz5gOX9FGQhWu43
VH3S8d4mzNJUx6pghHbIhP5SOP28jDCRh9qiD2TD7PPwGp2mdXxdCk4GxwSOMkl3
sAQZFOeRGVSx2c20of0/lPIQMzB2TH1BxrXJX6dqh9FEN4SIlKBh0aDoU/TBtlDe
ukrJmw9fvmuL6TlZbc0U2gjfxgfaZZNaNil2zG+DchKZ8nhqLq92P/okft34ivB1
KThZojQ2C8CRNTMbUJRvJgpiXzkBeUuFa/yHw5QFFR0r5yGItwUSV+YYE4wRovxw
BT/6JQ5kGjt+sHjCNKXDZeqAu1KsgM4CexU/WMnABWE8F4V4P3bogPE9CvkAhIFi
EGYXIUaDd1VEp4mxopUWKiFD4BH8BTPKuL+nbAkGtyIRNy7QRO75WBBKvd+faMJT
SD+cmlxOTzi5ZtMA95Zl9NPTvKK1JVhNizcxF3B9SGWLjmCjoRguhLgo3Aab4+4I
/4n8Qsxs9NXqfoUwoe2t8hVdLIDoRTcEBwF0miPxkhq4nxLT0oJwxlENoaqg/1Yv
yt+LVLgDHXpPdCNJDJWKvKrH5uV/WJyUMvhIDoWikdjyula6pAqcvGjuopOS/gaA
op3y+WSiUJpsW+2AA45NZ0/xh2G5Sq7RWwDyqZJsi7+S3/CYAeuVML2fJMqel2Li
xUdoN+SItKH20RQAm1DdUnW2J1VJhI2RO2sAj5ynOEjy7yTBiV7vFsc4TGKI8jF+
v32POJTXigyQBpBh9SNToAaO13OVCizn/2HIf37EY54hfW5MjRUBe3gcxlvQ8K5r
72abiDJfWld7m7QSjVyRKOJ4BqpPtfALwJmTYhDjPqPW+VNzdeLXw23hNiXAgb7y
az0Ilr10Mej0LgtNk7LAWJcdlP0BzOw061U7OmPZsI9gUDW4dWpXq91hCUvKAJdi
y8CLBzs9wZh781Z2KzPBrx8dVrYzkw1yBb6mz0sNYQC+XUnN4ms2jQyV6ItWy9/z
vlRtwULsvf4EVpzZUzbG73vZAiEol2ouxFrgLr15gTegF7FwaYRWpPEyGN85xWI2
9u2pGNy9YE0Z0J6vz1QTVKsdQ8kt5Y82LK9bHdklGmuU0HSBXWmS0uBMatLfoUFY
4qfd4MemCDg6DNlw8j7IvhYAECL8YUggUMJMn7X0TRCljiO1n1nLPCjls1Mzwt9b
z1bpX8NnqFFxNBTvy3l6JyrV4U6tTN34wXym6DWW+R77vZ+Hbf7Su7h1rXTgxScK
/9gmRCjTP5oQD/CvhjRt53drrre8fZeidIill8sxOZT9mDB9ilgteb3njggeeSEW
6XoDvzMmD0iejTokRfSQI4GZqm6SQjwK1RsCsa1kwBLXnf+dDxtYsWcPaSMcDoV+
epjqt2SSS5LwUuTZ2+JmCq8Oyy2Ru+PGW94HyuNmeacmUbHK3TONR1tW40GnPCgG
bCJlSnObR+rjm8/vyFICE00Txxdl58UELkVeC+8MbMyQTFPq6YVzexQJ6ivPUjzr
vdemWxfJIi3EmoSWQ/CwN56+JeBe/j3d5hOrkREZuAszg2RPn/7ljWUqr/FYc2dT
TnsMd8YOOEJY9dytNY02jYARk5hxr6sg7ku7ZFJPgcX8Us4WALdKIRmecfCarV4y
DD9bOv+L64yfepUcGGSzE99HOhR9Ns85a9Qm2nS4NS6Nb5NyWdl7/PbnM59n5NSM
UmJi3ruL1esnttgUxv6XMBFK1Yij8uuPliYYwTVhokisZmaA8SoTOfFR3snC2UTl
N+lbbHDnFn4ZRNMHHeiu48oqBVll8AzQLav63zVUSxxURHxO8q4luP+vWfgAHMH8
z2nNmwfkGflqTv9/mIoLHp/1axkBX3FIhRJKjBitlK3NoDUU8ADJ8mssy9o/QRiE
o/LtLS8cMAalT86ZLjO56pvQPurDI3bCMXvSfrOJrtPqTAhF2uvUjJJG53Mne5gM
DKwSKK9bFBWshf353TRX1rrJwGosyErhnQF253IVrP1RoKMJBLdEiWY+Y/KqmXUn
u128Sa2291PLiRsQ/4V3kb6hZRLQKylJtNYffs3dgP4AblCBpvtdZt7LEgWmeJIK
6pCt0yUmmJekCBhtl8kK4wYBE9YLpdtQcY1CkPtmT5oqmcoNz5VIFhKhKaCP/8gN
8iMg9SzUiBXn2wVwuX9i/EJGpQwwcVdkHS6uwjX9clYBuJrz1P8Yjn9mtefot1UH
ItnzSYkBOadapEa+ICQzIj7rJYr9+uStRIZ5iNCpH2dwQf/RK9ppAiMwUBfS2uGf
++2+4y0IRpfCpbgkbWH8a9pIX6HY3YJF7aauxPA0HIxAw7nGgmrxv+UWuCi67sLB
SMQh3YQzRfwQ7DXnLmXhK9kMuVPXfFnwnYDaIFKny+nSzcdIxt+xjl7qaRqkUcYn
to6PePlu6cRWZpxRhBCi1k0OUOqVpHaYdjgIW8P7P7dcE1joRkwRpWxj5qc6vYTY
RP02a3ya5D5QG55+PHIPyjLmHrk+l6vAQyZf9CTHd78T0+eGmRsC/3btYRNE066w
t02aGtQ2dd5M5l0KFQbRmOVjNZPo/f0SSgjkNvEEw4JceljL8T4fMToNxgmPxdlc
Jc96XVsZHRwpQumYPGF+mbrtpY1q/fCWvBABpECEMZoOeN1ByuILWYjbka8WIseX
fRdFdyjY5IvxuHuVhzG6nwiqpLBUtkRJXaYmIo8y247LFIkPiMQqxxmLqqBXfi2J
f+J9HfqqZjFmCFHGTCAemIV6u1bvEN43cY2BoW+axqrZz2iIJ253VM/BWf0+CO00
TXaFVpA1jutHBpY7JanbqGjkadNPtonVqfpXuZZ+lA5n2t3HAV9qzAmyRBhJ4CPI
H0syT6/ExQWAFNvu+9GXlwtjf+g3diyZu13vy6pqlSPRlmCoMmj+NqtTc47nNlnh
EdwADOMLl2w85K3cXC9HlfMWOFNr+QkoTFku1Gd31iQmvSTerjpCQmiUSKf18Pth
BnPBoXgmywRnvyvdrh61jhUq23PvX1ZAajLoMFcQz1y0dPiFmYwEJxfElm6Bbr5r
Wx4DALyeMj3YqDa0imQcQuv1ZhcU51e6HkgEbB+w6nMBDdtfI5XRLCq+u7nmuDLL
k+Lnn1qdnMhPWTPiGHj8PO7U47U4QXLG5aX5WyAZmF8b4AV9BcCRa0jbFw0oHpkx
+SpTcPydr5AAHO93QXVvzwyUSZjx5HrrWyc9q/ueuUkYoiucihVsaHGfYw6V1S4x
JcSvURAdUgWOo7bHHmQNaqK5/K45eoKb8vPvmosXG+AwDaCA7FFTz9ydd7JfE6F0
iR5GJFD7EO8ZR1vY71u+XohXvVMYVltgydA3zRYY9o0=
`protect END_PROTECTED
