`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RF4wzIqPMzbf3sF4Tq/rDnOth3shIeD8aCbDrz7tnaLvIkDFpwdmtphQXw4ZizRx
UfkWTwYLfmlSbCvxwdd0meWKLRWmJy33CVGnBaqrVwot70hzU+YVluFJqKUvRTCM
AzsHH5SeIBpyTHZto8D59guRzR3seT6tCG1H+XOZtFbuGSBHO89waPQTTZ8Cxvle
a/XVhvcpKCroVx+yPsrpciLcmsbszA97a79Fq0LaHXxuqsodE87/lgLJAouis2jV
hj33dwmwb8y3gObMI7bi2IabGsDVDsdrqO8MN0dSRLuP9aTGSm0xNdPQhyRSX510
jE+FI7+VhC6qvW9+/4cYLOr94sS7lD5y7yYQt15wkedEOgTFkHU6+fboslkg57d/
/kiN0iXgUhQmtJojMzyq6RngLi2b82qcn7Tg1Hiyc6EI0C993+jtLSs2Tfcx8tBU
gYlEQYz49SbeJrrLOsCNJWvA47E3/g+6jp39QfzqqQzGMniDFIoJEIdALi6U08RO
PbED/BPYxFIN+NBTyVf8ZXoFp68Yg21QGlTD5Wg+aJ/WgCexwCOuQILevy7lvPw9
k2TdPJ0AlE131uRgOHrJWsRP3RO4h+jyVDarVm84Kt0IX+uK+QsDq96QnFVjibuM
VX14CaDFMc8KsgligxUHYN9hvFN6tC1O2QKoPpqoWccwmsH3kopWi5VHjQllHYdb
g7VaqJ5yWnL4bmsrav6J45ph8/rSOc4Kr1b8uoB5WD52GSsY3m/MGmLWCZ5mqoDr
0htXu7/k9M1K2/kWytFHy4bV5WHe836TnfdicW/9UVdyLvTfpTLEGtthFc8ihaGS
`protect END_PROTECTED
