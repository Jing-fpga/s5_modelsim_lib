`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/faZXdETr/cPuLC+dn43BUUhzgRkngHzZwPp/dwbbT3oqkw3f5n+wXG4LMrGQV6b
vP0EgCQJ+sDZa3sQQgmUjL8QiV/5CUx6n9c+YfLZjJkDISYrXdMeF4yxbGX+NTmf
CHevIDCvPTS4j79I8rHPJP3gqFQaVqaIH0oEFSQ3lvD8zhOtE+qLOEx+6H7IKS3t
KFyOe0hqmDlMBa/PUMRF7vSwbwB15MKsqux/rWWVShibyl1L3tOJTz3q8qNKdCw3
jkvthFx1jeHo/sCmgR66MGr0D+/oug7lnHCaVhrJBmSS5IoM4c9MXHb2tx9Ecty9
1KGhumaK1M1+7/346jGdSj1WPf8XOqsREszr1IDByDc5oeesjCw4hNJVj1GdHxNH
nR+Jid0/m8gxhYa/amneFy++d/N8u5qSXPOHwHDVNWR9op6Db1TVG81KcNyI+b5X
OuOAfpbUvP7bx97fr4oLJxnAvAFkGxOFvRCzSzeBunZjL31r6DoE8wCABDbvrqYX
DGeOaQYu+Xl3UfbkQIhKq2/Z5hgQNtvpRP58sbGkMqX22htXpU4YVEfYCi0KhY10
fSJYIbB0yaUnkPkSl5SDx2lWgOZOzTgjNBml1MIO5qF30OSrttkkSx0e78D48+Dw
FBi9m7RjVMExcrg0hYkEruZDSvjmMYGPKBvAevwUYalDOHaVK6KjB6gMqiQeU/YT
t06dQrSQvYY49FRMQ18zDpFsgyPD/9sJdClsXtn+aMvLAXm6mwWA8UIHU5gLV10g
OQ328bC5SPd9wucI8MuR+f9FTkAFg42quTzUhocO1db+ot4pjrteci546wTBykda
pqdG6vd0VTgu8BQvcKFrHiXfDipiOBOK9S4uNXbyyIdgvcTK93pl63QYYOy7VbL1
HCXMF9JVdShClaT2/pAL/YBc02mpLaqrE2LALpXTyPuDVlAv7vfU8mI3aXK1E49z
cepr4wPUrMSNwzRKStC5gI807at9O91gnJmJAx97iXxK0+Rh5aUBWqJtgrC2N0G3
13gOf5O/Vkj5MU75Y3mm1MqQUs7gWXdwGGOhnVSe2rqnFjxq/mUaj9ftUXucANFz
zSsctN5PoAOuEFtlviaGaGb+spjpwcwGEqvub4apz9UeAn1TPqTYecYxLnPrHfHN
w/60YUZNuvfoUl5Aiba/BEZKfdueGNPxAjQb3Fk7MfLi2SrEml/h4CS0b/EN9STT
HI0b4S8p4en9zSC1td6SsAXGflj1yF4hmf98778ays8wjmZ8fFiUOwX25tWi/Z1C
NUv9GST0We8kNV/m3bHZyom8TbiqcANwW7did9jOwCwfAYdbt8DKFPHrNcnjz8bS
08a/WIFBjNlbKyZCIngHqxNtCMsBiY8EO+rGPmAhZ3GiXGL5iCwxkFDVwfIG90oK
j+t4nAcPCsKLrKbYZWJy0+v8HDPZ0t1eLvs5c4ihFGGdaLwoRF4v9Zn5GyVk5AIX
AxB2FXxb0MdMZdi/N3PAu+OOW+aQqbj5nrAi4wl6AezZ2ZuSOHtB/3I9W4s839Zx
3zaLpLVIjzFSzNNpYRGXVKw758l+j+1Z3++Gw4wlVfU4TKlOzMy1hpgfasJyErTy
Zr0OfPtAIrY62URLCOwKmDd8QiHp+Og9Rh9YVcqXmuORF0dLj8Ft46Qljn1ZcTvS
FaIiwrFXSBQMqCvKf8q6UepkI5ZoLBTC5r/z0waWQyYPmrK0qusQSYbZlw1VCOSo
3nn7X7o35jQaYZD2FYv1XjN7pNgAInhSWtXzAS+pAssRxLqU8ITZ2QRuUfNowAnK
1YblUSK6Yh7Vv4fL45X8IdoHlQosQPo9faILmQvdK5kNzMq8UgVgV0C7JuCdtKAw
ijqHgZfUYFfXlO53JD/amozsx5v5TmqdZ5n5q8qljJP41xBHYe/RrC7BcZwFpevj
WrvdWYv5xZ0Tb+ROg7TGNz5hroFWdpSNvU4dJywoLMob//sJhlwIdfDU+PzoL4qx
fUS2vIOxKVkBBDUw5N329SgszNweq5Kv4J0MF22CggcemOjzG/x+kF3/B/Pqz4H8
+IdNLT9dZB9isLFu0s/QPp1WWnle00/+2CpZX7UtjEmQWB0hr/TdqfLjozz3paAZ
54Ug//nfgtUPd/+ZsGRuU33MRr9G8xhT2zakeLZDv0nlMAsSX/h/2hm2WSg5w0b0
`protect END_PROTECTED
