`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FyuArj/+UhmHd0hsHExAFOmzxF4iWw6izRDEX98VwDik66ZPpaata6OsGZsX0vcf
fGKG/yKQhyoBv8gzG4JAIgszaKK75y/sQfX1JR87JZ5SfjmG7O08usocI8lbIwen
Ykud+yLpmb0U1rS7yy1zk5+StS1KIBrLY5Z4sMQj+9xx/mOuBu5rIVkGQ5U3bAfo
Dv7siGvFW/1mGj0nU5NdaZYhtlzf1aZ90+k+fGrMx2p5lXSZeX9xKREpHUtDe70w
+lZifQQ/eeQs5Tmi0nm8US1UQXYWYVyWFG5k27Fx7ZKj1YaSKq378tYw7NAHjWA7
aLBThCsDgAx28nje0S5GG3ZHic3epellGp9EsHTz5cJe8+UmVxr7bRdlkXwE8OxB
NdkNNwoVv6JQhdcYy07YUPfYaGKVPMhF37u3vmdSyDuRq3wG49plR0m9dnOTG+MP
zvfwTowxbpxcb4acNvD5sDcNXbdC7/ScqjJUWJjZb8F55vNTtsZ8Kr5I88HG8q/4
ZfHgofQTzv0TB8fZ6FFTyXzE+Om2rc9fgmsmWRpS8qvEc+YSqZgujwVtf709lnQ5
ZPaQv2pJ4Tenq2sPUKeD2Q==
`protect END_PROTECTED
