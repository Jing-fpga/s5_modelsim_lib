`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JTvGQkNr3M56xVx84nubCjM0L5YPwhuMG0AWwoGfkVnO8Pevvlp5Z9Tqx3/co/bu
BIyykE0cjH6VjWLJ+QN2OLFl5RUwAqzFJx3nQixhZMJfvLVPkWjJHNKU5GQbZ+T/
NObM42dLT2fLHIgJGSSsXgu6FTfKpbcT5kfhdqzpgdgJt/16jxtxFZYK05h5fpd3
ndF5L1+dbrIRkr2Cpo0Jdl3X15EJVSL+kvI+at6cHkbVArwZjwO30vTF6i9Cg6IG
XJwV4vx5LXH2avBHxbJF5/Dh/rKveqZGdAFfHSJ/vHD0fD8Ms9ky6jtedFS77B8l
TzUsf+rmUowGefDmvfNjJmDCJNF+hABHPKrD2P1CwT35YNQmagA9hZEuKBYSIjap
zZWxLoevyTvk0W7+vHTb7oqxrWblVdpjKoAGUq/AY6nxGm/nSGgxX6cZ3YIyepF8
HodRhg0FJF22dhIFj7iW/hfZjzIt+KSD+utr2YxnuM0cdxfJmL3FWujz9s94L5vl
sWtTY0wURdjQPdMFCIOhls5q1Xvua7lIzIv1kJQQ9lBsYTCiBFhcxBhkakpiFcZc
FZtITbH4dTkwpNoh9tkC1hV42BVQtBkckLX6Ul1odSxJ1k1hHkYygABTwG6IjUiT
t7zAS++ZHQCQ8kWKYXSBs5289mf3Pp2AiSK/plBRXv7GiJaExgKfq5MJiEct2rDu
ip/0GQ4A85mfIFcT9IhZ7FEdLRYJ03vkmytKVyJABp29zzw3qPudAVu++kt5Zff2
4ncWoAP+W4GphqF7Rk7lOk7RoH0uxSlXxnnWBzanRmX/JavFh4Imi7KUAjPjA699
`protect END_PROTECTED
