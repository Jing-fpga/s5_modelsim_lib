`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ckyD+m1V61g8ftAXcGlA9cThGTCOSDnk1MPS9wJ6VW8XHjamIws2FKphYn2LhcmJ
uwiiZEysL63NO0Ik9rEljjlFoDapc+KtR38N77AFLc463wtU/6bjSrCK2MNjKXUt
q3JBGiMoVKg6jDt99/wrmkFXTOcYTFMRsJiVg0+oofzP/Ncjm6eA68Sp1xzkEoVH
fj4xsHRwX4Dv15htjERyMqWVSX+NJ7WGaAEHxBcZvjRgOYOFFtB/Olo0JTzU7slw
2Fqs3fJH/Mjx6b3TsuOt6v1ISNIne50zVdFTGZ+21Y5efCRjdBQSiCtA1L5wAf0b
08RfRygZxL0thrzg0z9/VQisdxAFw+x1kv0X2cVfQR4XQsdNxN6lkRwfz5SK23yW
vKs0PqZ4JrvABwFAuFHx2HcKwsSRVpGaokmWHLZec86n8/+r/Pn+vKN+VDtCyPq4
QAYW0+NGjl4w8/3u3gA4y/DQAvMIaqgKRQzXyigd8NOVbKFJkRj8EiPJgvVxcFYj
39fF79h6WyP6cWzC1nPhEI7bDOMIFVVOWQnW0tD6+9UQp0G2gN7fdooEOPEgaC0w
1GtrZy89fFI0BS1oMtj7uXkPECCzJ6NiyV00rK4O8jYnqGMNa8j6KcinBD9iUR/b
XbQE1/u6YJIvku5L06DNe5IXQ72+Tx8oZwnmSHChVwS4g0ONk8mplc95LCJk/09F
G6/3AvCdg9yJQfZxiRvSZilAzBxT43tjJ8V3cjqVKqtr+yn7+825eDu97vXutANS
BCA6y3X7QVOoWylX61Ef7crshIQdTPKfhFZuHqi5rU9mcQX2C7I+63rdQFcMPLkg
n2XVFJxDzjtQuVVOxNpIq1zpH/X6/9yALtV/rH3ZQrobHvHaImJqMvYtoW5IGbbQ
TNQGraPfwTK5fP+2bR1C6lBmMgnoCEqL/OMfwtmSL6pnh9GOJLpdTk4VVxcSdrc8
AnwvnhL7j/SytKZkoVceRJRp8YF9n6QxYf6QUrBb2ajO1+d5VO1diRQC49JGQlXz
a1Y8QfUrMht0h/OmbiUpBmqnF6G5iY+V/UQbWChHAqUjM6IVjEKCwvtPVCJG5cCO
oFHlvtp/OISDmI/448IGzyDk45NRvNibTT8yLepr5nGQI8SrzwnpFVfn9I1XGAeg
CDv2PThhzzFqEFUK/XHd8DQYS8jfKdyPrTcVX6lnk5q1C60Z0aabET6dwXbTuRyD
l6pn9Fj67pTRQXohPTjGgLP5YERuyPBf1H9Xp4WPeeAHK85uI4Yg35kNbCjVeyaz
ptOahkQZnMA+Gx3j/zpt9jLlZ6HjtOPo+odIs/4FDH3giTo5vNx41ya2jIdkuBAf
mUrzB6NyT+Oyjzrs3CHIf3DnpjJ43RG9Bs8l9+rU2KOPHwbfi3r/dE7QrQ/TJI8L
3MfoOjJvXpWBYM7zLkHwKzx3Nahcd1suyj2Pfa2YryT6miM/JsXjal677JpAiUAo
coa1bHuh/j+z8wFAhDKMPnkJbMUOtUu50DcSQ0hEu4wBtNsULKGHl6XcIOprWInQ
mjUeI7kM1WrQxmvlp9XDaIL08VQ9CgXsj3uIFdnYejabnDsI8KgL1LPkE4TOKbvt
fScWCHR9x4dIPvgONCTn+7r3GvDZ4E9bnb6wyO3IBMMQorI+WmL5IHKpk4cp+xau
w3A+83QLDeu3PUyKtQfqMOc5LOpVei2bG1QZ2gFiimxVqwGfy7IRrqfxbicfbebQ
DwbEq0WGoUV9ptV+iRgEbZ3FkYh+3qlQQWX6iZqvx59DP5/3nwe0j609u/wosdyB
CuFlNk1RO7cSBlxCkWz1EW6atvEjOGVL/6Vu9dRcfCC9TOIwmTrEqG8jB+Np1O5u
yTQCGnOUtQM+LawwpymVpQVFjJDxPeQMFCYc4oSjDAqzbqvVO1d+YxB8yaHtapkd
JP+ebv+ADuJh1ItNNJcVfmjWqv9vuSeknJQIvXAXyCtJ4NcauY9Nni56cpYagYJb
oYgt6BismAKhlSXIKPBlryVPGyj1nGzHOptDqf5EF6ZUxqPbfbcGlMk0PDoK2ZGP
p/JD/Cs112kSqlogPeRGWtnQjIIkWXL9fjt04frjAxB/T14hNkLlyyYxGrJ2nzoj
A0nqw7KvVzMmg5KH1DV1cNiafELCjCPDNcXvkfY0tjPgUlroxQKO2trFOEPdrDr6
C7IpMGL6YEm9zN6prK4PyXYbgkBDi8+m074wXYnoGy1KvJpjgdZlv+7G/9/kHTCg
yurqfiUm5vS60Txm1MYB8jfphbJEVXgC+Wxwuxi4KuZQuxavH2rQOpPVbnyjkl5M
jOzBZpyJ3ldIhWFf3iO0CAVcz6vPl/qfVGVs0XNwFzhWfbTladZsP4dwpaK2j972
VgxO+Ke3r+FFrsl1tTUszkozIrwdD/lSXWsW3g9Aey9ax9x3Wj52jcaf+pkgRhX0
H0ftPYRNaZZFAcIXARJzCo2MppvGbvS6RZS8tXdEZh6tpYs/0VLVIGyP+DpEqmEM
BBK0RkTCiMrGHc/s23rjk++yusXeSrKrdLDKL/2z34K3I4qkTJRfQEtBOVF+bvls
GMTCCI0znUxLEoD0xHcoPFQo7H8gby5EGalfaU93mRY2sAt11Kh4W80poR+gGAya
jkj82oVrzDroLlJKjpuNJaKvgH0/5Qbd9DlME9QIR3h+Cw9AiVha9gxGMUDK/EWn
lptgNZkROrRWSOjxJPxtDvyHno7yvN6GKH/rQX8Bnt3adTLoW4h0kxdxae9EJkj+
RlFCyZFgE4MSCDux6+j/tstd7Ee+Hsv4RAg2+kgSOfmjdETMaRMTGTBcqq1nneCO
KykDIHavvZwJ+g8veSzJu0PBsjLnP8qzJLAropZ4beB2HEzQVTRklPlbS1QkGEnQ
5jF7BhUqJ/c7qAAZWaow32BWrtcJFXOsmgM03TSiVpTb00nCeFFAnKu202dBmFHi
hD9Ni4GVW5skqgqJ7PCDtDjJN2jDp4NNUurE12Zbw1KkSl7sFJ8cpxnEM0tlSqLf
k7OR4dTnl2xv/i6CnmObU+5geD1SzCBDAybPmMhKrmbiwd9Gc2e6yQkFIHLhcMlL
YzMIkmIui2KuUIsG3ggS5uqFyvlJnvDmat5ENqQWf4kEDnwITPuQ1DrjTbqgFG+P
UjIOCYZWmLo+TDInPCtBH2zH7RIXpNpxyIvbMLWl4mcn+n9rQCyaOHoUjNf7YL46
0r2M9NgJJOwdazGVepb15XLDlMQdSYw3V3114TvW1CgiCUXGdJ2iR3ImybLRezDi
1PSC9kLrZXYphJiUEmXJs2pnfDrA/x92Bp7TVgSt/2y8D3Vlx/rLxFhYtQ1R5VlA
aRymKvdl099cmUF8MvmXWUam2O8v/zpDH1fQf0iALtOqbzhF/7PbGT6vCdhaUEb3
NOo+o5OUJX8qqdRWmEorieYnpc/J++9vFx/TgMFxDXOGje9WF4tLCoMDE95wahPA
yJFTCKvx6HAtad2wprV7RQJiIEnwKvdElHOH1uNx/DeJvOVEBvoue4lKIcQbupi8
h2HIgHRyBHaUzmjRMIoKfPNe+RqzVzf3seXVBtyLzI7H0sF1JE+l/8XElWti/vb9
Qo0vAArdeXeBbAm8BoFNWY6PZJZ+nQqReLdad61QEpo0dBVcag+3SfKT+Mz2u8zo
b4p1hwLdWDwNjoGyIL6wWMI4HIMt6x7jSY8b7tFXvowCthZTKtqGbzQVW/t8Fwxz
a5xQ+fY1/X6pPyfirbDOlQyBAOWPE8dt1GTdUi2+kroNhDN1BvtATwJFcU2yvo3a
LwA8UdEwh4JhwiBOIaKxnSWZUChTwJdcIAoUaYD8ySyxAToauC88NtGObc0CYaaY
f81Q1HiD/9KvBlmBLAZYnE/siibFx4/yT/wJnCfUm2N3GyyhApQdnCU+R8PPdDqC
kYsCJ55AoIAkKzo76hpmzE1Pkoc7ZVaVl2UeZSeXxX4hqlvZpaZCZgcBTibNR29b
jDIoqGbnkO+BzcHvEXU98m7sKz8a6YhMOpJiIJ+cGxo1GybwuyiRLPaX4BWaJTwv
WrjJPTxWn//nNWUOB5iB88e2QtfoEEZ1zUll+frd79mVSw8OktNZWRgZBO9sC3CL
sGe8wNAA0eRLb+GPYkbpzpb1Umn5C4lmq4W2rwk9TL08iPrbcP52A8Q+BZSjY6E2
c21L4f3ttmRzku+suFHtFfQsAwD5QWwM2gGqizvl/GQ6tUVacKeA4EVULiV1uLMT
9PJV1EkVil8eYA2WH0YCog==
`protect END_PROTECTED
