`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AffTDTDwhYJF1Y8UEocA5l/zJ2MR8QfiGYw2E/e+FiAu++askFTx8gSzHeOjZCC5
itb1Ov/ZSDFg4gIa2J76DLARGxFj67bQ1wniG079wcEFcGxfnicL2RAfDbUbH9/g
eY7c0mp+AZSTFVnG32hf08ln2r8kM5BjWKarNLqo22IlAeyEWXelVTprMJSLODth
SG4iwiD2UI4TeCO0bzAZo8NBPgjycM0033yjnWRxtj8rDLIeW1abSLnzyWweWcJQ
DrFrxjl/afbj2zn5rPn+cmOArkL6z1t2tn5xv4NP3pb8mnPB8TwMqQt/Mz5RNhT6
w8cnkxep8Cgm9c36fggLeXqWOz+AYsdyGPtCMv3uJPXBd0In85jq6RrTgDzuAG2d
t+zDDmbzAoZakUuVDMXk8kon5coH+8bu4u8LqagoL66/9+dGkvsOV6ET23YikWGC
NJ09DzVD+lxHtutjPGEt5Vtj1dSdxnN4bUpxWsvMvuXSlgQRf6mQswELcdnRQKJU
1gzoPmPwUQDGjXendH7995iXGqU+IwUqBZbf08Ud95PNK6JpT8Z2J3iWjN5E+ogq
AJmA8dO5OE54VovJyk71vpMDPhj1ci+GJmccaVWegceJp7kihKdXMNaaphyW9Bv+
aLr6ZUHlsn5ImD01Z6AnZVJXaO8Cw4+cyjlkdUkm7aduHXWDk+J8izwf+7emyBg4
pEff7pYwpIsdNVtScIs4+nEO7zgQq7szTn/doML3pDaxI67k38RuzmBVcYsbGFVt
0aVnCdY2Nvbvysaha6s57kEgRSnU2+oYXluq3HofOBRgu5L9L65aBJGvroerB+/2
dXNSEPL7H65EtAwR6PVzu9sTzhV9eyaXxnGjOZU8DOZfR93yhFBZ8JzDQ8k9t0VD
ahM37wQBp/dgJcVFgwZ3/ubqylSuJUV+6PfCIYvR+QbKOlUlMsdQNn3O2jUeP/mt
AXPyyQocVUlpCKu2mWObI7tympd+ASh7joU7aEl/0VdEp7pi6O7+5i3ZcRzPUBI0
7llRQCimpigQ8Db5TpCmHg==
`protect END_PROTECTED
