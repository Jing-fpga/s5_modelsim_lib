`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0aWJQ/9BiWUHkxqfCo77nLzxA3rorn+0/fRTYwEyD69/a/BFrGRdyzexwS2irOLV
Ic9RHeLjal/jmg2o+0bszuUNNiDbYc98uro10pbhAHm5lJHlxSfhDVVmMCDlrFBr
63owajModG1zNcLscONuiptlf9kBlUnM6Z/THk0DK3qrIeyjj0MHAo05ds+QU10P
UWAyUswOFAGWwqspzu8EdHUnuwecioHbgD90sZncpREImJjErRkPt+ORUhE31dUT
N0o4Fj/EfpNhjdQ6VjyJnFv3hW8os8h6QkSZ6x53ZAYrB6iQgMOpCjBlT3NYW/vB
qsCX5Y22K661QGQGl9h4YVUK35bnVy1FnD8O+ken1dfA7JQxrJXJ04rUy6q01RzL
MrKw0vYnEAuDBThJ5Kk5tC0btLvyhraFfyK7pSyVem4SChO5NjIoGnDDhnjKxbzr
No7C1JfaGu4M0uyFkkDn52dN8sWTgbNS3uA+zs9tnCD1MNJcMc0sKHWL52Uz5Idv
bpx+nbkWlUXi0lm6bJi6ND/FbzHW5PuYvvho1hxJ/ajNddh20UldX5jxCVBE7WKb
7L35ddeAkCUoosaVFNVF7qMp42VLkel35425U+ntUsZzkoVk1aIsAFaKM8zaeCiL
QkiTr4GTYNUZPYVHqm/yK8lMJMqdSYQWy4IyPXodRG8=
`protect END_PROTECTED
