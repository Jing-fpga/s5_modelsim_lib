`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Ni2fmIbVWucn2TN7QtXiXtAe2qu2ODmZAS/wYeG/WY9gRAccE1DqeXmxIJkqBVV
5CRrDpkOvWHUXt5DTuH/yh09RatOeyV8VgZRz+lsVXbxhN8GZrW0Zm0a0G5guzZh
ZHNSr2mTKl3wTLwnmdBUTlMUwX9TqVBW76kP1dXrTdow1OHYvKrI7zyGnYZQtCbg
xbWOzoRIKRlRzjzNkcXHQRGZmeyXRHMDuj5EQVQQTjov/AL+8j9joEZJfIq5ReOj
3xDs4qNdFbYlpspZVqvBcEQ2HwniWDtLXQmsfimWQglWsx7M+xcZJj78Bz62NyLo
OCn47/Jrnq/2xFfp4JGmS0nFbrHfFWr+rluTQff3A6EdgrkUs59tcKHwpx1S8kmR
TqoMUcwcuQni18EA4gxpF1+sLhWni8AWlMWOMqCJTBkkBBjh+9CM2dJxXV/HGIAA
q4bCSfFQP/R0GfcpGPjqkJi8c2qXams71dlXqHlt8gjhtXi/U+UktL/o0kxgmQcX
jR5O28UYEnNM24RKxJL+OZyl4y9wBZktYtDVk8Zh2o+35kL9Xtz+/rs/f5QZZCWX
MBR4vQmq8qm1gwXY1g4l9caVimusokEc6A4EE4HuF2PPWI2BVIYM4SbCknBWR5VT
LyxU3qOZZmewmRyP6wgFDq1azQdKHz9anJkJbBjY4y7g/U723pPoGHSERMhQeCkJ
eglwB1EYjZ9yY0iM1mnFKt9y/yZMCRwz6kuKyZW6EGKnXJCoIFseKQbK03nvdyq6
Wtq7D1BLniOUqX3O8zwLou3z9DzmFBEwRwj+/TDX1mdV86iFYyoQP13omX0GyC70
x+A9KJG3Kj6jJ8hoKaGUl+edbvutB1lqlPIvOdQiSbfW5zXy0IYDJdXKshkiitbH
bbAMG4X9tdU6/3zNcMnzZPfZOYSh3Jku6o4EyZVmznQytLb7Gib9rvNP+ZXdZXrb
2plrZSu6Nt1X9W4OwjBuWcR+cjhkZI+i1LAgVZXEhTYdgJHbGtbm4H0NamNNZF8o
knt4jR1UGPOWFeFwHgM9418heYjiNJqG1Lf/cD3vw/5dFMlW3COfEXY5KTcnzZfJ
fY9REl4aak8ta+MkXDNp6Tt8UYXWI2LTL8iteojHr1rxQfROLW9iyIbJfLwgy1LX
35P3tesKPqLrLParbiZ677tCkLu0GQCdYS2QMmq12ThetXQdIzRZMAXCEHcjhkIX
u3g8O29vmIWHxmoFzXHzJRlkdOzbsfmRB1wPSIqTmJYxV1L2pZwSwiCryVZryN7d
GwT2T/kJceWUUQUAiEMv1CHUSL+1xMTCyT6kvRD1GI5CrZDKkgn3i6Hwgkgowjn0
USXtE/hG7BpX5l4fS34n7uXKWrk/gkzhY30Q2iuf1oVxtK7xslNSfGQV4+AQ0w16
rJ74KzhJzIq/H5BPqfaIszrmvprQaOR0xbmFYPavHHwbJFK8iAB9jty84xDquJo7
KuDbx3II+o7mydcJKkihaeW8ID+2zm6alcFAa+X6s5nsFnJbDDB3Qlbd0LmolMiw
RYa+e32dmZSmzrvs4S5L5KiyKmbh1tmX2H2PC/5KIPZWHv7cYelkPtrGPmxKwn4w
76KNRexeStH0GLLacguX9qrb9p8+orNQ6HMgQ8VdOa+peYbtKj9QzoDPlOarFR6b
d+s6UnxorRbTGWMmUMPCKNtECU7GLmVMlZz6vabef2Vi5sU9dZQLbc0s+QIVQnDb
xFFQoIOb0jjnOA9FdFIuGxiS5+PtSW+n92ePxWZ8kzEDW+L5eiTedfGVv4dI9Cs6
P20nveDZ3ULe9p/sAEwveXZWT4RDDDfWHulPAgIwKvqBzacFrqcCU4L1nj/HqoBT
quQRvcMTp2fZmDJ8xGfisNdWzYvbzQBccZ6QRSxb2pq6SsWOYx+/6qA9ZdA59+Fz
J+BgEomOMx+JVN+hEZoVOmeVNcFHeT4BomC5yWBmfOyumjmvmLT/ujBg3B6AGz/j
V3Cj3MXmdgzO/HoldGyu2x0I5HN2GlRePzIxUbgHCY62hRDYva3MnZqEkpsr94xV
O58c3Q6+ybQUX4GIK2HzijjLF9bdN1arTEj90/L+X0MCWtUIPkU/n8ITdzX/UXkA
LqPMIOGdfkd29mUXiub0HflrfFrEGRGqGdbH27hQuuJv0VBSe0vcMdPl7N55vkjP
52vc8XUYen19eyJ/pw01oSvs43HMbcO661L/eWuUbwg2pxQKBUiujxUXA0f1KwT6
HuN3lLiaywlhrQK3SO/gfhSz5VHP1DZRgHIHzfZpNWKaIeHgaPLv+N3wC088T04F
YgJkORaNgqrVj2B6ISdC0XK94SKABzn3UagJM1iNHrAYQ6xyZ470eaUgHHPAiBKB
MNwWEP5jAnyNzB5jX3Xgov8iX1LCuYdZ9Ao1NwuUQU/gY32UbaZcFX9qQDbqzqHA
ejWHqTJ7cAzsCcvos/R+Seda8o6PNiF444JyeLuZSjMH/D+aerkKIGpXoM8ImraV
0HdugTPn1niyD3kz+yxl9HJxwQ16TIxMR+O22oP60i9xmBzBErt7N0nYFlwo1Cap
+Fn9XW2S3W5TC38OGQZ/o353upVC6F83bA2aIjuqFL/yNSsWzneclco6nKWIfyJQ
vUcvCfrCX0oUNQhlQC3rRpYPfgLMzQOYmBevKS5NgC+fxQKalTa6HvlJnYtkvfZ5
mhHxc8u0D6e6yxSdKpmA9byWXQ3sg75A0YdB1PVfZx3qqnfE7uBF0bEtDk1MXKDz
EEYrX9dYOYiYazjojBCZQ05GM61R/o0s4dL4ADLhTlwh6OCRWGnZClfUAu9slmqt
wfTXjSxrQhF/FMakK7ZVN9n/QzsHaK+juauzosND2ZLyVY5/UZ0fxkoD+C2G+IFU
8tCuQ4CRdgKTuv/xAvA44uH+81S84J9IRp2/rwSkUGl5WW1fbmKWRiCWmZcUnrAO
EIi2anx45tMgXU6t1awkw/tU2MdSzteUB8EltzLkHbzLfOxSN9XJX4AdRTMA4P41
FKOxGmnL4E7Bw9X0qJEDN7Gv9KzVo+/AbucSA95vTawp5kTPnQmdr7DNnDwA1Bg2
+VP9tAqt/ZPykuwqK+btiq0d4+I5BRJC48Ni5i0CUL9I7Wj9Yo/q4hSOx/LWuF7g
e9zBrHqxGfozNnHYhNDd5foK4mrVyUZU1DDOGQmNrqCQ98mCwHLXrjFpqeNMwpxU
InSep7e6w1WYARNrVvsewhslPgfUaf+ZzTVhuVTLhpzJAW8PT8fUum7PZdzicQ6H
qNRtF7mzSDMfcAD/geSo01Fa2sZn37rkhJCuzKFCWHuO346AsNta4Lyf70+HG7hQ
5QI/OUIaKHN9J1FfwUvAE3XGTKSl2LwCk3Mjx4aMZUfce1YfDvUIfk9JQSCHO2wB
Qz4mieLpcX50fqNV0owQ0ZXXtUv9cg/XnFIZ6hoQoB4jOlvAk4ice1JCKeiV91oh
zlpZHfpgiL08yJbZDNTxgLKko5rwCjnBRrBaY6KjL5vNWW9R0G7APQUx5OCswuZJ
qfUqeDfnEQPpo96lbiRbBRxWz+eiynjs/cGzr20lGb+AJDYEpY4MUpSx8aZlXadr
J3NcqOpy5QBj4/gFKlQmcdX6wBkrRJYyBaSrz8tvuxYOz6ZUe6x3Mo2A4b55pFrp
p30Y2zJ+oiRBF6XvoiHybSccp6EF4e2qUcXaraXsgttESuInbOmid2y8V6zuVjTv
aC/3zdHarI3cgq34iXR5vQQKY/WMnM0LEkG/6fZliCG/kgySn4bcN99Pw58IO/n5
MnugHYb8ILj2C4zYeit+1PeH2XBuAGnraHnsA9pVtNoYJYjLJyUDR6x61+KZmKUm
s1ieQX1rEhZrRdYvIofbg8KkL3b5hwopg13HJBbdBEZIC+KaOhTV9n7vgnqgHyqx
L6Ro0ASLSXLDETEQef1UB2ZsTR97ZH9bK4i/F3HdE8lFFAwo9cl5UqCPJmh2XGoP
nHpxyFN9PheGJZp3X8xYi7Y2rsWwbdbwuEX3ynhFU/zoWHM2Y4Yf7iu5q0sH3X52
fZSVFsM5Rm9fjPu8IctBghhkD+a4j5NHCJKJfQIzibTJcYaUdwqnzqoUw7kJrMGQ
edU7SOxDRTqPbNcagOa0jy3CkeeUqKqhTHgEo5Knm9vsgxjnFWcfRbzElwXSDjTo
0tFBLJXq52m6k95174z2e5dgNro4LaXbLt38WQUG0HgPSZSFjG+GgAdiy3UdjdsT
eYbPN4j1+ctr9wZviAxVkBZjI8AoPGnDu/UxPq44RoqGYD6Cw+MsfWuDd06UVana
eYU3FccioQiYBjFTaAD7ElRHYIggDYRb2612+HdmTpOAlTgHKsG3C+1YtG/zTik1
vj3hoCTFM789SDLnX6NdX4auHPKPPYMpj1SKoBSlEaiHMa8akzD9i4MZ1lNmY0We
+j91/q8bgSp4drQDKPbZGzQh0d3cQQG4MmrghqFpPfI53gXY+MfRpTzRX8WwKpMY
12Mr0yminZV/Fo2aAD0xiav7+imTwKabyIe8xK7/tlzSaRYAoiFO4x4+L4Uw9/eI
GBcik5ZOsNRw7fvFSnZ/wLHSTN53gwu5R6rf67HGgi3TIneAv3dYm6joHlnNyD0l
UVBhLK0/TjpNs6hvRB9ExKqMs6U2SmXSysJwlv2BC5NpKszKPDvRahaFmws/HeRv
dKxcrrkgpEJjt5J/EzryUijHehAuLNCMDIceWJQtTAHSYbLMINzHodKOtz7IIYD+
/EG7DsBmS+PSGZ+trHyMaasJKXaYlln5z7GPn9wyizAwEg1LtQRqv5S3IeNOWIZR
dtN2icFPwVBJD8RjU/r7/0bfm1MCo0cwPoVGmqwmP5481ODLxeJGAi7kRV0i/LHb
ZTXkY8JefK30qq5lZG/3V5M2Rv5uw4vYbHYcuwopZeT+NK3JpzTxOMUWJfSELlUV
6FmuNvRDSNjxwsi+E/I09PBukFRkiCkSFLJjKStn1E3KvoOJb9byrWJHEzhKdxq4
nFXKsnt+jfgISgiGCtazzxhkdh8DNIKafxJt/AUPROvvhod/MondTY7wlv5viEYf
2GO1d3sNm+i1c02RT/wepuGzSNmv31IHPr+DI8QnL8GqhrXRTytDpGRJcIvI9nXW
68Xl0bJfbV2B7K/irX9U/UAwcNAV5N78NwOBFZLlnv3OmUdPEi75OhQvpFrC6Br/
kp4Rj646EDmpCzkLbt0uL4gxf7Nm5ogOEoddOZgrg4NE989PAIV9rTg1DG+xTZ8v
mmg9oo1VWIIYLyHB1273ESSwRobjeQvYEFjC7b/8/x8Hi74NAQqBZV/msdBIj5T2
bQLPme8Q0z6KlAn120U+dTE3dVJB0SLrgHC0rmRApHhJ88EQEQ+y61kWnSU39XwV
CoIpA+Q+DSxiE+x3ho9Nc3zNwZW5LgEDPpGDyQBP1+orS+splz1NIML/GzMT6fht
NNqX9E7sPkRADAOLMX+Vc9U1oBXNSfvhTAGlCjk974l1ELGQ7QbtlIfGgFI/ZW7M
bNl1OB7bQ0j/BginJOfRt8Rie0LsY6pvgaokTfExJ49CQfw6MpJt5fxJTWi8EtJi
JTv0Co5jVcBWTNLCnXYKv0j1d1J4gM9xQJhIJ+r8SrhQD/sF5C8023Y/zU2zfq87
S/GIcHo0edoL5KZ5recmj/cEUuTy0ABhC9o5JyxMi16kKSsqUcyPWcXumDVHKldw
G9CGxcJY7C4nVzP5vwXspswIcsrdlYamuqEugTHhAE0Uoude1IpKzCn1nA+S+oZw
c4fvquRzTFRFMjROeNO5WSE02GZzmidjAB+pNBnxyeVb2PeBpWKyOaLcI+FWD9Wn
+ePMeDSdITMUeHRgI4xZkuryePCBPG2A7M93f7vTAYqXjsDPBJgobadH/yfWu6Ra
oYqtA5vN3/qHxgXeUeyBzA9RefvGL5EH2JnyQWL546G3F6wUAcfIg7Ywh726jEu6
1mbgU98eRee7Dlsw8xWb5e38xm3KI42A2VEOqaSwc/qk+n0UutV60hj+BEAvJRPe
pifBqmBZjq3guNMwbUbED+dnJuWb54biZ8hN1YrvT93SsFafE/fz/DEqpiQfsPgI
9ol56mKo/FeZ0JE71xUADK3lDUDxSFo+Pfo/IUTDcgxcGdi6jDSqgXwup8gplaiU
xHc8PrDYypmx3xg5iPwjRRbMtCJrFv+HNJTKh27Gxx+c3b7r7r8kbli8GkAWv9C8
pZbB0aOiSw3R509DvnzVKPWBhRQnFv6Ea+plmVLgCrHGe1YCD4YTnsLIKGNH0Yb0
oBFo86nqRIFyFpJO9c2MWrX3z7G3Qq9syj9LtVMI9dEKlWEvW1gJ+7K3Pf3KLjFE
dmLqJwXzXQTdJeiAKIy7woy6Gwy9FiShupGWXSdkmZNw4n/7V6DJuATzo2W+gnpu
/2dSzoaLy3R7D+Of2/9CXZsBlcKBrPcZq+NNAkOjnmL1mSluGTij10IC67TuDVQN
+8IQOySeqU5cl9Uyxj46xnaxGTD9nh2NtgM9hwz+9EWqLRilNvpyJto3MgTyMNC/
YIcMDk5QpDw7LMaghT8rur7DQM4VSY35IHJyHgbB+wgmvCNs47ow/kcf07isXsz6
PY3b0o+jPRT5zUTNQWphsGLJ0i0+9fY9dESEEFyOEatX+Bi7G3V7MaBK/QtymtHH
uX5SJfZXhMTD7D4nOT4dDHOHqs0r07qnTzz0YGx/qxlaBcqch9AH5C9rzurENkPz
uUJmwu4WxfLrJ3xWq3TyTaWL+a7IUq6bh5uk6bS0N5/BiPN7SIfXGuLI9aFY2a2A
11CNXT3hACLoUwhQB67leDVk05/+R4lEetN0BLMrukD3XZQUlRi1FJUflALAjEQZ
wasncq1Kn3WqPRRY2zajqnub6gnJe/fvpNg2eBN0NAk3PA+/8Gbbcpmq7NJbBXUD
8S+mxjrGKLIy3dNP7rIA3NFz/aT9QamWPKMmKzcQxE7lIAwlU7nANBGbPdc9JGrM
LuvoFGVteB/PyTBqos+LoSXv1tjyJveFErjqsvBX18EIAdakJxGfCp6la2jUbdsw
xlnED1Rn28d4kIJ3HoxnFv7TQOTPlB7Mts3/CdfUHPDDwiA6iPVWN0B9wJVt24Xm
CSNC5S2/YUVLiNRgsZvVgYG6P7KfUFKbTTQlQxq8qDsZQzDmqOT0rCotvm1o4aLV
ovMfmg3HeK+3F9gA19AAbnmRmYTW3TZWRP9uHr+heJExLI0mVIQr3wB0Ryy76V7P
xNtn1zhx4uhxF8E+XiUz1HGgRDVT79DhknPODF1HDyU+6KaqJQS2oelkqHEbBnxU
ccRTft7YkN1vvxnFpVVeWBlTJw91IE49ALpnnum92kMOJZo5T8V+zot0qnWtgAIW
IdGPYf5Vs1VtOyP+O1+0Pc6IAA9SJ0JvXvujpmHg3xfDJLVSqDlhTJgaafZBWA6c
LTasegP3A+E0GaaY5wvfnBG/YDuLiXt1ebY3bw23gYURe+74PMT2o9XO+kLAp40d
LSbn4fmxtd2z+4q3QhnRbQ==
`protect END_PROTECTED
