`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V0t9EwRzRfKqkSPds9RyNImMh/bK/8nky3kSb6ef7hhCPGJGr6/PsLo8eF/6u5SC
SbdELjpCUeifK8fjaj2/3pfN2FTDQa8QsIwYui0G2ALGi5ryA5v9YA176P/3IuPF
MjTx6pum9uj6g3XXbKL8vNBeLsF8KltDZqVre9dFrE5AX+uCLKTUxezq/CblfgM/
lJUFzamlRUyJtgSwDjGwgESyP474txWJFoVQtxwQjJaloq59ynl1daCDhFodIqum
qhGwsKKuPq885YcbYeY0YKI+Ibrd3Z4ToYpTgZknpOqWT5bzjNkCzb6jBWE1SNqk
FF5Ucc02fTVDeLMVwgRpAEpeFemwWjXFQGcJAUgExG1G9vCLTPIejCJS9UzYQ6iS
KKdWb7JVA1OBxDjjvU8UVajFDxwyFaGlD3A2Uvy3Q/ty6QrlE4aLUHUITJk1yfJn
cTYdOtIPMcOLZ6lu6WFLVaSW6DpH5MYjzTLk7h6cDYbF6v6mnyX/wyDFhTs1g5s5
ByZhpHkk2QNO65yJrgpOt0eRUWaGcQ7MO96UcBvyIG2JnnMd4M7r1x0dlctJ9who
ThPsR4MMgpp2wdQpe6ngT2IXCRB2P6J42rIHRZJMoIEJ+4XSLSt2VGXONq1wSpDB
Mn6m6j5YKcSVKEAafEUx3nkUa1EBqpGFgOvLlR4A3UTLn38Lqdjdq7Rb5dvfq851
t7+mtj9q6Y9ZpiRpTkPuE3l38nK4IaUoWfNFiLp4c0aC3Ap7iWGpcnmqZPpSSoHB
V1s1kLVZMEKTPnqqH2sfszXTB8P5ttUQAu1ID4ToljsWr8k49aPNDf63e1W6TwGK
pg/ATSiSnu8z0RAOV5rzZ+kEcC1pOJMBbeCkCUuo+WdsOWymosuNToCbn7wX6482
o++FgGRSlHJOCbZ0ofXytMTRneQI87Ce8YKkIPkOUHd5u1qcbzj3t5MgFqN3MyHI
XY+JbJajea4RbcR3LyZeQgr0XhniAINvhppDUJr8jk0ldr9rKSKvOAa2zcf369Ei
9mtw99IqVc/RRglNo5LvsflRFMQcXWMDo3MyfhVpJAWcUYOSeMnJs8ijsQUcM4W5
TqN4cQpT67Wqw0uUlXjBydloiNot6QZl6USpo/LrxiZB0b0HsD55c+35Mzw3L6mu
pvMsApA23X3ERFxrVG2hDvWHn3VSr1VokbstLTrfausWfoa5aXHhaPskfQDwq2iK
uxxCxKCcEV3wOPySbou3Sp5xrCdkXJhMhSe4sI5Ccdv/Bv19D26ieQ5yj8zNY+0u
Xc9eIzr6AYBG2H1BqdCnySPKeyauuHjzKRx9tAmhWo9fgAHIX5RLyF3aBvbMNNNc
geNR+IuHC+HZdk/UzXrFhze6iEbFIDqsSRGOZsuQ6Yw8y3E66rpxQNczPr36WiXO
vxvK6dfsi4UfzrfmMMoxNDzGJOso9/Z707yeGfHyC0OdTNV34yu0aN4CC0xdjeVR
yhXzgiWrVtPmoJNWtbzfAbwcDn6n+SOAxHvi6sviha38QEyaL9NInSgLPercBBTk
NuWSrLbW9W+SKDPIxkjTFo+L9JwP2pYpxZ41oF/XCL+f+giPf8+k1EtdjlwQWutw
yd8gqHHlp0yt+LgHTDJpxk7ks5onbsLxePXGWwfyX4aA0J1S9xwx3EC5L9tDJBfM
sI18SI/x/hDDeSbDnGDOQnyzsD5O7P5Zc+FvtDwC5bLl8zr4mUaVK9zVqeOHGRmp
56+Gx0JYf82fxba+TCFd0A6ZM+k/r0LzWN1bCOlYjCDe0t33efxzzcdJeLLyHRfz
PYJkk6rfDFiM0gHZqgYhuzzf2EEUgO0iEXyM0zFLZ+0pPbErEmPMU7tkUNLmcSmI
HSfkV98Qv1lJsiFrE9PmctCfh9ySTOE2TbALPvweU0utr5yZ/jXwk32NSqAHRWMx
7tFansdAJaX8N0t6nWh8H4JEoX5NlmOoxYQotiyfL9Zp1f8xnqNjKeytFvMTl0q3
adeGeNLepSrF8dpHRJgrrClZniId1HFJOcswb9ml6jslElBv4peDYbOxwV/UpTLz
Ic6y+lGT+i09ybFrtUQRTUC79QO5k6laE9l1w32VHtkaXYp1WtidfDqRXwH1mMyD
ZWUbkBMqRTaMcKfCleZnfsY+4fDjuh+8639K3rROMqLA7U6/j/ehnmXCsSzQti16
cq4x57rLCuh2cxb/wyIt0TZZUv5i6XuV9t25pQ+eEUL0Op6R3JXe+Tk0s1mVbHoi
AIsqbMSK4dN5F9bjXtCed2mZXEZ+ca/hGAxe804g+ixLf1HKz7X1s1R7xP5ZlR4n
xe0e1fTtQ+bZ/VjnyCKr6FqrHF4yT0VjuZiarQTuUThm9xC3r6UQkG0t8E5sxYEw
f5Hawc4+9agfBVWIGSziF6kS5/85jsrThdV+rpkEfj7gRffROSJ+ZYLw9Rt7Bh33
wLcjIPQJC97VQXi7lEviRQCuC8jIU1LsgjOieaSg44FqHLuFm2gBHB2ufsdu0ZGH
+Ir5ocNhDQzzH8R5yx7kw88SndMy+Al9mCIhzBof5MOlgcrnnTe/D8iMIDSTHoOX
lxvwInPfXh1fnzPCWnfTpdIm0eFgksQeoi2PyCvMKCEZhMOMjDt8e6el9PQ98X6S
4G5GUltuIcUXmEwJbXi0eDYDrCdWSpeVq4EjbAxDarWfbI7N8+K8JnrL4txKsSNw
f9q85xM6MawyjLcF/4TAEHOuZ1ucZqmves1jNAzDabcwLLTehPAgJzu9+PYISMsi
8cekfE3CqENm3x/JSkcfeCaOM0XaKH7uWegOM35GTPghaqHHTd6ZGSfNE6L0pOKi
fD5ng6VoV1O4jzUeebKjbGlv/3T86rSWFtb3vQvHTwkEYS2r9cVUupAu6qmrLbR6
y2RRXBm5mxBjJ+Rl+/NHed0r8ZtiwLP1FtSVDyFIP08T+fu/bjKCJr02SzVFGCGa
Tpu79I6lgtIc4WkTIgOYGqaplVBaEi6w6Yu6nrNGeREwqjZvQZNrx4o+wfWehyI6
1/Lbb1spaBytCE8vfTkCg4fMZxkY2OXdWwwqUvIXSWRPR67QsXHNdvPS4lg0604h
wqt5atS/TlayTtaAwTQoyGrghvoZM7YehBpnNn2Lp4H8CQqpevPycOEqUcuHb0y4
dVwmQawIhtwznBrYh88Ga4P4b67vqHYv9HAtdjo6Acoec16O6vaCfKd++UTeBkB0
4HmVS1uz3gM/iSCv/4jFanqHcCv4jw7Ud2NEexAsJA/LqBiWXTxo+qH1GwJV0Hg5
s9HFYUIKgtVZa0fayt6wYTRwFNfBqCCqR4Oy5p0DnSCl1DAx4pJ2g9UWO0bOd03k
26gwB98n04dtIHqtIOy1N3tr8EA35ZXbfPgJ6shaBOJb9QKY1sMB0tp0tHEUhKYg
gTfQ+M7K8/DKsZIMVjeXfbgg+pN1A6zNsRorVAHIvwPY4WTSOy4W1J4p1Zq3Y0m0
`protect END_PROTECTED
