`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u89n6D4wsAWxbD2Kkyk3asVGW+FhsD4rwzu5iX2X7HV11NnBkETZ1EyS3pZA5VTa
hJheoXvPtiVAkfZJhWzuNblDbyU6rMXcnQ7QG4FOE8pPyNgAa8xM9bcX9fmnl9ye
cGHH/mC1yOWCf8B+ZEW2FEZviRNcy+QwrU12NMsBsaf8PyhBA7t+2vszS0a546ZK
qQ5t2CRO/muvl128nJ1Lr591MeCTMhHDEJI9tjAoUGqixwsnGPUnXeYak7ieGaW+
FShrikKkarOPhNPE8ROWIr1w//hMz6TMTRrI0h/QBMHi0MCXjxiiNrscRG/Yqsn/
v/s4O6NTq3g+HobsJMU/w1Dj/fVc9CebJExhb+3d3mp4RHZhj2JY4v/k4IM5oTmg
IIpx/OEcgWWqvPmymPPCZAVfE9qXJ3reP5GYI4Fp3d9h/CgV72K4KDFCFo7jp3RQ
NsxPzT8MRHg9+uzflhw7ekRPuIt6pFxDSJMSvP99Rd9YjXec7W0bZVm1xRNagJRg
jxdposGpXlFnAWMH1dbMFcOpkRPTF7SGDKHi4iE9ZPKT/ojUB/HyBlmZNHTYlXaG
LA4Ini0LPhEGnbkRWD2Gbu7xE6mIIGa2etRSjPBk8uYN4bFlsL27L9FNN78REsS+
EwcXHMSsiq8QG28BzwxkgeeFieukKAjtp5Q/c44KpTcD9De7crH2ZfO2uCT9K+Y0
7ZJbZZfB8c51NMfJCBJxBfPDAtgx1TLn2w5wldFih5qyWx/oiHIQN8ka1uRLwPGn
aNqu0c27oTOTFIekaiUCoCqxMVtYdURwlFT5FsQDcHGo/f4U52emHcmgPrGf9u6D
l9qtyo1CP8xQ+U/CP7bzYtprS7L1mFygeCLfCwQluiqoSQs+MegIqvix88nu+d6D
LSf5LyZI6f1YcMgj5PWqKZPwVu6BPsrRU+LO3UHfbJlR6exRQlyK+amVKKNiStaK
vVL0e6SPpSChXo/3AnT2rnfuUjt1ucHl1Q9CDDF90JicW0DjJYCKSYTfWCUoBNv3
DYeuNHNCZofnjp1g3gG2N6/u6zmcaumrYP1tAAEXMr2zLiYL2upzAa7D8SLKAdcv
/ltdftT+TYyTjC7qotlUisuTGVRVkbJb8f+wSRPeTfCS2sRjh7vUepwYLKEYYx6D
yEWAt6hhldwNRCy6YoTqjQZuI1NKg/R1pY5GJyJ/KLih34NNBswH5N0lKm52bUlh
Cu4DpqIbS8V7d/Bx+vKv7gdGj5+x/8Hc1qTqASdhR259jVK9TuhahA0tim0pW647
AjFdzzb08E9vHbr/1SDmKqVBs/+rO1vaI/u/s0Td55+7qRYXBaUY9PduZmP/nWn6
6Rehnw30SKywdfPXGqMbe1QPELkVn2tm0fQA1VgHMhMfRPKvuZmMWSfV3+9g7MJg
cu3cx1yH+7CuGtYe65YwMSaLSBfAt90Qu4KK3k8fkuSEdsd3BO9GoU+RaCWKWt6z
XDJ7B+CIkQBKj9n9a8w9xGysfYGyikcrxEl6lgo0mlqBAIqodHEbQj+eq57KVtQs
6rf27nS6Ms18JGwgtGs8unJeZFer5dhDXNo8h+lBkfq69Y38RhmXwP+Mp/PF63kr
ADHaUEKP0d+XZEaq1DnCA6KQpPr7a27JB18XqEtJgLP2Khf2I775DuxHTFX29JuX
iku6HzJOUEJcD30YZbNEIZGFxs+PpBQTZaigs+IZ3xy7kW13NcQwrzmytwlpf2eJ
t+ojgDtnr0Ss/cH51zzS/BAARd1tc1nM7rLCiFU3k8MsaEfek4e3JUq//I7JrOqu
EpGj2o0RyGT78Clm1ijI783d4IAm20O2KSn1z4BigyQ/hgkP67nGeJFlBMTB7adV
2/BSB6HdTVTc/IneBE7CTEUH0YJWch9IXVmv0Yl+0IO+o4456ijqvHFW96tMw6pu
OjyUqx6NNEBzgxw+RRuvVssguw7qIjAgImDvDRiy4qlH5Oc32bqros1mnBxzDv74
MMRBV6odE9+nM79H+HoIOEsBUGOUHq6skSeXCqQhuTRJ/SYsARnqLC8ffwu08hEU
MAVLGC0DuXscX3B8ecI7f3sabbAoT8gjl1QKfz3cEKajQ9Cfy0mNOimT0G66giXX
rABdVH3Ffo9tFVR/Sjzjsf7x9gCGcRrJlwvgXH1AgL7atbqji8Oeg+zR5XStdqKL
C/Os+Yi+M4J5hwikLkHEtwKKwxoNv9pc95uuk3RhA3EIFv+j6lDNLBQD7gHCMygU
4geZlKx3BUV5JUM4SrecsqzitL9Cbu3V/v+UwMizUZjZCM5GYt8z0Hg9p0e8oM+P
QYN43ey5uYSZju2DcB12Eokl8eNckTrVWzAnEPRN1Spt17grGbBSliHstcSkYBFq
N2AGZcx9sDWKiXJtDTyYR6+GacVkc1nx8oGD+FqfMlX5O5lbunpORCITguJzIU//
bg3sC5u3qNji5oi24d3LOx5uTae2Y+v6x4s7kep4Ah7h3i5DnKWtyiXIlw6PL5vx
HJtyWTGz8WAH2ykWRX73/r2m9gYMb1ini3TQIzYxqUBEsytEGmEdi2vAv0NfsgZ7
6IkphI8O9e80lChcf+69u3Rg/nk0dZY8URECkeXtMo25DBiTnTjHUr+D1Z6ZkNSh
yGl5h5ZbT9t1SxYwqHUUBe5Gq8W/QKoPJhY/ICvatlXT2VFrrGmo1/5hE/KCFt36
C3AevhXq/vGPdS6gjL34EtjQvzBy1DtfOrSCv6qiRPisKNIQePwHqand0vuJNEbv
r8FkV2rM2hDp1iVQp+nfntSiEql3X8tDysI0IGg4tvgYbmmUnya1ZLEEWgdUfQsp
rtUgX8DQtVxtFH1BfZ6DfD9RN3NlzglcgdfqIbi6X7szRIbB9tkdHagNm/NY6Cn7
9IWQPujvGrkqDEe9camSh8O37/rimPRloSFm/v6Qr4UNU+JdaVN+F7Ly3Po1NTqV
qGSHXEacxn539sJQMvGi4iNXxGZ5SxJt4y3XxrQPrwvdH3KhzPUvCQrfpwhEbf4G
r/qkKMIgt9Ohk7bMd5VdvCI4gKQfiC7AxRO5XGzEotNe/hh/oMtELLCVVRrox28S
twzb7ryK7+FXfthOjoKnXowkVqB86rPw/W5jwUrJVTNzwDaAb9zgbiD4cCum3nZT
o92cE5ZV9Dzlu2gi2T3NCIGrqkFjH+RSlXKAuxvK8cBqv0vFgzYsXQ5aSl2DdjM3
lAcLyW+c58oeoRJOfZMXQAikvyry8ONTfbro5K4bWRo1dul2rnQA9TgVsSljRuhm
rKUBmBYIFsq7vq5bqQ62pjeK3SXu2z+btAEEX0LsbzwOUM6F1np3kUftLiiwaC6O
TRIFuOj3qX9GVPf2z2A45vuhhQGQhwTgOx60P0lBBmXH6K07K0k62M9SxOEcQnBs
FSkfen5oqCr17kRuuDHiPKf7CX/iUMyqV+7fTpRSwlMtN1Gn2jJkNvOQU/9ZgjVy
khsvkPy1JqfRqOihplOb20cVEcojxjGjGzZkkZjyztKBYHba1hqpjo1Dizr21nHY
i0m4QQTGNnigRmCNkZ2r4zXhmQgbzH33D0YxovvOJ0+ODKzh8D7v53XCpGI5HkLL
1YD2/sncgx1nOzqrrCTRRvFhuqvLmvU6x0EpBIZhHsLAFhhdcQ6Zucrwsk55OkzV
bFHaHcZCeje5pOXxmuTwrpbRYhIvg/RbrCdJsbkK4JI8gynGH7p2msYxrj5NpAHc
ky5meVMEkULPrjj+ksR/kKxu32vJX9vtL1XCTPhYjTkz7YYq6KKCTrDSxa//FB24
f2oYvgkxB9vqQxaqMIPCQNLsZm5fm/MAWmUCGQtP746S46PPopg6/fuPyvH7WcXv
K7GcGHhot7EMnp6+fE7OJdjhGv2c56DesrchKywTQ6+wp4O/pYACs/YnA7l0hx2f
rrzIoUrWzv9b0ZM/yQE1nfQx9kUNBdjD77QzzO98kuwuTzf3075eYDCoTr+e0gfr
EBWyc13j+xbbOSRwxPV/UB18MoKrll+7SedPKutil4bdn8ELbTePXq9wtIfdW4JD
zznRIh+MN3IZnxXQ72AmyzaAuUqFwL1NlCjq8rOOIMREUbjBuIWQmjUS6DJBd5p6
Du7fJlKCv1YQKrrBEwj1iNsW89fyQ2LuBHW/6KJo4Rie23SC8yH4NTDNXtvEO507
ascE404ubjOu2RM3bg2U6OVOUqqDP/DDQrfHyeRvJNaDlhsEVgE8YC82PcMGmDZ5
R06UQ9f10m7+pfBlsIL80o2r2QjH32JWN1z1WNjWZGHXJuzwtJGSVb1ojZxv7CGX
rgs4KxbAaQ0uuipI9jwQ67Ptc+glNWW5okteR1aocEG5uB1oE83M6ovNndRq5MCa
vrmPPUSZ6EJ+0sy30Tf9/IRqGb5jQJa8Go5DLo8maAMwnJXLiU/U6PW+sZA6OHp5
0qc82z6BazbKP0BquhDKqaMLHVDV6+VJ5C7jv4cpi0T+yyHaZblMzGeV5elJQQ8M
4On8wDjeI78+UDzD2hEGfKVleXDABr54FrcRBqrFxnGFZoncGgpzwuKDLd6OVjk1
3bwEP6uJJWE3snRX2NH8RVORNWEXoPKOEBz3Tr9hS5ZXhXJqUm2CyBN17GGOVptd
UJ7ZxPCojdOUOqCnNgY12VCz1vX5dahSSPaN4Q2DoGrvFf2K/GEQdhmJOoDkRqv3
/L16wmN8RxKYnTEPTbbLD5T4MxO1R+xQs/FcPliJ7WwG6m6LbHzrsG/VkRhgFiHZ
A8tVGz8ZEz7Uz5Mo+I+JFNHiAvHM4GxmyOrl9vPdaFUfVx8m+YZHgbWPtKWNRmiC
dabdqSuyvm1LmKVpRaSwDtW4L9rohe/Sl9H+4fqehjfDM4tRM9SwDEMcabdgCzWl
SaXd+yaziqmfylMEh3aoFfV6axuWl3aUEPpBJ3IOcHWdd4MWuPWUeTmyg59Xv/a/
h4NqQvnZzcL7BEdzK8c4ZCFLJ81N0r69pfwnChrcve/k2B3EsruHxSbYMAZUiFUg
k8QJ/VeTLGRApcO8xQcc6ObjLXmR5aS3kQkYNQMc27PIraNRXnav/y88B6Z8ZJPn
WG2hhVI4qrBTilFnXwO0ajL8F8dkF9Fdp/3GZHQGRLEJRpIfi/9335D+xsuiTmmv
DtKArnoCnPUtYu5oUStlW3r9WBrsi5jYj2lEo2dMtnGm5v1ITXe8xbl42x9fGtJH
duJc/LQMrA3z9B+p0RTLPAvxn4kaWcKQj0cI9vq1PALXBg79T3JaFLRiDrqo0uMt
cHPJS25RynWBBC6rUruD9bR5rUqcf9gC5X82Zt3pEEhUsQFaSeorD776hmYPdUMo
RC0vBXgiNCfy4gkc6bkQD9/O5cOnTdCiVD6lCj7rCXdkzl7neEjuVFd3Iq7JfGyH
FZ9KoNW18E3ujsxFHekctzA5p3rpEIRn39fdTmxmUMP7Atxd0XjTt8fJsSvbn+UT
f2I1wiolauowRxIb9J4M38jK2zoj1/U8PBDmukzfj8jBHgbFQfa5yL8L9BDu0V9i
BmLWysJHPCUYadw2hRq7V50G++FNUan59MTRdl65Vppe0eOM/08GA15r2d/mQj0i
2GsBhaoSfaL9/0fcL/FPwPgVa/9e4tLEUShkDlWwMFpZruyGY24sKLk4ifdg4lae
BLgq58Ck24J3pb/XX1AF6VJkLy5O1JAwrMB7MHfg/LAAsFUP5SHgsnvatcNUHVtl
WCPVrbtqdH4HWBZ0REtUPOcf1Z08RMG1g3LxkwJQ44FJJPD0Q31XwhLDseZF0B8i
BH1W+tblC70labB+dw/N0cmnCZ61+OHYBIWX8BcB3pbJL5tpx6jOarZLu4NN8Kdg
lK+9ybXzx37CDwgyFdqpTfpBdxYiukEEUZU5GaronF5D56jyCKLQdIqDXo2IkWoF
VjkI2ZB0eRqIPO2pxdp/hGoRuTac5avqh9lVxy28wwyHTVxjUvXZsSpu5P6WUkgN
62V1d3NIMijaDYtzHkYMUq8kY6LN2y1+1a4rCOdHcUBRlMxe9iLoycx5RJqTlysK
eD8m5kq8+eoOSBIeF2IjWT84CY1FU84AY2/bulgryR+IIAd+Wh6KhZ6woyk6dQuo
fWs6BtXx8/OH6J+8zBF9zroSWw6JQ2PBFkG0VMDRbgaR1Wnj/YowMzg/Zk9QRBk3
5+gAnzyJMhoTz3oXxFsPQR+EwbstrwnQQYnrXKzLmvFlLFIA5u76Odk0hUx7Hu/n
GmXgrftUIIzTYKwdMbhbXeYadz7RXrGSZd9juDGoKJUm1Yzq8L0zfQ/peXkTV0Q+
+oZX9tjxHxohO+sqzG6G0Pyred1gX9sLw8+zDtlWmHDrMdr0Dv4KRPvFYKjrZBj0
7KGEOOT6iYNEHWqXMQeM0TrMHwii6oldCqD9gT37DmBkop+HeGyjWbvJcyEkiD/v
zhy6Vj7cJhnbt7OJFD7y2lVtzUwEzaVl5MP2mGB6fgRlJcjugOAb/sLMr+rbjI64
n5m2TJZRK+JEbWLpgccCmLEWr+jOC40gFiTuPiPJMsXpxyolpG2xvD5npkufnPDy
k3JPjYV9041SqWPeoMiCfPT2Kmr5JAAs2rjxebeSxeZ80fViZhdfQByoOl7W8/3s
PxAHIfhhvWmE/8NnNlmj29Kyjhm7foJC2TOD0k3dRtw5TKsdgHzf+btgCX0tKrx2
TCjfI4jVDBvC62hANVDY9KN/ekRZvjgFqbvSkqKmpSVKpbrBrxgxZ8vNGdFidy/K
4cDdixGdG/1KPDLdQiT0DhyB9HKwPVTqKz+b24rI01DGFZZLxrVkPQxbsQoPD4y7
7+OkuRtJ0CQL5T+UZqA9DQ2bS2tct5WbEFIE7+h67iYXPARK/xVjA0x370PH17eq
r8N7P56YAf3Ll40dVGRljHM+VPrRKZZmXYl94jNourCHwDhPhPfoI+x8zGWUE1Hw
qznr8xIG0gMrRLsHvRS57iR2NqD5uGLzfHoUGHpUrq9GylHu9+SelZOZqqboKA0j
sDW1IPFUr/qYDQEwHeKK8kiGOLMCxmkyv8sTiGIQbefC4ck2j20g72A21vJ9kv1Y
oHhlGDDULdNOKBRSayTbcgpOevBgSyjGDqNC8uIniEfVuxYOqWN+/1GlGoykeb0I
`protect END_PROTECTED
