`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IekH1Y2AhZaXtDl9yoEtk4JeOMSVC5QOnWgMzs5sw8p5+1N0zYOi6jr7zPejFOwn
rtx7jBmIpWVl4n6q/i8Vri0xJsKCMsaGzuI0pyGDTmx0IeG3inS/ACNB9PzJXkkj
Oq92gZKeO8uKdgAh/blPC1U47suLgwTrkn/memdO3PxtNsj+MopJkP0hMtLiW/z1
WfKwS/PPRIF+DxaEM9XlzMpRbg+HXQmATieoNuHTWqhwpe79XVWN0ahm6bBhX5kC
z1elD5ZMNb/CFbkcmWiJHQbLhUNCPIXKui86DCQmmVORNysCPQ1o8uPSh5c7Hmxi
lgMFr3rtTp44mX/no50LD0cldClTBmOS8ufwUT78Wj+Yd2Q3Lacb8vCILhQXQXIC
d6w1YCmR4qS5dV4KhycNqafnCS7IgQdfawH8ri+FEJj92XlJfOVJo7ORNT/G4vi0
OJzVVuETIFRczDQnQvGz37gtoPTKZtA+YUtd2sa4mk2NWeb8VfR4LNZ7w9FVJ8qs
yCxZbq2OqxXzdlinP0DRJhZ/YnTzKqaikx0SewtChQY=
`protect END_PROTECTED
