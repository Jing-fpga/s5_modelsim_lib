`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+NJDJ3jd+GUJk17tcn9J0XShP6h8k+jxZKqMLG+YTpgXBAfAKA12xtiWnVHW/uVY
ZQdBboxjV+UAkDA+dfhVHkLdZPebm/rl656Ck4Fd0LfxIIEYIHc+FiT5AwaQ43Ke
J9o9DayeMuSugPD7VdK5VSB3tMK+t38q8M711OSN7h/2YrvPVvMtbeC6Q8T/+38H
98Dub+f7EocVIO1qSNy4N7g0YxAAMonyAD7WUCEde49SUut8WzNJOwlsHTSNtMYI
YuUZqWuGVzUn8ZsiHxD9aSl/C//EE6y0PSpYbZv9sGK4mrVH5Xg04wAztxlRCHE7
WKIdrW87YXjMAv1QrU1bKVGbbwrnxh+YEn9WaT5SFNS3tfskigzO2THQcUhF+gtE
8jcpaYnv1Kua+poYJ8DcjvDDz9f8HBhqD39/Tyht4QedG2bDldAGRBkqnij95sPc
qQ2K+poLzrDs5cfeKN0TGv+zUn2P/WMbrmS1NjM+ibRA7bAK94aHZ1hxVdixslH1
3Vgbb5w22WZ48XnjXjD/JF6UA6i2SkQ7uyoIh2zbx5jwkMD5dHqmX8m42U1jLN6v
E3asbNuG9JZhB2ND5mhKHKJE9Y2qDwfXbNpOjZy9MkDaSY5QpvVd4TMOF6BsVROd
pxAoxUJfnDsWGQGG5ByoIdzjjzCS0JosvhIN6dP5qpLUL1SCs6ITNi2+PZwWYp7K
ugBQQK8teSDAfPR5u35bPgF/WavRouju7yZmmkCYO8RPSAmoMz7CJYFh56Z7AONN
MJUystxbfHncm6FMOfFQLFGWapXfSpgUDeVcFrbWwHX7cGku84S8acjcvuSwPdDt
kxg2C8IyNbDJh+cT1meizQ==
`protect END_PROTECTED
