`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZfFg24IYQMoDPZm+1vj1p2ZaFVT7pQvFjlMc2f8eirTe3/qfX0zpHhkRsRX3UpH9
SmohPwde5/CNcVnkfbzpVbciE0LavTz9qrUSGBn/Os2xftgtHBtM2i30BnLNDQLB
7Xp13ALBKQRlCtw0JzHg/xeI+0YnLzV5fEWW5vnBQmS6W2mKBEAHXtsJV/BXO/6E
0wTRUPWvb6bpH5xdhHqsczbx7vrnr/VhRO1QyyQ+HaE/ctXLNRH12xQE3+z3pEsd
DcoDo1bXW0mJw4Hj5EtbHgiwrHsg2+1D2l6aYtUjAu2yWx8xrV5Iodhycr55YZ79
i+QhgngRY+hm8xDJT3ZJAuWUG2nmr0HB5NdJJ0GObLCwkiR954Nm6H4ee3gt4ixO
30D67hMUUKP7PGbEJ1up8LIu8WPO78N0fXzns8KL5btTa4mWvMAo8zFu8hAznH1n
Z+oDyDsLzijvOL6mvOIFeVDYettVr1fOxxH7UxRsC53vr5Ud0shT+7n7zuTgj5/+
JzNJZBaY/TgOLo3WJsXijSZz2uvHWSvEFbUZUr3jqAxC+78T6y1JtNJeYRf9wj9m
W6tkvIfi9a+ad6B+poGQvdejE4xTmcR0V8se0C8riWkJjAdvacVSx5Lu36s488/1
i+WvyjlYPGknDngCLb3WXXRfdE36e71BHd2Zkg5XHlyv554Pzvx6byeCZ2aVxSJR
gfM59TKKlLQyv9sUhypHcfLvvNdnl73kJMAJHM4Dy2uJG5Epmvu+5qTFzbhpnTiv
KLe3eG/ei190VQ7NFpyVBbF/jveKjcUcjPcumyuPOWHq9ZgrlrAFTrmIyB/nwmuv
7QWXiJHd6Ka+NAVanxLfl6mHgaUG7xwN4zxSq/snC3lGfw6224kmyymSsI+Aq29B
JNG+aEYK7mCupPJ4pkcO76MXMfnEw8evYqKbEfFgH+oUoxPieXx2xgvkSk3toODx
t4skyAhWokyRBR/Yn7XPNiX8WxCHvs0/hEZ40ldm/VsOSvXkmB1Cv5d8vK+IpsCE
Xy2HxIx6Ji41Xmb0zRVL+YvbwdKDvzUYgmEXi0Fm0X57hZdSqCLc9VRJ6bMWu+Xi
oU6MEmVeOKsG1GRJfUCYxNWMGauqfGfsYMuQco6t2KgQl7sd1hUXgy/qPeD07q6O
xZikKTZI9XA/D9C4Y+f39NwwSD+uhu1woO65MTrEey3jAJj5tcxwQmJEgl6+V3lh
dLHU5lFRRn9MZMYfvMel1pMqG0wRo2x8Tl7NdFXIAUKbIbLItownTIJpeBABTIuV
p89EO2jclEWl1DHNnfQLLZdsvkIFJmo1QbfnoAlBBvnucuHLK+F7Vp4OWpimkEdW
hIATpaxi3P/G7ViMfYjSHd2Be8QcaPmEJ7LzDWZOU7CE2k1BWaVoOeuxzHZjAkxz
ejHnO3rwI+EEkNJAswn7DVQvtbcguxuPfXs3lBHX8YGvnHn2Ef7hAlb1Eo8jh3IU
OUcO3OI+XNE2XD/YdeKg7wydiwXDwXKYqah+Ws49jSWYbh1+VkuCLa6yxxKYvhKc
uGaq7+8TCAo6nj2OnwpbfNNsmzbUlnndsKGtQvDKxWdcPMpwkYhaHP3pz8xDTNlp
GjCbjeUpowwQACBOQ+bvxEVV3ewZzHRnc1hcoFw2tFHBjVtBeNZWrDy61ZSWnbU2
5OqZsR6K/YeQC9sMaAKOsn5rME8I1W5+1VOLbI2ygJN/oUFsyDY5t2uNFmFsy8FX
DE/ukQ4x4hfPLoDqsH5HUfHQyv2uFRdLcNUhsJTfI7FG6ZMSSHzm2S3MS6ssjc0B
9GyH707lSaLKMqtlDSFon3fg03AtQxQYayjiTa8yhtGDQMp3QLFbOYdn/CdX5fkE
gdjeQNnMK3LtfEU/DWN48vQWhRJ6xE7vUf12i18miQNU6GBLY0X0zemn7z1WacSg
DwaOLYN/+kbfWfdWpA4ai8CgerHwoSZpg6JrYLOMY+ydhJ8cVDBUlHqY65VA0WzA
pC6r8SNVC76jNTuxx3h+U08Pb33oAOm8GcTYIrGvBnKhZMjl6WPNhhxqCcsiTlKc
nmVp5Go0DNDkqVjrSBPhksrQpLleTMlM7nZ7hpoqtqaH497fL9JjfpchXYJBdtV5
aahIP6yiZd0hVopxDMBqD3UQur+aJNvUNBmEERT4WintJ2Z88M0iR72/oqnUh8HX
oNCmjNbaPjYvbknus3xCdM0puPhaL3X4rFUGVvZ+obqHJVciKdD7lxsiezVYSo3M
lWq3mTLuL/FXjY4zFpil32RdDhs5kI9qmGFtSZURhfFe61tJy8Ux50JpPmWoSWf4
MdVcZn/lM4bgV2wy/oU03mP/GzrFGlxodRwBqnU3tWlFcyIh86klhcaxkOpmGIv1
fQUMhZULs0pzyhsHZxkRRfg2b/FSbuceItsJvHDBeyK1vi1CXuAGRpQPSX+mPmhc
tZZYpLXyxbECCB0A/ZrHnXYm+5Fs7Rmt+ndFrrRsmaYy9QzBzjURRm11qBHsIgCw
hHpvTd5GL3yqfPbMWn8ZoW8pYnGDPObegnH4opMy/kEErQNrapQ6KxSqEDHLoFHl
+/Sl+XlZxSz5NmLBQHrAqTxerZmC/Q6vX5Tt1PEqdHjZDYIuRoqcL/89n0fH5ypI
wW2a659+sqnTSYQeO7fFbnqnnnR9KpkP3ozgy5H/hGLC11vEMz3hMidNBRQsbEhA
L0zwya6tc2rczKG9GsbdNZFIdMYgc7a727d9dP2HT6rHXyLFkkTIXrFuDdP8+zPx
xr6SbBycF+CZii+YF7i7kcsYRDxM5peD0yzcx+siDvd3i2Nn20+xI61g1MgTBZ6Z
HiclDmP1aOmFMHu3DLOvrfuLQQCJxyI+Oyq7RpBE3xW10rMZ5AW9K+rbVDtQz0Xo
JOeQoU0Oj2Hd87pmDCNq5iP3PZhxud1EP8xVpm85QJo5YrKYGCltY8bUjk4WnQVq
Zxxrvye0dUU00GS+K/xrntQ0CotqQrztbS6FS5jJDjDgmdTXN3sNqru+vEZK/rp6
gyiBZXvkNsRaEhBWC7MMqlXHjPJAdxh4t7/Uk7EwbOnATSaV9FsA2H1vQKmvysNA
ZOsDpyMA7tU50TIFNqPMAGMe4s51YxZ5582RJje7s9TXIVfHqKYdg/UNnoB43dJ8
ziT5WAreWHhL3Bq6Zc6s61rByG4b7pEnNrYdp1GdFqOfBXyUbYpUTM+SxrHYSWf9
HGPS/d+HnmAvqRu31vqD/WJwwfon9geGqT2tmVZXCCOb5j4MHkd0jUm1DF/6i028
i8uYhUrTQFVPOsBYyMAxIiRZiQ+694O3n/QenmYkpmT1Hlx5+qKSmAAYfqzixCQU
o2n1mvzVSyB8qYIavSH3t/4NUVsHa/jClxAz4e4uV5KRCFGJgK5tzGhBDZv5kBOZ
/+BD15KNbZJVCMBKZk4FmIWTExK8qbQktoowRAleIFbhcfXlLhd4QustoUclOTxI
5A6yclbvvW1kM/aeqMKzNoDLITyu9/mlkZaSZpxV+h5/+sZC7zV7ouOgrDkJhFr7
I5ao2CVK4yJG09yCLW16Gi5ievfERQnlulUTeLTSMdbBFxnhxg81ztR5/HeJNXvZ
2MAT/pDXhdfxqMRK94whwCD2IFNo5+emGLvR1JScVoIBulD0vQP8Cus1rQRmJ+x0
bzkwv539O56J+01LQEFQ8sxkcAj8vS3jhVj0V7W+WcsEACQBEtnWpSgB3Law9mlg
z3OZJwdgaaERTQu9OmpISYsFSZmz8MIajoBeZM2aJ7ES7Y3PynVRKA7h76AR4G8T
BNe+rOoOzEOF8AMczQRo6iE0IMGmYCGChxmsEsfXMg7Y4nHOm5sJo7tMsToxRlAe
N8eAqAEeDkwn/h8kl4nSwi14NGFX96940SEqXyOXia6zSIGUmqn0cZqObT3ql1Rn
5YEbyW/2t6PcFkJBXVZJOsg3jRUt+YIrW4lLW3o+3kjcI1aVLGKHXWLR2olhK3SP
zZbRl4g+LmXTxTkk/DbsbQ==
`protect END_PROTECTED
