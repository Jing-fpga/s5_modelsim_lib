`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rL8E/0VQSFYFdgnzXOOamHeOHMwFVBDNCh5ahch4fqQaAXDSC3rNDNIuuI9YRZuS
2WhCCoNNBuDxFmdhgi1yUJr4yjddBP2M2uiaY+2/vJbc5cxb9yzl3R6TrHtF6SpO
jHKP/dLdtRYMxi54a7h0SStzsjy6h0fUKPsgK5NIdIrTTUOmHL1rt6pz84QAHaL2
Bpfn8EQtwuIpL2OwG1fmFgoaZSxlVOeR0i/a0kOEdrJBN+FISYwhA42SO9fvCV7d
iT+NqLcu5qUW7EHPGYwX1odzaxjxdKXHuUJuTTFqgwMqmxJHQOitCtUu/uXRHOgd
FZxZW9u3joJ4HKEqI6prS9rQktz09FCEM3tJ5jW1fAhsnqTVamxxkhHN99+1yHEf
y0u+c17OdE2fJm81vTWV7G4b1vDfz/GLAdjacsFyMoWu67WkgfbUPAYnOEu7Kn9z
TKBFonGZyzsF5OzR7WVAZXy190d19+OgUrqIGviJsNKhm0RJIHfnmSpLRU3HNrJm
dpncItXr0DizGEca0MrRgWgBi0ZcngILuykagmLSUwgidyiTOJcuipEBRnGdaowZ
pYWGOsuC8og+PPWBLES8bgkSgIItlnVahN7gnaw5XqtJQXy4l8gkRsW214f3zPct
kZMIwMIw2t9ZQ5BdceK7lthOJwsCCubBOFd19/R2tO23g/aHFp9JHGJph4zCuh5X
9xGC80g3M+ozpoWYuXB+1PLW4EKJwQbaOfcTJGWqFTgnqC8JqteziKDQlWOS5ifQ
VNFwSkkYJYDJbzskQ/Oe+OhqoFBukn8EdJInNgk92tI=
`protect END_PROTECTED
