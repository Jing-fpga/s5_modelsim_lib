`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4OsKf5SNnyzYJX02mX0zXGu4Cy5Ayfwwgo7lSVOkQwx5J6loDeRa80rnjlaYm3li
8HIZ7eHxdQEQjdm+qnsgxX4zWycBCemOcE+sYeG5drcWfWTlU1in3gZEpSqW3mwU
PkQHsHMMMmTH5wb8iA4Ba5K6oD/87ApeFYbTKjqm+RBCze8SrottIZEE2Yi9Nl6p
YXaIaDHCiZ5b2CVKFpfPaxGM+Q170SKbvH1PhPSzlLDLpNY+3dzZhQ7+nu+/FYdl
nMlRkP7ZezCXWNlvLTCrGHNKqJU9pk8lrNBT7kk1qJO7+9Z6f8VLVWjara5UzImU
rskbdIfQu08z6Onx0Be0VI109wP/PAtvuA5T08ggoj7Ed79Rk3B4OhjjC+r4hgI/
zPIWMHWgI/ZcLDcwmTChVGBw/N8hye2N57eNWY6+IXxl9+4eeiOch58XhPG2EacP
k+xFPYHyfZ3Bp8pJ4ueUKJJfymAeNfZa1bcuoV2z4VGN9xJCLczAYAtUP84N64o4
xILEmcEiH/i/Ci7sBYZZHObnm0dJk0Vi2BeqdCWHRG4fs4oHE3Rh11EfudMG3s6+
M22qG2u7/pauPR8iJiglh5zY2ze+qNbm1mVH/Puh4Y+/J4RrotDMKWjS8L5P3WOw
TWY627fw6eUj4GzpPj8XoCCkTWv1TcRnjvvaFM+3rf0=
`protect END_PROTECTED
