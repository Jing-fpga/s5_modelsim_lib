`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U8+0OkhcexXq1L36g5hdF05DsuVnh52K8pPMsPw6g9WYlvNyfCiChBslVlxWf72C
TkJrnmplgTy8PguW2wrPQ1m2lUSNtppOpUx8d/WzTDADqb+S8kmSz3GpLFgzxyOn
byt8yVaudX+V3XfZ5ZQmD5LOViRwP7xndnT3gp67H9PvhytZrCQa4WdyubMaTOaW
NSf+3XbolSu/9x6Y5gOQCGetaPw3HqtYWLIq1teqZMznk42p9YlFiMImGF2VaAC3
87TfDPh84Xyiv5ztboHXlrQubpKcHiLVWDspQQtlLWjKNB9xTkjKE3PqNCAeUqlr
aWc9aFwBOImNxTtYGYftKMGCs+1htHjuv9mazfbrQlbceOy60Fd1mkIc0j4dgLvI
8DuD/nKloGR9k7tGOKUs14j3sQzTBxH6SsEcr+PZEUd/jH9IoE4yLXk2ge093krS
apt9uySsNFQsV8ByqhXAOrcgHKV9jU/lXEP4gV7J2l8OXe4BttV+2WfoU7izHCRm
LBN2o+3hWt/qAL120lrbdtgwDpHRDK2Xxv20uB6IbnDOuA9Z1l14EZjjYr/xS2nP
ZLk/MzWYvNzEGFgi6T/xAa+ts/l2XDQF3gD/Ke/DV71FlE8CCyNn6RNC4HhMTuOv
HDwRiQ7xvdTAaHayRSNFSoZbfwMBJKdiQA0DpYTQ03WskyZlDC6FFpnLQSFJvcBR
o46bJwn5720M+pBUbU2eKIHIHJbeQNG1WHA7nhNIWpeUYpFimgBYAV4e7pipsNf5
o0PorBPckOovj6+BvvyFbcZsZfpbQIVTVZO0VZfD1idk+9nJxWzEsYzXZUiHu3mO
IxqLhrk2wdmPFB2DhL7r4h632IEFaEeItGplrE3bVsGaArn3R341FZRCXF3KKYh8
Lp+TFEbJMEN3YAEW+uHgQI3lUt36QFlxqMl75UdSN5h2jNWK38Fsq5AGtt+ymp5c
f6sBfL8hOQpjY1AhHEj0GWHe+Jj56NGq3j4AGRARY7+9Gv6EMExPlt2puirpNr22
0dJWrOXQczxrGjF1D4ho49BEPYp34Rd8Ktn1XNWnXzGvV3vbPkVFZZ7JYT34RzEc
BQUp+pyC4nzIG/NFDhPRMbbHX01SinddOCg7IJhJt+HHjdhWYUpeJ4LDskLy1qQV
1rtoKZTESS0w3GpDyfcW4mHGVq7uplNDultQn8Ikz8yYW4ElPyYG6be7sAeA0kQ6
7n1c1g2OStR4eOXaI35+bhv8LmEtBEXhIhPql+07952T768aRBnOX8ZOe5+L3fST
loQJ4Hbu42x1juQOmsgggK3TEUhjPKSyjVckwityeC6RPyyY83y6I1zSIzRakp1K
+dYNSE/nCOx5pTnKiz0TgKWeokoeOku7fZUwA5y7ikcnTcA1Qsuu/eeI7a8dqnIw
ICEzy8I+NyV8Yyq+hsixOor9Dg6D4u/mmfi7GHES43Y95VqiMlmgD+LZCkaAtjDV
7y/ZVFO7lsOgFaoPUd9fOg9YIKfql2vkH3XcrTmv+8deqpncvCZgcUQWI1k9qsrm
zjJhbIrSk5ujbUCCrNElhtVfZBSgn91cAubKbQgtP1E5KPkT941BkzVOdk2roGqF
LwJYoSiF5Si10Y14vWR1xQ6yta6EZdEtU81KzOyLgQV7oYDtYZDUvcd3Bg5sQSyc
cxfvmY5SVWhJ2o/u7gL/S2flKe/9wROop+NxB20Pt+qmxekDCTFo9Q5AyU0dhLIG
RCJhqWla//Ewuf8at6L6fRzd5rkrLmPTNx+xygyPAh7vPp5Cxo4EllO8jT+1FfwO
5MUePwyMrw4A/jWNxhn3f06QQ9goTqbEbGWXIt+TcfP7e3iLLkN/xPhyV28aCCKU
8srfrQGXBYPV2F6UE+ZtG75G2rpB1z7NOqt78K1JyxDl6Vt6UTe/ZnzzsV91bsri
YDk50w9U4vWlkkK2YzIG+aZtf4/LvwQUBQNlCi80aq8uKDMPAliAiiMln8ekRtKA
AC+YLS9umfX0E981VstOFnPXb7rkgLupgVopoHSck0ivj7ZsKn47HiosFDZHXva0
58JjACpROCshlFCBgbjnR3iGubapPHabLtwwaf6OyySTOz4cDmKg9qNSuOpm0FbK
/Uga6lFi8P4zHE/Ez6zgs223BgGTdC6G30RT3iCWoyS7ifwG8TSgUrm9uvV+rXcP
7gEqpbXO8iUXYUe9VpTqqjPTmFxG/hgcJWgNWQfSzbPCcdYSMztIa6bVzvut/ICH
pkY7CZrMfgk5TIibnFxVBCiWmYE0YbkQ62mzp+AsOImpvg0YN4B55vqoPQwBN0Hz
vcL/q1JFyk+ov2k44LuqpjjKodYmrs0XbVrXHKeRq6lG+QML8bSUMAiSwUAGhmo1
zbPne4B99vYdSmFINYPzAQ9S9EFc2JtdLR69nQntZtJN/UwnFfFsPSMg3zlCw2Mv
EVGRjk4qovoLxxeMb7dFLLJrLHvhy+1mL8yLzs1cVPVTBs9xu4QT2KOIMLILPu+T
VCEbtKpnz+n52/Knda8E7zXJimNRe+6ennS4aiJCyxT8iXtRJTSJ2p1i2He9GllS
tOfazHBCM5Mh0/l3+4wlm+Ut5phAuoSpUR3DV3hwb6VQRMIyY1eczCZQoXNkmnuM
rVVV/OSV2UgGNXEVx+sJ7RDxxEARwKwyjZk/qPQgGoj755T1hVGLyQq9YPWXPSA/
ZFsUwRdbSmxaUy1f9aKPvETD5+kSNPurTe+CxHsprcx/akWaxL5BCFM854n1AqvO
n5CBy8Fv1cJz7TSmVXU+plnTVby4uTxuCtCfUtnSEpKIes0EvmQZl1qOZiW55hUv
+wYOUmEapWzgZ8E6RXYXZVMRe5ntz8yOvq67X6cue1inhX1BYX2VA4QsIkB5N3cC
i5Bxzqcj8xXkUAzZl7GkTs8o1ng1VdnVam6cwmfb1yt6PJxeWA9V9X/GUGxNFkzJ
7LAovNDEIF0IpwghARSDN/lOddrrM8lh7ESJqgers7EIWtIU25Y+BmYjPRAVb8DR
rk2ECcCMCInLPPo/XUPjo/EzUhoLAN/YWSGSfW0A3kjrgB7gVbM0lAishvY2nFaw
tMGSksd0AqDoTkdXBPwsERrwyChDt6yklquQjPEnDBa05bK4mWCVnCh+PQXE6Gro
B1B0srSblezJNJyh/mdjjEVPn5E8iUy8yWg+HalYvehfhZhI5tQNYY/rXtRFqfN4
QKc4qtdu/veXNxYMGHfjtuhoyP1c6LzwT4ioBi2cVfOUB6U5byH7k0NDriSTetQM
cxLk5gr6Yw2D3zz6jobVDld0etjqaSsTrWajpHshz5in0+3C87+zMmHyLE7fMZ2j
qlZOV+CS/v93pKFGVF8cXEOljHI0juJt8sUfBRT5zOOwU+e5YUjZyJTJstsyc7Uw
OiAsbuV8WXeQqJ1Pm4NAAFGPTaJYOxX5soTsWRaYcViN33MU+k5Dzp4tV0xNt7wt
KTUa4Gs/la4iihmkJK6ovqgu+nPjf5jMJWlRA6Ww/fyIDtRE27kE5WCi+p36KFgZ
eICevFnhlUX1DzvutOWVCYWYg2JVFlCwWnhfk4rjvGmL9EIDz96rJI7QGBqSRmNe
WtnVLVHfMojziMxYDoFFXne0mdpFbPDJRAgQh9X61R3WvvyZVfwA+x03dUnyWKZ0
zBlVvk0BXaOmCOJS+g4sVHTGSzogpJST6aLBGYSiANRJqfMhpNma1C86aSCAEfCc
o1RCbv5hHgmRri90sTlA/LJHhYy9/5HzHOXy9c9KOg2j5wVZVo77Sa9cW1OhyR1A
hYMnDEdUEGddf5waea5JgX+jpyUO8zl28wmYpuUhXJBLOQU1Rd53AFKrK3F6Hofo
f/jVn4HUGY1HcUow/bzSc0QgW2N1R+jG3DgvEtKlGXQYfHUFNxX2P+PKu9cyh69Q
6HT9lE3J0wfpd906vcOKCqobMFuBvnsNouXHiR0u5LFnsGTWSccZLO2BDh/PayFr
5Nubk/j4JKVBKigxAYWtBy7V3WaIm9FE5SaRHQd386zwL4afi5hxQUfZsgJzVZ+p
R4Wbo26bhNSW2a+oJRHCCAnPviFPa/REs7HXQw79aMktFDsFeGrnBnZJ1haQ26C4
RTJZCQ7IqiB57ve9bv9uJ8m66QpQdQmH8cEU2lep4YLxGTJRpisCEJ7kk4x+oND5
`protect END_PROTECTED
