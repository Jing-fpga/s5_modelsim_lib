`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CdnF+f0TgEUmBtv/jbTe3IEmoNPW17gPj7U8CPf+oteBl0W+W0M9RPGBYYFNsySF
tG/Djq/kU3210INJGW720UDuotaFsh+U4DzHxXWiVbj4uYWxCyIWg8yJCudnlE0A
2rJQ4uZPydhJ7+jtUCJxqGrdtau7gvwGfhNoLmK1NU5r0jh77Je8CKmd8EaYz+9a
0/VmUVxA2531uTRSfQnzpOMSWUNw0MnfKCIiH6N8vSsT2Tyzz4nyiVH0tK1J6r0Y
v38K987g2bpZE6/OovBMz8+y+PCGnsYbRj1iH1ll4DcdnwVqZ04jNFsCM9dDIpdv
rWlW8nNJkBor9d752ffGVFdetOmmlxFgrDkexEpcCjTz7YHblQ9WH1bQ3KfGsPA2
KciOTlbXEJo4dBDGuIBXkMNDvdFNh44rZWBO3wShs/XObKGYPb1bMw3+xg86dcih
aVohENqMupCPxcnZfm9a1VQFGW2Ba/vGlT0Cn2/2eMj4ocFuw1h8ykZL3nJfQ+ou
egd3NvpzRPdB0hZmthWQcyaltPT1BYMe5Zyh1+osB+iSLB/kTfafa5Mx3Vx2uozG
5C2xOjrOK7OltDcT+CK6HvNgaLBEj9tgSkki1ErMMLq2Lo+B80fuf6okd3yyioon
nH2xFJIqv/I7YdhbDPSQPVMlAAlkWpyO+FS7oK4kJhEy5p33vmf8NF1SI5Tfj7fq
xM9hhQ2+uRCE+vPOvBSY716/v0DrDHS5FsQ879nu+35YJ0tfLnZhKwxfuZhZ++ky
sDxRYQWguBYjs3Cn14zUuiGsQ+YIgaqrXTom6iDbLplvZ8asQstSoHx18BdrVBSS
K8L9aglW7UP5kLLrFyszwbJPO28gnvS2e+j6dq0eW4hypOMIst5TK9GGtTBdgoVG
zf/2tk9dFD2R5fwmyR+ObamvVxPc3X5zy7RkWYdgfoyoSCSfRUv90o7eii/tKNhp
ZZIJDabGfq3GIn6gyt1QXM4Py+/f4muSfDm/ctsYMZjL6WJSJhQ3qA8VtczkCniG
lghzWxDYxQWMdvqaKx8WQRS4xXZuJN+MQqhyG74pWoguHdoAluKByhXWEqWtRMoQ
xO4hOJYH4o8KUSBnnFUU5m7k436aWFOcASM48wXmaQcUixH03hzSEeBCySFDOUgH
hgN0YBOO+JWWKzWYUAMY5Vv8HA4zRnzJ0aavnQvd+UQH5yHpMr+fCF2UbpqnaTys
IlqsbNjjO9ogZuYRoby5eQ2Skey7E1K9cC5gPmwPJ2cACH9kcCkyN0kRmMTmx8iQ
0vq4iedmzH+njvmzodOXDS/0Xp+W/ecp/MNMBHxA7xVYVzYAgJDbjfPodXjdEJbO
hGRilvZkE1pxmz9io6mJyYptZgJzLNvgqtujnQhfQG84toU2b0r8Zl3iBMf6sFgq
yRdZdJj/grHZ4gLdrjofpyQKq8lV2GPxvVtqbtu3tzBSJaPS7xZWHIsimQvQAQkO
`protect END_PROTECTED
