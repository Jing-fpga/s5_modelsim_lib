`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uRtMfNzwJhU5H0sNdNHHCkehqSKxMg87R7+0JGXJNtIYEMGAshE8F9U/11ZU0gfz
qPCnmcBr5DdrL/vU9wg8A9vSKzj8tZIk+M/krgbCtou108reZKEqJHXE/rqw0nsn
9ADCDF/wDJIs5LmEHnR9Vk/TrHqPe8QmX6mEa5hV+/viBh6tfBsQ/M2CH2nxdRAr
dm33h/wCqVxJhq8hXNEE8BQxQmAq4sL7hLDE0Pg1Ao7ff97hwmyG1m3MUx5pDi3f
9iRI0h3OJRHeqM6UqkgtVYDH8bl5F6hrXuLnR8T5FDLSIVi/iroSSqeu0NCZPRvE
g2ECuT67jCYoe7O+fx2j1xF3F/utffW+6eiEKSXnj+dp9ZXhfqV4HZPAkTEBx7Bb
f6Nwk4pmEtnLrVSJ8kr3elXlPvUxXplFWAiBc8dCkvJRMAx0z0RR5VJvbBD6XTQo
J0EkLLOnNrXYgok8gc+swh4XcKLysYuyODEmDPvQRdtskjEVzwfT4+mIQTmSmDHi
9lYTVw21m/7spV16gQY7XTm2SXt2IujcfteMqONDiYtUfR+rduFhnRs7KUv9Z1eP
S9iG4xOunzCUMbBeZl8z98G73mC6Oxqcp9uUBSEtJTWV4onelbR2Mx/3d2ouvBXt
4A0tjraOIYw2DXQhCPNk7FwVUQzjbFtBr0p8uSQl4+UNAlYHJzUPxmJUBf9pFrM/
yHqtlTu1AH30lGmEOgmUgBN0XnrtOuIEPNUseKgdYPJTl8Mh5g8Ou0oVBN6uZ8tn
Hy72J8HhTNO27ntt12m82v8VZzW2l1djhsO9+tzsGRp5m7c3sqs9B7cakq8mNzj1
Sh6r4GY3Sxi+ULUfX+p55CkhZcvxACyZOBAfRA+nOxMRcGWgFaE2TUGKpKtRCeNd
QCgsNanHhj1gomuT0tYfYf0BNC2Sks6YrGuCAxa0l5lTrj0t6WISdVnQI/AG/t4c
fYjK5eGW7HUkNhTLx/6l/Cu9IKpuXkJCEG8ibuKkHXBWXHPwBNktTKkIsKEB+JrX
nygThbNr8YabXSWirJ0cgzCC/ictZDAkRRyf3bhGdCY/sY+OC73lsu27lWz24MvL
P+dpLyiz1W+rFbv6ODu1ckIpj3cchAZHbi/CqYXR/O+/Zo09EwHSfCDW49VwlGXj
2U0FwK6cXOmvhvSzwFwF7UivwsSxtLLzXmIvQhUaAkY0kEbjOnbp6yWC4o6a97eJ
EynkEMqj90qqSQkFJ8TqjGJWwrxwz3iOi/Xtf7YLEMSM4tquxllkLIru1+P2b7PO
oFH/LEQDVykEeRfuVJ5KafffDsbWtINWRg8MIvxYmiwZKRHcF7WJEIJ/d5P220Lv
l30DQcU2C3xCY66O3ujifZ9LQKOyLAZTgGr0M379Zjiv/Q7pTyGEElGTkfFr9iZe
mg1R8Z7Ev1dJFbsY6p4hIPUsi5lXAfUB9pk1hoI/9bwU2fNtRyRs4ZGPvLcRPeqk
zPr5ntSQ41F2azzB1JkkclEw2TAwxP9x8qECrPb/f6yJuyS55yzioLSay4MdZbFg
cj/AQmNfQwFANDeYIcUYbJ3ZQPbX6kSwrmIBycvNLAD73PBqFI3M1+nk1nHou2+/
5Hm1fqF7IyvG2bGkHNtgAE/1ccEaw1qBbcxVEwc/8L//W5lv+gsZwMA4K/CXWQZS
4xCBrqez/TwVyhT8CNC3/6yB9EZrBm2yXaC/7D6DnQhb1SlCrMVaw3oWc4H1Is3y
GFyGYnpoKGGnxKGhzKjlzY9zY4Lx6nbSBZohx95EtLw5bffBRLvK5uGwppcfhDNp
1qIO46qHi6k0Kwuqq76nlDxliMMKihnO8bIl536AUC2Pf3hMthZiJojilD9ZktYJ
glqMn0P+LlBXeWKDuRxWsGG4jDtQms16pUhAG2PZ6NZ/8UhYPbvqYbZs7EXxRyXc
z+RJ0i0lOf2OzK1WFA2V1DWTUA6ZysZy2zVzaoAbB56W7ZUT9G3RnZIfUQ+Ccjb9
YaglcDIN7AP3QYKW06zIae/XghSdYs9tXyTNhNadiDUG0QrB4lUjAGWDcRTPEcG4
hCLmEBSa5z1NHkFR+0iOszlZET99JxYmY7ebn+gjTK03/0ak430Grahb0LDxkD9o
jq2vi0LocVn2JHNSuTxBscEbqyMIKIQj1uvOH+f5oMX0/T2V3KpOw6Yyf9vvEeBs
MrATF0DfFmLOxcI+PyuqiifGChhJSOeAVw5YPSIapglN6puV/UBEJTqeyd55Vgm8
TvXCNzyVwvD2JKrl99siMNTC3yTMivQx18icWv8KQhSqOqFux4KMUfYtKKfZOlrS
z4nJZhiWTzhV/AdPS22bHM+YBhB29nbQ3G2jp5qrD+yYjSZEI1ZIG9dEyg6ua1+Z
CYvHcxQCbcZ+W449UmpkUW4OQPErb0kHqOoOy9aS1v2CSWyKZTEHgHqGjwGBZ48y
/NVtpTXsq1PddQeiKSXBwQ==
`protect END_PROTECTED
