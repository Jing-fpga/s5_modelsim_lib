`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qGGl4IPoo3REXy1r06ByEdPahX0MJEdD5/E7JwDMjYEP9S6AoWgCOCG+lEGQ8FiW
qK9T2MvB2chPatWREOoz963MMCgS0hG1rIAqVFyhAJsAhE3btvU/JNd3D+Xf25TG
W/zv0XaWwlvbaDG9YVtiiape/eObWnSYOeMMfLwtOPtJhWLdj2U1P/XzvJjOLZpZ
UEPqLFi9z/ZLKhOI263zFbP4HMbQGL6QmjL6WvpSuGKnzcajsL9f3jREOrOI8ZL2
mgv1bsJndUjcKpwGn/cd8uUWUMeJ8gaPu9s+PrylcekZDbM6NlNkCDpkZxnUk6Zt
GR9enpzDxogBdaxS6/aaU/AYeuSSHFg5eOc/WjkHC9oxlp8vyzV5s61qNBcelKrv
d3MP4oxZoHarVeXejd8pBqTEOhOHuTNaHDS0Hh/axqNM9pWBMis5HQxviU93WUAH
QIEDBIpDuYpcWK7gPEB3CGmWFKealVmIvCZbPVK7GUhDhxswWmP1a9v1ZvmrwtFT
+AmBDLi+/giahVTn2zaSfUq7GpmqQprITI20iRPyOly8p0omH/OOPyp+Sxo6dEJK
zuJ05LNXFFOY3CbUSGxxWwVpIchgTBjiCklMOn58U9ZOeVqGQKKnoMRGFiz+kvyW
`protect END_PROTECTED
