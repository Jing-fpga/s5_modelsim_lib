`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8n6E5TuifsbV7JCeLNHrtA16ACTBwBwll51orLCAT5jwD16JNQTfb3mQKkxGldz3
JTFO0DlRjb+6IjN095GYEdZAiEImQC12XAII1oEO700fvCWlxC2kRvJVLuNW5/7K
dSaaQCcyq6FmpjDnOtravfGvAUUVyFn5E7NjxQSPI/dGIyNEpAuYipU/M3/jw2EL
DYdmbHSo5JfQQIVHI8tuOVev3QSIqsmkZoII5VjHyFRwdXA48rk+Wh/4j1pfpkUO
SQ+acwpx5exwXRR6glSH1d3m0GhFuLZ7UuoTDs/bBWR3U06WD3wbl3D2tgST+B6v
Pu/ShUuyuzobuQFsgc3S1FxD8PsEqbALpU/HF/+GyC/i/lfhlHgO0zO5xIe8TNWc
n57YuV+1CsyR6ZJPIRGRUYMDyBo2aVPT6QERYRdl6QOZbN0/jQ3BrKaUNNnlHMRd
rAr6T6T2NMI/dTNb9NJahaeqgDamNOto3yRmofvJ3im40i7fM6PVxJYKiCo6f8nL
C/VJIg/fGCCAX1c1FvJZK8/YiLphWkHtAWRBtnaj4OdS+uifXtBedsLrDF/UjhPs
4T6IE0g62fjr1mrLw7D69i8rTfOJdZm5CtfyrCiuz6pBwkg9YiYOLe5Pnc05DwsN
AGlO4o++UXlfL6JnIMR9sZbHCN6/GH64OR431m9mDB4epz72VKMCwQP0+3DbY/My
kbhTuRkDukqVu/SRMZNocfAik9E86m/tr3Qw0UN+ONrdC4wbExPJBbmkp5Wq0FXf
j2Qo68fsCcpIqAa/0EmPSpFljQMC2eKmq0wRr1ZfniGpZ9zKoHNtpRdReLWr2f9E
dCRZi3JiDz3Z1czdM6fxAQPVeSyZAFupSEeomaL5MwxVjN1XusNrUx4wBC/6WfW5
g0SvJaYTB8fVJdjUR4w5Ng0xc/haAWNbUB9Ht6g7ZguS4Awgtsq6EqX5McmVO2Hw
DymGqR6t0tcEarN3yobpecfCC5ElzyZnGzibz8xfl0jeZlSrGdadC6qWZSlUPnT7
uwQ44mSwRAR3yrGe8XTyqbi8G0bJx0cmxW1c401gF1xpviOnM+2ic2yOg9YK4Joy
xAP790cQEYbRpRd3zxa5qySx0fCjKvwxaUN7EnX1TMNrGCptfxJzPIhIOiWWN55E
evMKE/S76Z3U3CGDGB7EAdAQfB1XB/dMv/sr4zdZUG0GUReVt7EZDF+a+/0s7y6k
gtPJlVOq4896QazEnumdsNcWKP6bJTgIMK+Sn0bzMxToUXAWngU9aZaE0zdaPd8B
3OV2wrikbJyybZU9TEbHr5ML6uMiT6krdQ4gpGKHueU6Dd/0uVA56TIN1BbP/J1b
rcHzkdVEj2ijKlHCyRIxGDWPq5udh21UlVOgHr+fC6w49aisUZS54UUTGXrGfnev
rtlDwpNJ5SS8oepEHT1UhbQFn0+wVBIaasl9N8YcCODXezHq9a9u8yGRfx72I/id
02/wY0gQkrEXgAyAp6Kgz14VVcgse2KX6pFdBLTt3Qm6zCASDB9ZucXGFyrapa74
SQ+lDd0Eusbqlb0eRRou8+hwAnyHaEcyFd+YIruuutAcSFs7urU6xd7qDSRUA3VP
zZ6KtUR/h5BBekFkrWUTeyZ3vBDxys2uh39N9YrgS0DtxsKrRtmpNk4ZV01HOQqJ
YQyiEKoR+y9jbPRniNpDZCyQl7FhYvs2krTMgu03ZXami3Rx0aTILYx+vLV7zz18
FjeXCcZ0hxXngu0jcAep/OVcrQgqJnn466eKXP4GspVWtwUcJy6hbhEbi2oY5fby
1fpU/5c33xT55WineefYFeMGmJlsGJ03PeFe82+OROhzqMVkAbhUY1v/OJsQ7DV8
MVznslT32kKa1OYFnrGOsmQLaNODF8+hLQ1VdAcmj9SIDAx5LBu2qRFDJEWM6zGy
IHvswz2GHU+oAGKwYWChK85n5xQbDE/DvsrR3TqR16fYkH0Dahs8MsE9c7+jhW2y
OwSUK/Hw7wRpLQKoDAAVx4RAAGqRmLJ/A3eu1WKDyA1VXjv1oewGXpsWK0xt27Nu
YkM/6h4ar4Uj9BFbK9ne948LsSm83z2IIyQWmvvG482BxCGX5g0968GRoN5elV/n
7CVCCZNRgBJvh1aHrOJor0837jXAXWk6h9BWkVZq79Hl1MkOriBexzZMDgagpwAd
wKzk4q5IENvAXeotXc12rCmgCOsbt+EgdG9UfmTwUeTy7Q/ZJ54O+ugAERv3HFOi
XqM5Z9qCo6wURjzMKu+zs21SbzoSABIQAdnpFz1hUuJPBsmY0R6SMgbpIbDW85Bz
g9h96RjptEH43nrYxQ9ohl4W51pjPgsoUB4ecxsJiwuPV5+vQ5Hz2YIyI5s0iPxq
IUbeahkgdnZyRRcxuEqyCu4QGPgsyLCpmQLDM6Vu9LhIL9v7dF5sZrQBGA6MT76w
oHiLcdcS/+78e1grkly8NXhQp99VUBDgchIj6Omn2KzfEgQZFdsNDtmS6bBVjhGe
QUr6lvloD2zQbmNGS9dL2j8x1d+LuSnFVep46Qw/UDN5dK4L+FMmPjRiHSwhxinO
gotTLhSx0ha+LXQiqKCMhSHS7nPAXrwVXjyr+x67+xO2NmU5ycFXujgp2y9sZQXZ
pSWjPQaVGm1RwtuIvDrm4Ig8Z3wOY7I8dO76igEKYps9qM/oJNFGjsLqv84WO317
jiyDJ6l5gix9v/XzgIMQOpJBJ2fQDBWoCmxcyIYRiDavfbgdTERvocbBcXD+/zDB
m9Eyd1Gi1rm3Wrv7y7ULtnL9AlUN0Xb24onJ2C93IROViox2WnAMPRxe4e9C3PLM
XyfmTUmw1LvaQzK4qE8iiu6cX6UW0j/F/PZ5UeP5loQTIC2t1q9wfN7GL7ViOppK
IiQYBZ/nNun7+/zRXS2WoD97BJDycnF/IJuL5QblYTjA1dFFX2dPor620m1bSt3p
zBtk/aYw6+Y4fQNTNM3/Q4DLN0Ao9rIJG7n96XwcUX9Rk/jQ/NFDqWnuz9+5HJoi
/EYeDYAkFFC2edhtVV3uX1j1RnllJzDBZK7m1dT8tZmLvfxKtLR1iIs2tEhqMSg8
BvnXbmcPCIB+SYBB/BvddvmmUgQGc5tL8q+Ew/bX7MjXi9dSEiZ8KHq94ALFyDQ+
DtTQX5Aq2FIy0mux9VXtbn4bLOoedYWyfpgs4fOhDBDOOcC0Ao2H3BBHLI8v5ji1
Uv4N0Wtt1WzqD6TpwbRW6e9C6HQUY6iTJbWaTd4kJyvG/eQIeX5rNsC5GanA564+
XqtYupTy2248pmxiic/3/SFVs/icuZbFvRFVVudNZ9vuau3RDC9k/V7ehHH14aa0
Z2P85q+BjUE8JebXfmJgof5Qh7Zf3qseoYJKNlnGezich7kzRMgXzHSEKF5NTTA7
OjK2vaT9JqYKRDE8hDfeND/HWg9M3SQG/hPjlr683rRaySo7nMmsdWYzyhTd28oh
iysfmBa+fy/Lcv4/vAyhBYq3A6fLG8ukJLgdikfUKymrkbyM8bm7K9S+zc2FvNu5
BcqPzr+qZmk/oC7EFUkURLSr9Mp0zPocdwY//HmKo7UgjhHj/jHxEnj1nL3fihtR
WZ9GhkkQTkbIQENZDIueZMt8e+LC06FmTBc4p+ozcKNYZTcabPPLkh/M7f8GZn2X
ueTk0oRwNBP9pjDZquSBZKLHhGC1MN1TVrmpUhcpZjXWfWEl5kT/0O+73lnuPsxq
J9q5NfwplksBKGCy5R2QVFvLHEGuTb+jeKNhpt0VwNZXZN+WcOAiuF8eklfXwXri
179UhZ1QEb0PYSoSLa1KFCXxrw6L8+y70wvaiwxC+wycdk3ruy1rHYXX+wC3kL4c
QSgsbUnwhBq7a195hKYUZr8STfOS1NYlZ8Y2B7w3js3q+UAyiqU86T+VCHhFwjjT
Au7kCoOGqw/Z4xmCHdYR+6jwx3yS5JQm406ezJdLoiE8Gz2X0x37agg451JjceB0
z64GyAm6dGzmBS8ELyjuwLmphzj1BaEdzvhwBLTnf/WR41soX36qYbj/QE6hkXOo
DrdJzIudTX2frMAHmr+9yR7Cw+i4n9QnVT2MJYaC+x0zPA1PkqKLunJQ0wW6vwm2
qoAtdSE8W6KbEJ4D1TBUZE0bdpWquNnrnFm4ggyGdVuDJs/nzdV62V5ZhaWTKg8P
3402Jyztj/3EQtdARTr5/v30+quhdpMJQzfrnUo7p9DxiDl8NG2TpXJ5z8WQp2Rs
fj1c57MsiZuCuDPm3HcXJBEvV0ppr2xbrsxvWUmOysJ9ctoCGC6r30IV9eSSoosE
+Al6sBmpGMmUCBYSOmG2gzC5EpSsNzhKh+TICYl/EmlreXYWpXmXVGw3y5sZlXOH
yBikAPuo2sR1Nq6z+QWKmk+NvhPvhkgzU6hEIsozylWJpMmuMxSbbgAUO7h93KoK
wGmp7C2OVj6WzXDr1Qq0YIKdp4NmoBOMPWzrVQrrtiawR9ktO3zC5Gato8okpUz9
sw7a9SshsRV5yaiIXMVzd+qAAv/pfy3NFfWbiDludP1CwRoCif9ZvJkf1X8HIlFf
8TqJsqSE1ydWP6PYkMA5sVpPx3DS6Cw9QnLJf6u78mL5qu2+2M4MZIahfzPkGucj
jg3mXRGngxbnoC1MQ5wb7AVxq4bartleokNw/YNtF7ygeR/XVcSnEjtmAdhzQB/g
Sm6va9Y2g9imdfwbqMVg9vVcDHt7qL9LR0bRIM1lH2/cBGY6q217Uqf90CjpWxbZ
CCzXswnFOwSY4bgaQDsl27vWkDPZlQt7Nfwib2y/9BqhLkwMk15yvluJI/bUHi3G
KtaiBS3Fs8774IFuvtQuP4ld5tqr6rt2SXY0A4VElHW/cUA/rmEJR51bH7z0GnDU
xtBGwBPNgiDZ0q35OE7EDzKhrpwFGWNn0ST8YbOawr9qzOhpclhfidjk/JJZTvBd
En1ni0UbYjLTsNk0lHN7hvdLgQObql1QAGu4fr8IdvKHfK+33P9x+2K/X49Hf3FM
RyDrCNGxMmvgD4K2F4aZo6/YpBYWaDkZBg6NzB/xSNRgdiq13qIYRMcaOaRcZ3YB
txUL4hLC3dqXOqb7vK2Yc5qEgIVRe0zbqQ48XmFAwhHJGmMqBI3JmQJq/ISSKKZy
cq1d1gi5w2zOhVzOJlJ7QlKHgB011jZbiCz9Hx/Ec29FLNYVnL97huWnwS7vY7Wr
ldJ9KoHa3Ro72d+GpnQZr/MpfCVjixEC0UE+espd3nBxIenAowSVqRBSLv72lqHy
7o8OUjF0RMBq/EqYaif7AtlySFKiXVh24OnV773105Hz8HhZztjqBH/XC9MmWkt1
MdcYo20cVIvoEZRn37EBK/eHz1oubLYyjq/n1ulGlFAgoI0Wr9knqzOMgKO9EODl
OO7itsJEpln4uhr+GRD+72xgr2cmkA4umuQYU4ln47lUn5g0Xc2gKP+U3TfIWtfV
eHkCAj1w0Ww4HgqIw95HFBR5jS/JTQRdo+XxZWrBNeyGh058w8lSLVlGnO2QJWGn
bsu5I7NY/cDfF2Q1VEGQLG9wjbXdbtNXwTtPV8MW5pSKgTvCsM6YPsuWhDb7KBLl
CFMsfaDcy3vNsIWFagJ/I/HZL4fdD92u32ST1fYysjkQleF5arMAvVVWrvYzu/C7
BNSIQ9CBtjr6YdZ2XrY/qTwG9lKJHfRVcETT+ilVUTzagE/JTJm2ySdpggIvVAyN
EmbwjI3R/ORbdTc2evXR8kX1RbVsCVKWtueSY1RndXTJyeW9lZHBEuOwUiAhiVVz
r62pRgAdTNHPBnfcahYYf2VKL4QdgptDVTGLmXkzR2yzO2H+FSOzBc2XFLSAC0QK
B9OIwNCPpOFk5wD7imMFEvsIB+LsAqN3qRJAXtPaIhw7z6OgwRJW7Nr3j8ROYbaE
vsMcUPtGZArwJ0GY3Jt9KbOJTY/HLPVIzpQD5hxS1H6n8ByrAmIdugWxMnpdq3IQ
VAyZucVk9ywgv2Gy/AuDPEQy2b/97LoLNVesB3PFfjUBRAxZ4ZE7TBtyUTyVKYIQ
AaWVfOBjWO1GAaWI9JmrdUml56hgZRhqeNxSDkTZazJ9QXVVVomkM+TryrPshyP+
JkwwimZqZjNTNTYzXNBuz6rNYQjFISNL/D046p97AOAWAQ8PxW+6N/BKg/0sUQ3o
+bbvIxvgURm74IiQaocaZLD/0PgnS6e0khouDuDQEMQsjjAd+x3WOxYzpHUZ1yf6
usgIuOcy2x9wqXhFQ9NrsFZTvaUnkz/H82+FcJV3kylYWpjKA13WxIhxkcaRRZLf
anSnFrs6iLjrl6BgjTRk9e/pceehg/orYk2OOsU/Olz9J9zmzzTRnseDD6LhR7pH
zHnlko+GWSc4o7QgZr54nX2W+BJsxuoiykslANphiRo12fGiutz9TdpWpyFKXLZd
B4Ho/Teps/3mTpXLsH3izBsz/VkNacaIR/sJR2L2D1Mmw8s4f6Lifl2SmJ5S9CBG
1xAXbMyEXwbdu1YJt081z26wAPnTZAXRyVJmqfNC83VKHM4v4pgaUXHI2oHhv4jr
dIBah1Tt2pzrDbgHv836JWOe8u2mgoArcoqkLMmAy4GDfB7KMU5FaT9G3ESLlFVg
FCsV1cAyjMxtbm8eYn8EVGvuuRTixAqPmv42P53Q+TkhQUsRH0aUYf9SbHBZdT43
lfNDOUHySpPUOs+uPHCgszR8cV/V3PlzZJBHZk6gpcMBQqZB4JT2lot1MJxcQOv3
Dzs787zy28ZKeVBaGIOjsRB0DYdq6G3q/R4FfGZ7Cy1eqMu25+8jsDFRutoiassE
eLtSlKZ84v5GEHr7g7lo6S3Xua86obSRho9XnO3SS1CAqnIBqb9P3oNYxPVLmEk8
7m8MD8Szht+QWoOOBuDzU7mZ0paiZqTYfRtNTohvnBZ8zHWd8KsjnyaAjEgD0AOj
8io85MgDMfwk/KD98z5f8F/sRY9yyfPGTh45QeAlCqexMSgQ/T3VDG22/sB/jQin
aY6zcfhdnaXm654alpMO6cm7R+SEwal7jI1S93CPo2h9n+em2aV2SLtGgtdkAJMa
g+VKQmCRdJYhRCVTYWzfnSoEiUC+03g/v43owqYNsYJlfxywDu8bP3hXoO1gCmTX
DqkDk98e8i9Qf7H7HmPbasoNM9pHn17thaULUUuUVt5Gtz+qCSQ8ALXjo0jIeJ4/
iNjxozHMGwJWPKzdXgKWbS3+JVsut9y5BoQzYj9uDzQs7scvaii54nx5R89vyTct
AvPsPTFhrL3sgC3V6gW4dYeGzrm3+YImwvHLiL/uNKyychoCylaEO/2srSuNxQ+v
zY14rgycfVwgd3SrjEqaoRE01LDFCsnwKRqk5Zd+O8oSpPhKu/vYIUh+2A1KDKkA
zXGfpbMRAmHkUYi2UAzCAec9NAywt9VMJcGGlZ72CeqyWy4MR7zPogAHxc+WCamJ
6RY/jQfM65cBytxEqwdClvNhgi/9owdvPh4vEaHn2pJ9jaFYpw4B8O9GadFdbvj2
vQmxWQoJqyRBHXXUhxF6cMplOg5DR89PLgRSDAWtGBgSZJqCjgcNC7+KD6NMejSh
fKU+BNcHJg44+eOmfxWZ8lUdrNiMFun0KWKHP4X7fVsV2qavUqZdWYWOKLLAIqZM
Tm977EcubPg5Ekku0RSL5MByz+n0IcENL3n/t8j4WaqcGzKux6Rq+NVmRNzJ58v3
s6w5WUkrZWLgzKVQHGgqI3jbDmZMXbqmoPSI9tJvXRvJy6gHPpy6+90tNMY6NAnV
M2Y1X5IX70wdVp4gBH95n1ofmqMLkc9u2TV7DhrQtQDcQVoGJn0220Lz8mkh90e5
Io04TCxHk+aOsWlEPHecKrgFFvFWol5BqJ8QuAPO7WX/fubHhhLKtKauvnBtiJ6O
4WvyqgvVm6AtgFXfvJcbOZ73w+NFavcONe3eYyG9HxL84Rtq8X0CnJbKqliE+Puj
WWDi2aavX8MUHkXv0eo5ShaIvGPiP0oVHiUgpVpCmW+jG/cwnxz4PL3Gq79LWzw4
2vE5SKX6nD2g6MMfGsEGIbBHLf9eCXxvbQfesABS1xsQzsjwFUUZbUz+vdrRwHcr
Mxd8mRkaEtQpz9ZpAqQXEne2dg9kv2H1HLhzjIx1ocW46tcKI3rsC/5MtV0tYACh
odIFE8ywrpMH2Q3QCLuQc4bWtQ2qXlWlKVLlkukVhVholSICMXolaAI7AEiKOrbi
P3mD1XQHHepUPXfjrVJU96GqZz0hdruLYHqTmiHmwEm/ocUJ/D9JwynzElTgpJ1Z
JWAFPPKa2viMp5K9uglBLMwXU/QaiDV0+jJsB8LFb25fM+hgHn2+s+8LejErukjd
TCHz19asokDmLNeeBp6+pz+2C/ofXURYBB9wsSUBlOz+BFAvCsHXLAM2pfrMwUwi
enKb96DfTJaaAPBr14caXuYjepgJBlvG62cjdJAaku/FEiBPuoFISbtzS93/tgvE
RZaaeYegJx8ccfMrsk2/VygTnJ4aj2JXw9rVlbFKGubJV/FxSer3CDDDjBR3P+YC
e59+bx9nrbfwVXJLdDxP2OIlSR5gkfXeNAsNEdRzOWO/X6JyT+YJ4KE5hZm0P40v
KGdVyLRptyVyj6mkz4tg1XXkr10W1eZmDfM9Dz/Ld/cZnVHci5AbmYZB/BJ0BMf8
QvcXI4lcY4LZO6DU6p0+0dD5NZIu5ermPTH+Myj+4xuoG31ph4JaCcHkUfyUKD+D
u22MOrv1cNe6da7limJVKeoTRPyUNiiCF1tjBNltT64vZ9ZerV0hpP8XtAIR3WeW
XOUxMQ7SRiC1457fuG/QXiaWPsvN+Jfmq1nFtBJJ5A28zA6Li7hykKRwDTWTVb/5
kcTqsBLXh/uNY3O/IED3EfUDxxNmTXk4vv4vHORqxLBdPt+QJLtWlgNKiKxkU8NF
TB9smhEypgv42Y9Qe0pSr7nT51DDFhphM6mAhJstLHX/gyEGSGI3SS9+5hNMsXj9
53Tnds4QO2EeAFTqN2p1H+ivW6phEbKofDxwt0xl+Y4qUOA95qRviG8inEZZPptC
trFMP8MfRgcLeBTb8Oz5rQTweUw1O38PZjVOKYUlSa0JjGJW0UKNRMVMI6wevhs/
RZgL7uvb6L4hEqmQZ3GFbWGmRYr6roaSTmCBudkUHXZxvc+nv5a3q+ytF4oRszDg
ik/kPxgXwq+HhsavtVf5E+UQZGYhd79DeJsIHObBmn4h89vOlAttY5siLbriV1E3
JZB64UcPYLiZt7ubjaSUI2n2nIaSXtBBdBQjCwQuBiC4Ru9p52tuIJNl5c2MbjEZ
IrLvED08Q0g5GSjTG5OzY866KnEqm/h96undyDrPq/bBV7xf3oyMZKeC9F6CzkpG
TLxSXCAIeVuWd7sOdjV1/WqasN0O3DTx137ksbQ88oH2wUf3hmGl6Fyxc781JnCK
`protect END_PROTECTED
