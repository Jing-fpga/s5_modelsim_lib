`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9slk9l+Dze/Mb+nf/Sj1ZMeUcwHpEiUdXo8+7cGluNxnk4fV2oIGmAC3ryFTXoi0
axs1f7hNwTlpokZTuhlBEBFxfvbeW+LqU6AOTf0o1X24j/kAeheDpvmQRgW+cHL0
LtmNZfnH8SsLKqMdVoAK2UTbQIeE7H1v8incn4kfO78gGNlgYcAyuwXx6P70i1t+
g6iO2LXaSuMJFU4qafDuxm91ix91JxtGLY8lIhclD1xM0aLCuPfXtGFYB4NwIrCp
E5s7vHF2C2CbdyYrJ7z74hjxgD7BQU2KL/vjvRl8xrSzsLB/TANFNeUMxxtaacyt
pjhpoVstD8NgSLuNSO9TZcv2KEiH6/Xn7EcTpM2M9fXDkRBwKHP19NiyRe4G/gRW
O2BvxNyiGQgzlCRT/IvdD1/FbYH4jy3hYwOF+YnzoUFBB0E3tD/edcp5U9pUL4pG
ZjaHvqDIZQ6j3rJaBXDjW7LaaGFXDpwIo1zbW2CmIpt97r/TyWIR+E3di+RfWso2
7HPGvdsrG8pmyhJd0Yly+Ulw5vwWk3uLtFv3GFumySJJCWSDidHhgg+P0vuoCYb8
Zjs0pM2DzmjHBnkJtqFuD+fFAlrcXloBSSTdx/fI4XaQxuCRf4InIb7zCSJS0CJs
vfkFl0GCGM7OwmDrx7x/jJAFC8/BOlW+rp3ZErbuZxhc6hHMMMDtmlDcnyUWlqmw
LIEhiR8a14Ixso3QEpty/fYeKl/mllwwD8OlFFnwPmE16qRCmeNJQE1r1dEQ6naH
4SoQE/SL7Dlm2nTH2wfZz2cGV29l/IMH22XKUvMOdDwuf/XjONi776xnP9l0YFFE
TCiDWuVgwnVDTJM6TvKLPtPY89m+703pL0Ut8HRvuphwfWzxYBprgQ8myuaECYe/
WlEKXHhwT4hc+cymKB1EuqJRrFOLygD5eXU/uftPchfueh3TgWa/o+gYymexpvLb
8JagAj3Lqzd5VpcBczdVHZMy82mQjMaV+2QrtxHuPUDLbIOpYM0WAA7mCUV9ZDPw
jAwjjWG/XNl29agcuaYngZ6nwEXMrAehqlcaOWIRaBWzO/TjVMTFF0A3W8FAEOKl
eB7gt+lqBnPVMkCS3Qh5hTiTTE9lFFSJKcDfQNlp10pv4HgwGsEdWik6wwBcQz9U
gr8IM5DFjn+NXy+NRQVaqJokpDwOg7pYkdQWISsSdv74D0rgRJrObUohZ0XFuwbM
0VEV4SDiL0kafsX1+8fslFO07DkYNtLD9ZdyaIKwd++PyxZwCc/mjiDJs5d1l8qf
o0StKTAuy7XmhqdKNut/qRPYo6F+P193x8r4blhn4fsHqPCdZiJ8kJRFtrS24tcT
xvQgEXlVVwkD7YK9ubIOCsfmuKS1pTLkpvc+AKRszzPXh7m02dNw9tl6SJxDojPS
VmzZDSRNdqmcmUtivfixdh5NCkwRsqkIUyVSWVKHGUBui5BGbiEiy2A5KjnF7uJl
I85jysLdYs34R/w3gE5G7GKors7q9wyE+rMlonwagjlsT0/Mzmx5wh3dl9iigxkL
UY2l45iOUjCd4q252fkEUf29wQgSCB4XCskCcoiTwzOYX3YZA3deA4FD/9dsx2F2
XsZ0EkcOdQyjYiSE6DWOiVvuj4imdqWC8rJmMFvb7uyMk88G0VL/EcnaiPLGA8TM
yBapPVA5EZPpIiOBNyAsaHoaA4csJ3bVqkEJnb2UBRMUZvMBblVszVtNvr7OavMZ
ARsz89HDP2yKDyjcxPMImJ6eS2m3qgn8AbQ+KTlRX0eYXrkdKt0CNvtowB/9m5G5
dtKgvUYxmakGeGmDMBB9KgYE8OuXkuEwF54yDKp36oKv9AQF2hLiuJg/QhV1sDLK
UsuGLUyqWfFt3Nr3dYJudp2/WXIojZxmp2dykDQFURyeR0YO7gIksp/Rj6TDVzIb
gl/kroNq4JX6CC6x0tt1iWRHKqed8ULE62ZsZ8O7NaM3l23zBDnAdQDCjYcW6Xgw
QK/rkxd+OBWBiLSjhmb5x9M1rlYmFgzLlVZlvF/l0JA0ZVVT3bnf7A9/arQIOgb7
NGR6pdGoG95B4vwX4Is5uMGFuC+sxCRSRSUmqSU3gWiXfquIkIGY2FoBne9MpJ+o
pgupcMu7rjndyNdte1QV2MblhqzSGjxMyVRY1cKYAl4+tDLrScNGUpcpDUZh3cKY
m79bJa65F/4s+WzyI/jda1KN2D4Rhx+jjDhIRu5lqOlu3RlUZSYrwXUMc8rP4JZy
Lo6a6VBAZS6IckzpKqECGBKHgJ+kmPORfe9Z0pbEHg0bPle3CdjkRhIIPXLZVU2d
EUBFxif8vNMlxA+m9xeZVpxWQoMGYmH6uS9Nuu3pcSY3gs+BKzJGs2P/QFbr5oPb
9V5YdNCpzlLW6VJ/9VZh7FzzdT3ZGWWJCkzMWstZCYhLQ3eGew9TmJW8/Sf+lXLi
uK4RExfjOSaaKokC9zxk/8GWTMtzEojPOf1RDGku6/8lAA3fjWUdmXLtvBx0q0Em
ywcYb39arIq5TQSQD1JXh6j+FfDONsoxeW0Bnsazi4a/laQUXg2TbWbLteEmKenf
E6Huu52etzhYstmD7CrrPae3DI+qh1fxV2pI5bpU8VIh+Rmv+NfR8fqKTGtiJjom
7BJPLBlP1mI9w8NOVAV1AezrC3YZJJr/u0h1Zx1DQwT3ghBFU2N+B/75XDjrZ0fe
0HY9RtXDUXL81wTB99yWFr4WBGKjX2pBLCb1be5mKE2QFvaiARrQ+fMIe+rO44/a
AyRsE+rZW97jBH2F41/FYjzplCib8faOLeOGArl6U1racaYPSKw+Bq5RhRiwkp9B
jkSdK0fOfmVsOJKzT4ZW9BLU4DM7Xtte+FBiafgCn5UiE9oeSlD/E3i5KrpMg1hy
UC303wVDDD0BRhgZndVaeNMpdHxdgYL3yaqbn9jgo4fFCdB9sQcSlg4SkuVfP5b1
wCtTxi2hwVTSGyzhi/JYzVSV8nCLd4t5aMJulEWWRHPUEEshJA9J6gpmdd3M8uet
yeaAYwdB1lQJ94500NpAnmZz07ksOomEOzau8HkMt2y7LwboAyWwJMsy0KS4WZZH
EOwiOGj4fHK1K94OtM2C1Zkeo426V2tRYv9ExZTlWm3p4Tcqw/GtLSAlefzn/L18
i2KTILpPE7T/U5DGST7+azHkyctlqnsDOYdGkr7ufkIG6iWDEJmo0z+XMciP2Q4H
XLGqueSga8pbmKkfehHYwY2r11VR2e9khALPuIkBMd9L0gAD9I1umUyz5Ka35KNQ
VotojerT0T9Iq8AmWqi7spnhZX/HL0jD+FftMY1uXEAUNPRSAj+ckDoJz5bvatfd
oGLH0vNVK0XFIf8rRInRqKdkhgP+wiVDmT9D7Y/FnByi1uGM7uvnalkKEwEru7iC
aS4Dbn31FZLrZ5fYZ6cZZeFwm0jpHOOD128e2i9ryBLdS7SszOSk7HrNsro1HWzm
mq1w2d+2qqObgRmoU23Octldk1b0I8z7kPkynAaYXR/l+3s+GfGTipTMulBl7bxv
I+ZeJSCpsJ/KqvEGSqypMal40NVwFx1ZEdmf18huWcEvbJElZEjGdKn9hXXbrs5R
yAC3Doi2jKtK4OKjNis3kidteLb8CK+afY83mgtDU0yBaHl8iokP18U1HoPhT2sA
dAGkFuaq1rjSQjUwQbaF8mJ7rKn8Xxz+M6xSP3wnUImHWQ5KtcbhU/y4ohSYkZpa
ARiuz7mpsTLfe7H49sK1HNhfRrqf9pVXWR835BNJNyvncbHug9R9HTJlXg7Eksnm
j64eWIFw/r8ttMd8mV+MPl+KmpS5HhqHLxF+P9XRB/8STvk+aXhuVnuMg1MENEmD
A2OUjYRn/faiOyFS4yqSYQUE/7FNe5vHGGO7k65l7w6juV2pR0ogGk2WGWBDN9br
SI3Icf8jU7ANEiFGInh07wHvpAlzzYnO5HyO7c3j/mHoQiK51GX3GK8cv4rX6kEH
hMM0eL1qH3p7mH2KeuqxmIJWS0Omhf50AXIEjyAWCDV/O3CoW1JkfbLLquEJIzaE
6vUgshOpYHiNqOcFoJy+c9FSDnxKQko3JKl7UDp89/XR5oO6c4MPk5ghN6rTAl9s
Sna/nAXd6V3naZxCelG2TyMBOVNxBC02Q1UEn5Gbg4rgBqXQQ9HTUMosyNuB1/Lv
T0riZN+U2JwQOG2GYeCksKLq8ZRdh//ONpAF+Si0YJ7oHzZaOFdeuUuKNvEpBVtd
hjBD+NRb+HIRzFzwJbMv/VrN8N363rWOfQF0qvraVb5teWq74xezNuGquqvDIBpY
P08mNcfH8h7IYNxBn+APZ3fYPYi6whrWDdE2CSPbQ5GnEIoChXWWumcOoEX0X8nQ
Qaxu7YgIoMW5he+ziNdJN7iQjb6C6irZm9yaxtgkiu7lCWdVPuAFunHHlqhxVJLe
Y4epYIsn+TlyQpxIQbGNggsv9n9cKnFdxWvmZ5bj33lWIAZt3LixcGtT8x3YNMkX
uXQyjm0k2Prt8jIGOzrVrDL1X2FvnqWxKY98mYQkYjWzH5hRu9x3l6kjQ2hRcgIs
iVh0CP+M0BGvM7gdrZVqFSJxwhYN8ZyFmQGmgwF+Tl1Jl6wDi/uftN8J3QjgjvFf
0qLYaVv3CQyRVumDnVT4fBhLrQyEMcAjJUUUMJ6L2GSRbIoh+wFccrGKpGezRBve
0SzSFe+T7Lx1gxLyBf4RF1fPfyLe5SFv7F1YBGahAE9NUHFef5AxHcSZ3RNHKwiQ
4Y9Uq+ub3VG5hNtYB73+uSkw9ef0oIwdmLqaCHdEIHjmuB/S+fHOgewvGbqppeL7
Y823XonoKr0X5jgIhW7uNT9Tk9DgRQwxlt0RNXzEHvj5SxxqjrCCklxlwqy5v8sA
/rOdacMIJrIwwGoV8IRe0chZrvn6vN9Slnkymk6LQp0odJJWZOi9JwfNvKaoGV9d
BtLMRO0W6yQ9smr+0rODJR40TGHyvoYCB6t80YaiDWPXBAW0KpogEyzBiQYd520x
KNFUo7vWhUwVra5Ym/CxcBb6AIFRx/bGb34sNmaLQIelC2D2ZE6k6kQffcmGgoMy
g9r1UTaReiSrUFchuUx37pTCnXDaOZVmkrc4dPEzBAE4F5ZHSOV1WETsnJKw1hZ0
DiYlb/uFSuAiDhDc+SKM/koiv0DGn0eZ5brszRQyb3Vy4TyJknmVSRrLhUCi/rRF
gG+lRg2nC8SlFxIPgPAlga0werZF3C3DDbhD+7N/s2mn0LjJFv52IHI6wO1Cfi1l
1sQfLg1nPj9ORBajoCr7zz31GpYYIHTAj40dKY30Wa29zy59VMC3fl2Cbj6ZiPSh
2udhckBDSsz/jIw/UUBA7+BVZZz9Lq/w4JfccJapjRLL6fhheiH/1ESrxiA5c5pK
pLbgfDwzD1nHynAzjrRRaMeaxgjSFxn3sg0BxvsrTIa+qpHMm/i2ppgi6Tdqki+V
29UBTBIp7TENPlEE86VF1S1Z0sRwnCoZfeWKXWW5l55JslSzb8Co4YWx7uyzpMFo
4HJb8pCSXEqtfSaHSnqecucUqhnxiw3FrRoTEQjrnmb6Ubc0YlCVTXMfUrIe3A9E
`protect END_PROTECTED
