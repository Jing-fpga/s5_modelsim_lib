`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eZt3xYFEyqSuhDiuFHUCdkbZ+jq23psCMtGrYrxVw3KkpgWOUFB5IfG5y2E2Jq5l
owv4lRj63D875CQhUzYEvBOh9znxCAxQ0Gk/Cr5+Wksnf4V+xWa1DbIvtyVkny0T
JPNzqAdZjvbLJhUqwnoBHpK6t1q2AVZvMBFhLxEAb5mhcORkE9UFjwO6jRJfaEz9
ZOevYBvPd5AW+zH0PQl/9+Nq5wpeENgBc0pUFPNFi1DPQuwyAhOIJt3CDZzPjDDK
M3uWiAVYm32P94qrVLLWylXYBTTsXlMXMxilKA3NQunLEsIBLwE90h+at8ApBufs
z937jsfCCK3pKJsd5ukdywUbzkfhWMJY6oxHMGVDUXS11a/ptU1vcMvhYV5xkRgj
oxvCGqVHJov1aPca0teNjEe7mQyEqn9O0/0bPnFZOM2VbvgN9qOKcszWLmuaM3b/
A4QapwzFOhuzi/jtSyfVhYxBvhOKH7WIhUr7pL6UsysSO7rgNNUc8uc6eHpDN549
GCfZI4KULEnAlY27JyR2xDjZlIhX+iDatiPwWadY/IL0q1rwLmklZbRnU5W8yG7L
dekBUdSR1+75YN6Sg0WEIzDSFg7PFro1PyUp8aixPc4MDjrw0m7HyX0lxJoOlK6A
CheZdMJ7sMEXTDrKvoVqwo1VzNwfMGEMvgp231TzcR4hwERFCfvHGFos2N2bXk5c
8u8R0woFEgz3nkGAZKMAQw1WAHVKw/T9wYOJuvwCBXHkYgYoJO+gYnaVb7orv5KA
9hWJ+OuOrzaJBSO8G8dzYugdBFlFFSeImWjRnuZwPi2gbJi7MzICBuZj0Hzld2Bx
IsTaxpf16nUmBFd00rNUxVBUNPVDJ4Wp9DxYYTc40x0hbiQsir+ugQXIt5VOw79W
4NsWNQjLOujsFy6jxbx2Alap/xg4NO9ygYS6GI5pHq4q5sOZ4WjNniISUjJzJeL7
vuwYkzP4xy/b3zkssgOdawO02hA2a1CRjY3YVdQDavmtBsNmJcfcLx2KE8XMB8Ry
w7zvWmDH41eW1SNB1jj8cT+J+b89EXTsuzjN2iRrDUZPWW7pIXY05jBTD87SUfCr
wgQ5A001U3kJKUykejDGtT54hacdnmfcPwiHQ6+skum8WsBRdWk5+dPRblS6I8Qu
98msYNlCMQHIW5UzhEhRa9AwpuinbRJnB0pDj+urS9Y2G5pjw5Hrf4OcGduaXuAl
DCJ7UKG1DkfgV8G2aFUvaaEDLuvYgqBATDBoqlqnWweHU1OcnWFbF96+gODhIl16
wsWcw4+dXedp3DX4Xh8Zsuug4Yf5Z/gOEDARCz4tjJVdclYXFJrWH549nGg2YWrq
Ed4winPGk2aqsd5Yss/OvluxuNASC7hlrU/TeVSd0CXeO4+iuKyVKWbHXudXvJ/L
QWGf2A+5LCJ2ToY16HVSBDGVsZtQ4ZHgZ7+fEmSZTCTzQJ07XhcKTvlgSuxj4Ycf
`protect END_PROTECTED
