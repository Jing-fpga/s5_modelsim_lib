`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5gj/8p4KMeyf+fwaGFAFfcA8NHL21wzntHsi6BWnstLP8uoeHhf8MC2pYZYho2kH
bVzWM0x5MP66FmZ1NOl7e8P8nHje8Ith4qvmftyyP5ANIbJiIgS1u2nRgJAHS1+p
+hjyaVu2wsOoplOrVyTy9mHLkPeG5R9bNXxDVF+qmjXk0VqayvpE6BdfmrC+k5BY
AjMJ5TnctIV2DvPTxhcAMo/CK0A6LWR3SUU6e51kr2E7JuHULehfY97rDzBsn2oE
DKhVj6BaZfemkRnAtaLd8+BaQ6jOHie8wun/dFwpJgEnA7bmWR0kfBbQd38Pb2Vj
XoW2kACPz1ZYHS6ALzKmEpwVeFEHGZKodObgDjne9HnE60Hiq8M4Sh1n4JYjm8cW
y3Q594G+ntICPhtoQbDo0iLUmmp9yGYYBARutFtn3qn81r7yWyS/cMgXVcktZ7sb
IatHT132+RSGwrDyOl1SUuv3LmLlbmOPwoS7FcM8TN1TLQV87vBB9fNjAypm09hU
mEawy6FSUnlWEte8I3SK1pacK2tPnBP09K8QiIffITRJQ2bn2sA8UZZQheGW63A+
0dhLheFbTxLC18vqWNO/yahcDoZx+FkNLt6Awn3KIWnRWUvtBmIlE8rPXvEs1Jeq
IoCErR8lNSaAup5YGV2lXVKXw/xhmvSKQkB+uD2xQmff9VSX9hRHS58kiZU6Yap+
zq4aNdu2AuSV+GEzwV13E4PaATZeOK2N0Kw1dbhTKqvDLsO9iAfKbFbLeMo4B8Sv
+h7FlbrUiIlk1Y9Z23v0vlu37ASzsPlgnpZkf3N16uHw/dX0WSPup3vnxuor7F6d
V5rJDdW/GkgsONBA1PreMA0po6y2eGCjNFjiJnq8yWMYHqOwOkT/DmyoPLrQJGrA
A9OcpTlS8n3mubGaa/KYZROtqm6XaX8OXcFAIwlfokpEH4F4h5cwQYXKY5n9L6yB
M7Ctz3Bk5d3SjoL2qB6zGQDnbPWDGQBoJFrkmapKxSkpdMmEGHqya97Ql/5bHJkj
xwGnQdK4OY3kxFCNUcvMoizzzF2iM6Hzc1hKxVT+qJyJM0YJrgqzx60N8cQ9JDiE
A/QzX5NGmqI/In2o02EBYxt2dQXrzkip+TMeovVmFpyxn/DlLq5PiIVhsmEl/it9
ZubMtZux2qapTqSlFhULmFk/mx1KOrzR9h++FUy0fLmzeBba8almik5Wta4R4JDq
/Z1xyO3gCaLJSfqAFjzk/6ieffdzMkb8Cm7WiQ+GluVsgLuaLtJmPO15UDqhWG6L
M0w0FKoN4O/hdfduUZN/O5JQmV8x8nlq42vOa/RFURlf7zqEphua3qeRkpeV5kgh
n+2Q9MBpRdXp5lS9V3XdSe8u860WfXv76XWJObR0Qc6Rj8c9741m5mzr35Q12fkP
9VQd7zqKEn5/72u03ST/BEafkx6KyNAHdQFszWntCDFaXWz3CbyTgsJ72KxOQdRz
SMloyX72NSy2nYr8WHdJUYoUxSZtz8IfVd2f+PsGqkK9M6tEevXspCLaTWixmpK3
5is3yxwyTVasN1lDrQjS1bEQs8U0mK3xL5ezUaQUYJIHPopa2KTpd7zsGg5nl0l3
9NW/ySTSH/R8Qj+JDMXVf7Q1k9qiysKtFjV9zJLysIXE4+XdajW21m3b1kop38/M
9gs6r1XCMkIHIlPOR/11zfu7plsi2613ew/9ENpdVS9+Un2NK1KcU3ikf5U6iySw
JCKsWTQi8ddhDOxHSqgm0gAJJuvmlu+TR2EHi111QIKktqU9dqSNbNNoGXtyUfgY
3x6IWv+b1DVxi6PSXG1FQxGqQV/skMEONG0IJKNx05Qh3q+PBwH3RUd1G7Es2xnd
XfAEu5qMVI0ZEd98kj9x78okNinnRmYJPMlfkLx/ijpImJhqCyCOh/5Zd+pYx3sw
ThEQOdyeOuoNwtwMz3cG3Ku7iy4SF3wVan4nXUondGjpkomaHCYnZITM4jctmLVF
vMGkq3cISxhWnkIW+Fa6/LbMO2Oo4onz7duL7OYsy2O/XfwTfh7z556Hvp1szF7u
WPpudeXZLmZ5cYulr385Lsyx9BGYZ0CnkDrxxPw6fhgysJ+JmcpJgmxMX6I5iP1G
96XKYpTfQMkyialz7VfoaCsUKltWh00MB351U2cML4pj4dG89fh7IrZqBiAkoimM
hGT+te2nC4hzMN5CB6Dd+w+YuoBOTmzmPGd0RSf24+FW7yc47xbQNYLRU0yTc5zv
oTo5e7ZhoFxpmD2WNZgro/V7O3wCN2vq3YSm/61g5FPFsAMcxvVqpkd05uidjQgw
1HgFQH6KyQabl5dEXuI4g1fGUmb3QXHT6z0XZlkmlED5BcY+PIOCenD+pf0N6Mqe
xIWP/htAUirVTiDlh8c6whpk7pQe7zdIdeot5vgRaAJpRw8LyTcllzOvCMVl45/x
wN+gWqxdO8NT+vMt1GwSvh9QaoEdQ47ENXclUwrkmpPZlxXRYxewmMXRsMgjlvka
nLPf/MEEXx14kSDjMOgCeYc/lm2WuDxLEkjbnZDPuKBNLj9e2cENIyFkEFBDSCuj
fANC86674kDTdXD4tmUThQH+RZLsl9Qvm1C3nf0CDJZe/3SB6YpEU87bIIKS3a5s
ZA1AbQqm/UTJ1LWLQ/wv5Dz4VTZPwD7OvNc6kHvsmFTtcFrgQPqmfPQJE0R1Ro/G
m5/mWXO/juSbgGSuDl73Mf8uf0SJYL0G6d9oCssFBseurh6Of5TQB/N8bRYrvXR+
tshpjoW2rC3ZvoQIyJBKml52k0gb456dFUSNdOvgQZGq2GhSuvNnDnzXzmpT9ohr
HYR38kp70Q+V+Yozu0Pdzrxi3tjkeYmzyZxRHm6sUvuPjtAhm+LulYLCGy5tlKT/
MPJxseNffNXIiYxGm4jz5keokockA31dEW4FXYYxXfgJOJHsTXjhp6c/0P9mDUel
0PKdPKKPgV7ads9bw69AXYiM7PRg4Bxj2/MJVycEXmdpuwsLdQCnXYB7oflNrXJq
EmTs+AbNHRwQ2cS6LXc4re12h9WlQn2tu/Oub8DCO9mH8rKZxZp7htMbMDel31wg
y2YcLyyj1uOz1Xvz3eKcFd92+5bzIeuuO4cV1qx9HPIdKi13IcTChykGuFEOMv8q
FdF8CO01eVpPp63S5UY0XDNyfHTWJJJTQM8M74fJV8DAl5K1wugLXbu6xLkCKhYf
PD+UM23luJvKwWWhjnVA4FlJXnwYv0FjnsRG9v1rQms=
`protect END_PROTECTED
