`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vp1ywbxzHpWlc9zJbiS4PFarYM52vJS8xGgW1fNonjxSKupcZl4+9cUIoa10wj6e
QmxQ+eNNvjP0iiVMn2Mja8sVJxpIn4kNDRrLI7ShloE+CCZB+8+yi3rteRiUhSyx
Ku8FN7yH7zhvN7M2xYbA9luh8WAYs0x0LeE6hdfcLcXmzMMALwtgZZnFpawMu7gd
cDqNTkBJmJiZC7xk2ucMR+Afy3aQAXNa7+EcSAtz6F+Bv744UGKxjGQyComvThNE
1WRW0DUXuCTm82K/qXKW615gKEmD1vH0X4usIFxD1k0WPF2zmiMRc9H5KvgI3uyv
Z11rhFtwpUZenfNhKkFbWjgXhK5WqbWbym1ongs7luGS8H8HZ/rU4lCqBMpgD0su
7X40pYO3+IfGUY0D26EwU3uSB94RkH5WIg+1Oo1PJsErj4kWDM5P8t3l/H0udOTu
r17bTh3BlIQmwXXelOJJUkNB8mSOfht4uiKHqr/IxW5g+/zhJMjAPy2JXMPMxNW3
qt6QI75Y6TAaCptXOIMo97UA0bffCkBA/jYn1xs6BubnBZKnYKR7lYQZ+F0BRf+d
7x9bRki+puDoujIrEupjdwzHVjpurqCAr5l7DwCPL8x885AzRIQonXFUSmrSjrgF
UeFNuV6snsEmL88ssMxDk0b2m42QGtqvAXCmzLFbYyq1O1OEzkR8d57sZihgb79O
oPd3YtFZwmqZ+i6U0jfPSxCqGVr6YwXrI6VT10sp6v689qhiEfvuSopQiNOldsUt
9fVS3AuicfRQVgw75FWlSVaDeRQodVucWALsbX6M0id8rBDlyzSDhy8ZCaRrm4A2
TbRqJjQ5cBbNaT4+3XZz+LaOI9svO8grdCayorNppellzzW4r9hqV/2kfE5aT0t0
055wqvReWwHJvBQ0jwn3SjbYD21AyUoZATvbgyKW+ZufFRPCBitwEJT0fhSRuBU+
2fFJ6YC5EU0mHOUzJhYeJdqsuFWCsL3jiR14d05mzgyuM5sDNw8Qh0EYhPtRSeLv
o/Bnt/xIdzXaACSgWaqhNs2YM0DxVIghLVK6p+xuS6uxMXH9PIuSgh+RQtpzLOYi
k6IJOqpywmy2C0kJLPueGc6wuw0M4q08hh9RtamEgOrN9l+MDEJdkaUSluu5+oXp
SkIYoJ+93wR4gxx2fLVIdkuuluaPd+OBPiri5aWQVrBbvbAR2fbj2PdocoCogLyd
52SqppB7JeND2489NGL1e5iUYnj1guw7eLJEwWWeXezGiJ/8ZpUif11KeLRmmG0f
lqyqY8hBufJAXmxbj8zcIzBwFFOaLb/r0BoyyPqvYvcstFeK2c6zytucFjQFmtbi
ftpqMpWm9+uEQ7u3HJ9gFrgsu2YFcjfq+guFQpWUAO3p4ARQBiag90GkdGIDE/l/
+0DSmS0d7z6ADtyq+pjDlGNROJPN8ZQ2lB7rwx4j3JP+0e+y2d8ajsMcSN+qTdXV
25H1oUaNrirCihgRprEmy3gCYjhtE3T1rhduen/NnHwCYQgYG3sRE77VIenqGhFH
tjizRqdEC3P0B+oANgM32Gia5wsyIUd+V3Gcs+4vGqjK6ZmodriZBAqMhCRI/BDD
2iZZtjT0dbP3GYntIppCN70RfQFOBfYNjBjWvoTU/CXieOoI9bMX8bbMA3RIjqMj
QeC/HEMUF3hDS8YPDSAJrerVRY1fi4XZ9uta15xDi/XjPDN5ip0L+rbtnWA1csOe
KGjekKrXT2L58gC/hW3ie5w3kmuNA1DHTKStAQM0pVshx9VXZibQMRm6VtgryRgt
0AbhfkQIU3PiDWg7BaB+5zWgW+w1h8tNu+NiMsyCzZ8pK7X9wx6fQde9Sfk6TqZ5
/L1KA7ohGCKpkyxIh74zwNx8cABbrtGAGt19galJ2CrV69nCB9MYN4Y5XUoIDOe5
RN4zRXS5Sf6quVZkzLx+nmfAbroJUOcIFEfB8BinepIp7MCUC7wMmEI80U/BgWos
Oeh8yuIlkiNUX6gpKZQxMEFrwfPIIdd0WNMcVKtm9qqUdabIwH30PcFCOYrl6GNX
yN8yd6jASg4cpNY9nq9lqbNJEdd6lzijiUhTUdISLbgLo1aI8xyh/9QdsBnWs7UZ
44ogwaZJPLaRWCKiEkC8ezu8s+S5RAKvSTHm9rQpiahYwBdTajQvh8KQcGqYgzQz
JeXLKMYAAA8sIxwM82buW8G2/ri2ZkPLeFEdv7okDkyr6zw7HBOOZQKrvuq+IyJ1
sIv6FsFKjchF1sGXmJAypnl2fUksNwmuiW0Yu6KswaTwwtdhHcIOcaj3/EtvbpLf
kmgvSPDE73y4JpLlw13p8kkridkr/hYndtXD5od8quTY2jDdHYzwj9DZ393A2Vpr
oNFlUMtPq7btp8w+scDOYg/q/IulrD5WiZEEr9yzU5vv9e5fsh7x9sOpjxn8gvbb
rzCxtDQerxbjqykmiq41rRfsIHB0UMBVxCpy2fopIkY7GdHE8Vk0I+HdDo7o2t0K
ADKQAzDYDsdp/3RkrNWvh+JucGa0bfpYQ/zds6VXocAe1+YXy2DwjZG88QJl2jVW
VQmr3lb91JDuf0nrxNgCJg7zUGaDLdv7Kgn2FNs2BNO4jpDEcN7dzyMt9Pn5hRJ9
JHevIUx7xxeNZmGolqqDuO0J1zGmMMJVTtWptz+lvgo2BZOxK0iDtD5eaEQFexFp
4A3S26shyK/jacG/L1d8n4+LDRf0xw9tMX+dwoy5+leH9BQg/HJJGh5khbCpVjip
ga7puTLrJI3m0xxfWy/mfeXia0oLxkRqARxkofGF7rXnYlnnRmhAXbpPJVe1/rK+
QPgPgo2tktNiu89EuMwovkTFy3mo3T8x7HtPWamy9VJTk1LmyzGU37G3tCw8EVPE
h3GS08+1BSbrHSiurAqNMd3PgNIXMSlADK+1jR0+EH14t5pUYV4ahVyKI+F+m7JS
eqowLXHrofblvxb+Xni5V+QaiHhPG5H6pDseyauMeEWDDL2kAPtkY7BFINUfPlJM
7ZL2mhJdrTQYzzaA42AyCMFbFC/WSIpDg72NvfE9400KA2gBiG1haKDD8ciYQNGn
y2p1/FRN3YOeyq2a9MVljb9Xgx++JoDFS0giXZIn+dnmhlkaQBOIv0Ydc+F3WymC
Is1fs9R93dOY2p8M8H9GFBITQKcpGoej54U95pJJvuquXMwaDUAjfVqDr1FubNsI
ADxSZZ65+XCT/nww8ceLWMpGqMkNVyJ01LIOtdnIqEcLaiZLiYDPB8JsgowMsHQt
3vtqJ3+sbs6/If/91r7FcyvMRaaQl0jOAgmc/QeFlakAwZFufYYGvmq5k2Yt4t1j
evZ4+00MpXJT7ftr8VBYSUWfrTDEF+wio3gEVYIrrWCSbXtTL7MRz/n1mO5T8ypw
/yKUqP2Qu9mIQ6WapmVNgWvqwhn5rNSfjyLdWCkPIvfMHcEhIQs2V2bxzlDxTAZP
93mSSC6LjkigKT43grrYEh6692e+8TGc2eZnPNQr1rq3rJuekVrGRGuUvmdWl9Wr
7Oa+fA1m+TdMpn1C4WhAfco2KSrb7UitIqT0Fev2OvFdIdn3Gdh/4E4rEqx1EEAW
FjYAkXFxc8ZVOa97IlZYRWM7UwHlLcmuHWQ4JMgQfSGtLkBkUIMzTT5TekXmnOPH
Aoc3JiWA/86AQT9s2cO1YyMoJdCwpWv8+QFZovz25d8+1R0wgGytiFtmX3UiuszD
cI5ot+LAmJrUKWL1amdsVaaWxGAG7r1Z9EckyOE2Cn+5RZ2sI2h0CIiMk4xuPMJ0
rfg0C7qMsGr8UPO8IaWzf9ac0G1p91UIVNF5PqBE3WWPxibu/Uknyll8Lv6EVevh
9G6CdZiXReXaZq+nkz6hrrilD+n61viVgmfS10bG4Qf9BQXJE4jnoFMcBj4kpWE+
nuXcrVn6Caf7R7R4cTQoygbO2vriyOwT5PhHQwq9I2stbu4ur/EHRG9FrjLvPrg5
P3E6i+ss5cACaegoGJNWp2yiHPK+gXJ42nQCdkXFPzDPPt9tqyAKuEYBexuupL0z
ZZfmQH2detR27yZSMwzpJ2mARGiswhgGzz/ISkEABq074CFj8oJNUFnLnDHhZusL
CpxZEW9+B0uUjJXLnHvib3uuSjoSw9kNwUJzPToclOXl/XJVvx/5UW8iV1u19cD3
eu8sVG46OvueVw0CtV0TYK36xU/rZcCuzGUWYRc/wp46nNgoYSaxvN7IYr24jNGl
wauyBhoS9Y1rPtEIQ4QdwGvz1XtOYxxCo1hovFTUMCbLVWtP5g78w2PMdLV18v6U
KYURhrBGrp98rA4NvmKfzMj8R7yrbuVUeN7g8gyMp22bhFTn+kQJfe9gTRcSwNXN
YRmicaNkatBpRgf3Aehl8R+4TlDFvRKxUxOqHk46CWcrINfxSHFnRSJPNeEuusEN
D61bPMsU2glun2MeAcFNgSrPCrqOpd7ST2yN5DV62shKXPan8aayIqT4yzYR+QqI
BZ84VsWmlCvaWUyehdfQccabid+Q7ddAcr3O4FtnPToDtEY5MaJz9WPrztUv6+vY
dcVIMa4uXspkVrv1PNzcDITwdLb+K7xEpoBM1YWGtSAQw5kMirXyqwtp0Fo10Nfz
pqNPNygHrWTws1K7MR3n3ZHYfT3pUAwRfxSomcROsIvK6wMX9aMkhhsyHHzAvF4q
3pffpXkaIBlU5SXlyoj5VUvkZmq10iVSOJzKOeweyD4rWJg3k81nWjOxct8+xjPM
5ix+DA9lLWF+VpJvncMmUtvMbQ2FGvsAfpTD4c4vhp/Wts09a0QCouBzriBWhEL+
tGnHtQUDbzWGmXLJdQObkw==
`protect END_PROTECTED
