`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fg39qoqs5zZNo1i4b/EMSyvFJiz/GY1iHcenyfPU5KLy7KerE4GiI1ho3kuqQy8b
+Z6653WLDwqplaWKHFIKyNR8AcFHVVYFWgarN+UBNm/9QhIMyLtu7EvxE3GGqFQU
WSI212GrKi9lv7F17LXHBPZDc6d3/prOxB2wnxeGgWBWbfqpAxJQ3C+6A0G54opJ
8QqAHVTeY2G19wLW9Fejr+FLLD5tZLtzZ2PVFXHtpd6gZ0zQXP+ohMIDE8my/2fJ
Sh9yyH5KzpYVWKMJ1u9Ia+WMRs0SoS5florg/hNJ2yxeFCUj4IZi4aCRcQ9Gp9Fp
9o3aeyqBT8TYN1ARffvjldwYxeWdebKgpeBqTXY2zdWz3HN26tJhaJd29IKJ7MEt
bNfraTYSefqGA5GwLbGdLQa/QyV6ADlN0sDvCgvzTLVtAt2NKy7I44gmdAAwx6tV
IXgjKS8ke67AyacFPyTn+7Y6+pDyumCu+kvZE1TLOwSgHBvq9XEWYhv74Ps+ChNG
x07nujSTzwdBfiBub7Wyn22ZoLcs11oycYGACgUmTl7816smv+SylnCTjEx9NXEl
dTnIMICZ7lue4C5FKYlWIvoplxIZ/GQiRS7iJ/wEyBfF92WLyI1i9i2e2kPfo0jf
te/gIj3whzZfgun63wWJkeMWz26dSRU1o1vdUr9rGRsttGSZ5klSXKBSdIxigFnC
MuZSzFb7lnc4b/1hsE3Mkk/7ldCPWeJp9xyVt5j586aOghV53GTcUiVK8koTfDMT
593TrXbw5vuVRgTIqH1o4EQ1PUjCek8qGVmURSETUmW+6bcoMVAZjwH4yP1/+qu7
uuLtFfmXW8i/L4vogUyordSDxNyQX0lmho5aDEEXFt2gssHGtIzEGjVjS5AnbdT4
q26n5+BiBi8LR13EufTnv769fCa7zKmbRSEdAXsOsIgMsUPa4SMSCZHjUIHDW387
dxFOweYgbS049BlIdvSW3SbgyRjswH/MeWMRzTqB4MKMYLgdFXfeweeccjM1sR3b
SOPaz/7rECCO/KZixJZfrckbAI4h+i4P3ksB6eYMSwjQkvraqWPAnryMCVd1QgKE
3MSRHxBvN+P7sX94LQPY998VnGcIbrccjbAxWHTUZDu1GuJHYYYud9sUgLBFrPUU
BJZTIaV07eoGP14jv8e8qkMgxoRJ35fRr5PqmyNopDDteYMipFBQGgVVy7e6H9ru
quhEzzC02XmZ8CDLA4AzVSFXgeBH2NBAVsU1jz+dPAebT2DfblHjTVvdSMHFV4gA
jUHT2Cx89a9O1WD1Qk4zNczAoHtrXgFQtp3Lhy1yga8yw5vOdj+a161MBZVyBdzl
hPnYMX9jlZ4BNh7CZc/C15ENfOTgJd+GdMJRfdwnTL7J1TrkINUd1/H6YUgPF2wh
Vc1zNfxji2o4+NmCghvmM3Yo+EgC0HvXaW9L7u39Nf5VGcA5xzktR/zCJpon+hBH
vVifz0rQoOGsDzCIYP+iWeIV2F6p1kM6+DHWjkzOiDUTv3xegYychsFlz9uC0A0f
dEsBkWq16hxkzRZSpI2UuW4OQPAa8uDTnvkQvDgv4LKOk6YaNhqZ/jCE8E7oowjl
4DyRlQJhw3x259QIw4qAwS5X1I5BbWpd0g2odcC9WwtFPHF/uFp419LnoLKP+PZC
n64IMq2QcxQMFqJzuW9XlwrmN6OP69TmbzK4d0WGVEksTAWs9uKEOCCRRgeGHbgM
M+V588T5gxvO4XiooYxt9PDMuL/qW7fGRh8TEXd6OaRQ7PlkdAuwwn3m1CoKF5Ab
0Q3Z81b0Bl5OpG1LFnCRwGxW+/QnTTprJGBucxPt5juk+qdKqImCWxJA3Qw9CtKS
Mir1hLvTuhxT0goEhegkerCtZ9hKrrLsJCj8XZD82+75FCw8LtsFSiqWlocvAPRP
EcT5bqsgPq0jMxsTuxw9/4+YM8VSQE/873RBILkqGeNJ9rLi0HwOBuCDa8crTRL/
tsfScsagZBlY2NvQkvl6/2KCHhMwFbFZCOU7tU7rSZMlYtH/ITFt0UUGuXis7Z3+
FgvLM5PoMWwJsZxWZj8DOTZQuv8Z2FH6N4H9zFy+/x8CS4HHV6YE2o7vBHi/iI30
qoEKuvvIjmwGXwAeEsO7QMxTV4QonjF4DIOoJQZwWrQl5I08JrTCJikM8XRc1EGy
7sgCvuZz5I30Tz2NpMQf4DEkUh4r23Nwm0QotUJQI8SEwrMxuXq9/yNWXLXbSb9Z
PChZICVO6ivYE0VV0jjPfzHmJZPIxzdIpj241d+1nSunzAPw3oOwXVdsUGsWgscy
7cs3yIJIDG55lSZgGbgpONzUrgtSQWI0+8odqk8n+FIsObhX7UM1rGW4QrIAv+1/
YlTtrUwpR/crhIie/Atnd+V6Nxqf82sdrI8xtyWEow+qSuCsqZp/PdXeCpb1NMUS
/976Y88XWdFeFj1SzxTZBwxl+KS4YQjKnL9h8HN2UB6RqNzsa/F/108bUCNd8xi7
cmFyqa28noAsHkfhUhwQ1XZ308BjSBMeE2fo8Nzsx1P6T/YEXIQvqsmqUDlOxpB0
pcSn+S8/KjB6Tty5TnQg9awmX1ztnHIKGPx0rKHmtTba0qw8JPSeNaUhx9fulWju
s/sdV4RMXPYojZCZ+mtTf2AtAMf8bZX+fmJqX8tqjOCTn9PceJ1Y46rMboOmp7ya
I/NsJjgLcaI2AL/Fxup0f6H2Dld8EvGfqwSdJ9omJk1ci6hnzUAxttJeE0qoIkX8
nLVoSvEg7wZSpPJFZhxmV40a98yO1f+IFKHSuxuUjO2ptzh6C31Zi92uj26Ur/VG
Qh91bAXES7Keaw6y5ldf+rolpGJlbOEdlUdml4HaDbzh+CYE2ShlhA2WCMfJazQW
xlgy2HDi57oTFHO79VTuMqrDC2oh4vOWp04M4ZYq387amZD20+7m0c0DuHym88gI
Zj3JKOfHkWteW8aNuTrsM/DXUqIDCVGpcf2EmYh91uo1tL1eHg4UB4l7b8Vg0vYN
3PHT7ktGkWqoxvBzV/G8mBtdhqzf7Sq8JkcjwHLMf4pOES7AZZbRPspLXNVSKdGW
NiwKZjGSGVWE/wItLD/FeCuW4BfhNqNV7OlBFHjFzgYpy00HhkIssPvH6f9Op4cq
GnLN6bJf4u3dLBc86AenYKsMGiAB5/BY06g0mfgDU9p0gM9/D8jEsH7iBRXnGjPY
5zkZd/m6MohxQhFWkkV6AANou6934PnpVayVhBqf2TOm2E6vY5rjpXG92AHbSz72
zeL6aaYpdw68CqNX/NcbBwdspEzJB8ZfQR6NAucIBkMqD4BCCsn+tCPmn5i7TGsG
8ygkSShglVRhNWnqphXzsIG3jX1jZ08mPijunbq5d4XUXE2r9svj5OgLZT/CBnru
DZleUXEILC4eUkE7i6EjFkT4e1i46i4nMM1spWVUIM3h6CSvYGNXENAaFv2jikWg
/zE65HC31Hz9/+4SkBBli0v52ghJZ1afB2HqPRX6ZdeZpHDWdSIs9yPew9L/wv9l
LhkOSZrcAyqa1DPmJdsseZEYw37QYQIWvspIq5BGm9rW5+Gd9Fs1AkOFZQWBb3YE
QtkSaTGfvNbabWGHudZaO2EDcCEpeAEUkmBi5934pXcigZSagM+IJ/K0mntKcU+0
fWd5rfGCPALrLoDMbSvzOzTKD9w6vwgb8loWSIfMaywvpvR7eNsEL39jXkQzJ6Z4
3WKYU/SEWHQYjWJ+zhWBjwb7Mi6QTt6f53PG+61EZ3v24YYhJLumaWLxLCNhPV6h
LFCqPTHtHKeI+DL/icG4LQ3fILjTGreIWOAhvlm3rHEXc03rbjvHPwl2gUDJ4HtM
GrFhxg4nl1F1Hz0sX9m6ZaAVNm0loBRW1POrM0KuJyas9GPB3sv+ruirScu+xIWW
CPT7mhXW8aL5+x5i45U8dChIxvzGBZ6QHfxGSs0w9IUL1RPH/Kk89j8ALZ+RhKJr
NawgLCFPUmixeJvd/+92xZhRLfGyLHkmWUerW9oH182xM1zuCiGF+isdOyFXUDOg
z5eDF6LpREc6P8gurv9EURB7hWYsK3uxKzvafD8zqRlZiinaNkTnyP9G1A55StEB
CeVgQoUAsgwiWAD3tSXiSuhv738C2Jg44nOrenHBXYtFVe1mxzW9nHkBacrnnQJY
oxvjdiZQLN6x5ZptUdcw/eUL2rQnY7wCiQp8I+yC100YL/WJWBSdA4FxYN1Yo07P
xs9b/gxhmS/9Kl8pM1Y6qqfbz1J06GZhez0j0/6f00XD1f8HUl07S9eUuOsdqZQh
czCvuN2Sd/yGzafuW2j4w3Cc5abheppPJQOXaGUhYH7WPmGOKlNGlfnRd+NbeedS
fAyvkgXvQb9owP11kDZHifefhp7c0dHBUKNwQvxe1vabp9kDtS5XHZ8dNwslJBk2
EgTA3CfJGGeRj7J1ewBPlcJjbRU/Aid6WYrSCcz9bAUNAERkHZ4ztHyjn7NRtxl0
jQmVMT6KY0+5HoiezsY5crRA63/RYjb/D7hpwQEWwjDUA+PdnSCUW94DLBWOE3jV
5HHYfMVj92yo5/QQximNTvuQL51FzpQQ+7aPrmsu1+jHyhkw4OLjeY2lL9TFoIfC
jeak8WBfK9TlxUu2nmjDDh9yt6a+9sDqTnfnqED1AGELP110QNARCQSq5JM5v87b
Euy6xgfhrOdatpRECKUnPPfDt0rr1FlRBfF/J+AD1sGSzToMfM5eR2pc7DdKMhVQ
CaoKRx0yxzyDUfVAQt+rpfmL111Y9lAG6a1utpuRgkenCTsAj14J8l0I3j0z8cSZ
VUk1G6NdbSQVK8GZZzgGc4IpuVyK07so/dgigCEho2hCW0hdMsOTfee16NnAuCP3
X2oBykG2J8udI7LcwVHmOGyghMlTiazGz0CYcHENMskcPmymZxaSsgFp8B0UJcGM
P/j/GYLV2IF9VHXyxwg9AfhDRLoOieUGPuYf5+qWfw6LXj8CGqRROf9O60K7fnmo
ROAjlKXxksjh9TtKdYLMSLkrLaJtKQlS4rvj/EDUzZcA6bA//MXQEZBO358vnT7h
dPX8Qy61Df5ZyZUc7WZaS1aD4MN3tO+b05lM07lJ1GB1QzWaru4THQVeJadf2sJO
GHBBjz5lcudWncZSQlJBM1DBqM6IEqMvunPx78DB1cjPb3tPk1dgZ3uTyUQ+VaLD
sUiAHsTiA20Gp7IbHJTfkaoov+6L8xNRgdNt863QXMFjaZno8RTWo74iW/LWa7Za
H/5PDIXenGtgS+jaJt/IowVg+eD/xpBJCxw+I1Qz1zSYuGMqe9q8kRC0tR8XAzpb
KPRaulUXF86rQRzQCeWHYJ19NuF1qv+itvjiM7Qc3tt6JzJE6gl2kUlgB9uQozlv
eY8NOUV+xiGu7wBo1jlT00UIfnzR2rmynAGwM/hgp1P3hu0ReP9XIwUWhRAx9NBU
kw0ItCU9eaDFQe8ZN5Xl6HH4wHUxZWuv/cZu2XS51HdtC6hCAYUIdY5WhP7C+JQt
lRj4vY+qZXbLouXc7rFUuDafIK9pTNlDE9zgrG2FBxrLjrIEW9HJO9xfcu/J2XZj
R7wg9TmDYC23rFeeK/PxTGN+A9x/5PQOC0D2DVVD41uShWj5CA1I5oVXiVi3rCsO
Tt4Qu7Y3+XAr+YTuCRNneR8MtjpnTXRfTxEV1EpaZWZvFuYje8WtVz8jXZv7FFSJ
gtPJOttE4sViMSTwjlpF1F1Jh3N+qXpDvujq9tiCG6bNQV24EOlLZNiRQuyWU3CY
2KmttJziCVt5pJHdDuul3/Zi9KjsXTqshwar7xV9+CS2Gy59Amw2C7ORhu/yvnaO
rLTiveLIFaXtMzZtigppF3Hnh756FB+R7RfZb6hl6mF7I0N9XUesyIcoz1kz4B2B
J03cQiwGAjLD9j/xdiSxEKIBRvx4hT3n8NwM/dHq4akFyAOn5z3m9WIuT2+dLk4T
0rAl10d7YPpLqqOMR4Y0KG3Iy4D/UHfpopdmwNHpCqRwx/9czkMmwDLAVMxxeu8H
HkhrL3iop2ZtdxGUZfJukYW10gDrV64PDySDWk5x8BdmjMFqrC8moLdNLZHGRqvj
HpC6hwTQBT52mus3RqlpgEBuDR1XBWBGpcUCnwys3r48To1hGAV6l3gwzJZM1olZ
eDOCwndR9mKae6olEq03NQfIMCEY+YRNL171Se/S/m6OexAATNHWF63lGvKr8tgB
if4wt9wgaQgZkaSN76T7jXr1NDjhwDieO1MkMn0ZRvUBtSQjRFgxEdvQd8+D4ZN1
QsHoXLxzE5SCsZGTAsKBPVEAbGpgdxtBB/newiYsa2rRnuoEo9L5Nq+4cFuRoae3
HMUKAI2P3X+df19vEkGNa2oUDEXqXS0T+JklC9e83JG7aY7kn6Lj9TRa+ppK6v8U
qSeXrmdrkF1a73AMcY1U9KDPpc1K808spLisigCJBhiF1BNFDS1CmolxJaj/CQQP
/GUiBf2RDcLiF67KYYK5RdzJ91y8+TF4OEmQ3DDVIYVeYmZ9MbPekVcUqTD0Xc/U
F4M63ZwiqHIlaGfwORD//L773mYKWyVhD2zISNA4G3LWdtXfNVdvRI6XGNNuEOb8
OODmie7YOjaDPWkEYsUrO+BLVM/GKB4mcTI5fVx9+9HsbL2mw3XzJGvG5dXxX9sl
4yGVm8KK+jMTW4x+hA5a6Jcc3yn2iXrcyxQNBzUn3RFxt+ROL9QwNuzHjFFBlbz7
w+YxC8jvh+sE4myWL4KnBfCprAPkELIjCVgfRoYGEgyJiosWggxVVWy/iVDMxOF8
T7m/rJi9Y7Q4hQsDRKsAYQ7n6BxFtHcXtoz1Exq9ZiMddSsi50lysAsxT75PcahQ
6IbsJgdEP+4NzcBD5ddx0mmbASl708lBRB3jNBCxxNjslj/SD+V8LhTNB6wKc9e9
okDBRHinw/dyrqHEUaDubITV9u6+d3Y73hOy9ooPzsHp9NhFSf4rxXL/Kk4nXsTr
S9TYM0iM5kKAAC68mbAmfCZPz3vnu2OIuDHWQeHZVuU0rO6OZD+jn96hbsl5gP4P
ifcfVV6E1LON0DX04hbpGJppXDc4esQ+yM9XaC/poQfD47Vlz/NJTpNCpBWMJ7rS
SaaC2ndDlOVQANiomtRVsOHEXRSMg5t1hlsaI9pZSB1OXEDotbCY9rWB6uw9te7M
yENRWhuodPILYtFtrbYZlh6YOUFkQcJcu3Dc8M3+G7HsVioBxOXfvtJJ7S0mSEjR
bsH/Yq6C/ae9o53dE6JVozpTUajeRkk8gmsRaYZx/OAWv219d+MXWuKRF5UrgV0Z
TVdZVMsl5Afm3pFIcrILMxb13a7Iq3X8RRP79RpDfra2+9PkZhwDFx6NmFgd1YoN
bUNYNx76V16wR4DNAv6VLlj0E70ZwywARHm6DXddWeiplEqn/Xyw9a9hxwKXuE6P
gewm8+JzkYgyr3P15NgisLmGhu/wgz6Tb7bkbYylTNtRAO3tUfbnPjna4TQtb68R
aqozkHVArVdrE1pc5k6wYNDEpE0ULpCDfvsOJ5TcaHGswwQAupEOH6dpzqAZ2etD
+xpDtqGgv8ti66GlVWNC8ULOXZBUQfQ+yRThFomPSafMdc5+V0k7BqcBVOMO7uwx
DlePP3LkuBxxpL5UOE9KMePwF/BE1pDhUZRTmZ6CK+o7Qpeylafbg3kKLgxYGs6W
Qk+s2pcqBzOLf2GbBY3T42+Ualjh0nQrThq1yBmKrwJ12oUOqwJxvnrPe5zVDC4c
rAl7t3rRDX8tamfimpC+C8HEaWhuQZCBN2vo7jGMpKMzjhZ3KYGh6g6DuSG52STV
OkxA7U3bgKQp1icQ4ELSCAS4p4zJW4kPNlj3SKvsWK95jBocSLcqFM0SyeplFxRd
183PMIR63G/cUWI+TjIjNUWZBhTo9At43YrJBdKT/XJjWzRHWL+Y+q7eTtLnFdPK
bUs4cYseHL6tPnPbsjupzf5rMWhkV7+c5si6qAAogdBunyfTZrMzt3VZaI1xCOUO
SBgRI2A559C/ALzB4svR2WnIgKuuLCnbKaFh9QC4iPv+woD1yOMmjbhh0K3GXMsP
L++ZWk4VYZr5Nhmyh20YMPEQdpWEzszPY1sTu+d5V5R+IHXPtOB1nIpRuancmZqC
OzSyi5JF6VAR0CwvFK1M0GyYNvVkHHp46SwDtQaJppgPB5dR8Yj7azEQKWCVRgFP
vZnVPFDzAE6ldLSNFk2jnj8lJ63AHIgIhrUKxYftOth8j6W/FfbctK5+YpoTzQDf
mWNqLPWt9w23KScY4bTWfgjj22LtVeqq+VbM0baM75tVwSiEPloHFDXQiMrJgBzx
vAB0KEv935XKOn5fg4LTZX19UEKz072aneWSA9bpt1uwdAqkcSb7e8WyOkdzxD9u
/VxcO9Vw67CE30HAqTD++JRYBxM/jWBavK8Vv8e1y8LpTv3i7/QMBqUMYtKmnkA+
h5YqtXjOcF8XHcJex7msVH/otT0R8jZ7VdcHPnF53pYRuOAei2bFxevOhHsM59jE
y/pTgZw75GqvQ4E7PODeP6l7wdWfKR3uy4SEY4afFF6MK6EPPX3D/I5oEQBD+ZNB
CV+BsPWvstPxMTJNOlxExMswPnrRxk98iY0H4GWLR32IEit9MqrLsmqBXziN/D4P
qeYSp5ai8qDrUpA/y0X/k5zRYny2fhfk04YK41hmkNTui8zWzenw66lG1PzANG6V
F/VboaNi1DP6DkbMv2QnMATO8mkdf9OSHCcYL5EhwhBN7djW8g1bcI5lgG4enEJz
dhKEAlfvo73FQNGfHjaeLpEmKVEsRabRp5LQAR32kOvEpEBo+xXw6ebY05LBmN3z
jZhw9sEOWN8i3XD4kHwaIboj8R5lHoz3nfVZv2PAEuhksbsZqA1ZEZsKd0J1M/j6
/j5ShJjaN9zkasNiLBLZhpkjArxPkvgzCrjBTsqeACD/FPYBbpuwv6insf+ncQ0T
adh+o+9nXiA4e5hNdIhbhwD7Hws0A9yCeFPE0UmcfBMsOAwAoSNoi5miReVUYpml
kM2nCd+/ahIunIccAu6rjaD+CYVnYG+iDubxEnn7AJG+DjmJDL5Y+hrodTo0GFbk
8MQ2nIHjO/dwH2YCvvxNO2ucI8QIUsHUSdabh9VkfMg6XJl/ko28DR/kAmT1gIJ+
OzMLgAlfPntzDRCSM1GDHQL8qYVUkpBxkBFmcGdOiUUl15CfItGVmvN0H607B6fz
z6qhNH6d0PQXcbKo0qeYN9fuc0BuHOycpreCRcDOLYc5RqqLc4oPYB8ae63wWYNr
YKO6QttL/PthdJVyq/I5E7ZAqFnJyBxQMDr/FuEQSD0vFYYU/WbTW01u0sxNx0zN
d7Zo3pzOjWvdg+srv0bS11Ak2f11GEVzn0DcXm8jEuFu2yxRRtGweVSWExhJRZIf
`protect END_PROTECTED
