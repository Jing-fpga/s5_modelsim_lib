`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w8NCIbLGD1f61FNlWwjKejuon7yjUO1q7TmRwEODb5pMNtraCB2TN394T+5+0RRz
JQR3br6Rj5Nzjuci3xnswnmMOBPGbCliPiEWo0uWZtWZJRdpDmgvYNBzLb4wfNXw
XIvjX8UL/2OIPZDLAN1v1xXec2cRfaAMF2g9XyxBunWMKU/EUUYn6/W5WiXlQ4A6
Hk+JnGc1RN2Ce5YSaq5aaRAIUscsnxNyfxM42avTg/rQ/+ZS6e6EouzD5Zc7lvu+
Xg+cm7brtnzaubOs2mCvgTS3fUtWhsgXu2ZuLEfq2HkHpxYIAPWo10dbDQDOXShn
syY3Od9gXHJaGtsAyBLfHpGhRD2y5yHmHD495f32kTW4SvLZoouHdm/2gGQ/4HTX
6cuIU5T8l+NMR6kutYS8qKwUP4C98sRS3C9MlXWv6zDf3mhUEGsmMyMABR14jTO4
onS7K3rGo3qoSsLQh1U6rXLOHz7XrRkW4OLumamYYW4Y20ISi6HffhbBb/at+oxF
YI2ZBpDR2eGK/pmFuSm6RHHX/VsSTgr8yuV4YsPj6D8/UpyWCTRjOvuZFnagfK8l
EqRP8j3/bGkAT/tr4v6LTK0udE9p357lEihC3iNuIHM2k41G+R3biRJVWBZCLC50
bkK8lbw4ZstA2YcfVRMtC/ZRqqIfjE0+NR9AlMzsoR4RUI36HQ/jtTpaVFtVUAqq
WLZi8DC8OWvJdwprz+lt85ZMmdj3Q80Op7Uw1xGCptTDDNqLHdWoTW9Dp0xRbmmk
wub/GxZqeZ4VFkREkk3BqyK4FXJPUfP6lJ586kowzBfoKbRPMh+HZm+PKoLYcN5R
uVVY/qInoZ/Es7FOro+pE1hKN3T/viOWAJmROTKrda7vr/J1Wdeqxzd9ULYNl1Mc
OSAS7LTbTISoAkFlVuKlEmcMZsAQBOYHt4kiXZQbIUxb6B1HiKuOZeHczzcVSGM5
PGXt4/aZz+ZqV9i8m1RCRaXqydukUECwhVnY0xr00Q5rJtgi2QeOO/LD2hOxmlfu
jOGtT2WvDufiI9b4HH0va25TgDXm2SjtSyHNHiLUBDqFl5p6GPf05D9K2GuLwl9u
ND7eztRZSNRfQkJ0dxi4/B8s1xUyC1YzhnAxvEiOZtn+7yaala2U+svcFRQ1zM1A
C/+oG18w+71yaMY/GUn+CqxztVgE/Ietw+KYReYmaDoW3KlfZTvLCAgt+Ci9rNlg
bInKaFipvzwYNQ1BgRW3qp7aiMSbuuAfj9K3jwtC/nU1Np8T8rfdtiQCZA3Lxm0I
Gq0rfkm0+g6IQ7shmdZbJedkZ2dl0uK9wwK2Jja3DA8PR6SORJaudgOToPb1Ske1
s/PdbC9k6kr+Y6fzyBDd9NZcg2DmKhpmR9lwu2QFu6ENfxXaEB2gzCwNn2pEYCMs
mG8ZY0ZOT2d0k5n3RG/5xP9YGQDaGpAExJ2HQM8I7fSer6JJNlNfzzLvS4wBLfnD
YH1pzsQtRJaRycgQEtEjUiiDWocSk0U++9Resw5vP9YjdOOmtQlFi3lrHFVjG0sF
6v2I4NNUED13cgQ02NtOj5TsjX6s+dJOA3yjO4/AfZtnJIPscTbosuQEh8ZRdm8I
ucNQiNY5NHJiLW0S2Z2KN9Ibfb6G1JYLgX9XrbGc9Xg2C8eNfVyt6LXfQ2ilypAV
nbBi1nkCp6pFElvZiVgklI6DlJQOoS+SmMe+v/tRn6WMb5ila62XgF/4ay2r5KZH
1Ft9RATHJIbpAlUFCTEEiGdjg7iPpFDybhzeKfqws/8C6gD3CHrTrWfFnxZzxo3b
zO1wfhvTRL09Z5a2WoiH51c/IlrL8t0quKbwpRtYT+JkjsThz2cQMBGfIsWo35Fp
JHe3C77Dg/uOVO41r2SAkQpCsqzXaGfswqtvNB9ow7tvvzgOKphpJWm1n+cvFN1x
t0Nh4xIpRTMOQHnLTkt8mD3xJnsFunFfM73DQgf5HQ/KjWIwuvJmkkfPsgdDQcYu
HIBMsvhJyfqFcltTpxJf4aCTB3i3T60D8s0fljUA52Tfhc27hm8blh3qMrRUO5vd
6kWJa0YYzrCX2CUMHM4KMr0f2h5KLD1L2YWzGthEC1I8GF7uhAFKy/fN02URCWYm
4Eh16KDpthlropsYtFLkz496Y676xMKUruZb6HxdNSs2Iy4JxlzPUuIJ4wLV76ew
m6f1yW4N/HlRUNMCz5eLHeiq0dW0SWwsb87db4ODpNxVKsbByQyUesjf5lThJ9Z1
xj9OVIehk2eRIAe1KQ2f8ptLUBOgZwwHlxQ103yaDZ3JZT0sW2eKeCFaLrSsshgA
bc59LxU1twrPMrJZe+L58A==
`protect END_PROTECTED
