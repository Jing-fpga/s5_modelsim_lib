`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ex32vjRNheukhNn1yxWT40l8EuDuQ/q/mmqAJH3hvlLZ7oloCQJhwMA/iaMrwGR
EBQxOsU3vpLHZmWJkJLy1RHBkNqx3ls8R0OzoADy7KBE42+yiJYQL3qnObY9wzp0
xA8k4HbVXspsLs0RZuoqvOpt1Ob3IIcyFDctRk2CBmq2JSbfgflFwU1X06LhqUi0
uuE4zWooGdQyhCEWMnSZdigABEOTcNYkqPp97Nz4CFkAmRx6ek40XjX+bwGbXzGW
q/LaUlhqTzCBohCz8CKXHRHFN8AwVdZkJtyL8M7h2WNUND4xS6f/xAhEkShByBr4
8qSth6sFSIMoj908mJaVnvFHTK+5Ea8EEPy4ycQJvLMt5s7CR6FmlBuwhvGT0XEr
2210XU7WXw4TbH9wDzy3jx4JBNeFt2/ky1BIPXMH7nDuKAYwn9AbqCXnUAHf2nDJ
DMqdE9m8yaf2PKEjmqX1P95odHh4Hpgia/TJDZtZDRKGfDfBW1cIa+U8kxgCDOhk
CxwfJIFpbPY1clVcweUW7cdh420HX2HcGXOHRxFEOL5ccdvR8+I1UUGrhTKlmnFH
jqfMgFFNb+HP+mP7Et9iJJtNX5kZIz8btAOu6ozynzLqKvn+cnfVW76igltrCTtF
L6GsNuVwhIq6rc+i3rw/biqqmozak+0LyZL1PaQNAZaF+sjxEGXnA7o19hQrT1nR
YI2pf95OMRF2aTC6zAggYX/C9raDL0lBfFgFbEB0c81aASPzA4JdV2lz6yT51RbU
PSl6gNhSPoIWtWGc+zzog0bc2B65fHg4jpxMv6Fwn4LTBy8/uPGbpdPjVzCZjbCk
Th/jMp8PDbGB8pMJ5NgCWFrLHcKcUlb9qtr4Wu4Em5vH5kH0NLUtD7kJzNCPjwL8
mcj1QYD2rjJQlhFKbvvlBNslnnMbSCMi3PVFHbhl51vXVloygk+JFbpkd1AMVLGD
92i9u1c+HBsn2vI6/9ui/6fk/Vzs0v4DByIOn97ydRgQ8XJACNpMXx1FAvTBnR81
J9VJsHyNOQu8tNZQlk6vTllYKg94/bRjsxEhSaqa5n4pn+81TYRAiUUDdVpKhFcm
g3PNjh3hNd9B9B/ZXLm6hnXDuY7HsjlgBLeLtEx/qeEMWwVEIiOYaYC0cf7A8eiz
zA8W9ujeFGXKwmUHJaWMEl59EPDTKd8OfoQm9nDv2tgQeT+DGtJVrgZ9Vn3sB0CS
kl3wZJz8pxxVbLICw1nNaghGnMLFMWZo363Hd7dJtpZKYFB+mLqQ+JbfmmrHf9nL
FmeLVRKNgKomYryutOLmYcYvn+5HI7R0sbB9yUxCC9slvAemz8YspWaDtj2RLbaq
4oyvbTimcjj2hHaSNC+tV9PnXJF2W5xH7vo1R/0IDm0ntOYj4FsqGZDYm4vEUZiA
`protect END_PROTECTED
