`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OHoj2ycet0SzCgST869Bw67snyojCU9/BpWi4MmCtoKBOhZGOUYxG8ftsTov1rIq
SWB9MdwJIixEmLrMDV5PjA3PY7TpPaYNlVz5rWGO9buhMGMTLC8BFO0deOmhJ8qn
IIfGlV/TANS/b49t0Z8sGqL8rnRNix/tujLQDi/B+gYjFYw1a9x9oi5m4m7LeEhv
YcDrYjhVdnib7t+4nmVJCnAoy2Yd/StPxZiFvFDiGhChtXL2LOZ1hWCGB7hPGenJ
pv0YwjN5If1qWaX9+5ni8Ph6q8nL6Xkw9OjVyVMdhh2vaV1rvmROEDxJ7EfXthYr
Y/xdd4t7yN3Di91HPcAE1FX0DGI7pnxZXoxM8Svpk1uZS8YS/n81h/PBy2+knUdk
QaFX4ctci7ddyNThBkfMxhfmAX4/OjbRWbBtiC+AUFQuKlcj077ntO9LzWtgym56
hO9HnlMzMOkq5VqoGW6BwdtkVZNrGEOJYKyPFdl+NgFxLgkKMtYHzk4Q1UmnDF2K
sK8KRzLsgzvorS3XG3u0tQNkvGTf0Nkw9sDuS6xuM3lHn2eNuV19kab4kiPos/GF
TyahvZF4KgDKOAoa/3RYPphCN3imUKNxg8IsV6mjpWwdPh+02gONA3BHSM1X4872
l7+oU3hp8qAsohq7gWAOdPSvhbWc1GLS1qrAulYsdcyrvmjlwmRxGmMKtctvWVwh
gGHJq5v2hP3i25P10kap4A8EpnBXsWMxmm2yXh1WrKPADuWgeJZ/QBuQUPknp7cR
oHWt7HvcDpqJQKBhZWyF8HUCXik7wrHwxUn9z232OmyyhTQGEsdU7UT/Q7fiYi2P
KvsUzfXamqw6yyebV4El6zYe3FyTM/oTltbISApy3v9Ja68kp9r+4KAaKK8hOR7J
2WyvuPyumNlJCFxL7EoGn8vmCsAJ9l2oNtUgF7y1hN65DD7MWNzI7XxIbuWqLh9E
FRbr/VU2rPwC+jSkzheDFA2KcU+6eKxOWEvLdtvPUR1om+lNXbrf6fx0xnvYKNs4
zX2of9yQ6wqCzhs15pbXDe9xfjauqJ3PE/74ZfrPCEI+yntud3n7sQYTB3QxOLKw
gJ9y+PKO+eJpPosUdHybLjPgG2UiZj8oGHsOowUENjEIYejV1fPRzzcSlIG3RiMT
reajK5c9E/SxrINbA0757dXoZSIIhVncOG0RaY7ciwRJxc6EeAdBvTi+OKZIar8P
dUbxaQyIA397oSMGMJHxyZszXocIxtx/c7WxSnq4sQ8ISPte6JH5zK4hOfpwE45u
RvmsvcE48sWnXFy1Ums/M54W7LRw7uvL4KCS3dsdk+DR6nQI81HIGk6OkPeLLy6t
XeQFhR56kV7eSjGulj+atiQjJcnwUh1ZC+K2pnX3im4Ihq57iy/etY6rXLgrZmHV
fBE7xNP0YnOCahU1W/SZlQfOHdnakDgDphipKgMagkUxtrBvcopxOVV509RJmuGw
v0eKO7xp8jhQY71nz89LFipvQXwZgxnHQ+Ja6DrbOrghlftJJiVO9tOyTa2P8z3h
DFKT9Bh4zILr8zV6tKJcZX3NwLy6Y+4jnEuadyfgUALuvBKtGylpXNLjZNNQR3jz
ymUFbEsuPTFKHQIaoh9zkQ1wq3VKtaH7X2uRUI3OmlDgrxtwXvLgwGktIjUNwd84
VvZKUGadTz23j5j9wmRYuuK05vVZisPkuMzg3tZ6r1ENQ4ewUnINCH/lsYocCMNa
xErJ4daxgtqCSYwrNTLSEl0QC6ZdqZRbKUwGpF/eS9Vaoj/lSJsTsN/ihwt/4/VP
7KfjadVyoJEW9LvTUkWoY5WMEZ5XR5DNb46cEIHAW5af6WnyEkXFe72wmdiE0hEP
06jYgWJvfD8goSWiSfF7AXmNKiP9K54F7+0wiFP0sVeaftcXwcge+piKtdhrv/AQ
KKfpEKPjYr42rRiql6gjgjlRvEmKlhDdsv/xi0noSRkgKbghQ1RAhLq9OJlTetWM
FBZkOC31/ffoChYDWbvtqXrFlpRH86IQAzXcf6hu8sTQ+9Wp+EzwDJS9Ur4UzSSi
6GLHQThTwvlct+5Xe6e+q81fFJazvRamrEdw51zXm6vZUTFZChJgc2BxpOcyP6u0
W1esRGBWPKWEPHcgHflyfRcwBisXBrOJYUNkL4uUb7rVpWYr4ATEeVGcdNS+rtwz
gORrKPj/aMGNn5caTM/9inkMi9iefuYfjgUP/CzuA/vwiOSMQRzqQFL9PJCI5Bxg
RNqWeWSLSqbteraOke/9MyFdexqHcnposBhESnYuW6nYyK8CReUmFH10SbjZZHIy
sPtzx3fkBZrsMyYZOPmUqonAxvU/WWiCg31kAWP0vh+jX2sc1ATrAQJuPl4KPUiY
xcm8t8Hzos+MPdyglEihDsAApxm9wjfVd2pbbPRH39kkuM+PHkpcSSaGX+/K7+kY
CJe2MbvgEDOZzjWIu1cEonH5WOfhgl1JbKZOn+aqEpTZjr5Yy8YN44enGHQogOkH
ZIcezcPClRSvx84fFA1fn5pEZaMnwtHKDnjKCD1Iz0l7ZVi90g4A3r83FUMTvXBN
SO7mxstLiXFfXkV1gbND3mDMlH3wzUjCFepEgWz6wm4s/Rr6biuL/fYpjL6QdEjv
burwIFKK2KkNcpOzFhvnvFzws8F8FM8e4IncwbIdJb0p7ewmPr+ZhE/7+ZVu44wz
wh9b42xIJ+OInuvDKcqHTYnAfBo+ZHtAkFZL1NtdVkbGLMJMiFB1ALYg8asC1Gq/
W5s0FQiP0wpNlK5YpsDhBw41KuPNh5wx02JI2lBM7MB7IODH5x4FkuOxlrPq/R4O
9raFAR2EpwnK4Zv8sF5TiLw3le+APr1oq2i0gEKHwZbXJnjd5G56+G2mYg1YwCrC
RWafvJk9nwk39wj8Vf9pNgHaJgiMfoS/Qa9utddkVegkVmZ+R4PfH7VPjQ2UepkJ
vbewy/MJ9hz8+bHO7SAesuRPoQp6AVBewkovvGVdu6GJ8MiS597B6BYvVJC1KcaZ
oGHh2H2HHud5brnAkBbIDtoCNah2egBzpy1DcjCNTjFR6YiE1U6IlW960oDQcJIb
/SXGyNZrQO2/2BH8B7sqYctAZBxbm9CY3MY0E4G0mb1zudpBiTRrOvMyeY4aNdYF
sChKfX89m7MAH/UW20nPDbRBCsaUrdnJ9QFZXn6w0GRmTmRqxOcXNfl4KT63/HT1
Yae/ER4DnQXV2ICzOcjTPdqIDQgxk6jZ1xmakRs6kT+g+adlztukIyND9jxxm6HB
dj/fuMHZLkuWpvpiDA7WSamJVxKJT6BtgdgXdYsYq/USjIRImVvSGNoBMJ4MlHxz
/myCn8FqER4k8QTfl2p63pRSnUPVc/tnt0e4FzBvnonMHFFJlCHekBFq9VeGF3P/
M8G3iwyIG1/AxE9LhOVDaFj/sNkYpcg2zQLB7lsK+/udGTXYi4JWZiJvIG2V5WSa
8KlwhPoDMxz9cNh6wC2zHcAQ+rvYrsDcN/AxCtNYTfHBbMK7SvYXSUtxCVfRPIw8
udYSnMuxjfaoJJ4dIMn0qXN/N7EGKKKt9KSzMiZtlBhE7oAJvmC35Ah8Qdttpar3
FpIHI1zNtcORcHWo4NbF0093ovV1ZAC0RBAIdmvfy6hRqUath8IQfcGDYghJFAVP
GLml5zouhhFpSYhk/sZzvM2OA5t6QuEiNUlEi+OGgCrqteNeEbZVu25QTZNYMIkr
3iD/V64ZKbwVJDmgoMEJAHv8PoEVKSBiaDNsi6KPT7tDVLY47tCWyabkhXTDFkY8
V7DNxdwpo9HLL/0k/TsRjZ8b3uv2wMU/k5+mvugMSpyCD3yS/RIR/QvSuhBiUpLA
mopupiT38K6NCekn3vaiIADZFSZw3DuPxxwx4w5d0v/OAD9KdJHPmV8l4As8wgmg
UILT001aVu3fe7lhutlCrVhzf2M4kmvvbN52Egw7TkwINs//+gu4vyqVPvRDq4Im
fgKgZasz1Xp48d7EpUcmlIase+VBy5dKzyp9EdzcBW6TbrfjSr8ArMO2gK5flUGS
uEy5S/+VeZexjAgTwwxVOzg6FjScktlK/Z57vpQWew97eBGq13U3hgefeKD2Px4q
awsZUgjf+Kt7hB0jzsXbEhSgy8LS9h0ECT+TyZb1nSmKjOnslpSme3Yf4Stz+ltn
DMFgvoJ9o6OvqGpNsshKlNRtnX5FIREd1pjk421TKmSgQsycALa2xk4PE+RXrH7Q
djGba6vFEBdtKK/jJe9vV3tpUPnZFKKBPl81znElbluKhqk0EP9ab70UXajq+bOz
3Ur4N+AIv/0hUpsToVOZTV3mzEuhvAC9rDoIyUDfcRSSJG/1JJsdaT3dC/qais2a
1dAbEvlq43ScH8d6VBxqpRG5OJ3pgSvbojdAwiJW9TEpa1P0J7/CJw5QSrFuaO0k
wGWVLp1KUkMaK92NqtlhcMp96UepApuCccP6KwbHVmUR2T4G6QxMTOMQ4sytZw9b
K8ycDHp/S+8Dk/Vd6fablQ84Rn9+BtxI4rfuHxCC/q1NavCaScYoqW8B7d33Vp4b
NIu+cjWqGPZTk29BECY/xizNLEVu0n86BSICCNEU5yLOFctflYvDQ4ykKaJCK7LH
svxxnXCua28N0K0cq3STo7ULL6DBdf6XbzoSEu3gNVDVNbDIVWXJTOvgp70V7IgB
GFSXQ/d+/VQjfj30yTMBNGKMqfhyuCFuvRZadT9n+w4N9zyveEEV7ptueDWUVSLQ
QZqxg3oRtFVb5xEv96PmYCsoTGhY7a4snJ4c/vLMYFUgRf9RXEAiOTC/85+1vKzt
X8JpRGB4ZQ8HClZGKlne2gbbWvioHt33Uhi9+opPg4FwAnIq+WT0ARex0F0PpO2q
DEF27D2Yku6RIB2dTzRiV1ZnAmzM4yUEdV6GQJWMHm7VkCd1LHvpmSXzMaCPgsKG
ieNb8XW1EmoECpwI4YYIQybw87u2guwz8JLE+RjUny6HHGWUb7WHV4FotrWWYUO+
poRlp12VWlmcMeJd5/O1zCISIOShJ/dHjZVKVOrc1S5FKYEJFt/A1ft4gzoDWXKL
fxKqOUA/56k/HgKeStW2H+x3Cy95sRyb4lPTGAP1lt8iswkEIoQsGUtXmLWdSHFX
gFll1vNg+pW6nerTTTPWwwM5I+PZHR7BPX5szZGXaKLBltshsfv1dCGKyWlKviPw
0N5CgNfCjx5+8atkacyfo6GaBqUDrw1RhxFcVmQvVD1f6uHxf2UXbPHzsq3IxqrX
lzlwflYkUYHIXBDpiAUJ+09/HEruUwNQdRCILT0y3ODbX1Tx7FOKfzXmKOXKBugc
sl4XQsCsk11VAGEKMQhTLakOixRZO2fA799Mu6saZa9bS0sWtGsCLAnYfPdS05IX
Yb6k4qTDyo88l8zXSJ7cBYquNo5FOn/VgbxQRmVtD/bCtKPxIWYKpQ2hRFp0Y7xj
rILcjG/afR/W8KEjVgTaqgbbiLuczBnb8xyiAHmoBSskR2kEM9VzwhCFGtL7vY9u
ztFAZgo+PedqDyCZ2RMUaIzx/56teFzVoCJ/sRqVJJHzXRK8KdL14W4dv+F6dD63
3RQ529w6wXaVqJudS4VOAEgxyzb/qroncUydBy5YsF4Kl8HtRqPvpboNd9+h1zpu
nKHCOnj7HldenjKvJu/x2cqJFcDVdECLzFla4+PWdAWvjEGlZkjubiSyFhnwLNyi
oWX3acAzOzNaenjbQPWnrYEq7c79Nt0TARZ2dg7GoEJmWRtUcjs2ag5QTP1JxD8F
f7AH8GZnEG5IqQQzTDyCO1lwSTOy3rR8cyabFvaRBb6/bajI2gc6wAGHKWBzG0oz
`protect END_PROTECTED
