`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nxQq9MTG+iINso0LBYQqXJX1IMi8HIWFd/ah+tu18CPE7Ijl4vWPoFcq2I7fKtYQ
jtuAanEvnxN7OviDYY9nLl6lbydlbWVmp6vbSrvkIiMj4W+U2zcOMv4lihwg3P17
zRf7B87QmGclbla73IziNciFkBh0l/Xg/kV9SeZ4FTUZe1HJkK+9Ot7mG6SKr4K7
dBumZ/mCIeXTDsjJWEG/9pWpxXSRz13ftc6V4l1cQxec+eWQxmhkzH5zcWLPCWRh
NJUjjhJrvxKuwNQ+R9bQHBI1Z4+P7ELy0eACjjMu29/uNcBj0+kug8GdLZDAPT20
q5sMzx2XZ/QPp1J6A1ZQguXGqAlV5xvuMOhbbixUN0J/eVN0IO0jQ0M8MpBBDzeT
ltrseo4dlwpIM4vmVgRtJznw0zZePwFfzXnsL/fujGO/ADefWMADrvNLOI0vFpfb
okDrETUIP3lq29zTNuEbSv8uHn+EX6UFOrII4h3TguMVYsUjQMjN4T3n5T/vyr7l
ZnEZ4UEoHVmt++3zSdu+6JXYTHqaPo2pQOXqz/P1tOUawETGts4yAYRsipORFRPt
uuIiqZ9yUGiTPvHGCZ1jIs/A8M2eKVG+cgJY3nXfGEfhF6J1t4rGWdW561bLRdnJ
K9hwlnL4xcFoqbe2CpGcG+5b+kMOGoFrUVAGLztkoJRZkghILKbrUawvlg8p48us
zv3hEixhnksl1eUN0fqAblU6eINs72Bizagy2puRPrguOQCRlyy0jnbUIcBxDld5
KaLkcH4GBWzCAqHyc2VzCTwa3kECGaJunzCA8trP4sVVJndjPzgm7tvXhgsop4i4
fc++srbfl5E+7DLFA8pUNqNXVFkal5DIOLKqUD3lbGyzRKoxJxFFQ2cmK5ZlGLC3
6acWpCynqwKktZx2R4rPMvZ+xg1pVAWkq/BUG5kDHZHbwa3QGaP5aa7aIVGFFXty
8NynmcOkpFSd9+9MGROOmZSqS2lnsmnCLR3r36sde8zO9W/EyjIVk4EZmaoL6yn9
IXVBU8BgFJ2avB+oMj2FKYMyiHpRZkNU9K271SFG0tIHKGAbNHfXIuGA7FP17RKi
OyOTG1jWmi6JgKM6Rr+tXyeVad2YzqwSJEKuhhusUGZOy85E+ZzCNQwhA+k5cCLQ
/RARjOB+xVRBMrlwJbQ7MFpQBHfm5fVWKBrHoCAn00yKQ+POx+BXqyp3ao7lLMnT
qEqY/88hfk4HbFsArNU0SBbewqrEJfW1Dy+WmbYfZSlQHdURKX3tUZ00C8dAFWaq
V7LvngMnWsp5xN4TKunxDVJvaDjDRmk+mPzM35tpGExfdilCwzXxtkIgh8BSNWz6
c/cNpkTcjCAcU/Wrrn92gvpGfZxuamrxIAU3cBwYnQn25t9p02C5tJhMJT6z3gsg
pSCMEdNp/YiIkOytZ2Ebld6ycM4mrkPLw1akQ309VNwA/jOTGSYLMEs2IPqQbetO
TzM2I+/nhrUIjzzEQvUXXZWkN6fqJEU/QPvI6LHmWgTb3LABc1d694Q4kx5XuGcU
/EjfvckzoWG4MfuXMiTjrhE+4yjzpDLTXemiA9rnF5kKROsKE39/HDyFNj+L9beP
Q16//72ZX8vqVM2gn+ycwMFUBJ1+r7kfotykOhLkX++aj8u2o2yV2mbkmWLv3dCJ
uTqNH92ZKi8P4Li7PxYGnnq3jlzPfmn/xblLUvOm4GXWlmPwEwCS3S/TTr2+7LLC
f9OGaqrOUfNkqiKPOfhcsqAQDQZFrfWZKCU0SMp/ori3YXiZl4K2XnZrgyX1mVFZ
/sXONrnEswCIsoBumb6zf9FSxP+xOSRs1YEMbGuK8v2KUS0aK0N4sJsZOhr94un5
JDTxe2VhrEWZQttK+cQkf82Yr248UTGpsif6w31xIU0M2MS8e2Ck3/Of56QddMNF
wC8MewvowU7fx7QMj35DqsrS4O3PpCNL/CmnkRrkxxYmsyHCYbcSBRLE3HXdOX3p
8/5ca6BYMrsv+hs7JLfBAuH4Hr/42gn7eKbFphvUSz+ecFk81Rq+/EUgGMGVASbz
05LkKGSCptJZVx2I8l9nNX7aoSJj9TRXdQeTsoTPqC/uKMw4KxuaTjEz4MF/9xPP
mcW3uxhqkdhz4t7523fy8aBMrZjXhF3vWXJiAq6GJ4+9wrKgPrcEf/PxMYvgGNbV
Sv8Xi0gdX8ulc+5CjdtBybTzVlbASNOOxacZVuZymM2jwgD/t4KycfxGORS2sbL8
0jCZyVY5AB8Df2NyP0383nLlAqAzsutHA9qyfeI/3vpCGcJ6hE51GsHtGAFFb0Ti
DBO9DUAOMb0TFNWjA6Kv6/tOGgi29KfKMwRmoS8gjHCa3rdJdjJEuceyn06wiCxY
DxCSnlYXPWBV6lCji2a6jO8upqv8sA0ZCkYNQd0kDSbS8RQ7kW0uG0qdLzY0u9Rr
lVHNOFbaZy0oYhcZs53QCyOQJkvSauPtg7YyOdLN/K2+saLIVFvZ1Nb9o8y3uNpk
JBvF01nTvKojbAmu/4SGY3C+nua46/N/3KQxtkJgDFG/adukVNtS58811Ev1xVIg
3JgmjqOh7FcNkMFpvzCK5nO0J7EPLiJRhQ4oFMRWXlFguOKsb9O39oU7ZTpZdeYg
zLSUkdfTH/3icMr1Ey3z8TY30Hvk4ibI/3ySo2Mh8ky1LOcDsft/33a3diBsnse2
CrreedwLv/lqs0Qmb+J+ehX4sfyUYzoC7zi34jHRdl3W3wxju1d7yv6oh1mxPBOe
dNIfq9U5yJ5VMdIC4nYVgT38OC2jRockpA06t4S74U7YubivDzetUzTXAi1BvYT/
fqj3/R2Ckgo/3OQ+qNtrU1hcapoTXcvX8Fk4hTqqA/MIKsNGLnlJriLqkb40z6/n
Ve0Y1Ir7AF1ObchR5kEPQ7eOZFCJbPZJAZzn8TxkT2TKJdHpSfZd8lVSGqGF/23P
xRYKrW67qgXRQP7E/c/l640OMhRcGvXZRi0H5Q/Zu9e0j0BJxYT90/Ev237Y9v3O
WOXaUxIvdvTOThV3NM5FrWq7z56tLx7d684ITo6VXLk/pM6llwpTwTQMPvhQ4Tu2
f40XKAtG1G+CiqhTVuoiASlpFFAUHBGCqEmkR2vnI36f+3DSWInA6DplAPErhJFd
gxLGseqxKvDHZNHlAJlOcyI2ggCmocfc+ZwNy023q/7TSLWalnd1F242z1S+YPnG
PWu1TNwU5Hu10f36EKnbgnTEac302O8kN1jxxH15DXESNN1EHRWcxYU/vnt6/4Ju
TMCzFob2RS2pul/BGrK067wOriNWKSM7v4ISp+wLamynF5OlbCOXuU8c5JAB8vgJ
ajZPd7mtyMIsmPaOBlXMMw/Ks7YtdiHTfb4LJCigOC6lrZdJaahs+Csqs+jitk/x
uPJG2JCIPiOa8HNJjpcpMTTb9IpjgV00iqL97o34CUWwcZ3T6Tp2U5VqMviHJkSs
ynqRxqrJnGPvcmcw9IlXavPfYPK9BuklqJsiXy4KAv2jJU4l0vk8/BtiBdhgnbB9
qL2/E1Nz03OTJS1M0gdA0t3vFKBEM88grrkzUfOQ0CrEslB72+1uvzU25XeayjDt
y12qtE3jeTm+KMNHr1PvBhJWvkCVIRb0mlYJXPqR+FX0Ha2O6dIVDRdorPYwp3BF
nOShQnADw2/OqISZ8kwUaVmDe2IaTNP+o/LqDLDdTCplNetdCJlq2mDM9E1HdZWr
6jpeBq2ItemtofaRfZCWCb98CVVtitqjZNpy8EcSE2yAC9xHu3YKU8/nYB+gBlcY
YtL5BR4IA3USR477FUIkGct72e+7TpeSv0YAQswKNJNY7MJFI5hrXlLe2xGd57o0
Rzb9ec72OlVIPekXhDWrS2dBiC5prb8xh7gl0AS/SOHjUNa+uZsVE6Db80IYUweX
jON9l/divV9W2lPNhyqWupl+ZFDY7dgLPqpdneUrWARaHQv0XEARZkeagV8ysyul
X/h8JEQbjTRY7YGWqGK7+9DZ3JFcLEoP02rnAfkPCW9ieP7o+sayXzJ/99zVlo4R
NZXYysYfMLk0vhNhm08p0WC5GHne3lfVNVUgzFzQikmUaIcct9bWeNCP7kFmZ3Mn
qlAOHHVFgMTn3kDv7NK2PmOIE9xOpPpZMoLkhGbii4gScFyw4Fl+7dibWQt1ehaL
Phn6fOPPEB0hwPKvPZuiByf+llki2z9mEePqknncVIaTbt3IfVb4hX4NjCfnyfF8
HNDVYzfG+h+tnADpZdv5D1Jru85C9tsEp9JBRMuaVyBZNHHwcZO9hsErkqam9HsF
iGsSMP3MCYJOvpDknVfr3LwBcoOFfrJH87Y8X9vKSxk66UeP9lzHmqoh/kCH0a/A
H60JhRpXGX1fg54QbV9BaQ9LpldsuKCfT0INZDlsU5gcV6Ozp8tpUjBVVF057zJX
euAKAW1/Rp8Br5no5ovfgh4vhDOmWPk7z3TS9iGmheG9Lqvj4nPKVtwHmYojLQ5E
gxkqUjA2Me52K+hZQgKAPxoFMXXU/XyAcZk+fZN/sjGcgv9Y5iDCgS8GkTG5TTBw
V4SDhRR1h4CyDPsOM6++ba6aOYR0ta45fl7mzJdwLp7qL4hq1V3ou7usXcYZj721
OsWqFosLn3UA7VeLfGRctGhV/Z3z3joJ13ZUYNlAE+AkqoFfOZ8J2rIa+MQfRWq0
7CgTFReoA2sUiQFOi+VtbVsDKPy4HZfTxYRYhZKfcAIR3zfT4FEeCburVIILMPda
nnZs7ZhZEfiS/QfTIbMvUJFOM2c0JlKNKR4goqfgL+1Jf9g0C3lc7RCZeV4q2x4H
1xIUJMaPBUautCLoaYBpXGG6tBFmg70ciLhpjaEujOPV0d8msxI9Jgj4aIp0XJNF
1l9QIcvnevWwOFn2QxlAriFJ14dkTZVVLX95Sci6M1NiMIWdRLd8yNT/pm8rcwLg
8i3wzwWH1mrFvt6m5A2Q8eHXIuD5F4xORfLRM4gKBF+nxGsNZ5KSB9T8KpMzAfls
u/2adrT7Fuw2tXqhEij9Wkf5BCNBqrMEL5ZQXi3kavLsej3CLM1BK3dLVJFabaIm
WG0RONPEUBLoGsOGuwBNCgJ+3Tg3TeobSNFd7TBBXkJVKyX3FoBTecM1OU57Z6t0
HEb3sxghjyfQZFmNtQcyk8D/dtwv4xDXkPo6h/eWsaT8VfVjrcd0bkVrbyOQg9Q8
rNwwCicg4t3kfJ/GB/YQWDjXp8nFlUeHNAeiZzFsoi4dH5+N9xbhLWgM+KTl/nbj
SY8ogYQAK7ztJpMDc59kKXOmJykEpLYZIc6wF/nu9p7kN7m2At5JkLekhkmiAIU5
wgliqVgKfM9bxd6zAzfWLh/oWDuNlDysq7BXGZhe87Gex6EEqko+zZlGLJZFhV41
WX+5aOL2wHVEjPjYZrlgrcCX32CXTCozLpaM0yKMroJGwaG+0f3S0N8UXaNI1htB
uonMZsb/a1w6A+4qVX7UJ2D8X8yFmnE9yMV8cmzoL0pgQ+FM8EAcikoY2g6J/DCF
JIwrAfkdXTA31J5m3L9N33axtwZ3iYrJTjIzA0zhCYxHmFI7YzpHgR42q4It5hOR
MgXJxscV/vwLOA03ON8843qDFO7zg9V9906S/kuso+MxwZG+Kg7bb0FAFEAHLCqd
6XxVHu+yixziI8O1dqbeK5lHb4REQSd6HhQxFRfaESLE7Rvvc6Z6fF2eAcGHJbOY
oCkHXCBY+0rP9lP/d8g1e5eBiJ65tZcyTyzcLefrxVdeqPGmP0nHod1WFjKg/H41
jYkB0Y34CH+1htBZT33IKudbqy20XBmF4/88YVWkJyM9CccR4UlyfNPE/HVSTn3k
O1Kdv3ExJSL75q1baCRQpvuP2tjafYCPzmGJ+EPW596ql+EAiaf0tMrbhziZmxWa
kSnmTX0NQcwhq/MtsNWH0pBHaare25/CCB4JRVUj7pfKjoLluyb5pk2PnB1toMkI
6+UJYR1c3oTY4Xl78l9xtc5cLv1DG2rTXDIZVw00CR2964mCWSb17q/wz0WqJ4yl
wrmlsaKrGTDCDprVESxZQBsxGBns1sWp6pIlh6wy/cUW6wkon81kiF4y+mGRPl12
FxjNzLIqlMdzdw6JRQ35hwSaemo8Xtf6jG2uBISp/gANaf3PmDzOMWUa2DDqbEfw
hp43cw220Ibuk+fCNdRwZDJmRVfLfcA1apUEj4PHXsGYtinrjKGfWv+fjUaC4NTY
k/ttUtrFDvibd4V1NdMr3ES2kNulH6LV2RyEH6280TZLjADvzwmg7AWXU1IOwYaM
MDwnUB0Y2El5P+X2dTD5ry0Q3bPj8lezgvbEnRGEoX4ccykFmy303ILN5VsQosRZ
7LQFyFAWhGhQGP8qmp2lu0mtav9ds2LtUggvOjdlf41l6h8+FYncgLfADpz4E9v+
dhVTjcmcSHBOZJavJxiNIkXZALg5jLyrgzWc0/MmHq1p5n66iY1Jb+Mpbs0SdFgM
PYEp9ZGaaHAkQTeZNvFHvB3mNFWA1aO5eoNYM06miEZXxTiATdon1FQnopQ5tybr
XGv3aWo9fRsJsqSex0A8Tngo7Gi7cHNNVPi0T7WajiKOxmg68Dyeq0wEi5i6dBsB
FORxNKEaaXzsUmMkIy4BhEm6RMLgX/S2+GV63jYKolnTll4QZNbCFxUx5MCEVHTF
XRs6d+I3V4H/vhf1tst0m0ojQbFmD8e3IioYUS3vFq3tygDcH1IE9HT8Eoam9sWA
TgE7z839kQpk25SiYbHJ+9/yexHxutKue51nCQPGuccPczP6YHpSmYL02POaFZkm
bCC5YzhPbfMjWrFvQYqgdwKH1YscKRTaURnZzaK3pm7Ue7/XNr/d4tpIja4onQbO
n5PPgMW3oRP4sqlJyJAHE4ucc0JjCDWwhNFIJEXEJg3qd4VKsmgO2VqcBIGgAP7A
`protect END_PROTECTED
