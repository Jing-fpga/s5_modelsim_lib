`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eGS0gGO5fElaxieWc8jvO/XLvYQ6frbKUXTabELZPea7axf1AwPfcRj/bfnarAuO
yxLnjBJFg5YCpxCzpmRJ3txq0xhdMB5Xqm8iYxisf5Ne2M1vQrgoqQ+/TXKTna6n
zbTvh2hV0OhhyCG3uGAot1ZN38ns7OkWz5zwEZrq5yLu/A8UihdeaRP+f7E+7NvV
5n7V6w/f+RFd5ZNWNG29SxUWmSfjyFJm2tDsrO1NvgShxmqcULEc/N1RTS28fCp0
HDGnoRtF+UdTS1MwzZyxz/1JP0HqsyYiq1ylsJgiCCEiU/WPHmuxbBswGUOtRMc6
ZTDnJ1j5R6rYC/nvJVVCoWamIBbRRi+qfDCm5OxfBOcaCgA1sJXcMWccK/5g7Q8A
3P6gDlj/p5saJXGbr1jvx0KErp9WlGvuRFxJkfgKErfs/EViZMViYtzWXYz+h3p9
9NhDrY5eOeD85wfkFYBgtxmsmSM/UqpotisXQaPy+cwVfXOer35Dic0S/XxV3FEw
OnKdN9ebdTGtc8Nz2ZDMALTlCBlsd/ZcMEw3OCpGkkAu0CFRWiF69ukvJ0aYmlTX
fcq58RJktdPH5sLgU+CG6JVe09bPdnhCWipD6uQ6p+/LkwMWiqmsh7XS9xV1tPsx
dGCL2CQW26/JMi7FjiuFVY0m5ARYx7gkiAedj+KaYCfoZgmVnrs6KG9A7URCp315
G9Og+qHchbD0ONJ4ZpBr/BkQ+uo6HPuq6QPnA84vUnuI7Rg3aCaUtiVNMNJWxybU
j36ZiDRl+E8GvERgpDv6makznfDYc703mKjpsVtXB3W94Y5246r2qfs3ikInqNw7
aQ0jvWiIs7IjR5/jMJsm+JAcADrHbV3MSh+ByRuWFir3pUVHqt3IOk0rZrDX+Rjb
FeCdxjwPQ19ebghK2tZneosLVJhTlxCTMDbsd57D+py5JO9OqExLJWWJxRUsmiBD
+mLtR8vt/UVdgJ3rqW4/PHKpWuIxbq0fbyXZXmyg8EQTmlj6K6ufiax6FgPpdals
+6PjPJybais54bx7lBRSoDZUKDZ5u8h2mOxhIHCx0kyVDhsuIBZ+FCOVmxd4khYQ
ZlVWGewr17j5TVFH6BGPb8qyXFm8Xzvu5ov/wpi89pKO5dj92LCgn1t5VM+GfzCo
vD+YbVyVCk1GCT6g/B3c8mv+6J1uqp0rgVUXOpobTqwXkztnKPGpI8trkIBsA+WQ
mSwyH7Qsv9d6ZEFXad92flnHgWVWWXx0YFLrJauQR1C+WQt48HtqBS3yWJHK5Rji
iaK/LSkQIcE1+z1UwmVw527Ki7Ba8HOQT9Pcot1e9rjmJUCwPB42J6b1MAM+dUAP
mBzaZHRGijnUmgjYQJwXzRsbjFQVlwN09k+3FmShVKMlTp9ykui/DSB6qFxWBNfE
jGL6OUyuzZwZ/ooywUOdaWG3+GIy3hR9ACtAM/otRj6yQVmwSwmqhn7WgbQefCO1
c4f5mTtEsT+Q63+gngdYnW/5KRpa5S/lUDmqaG66gNIIb/r5THXWOQHPYTgcyes2
8+ywRHKQpJccfNMenFzkw9b/2LWuBsULVEI8e+J/statHWWZ2U/tb5Ir/19JzAyb
1CsCEcZkt/8r4OT3PlJe33tE2DAmuw6BJ23pmop2Z9WPe8oTLV5KLGGW3O7n93+8
IWpXzid+ZCeRxxnLhh6n6WsfNxRD167gKkjlz3MiWFlDi7VkcvvI4Qfw8IrLTmgE
zJgzs8GpZkEpxQtNJxw4mFS3fgpDW4BvnGU1zSXhojRhzFvBJJecnOElFEwQhkVs
nA9VE08TGlsuk+yGv+1lmoxLeHnknoFBq2SkErLxQ1jIjlU+0dDUrQS8+f43KN+X
LiygQdcljna/AW3/cXjSSXiLuzKIi7b+raBZDS49Oayfv6hb7RWZ2GV28TuajOgR
i/dOkDZqWLWHYdzXbB6a0n6ZUmF19xxZQqtZWePJUO4ZbxDsoNbUUh6iImEOynSl
wdTzmlvwouXhwG5t8d3IE6lLJr3KFcu+P+C4GFTPeAFFTuStOExIiVeu68hIFo9G
1ec+FhNIm1/xG/qzoNPS15yd9zjoySY64G5P6Q+r10LrjSsYKQmp0gtAN4wZ5tVe
93h2s+nn6JZnR4yqpIpRCOB17+Sv4oOgdh4NnxS21cpP/GDXaszvJHA6KsJw4v2h
0KE1AU5x9shQF2z0IDyCXcFxqQrydXRMcN1ty7ntDhHIlrSzrzwCj5L4rUQ8am+d
oy6qWKzxs021i/eWB4gqpxGB5KYkpU8s1/gk4h8jGBRLlb8UKRYDWp75Q2Pvz5+s
bZo45Cqe8D1MzKqL7AOCnNgFk2MRG0FlZeHe+EQK8D60gQ252Wks311HNCpQj1RI
ILnET1UdvZ/d//M5YHTLwyIvxfqMODjrYgutQKGczBmj/Rue9dUNFXjT5zUhC3BT
BiGIaZKWLjV9R6roKQT+rE17e2Advz4ZeZgBsOt+/Syodavy55GLmvQ7XV/XeF5U
aYsXxx9bI7fuM90tq15/XSOx3j+FiY1bueoGs01ZMc/61s+uWcQ7BhMWakRgxyoB
SeoYlLdmw74V3Jm/wuS206TyaCedGA4FJRVFyP9uisvX1z1gN1KBkrHg3AoH/ER5
B4r0R3FEDwFbsvtI5zu4Ga4UGJFUyJbxnrstD8bSVcr5ukEOVO2Nf1Ps3Ey1kIuH
JmwV9YyKSQ3ROrhxLgkMPXTcHb1zz5Nh+bQn5JJyEJXyLzJBDzHRUNHiOkTgiz1K
3G470L8z/AET9LODo9pqOaD7XZRzavZJhfcgfV+fdoOtsOQqqpDJu5Gti+ogREWI
AKNOwUUCfdsWs1jue5GzpkTWC9S0OqkZOKB8WTHL43UBoiLSnJ2e0mXpxXuhygqR
77173s9+mCpuf99NfBdmDTkXC10QTw7TzqZMKAje4zAAdqOWRyVEgZA6DfUi4/Ty
n4bqQE37v/2bE5jbhwyZ71Gc7Xe8N1AaR5lGCZfe3iELl8hfKDwmk+so22g6/m6p
HPb70fxVBdoMj5heIGCymPBc+5kEQ411dkaHkBFS0rtOBRG1FF4LWS+pjmD7thKG
NcwEXN5CUhP3/v+/1UIFtdbWs/MT4I4e6mMUapZwqysZhUfhY/CVOrbEhcySFrwN
wb8NZLIUNmFdRiDVyIPulCLhgGOG77k88WWko/SAnICP8FzeUuSlGoW1nNPOL4H6
rTwqlzdq49smscGvRGwryQ6nLZVbr+fUItHfApT8gk0AcakGcsmCBhZKrz7ZPxpr
gjTHrzv/T8tvW/QYXR8SF+K3KfJB2HobLo47rlq4+lNVPWmwi/3XClTY1oKLpyD0
GEF6fImbJAhmvJE8oQCTcP8lKf+y9YbnXf+ADRChZI8yWKjn73Nt7R0x86LaHKf3
UBvIxghY7RnHtVI4eUf/8yKrNl/rhmW3dGXkP/jwdF3t5D266d/+X37s+cPm62sF
4jSGb8dv+8Vkcpffch1PjDKU5wABaCasH/gHA6z6lQ6w6UQ84ePCshWR93Mu51jF
JRwN7Ww/vYktOfFPzDkb//DNcLFFUM+SOauskdSlKbT2sHDYeLNc8I2daDwE66L6
z6kT5mjvkLSlj8hPjXFEhngYDBjk97U3iXL4MGinqoWh1BnbWHTSpk++4qhKUXH6
87XiOv8aGgvfMYpP43WckUjWwDOmhGjpfM0P4oe6/d+Rt+/gz09+6e7y6ppLv+Bb
bqNt0WrD6gwPfBKX66MZuW8TK8Q5KqqJX+zEWgzQx7tlHsu1xvXcnKiwyLVh0Fwc
VaB6Z0nSh+M3fesBit41QLWafmYhRU5hpvB28DX+TmWD5RzSgW15abcy1i2XIPjA
SOwCGO2bEyowcT3Vqwz00wD53EwESztmkveWsH5176MCqGchljDuebTOTi3i7Ml1
BSC+las6gW21YbZVtAjKYX9Ru9qUP/64JpBA6EoMFJBYMPQQvFQj6eIhtWoOtZIe
Nr2ZzHneNEa/HAS/79z31Jknksm8qqznD5SDd2OYW8P0qXC14IMD8WQvZJMU7BSm
Y02Aud0WIVNG7TP83AOpqC0AgorE4k4lEbnDaTwtrEaAuBJoDkrOZe3JWVCZeQdw
/9hMrDE5JImyXp3RbdBcFi+iH6IwTr91mhb6VvlqSAJtz1JLn3Bl1ld1jQcLQk94
J7ql2EphlD9SPPzUOR5w12QS0lQHMU3oCEu4QD7u83httniOOVbJtXXBWQIs6QSI
mcGlVUfKOMecqt0rdK2fTjlh9jxfVBdS4araRnS1+In51tdnarGSUy3bP34IqtsT
MWTAA1a39FNHsZ6W+t9M1xNa9L7ErwH8Jbkw2Y9RS0hplplu+COXWofksPAmxust
mVFs7NTZokcrmevjBLCuOcsuBFJ4fExROZ9+Dz/QMMGSM91773I187Y+ZM/Im4PE
g+Iw0ntRVAnFDYjB4BnBhvN48xs6sBKfK7fss2sat8FYQ/nDFkOO9irb8V9JfsR1
fUvztQHBdVoLpw8pX0fyQs8GLw2B4aWP8zaiKvuseix7LbWbhovxY48sns/CPlyp
B/N1uqkLO9f/nCnbUkVKVr0bmhtAlfiDi4QObkyp3iMlcrDoqpkc+KTtvV1ITzLB
nbY5GmBx4FCGb9aFTzDlwhyDtC7wA81BrOZiqob2Cad4rqQWvgySJ67zd55dc70Y
h4LNL1l0sm6J6mRK/2XLbXVqVum7smEgj9WFemQi9dPCv93jQ1U17IWj7v0agxRv
q+7OQa3tNfJ+kgptEhPff/p//lQ716sn75ghtWLzO6HrEOY+mqMz1rSczOglOw8l
pLbTxb8ljBYS5CE32ckYPTt5W8rGz2GFn4Q3e9DULR9s9pcYmw1uyKz9zjiIAwJG
4EjxMDB9bD5Ejpl0OyjfLttXy2Uh7A+Ut7xo5zASf/rmyBjhms0gYY4SjvacDWQ8
92YXkDfQGbpxyIDVvOBpXm7vFLLoakQiQPlb7RsjtygXf0bIbFOnjZbFtFxhRIhb
yM3GvFsVhEe/LiK+eM6BqRFpG/WLL+t51Hs1gXH6U4MmxLPR6Btktsk6g967Z5YM
hsAxzEIGHEOrVh+Qct19hP3o/zxUVHp+Yjoh2ZEIUXqwHW/sy8gUqm8vK9bx4NQY
KWMOynHBPqEuvteOwBRPlDGjUOu7hebEgIaf/rKoaw1TNkbhoU6MIHmD3wc2/f5T
OzroD1sOoJG2HS/q33UtvmuL47oxOwj8juktOoODLmFlrV8/tV31Slji0GYV/WRH
BG2GGGeKQupw5XJTqcvZuL6YdHdB1Z7NsfheDWYyVYbXaIhEaMZQ0ce7QJn1s8TC
Xh30dxuyzau9gztBKQR2qus4UiyjF87PXJ9XXV71QiHdtO3eUZbJ/2zUo4eovQ9p
vB40o7llehArukSqmciL59xjK8Ozm7qVU4OA10poOGxX91RlixMVkJlcReNrihMd
rAHW3rC8/DojKJTDbesRbGWMADaXUvPl5CFwGvNtx8SYrw5QWFPv6NKYoYrYX4aE
EW3qFYuCGBYIQa3aHepavWrCB+chNhDatpDMaVfjR7rkvnXKT/fBgFpvsZq/Hmo8
2etekGiVcR9/53A32iqS4yfy8Z64+0OOKgmYmMEH6SUMBe2Mo2/szryihptX0w3J
2ijQW7kq4aB+MPcZgbD74rmVLqkviYKs//O5D2yizVnTkmsrMMSgaWqEu36qcNMG
LmEa5UeOm/6LDHbz/OtuH7HJgOnZ2WDj7PpwuRBIhm8Vf4SFMR9TqoprN6/JpyYW
gOMZRhTxGfQqlBqHwRbm0T9Gp5OBCfi+cRAnvD0zGg86t9bRD+9ok7rm5oGFVmML
nqu/djSOoxRA4GVM9RavzbCw+Osq/lECAVY0mzXFePFwJu95JamF0J3YqlNKE2Iy
tX1SztCWIFnsC/UmYcoeaBOXkm2dr2A8xeoyH9JW8FCL/Jpy9f4twpwyM+HUlZQr
K4IEARG0ESoQ/LYz9TNCg1C2BF58iFzoyvUlLm1Bs5gPPbXcr9StU8M28XpSppDY
M2ARBVVpX1W3DfKidxo4g2n8zZT60Q6h72S4TOo2zAXpJLxGmTdogtwp11wr+7sR
1DQFFI52G6jbuejSXrDwFBkOJ4F/RUXRRES99WiVIHJivCATzcLtKNkNFOlHN6BO
nTGPBN/cFHe4Qei/ADP2qq3N3wfTKpZxn9lzL9a2JsolNy9SJmFqB0wITuMbpr01
eqgQOIULycPH3/NsOJN/BWGlB9DwWKdwErI8GgQw2VCXU0aSyAOTgNqdfdKMGd89
Fv0F4rEepJj2aSD35sOk6o4qT1gfnsy4kyhlf+Mo9lZjrO5ijeZhBOxHfrli5w3G
xYfV9PjKl8KUbIT5MhprWrvkjEvmLOC94OJaRN7Sa8Ohr3mosVEgh/mqBNiFLkPO
hXQlwuwtz4hWcGU8IRMzim/xgh9JHz3QKYCInLsn5dQ1iGfuJ6lnVQ8pWfWNmlky
oUfMpYKlUuwmQL0POx9Y+asT4vTd9gYB23iRXpSMMleLzV/E93e2289N9u1JZwXZ
FNpYZ/kRNdXtxoZupky3UWMpxKNBP/eQ9DYew/GSJ87y4r0iFXkV4O1GF5GYbRis
7ihwIG9kaPdXRWB75vHRN7d2Q5P8ocTBxdoRStwkuWC/zvr+X/Rj3Wp2VB8jGXfG
X3igEFEdq0ua1dZgp54ur6caxDeW2HwD4THlmJdUQJknniZi7rPK7CFYVT42adsv
7pgLiSklxj9oLa4T6VH9McNu2O5A5cGdpOReEZtcXjyuCPlpjmGRG5VW/J4yKtXw
yZ5K2+wJIc0T/txLnz91QqIRGo3vo+KjjFj4JYzWzfdwMW9GzxXrE9if5kdgAUbS
e8roWPdFIeUiTeWCTW0WonbF5WJiZkOe68BXZLYeuRS/1wxuOVlZr8FMXSToD6ZA
06+081AS0YK/2+TfCd5pn6Ic9eZ33sfwhmCCxQyvvhkwqPFix/uJQcnH4dpYo0uE
MQkavWm3gL2kx1GAtfS9dPdzifiHT8kT9gxslnZGBNWF2nNd/dX22zRFXjEG9DU0
mwJUG6RcK0uf3HbFHbOZVlA5GNkP3vocelEeT3Apkqvb3/A9xlJKOCITMOGQiJlZ
`protect END_PROTECTED
