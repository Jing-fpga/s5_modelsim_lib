`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9xZ2Ef/thlLdtPFRWWNFC+lK8TChchjaR+cZavOs8HPZRZ61D0P1vkk7ADtS5XaP
v3Zw72kSjVHRjgsHbfjNqG5D7y2I83FV/qJVkaAmVBbDvrPl5E70+RYI2RucOY39
YO7WM7ZFmdP5rjxu4aehz9rV2ow4hYZQxuxM6I/1/GqEhTJ8FRgeqUR5KvrDZfp2
txuv5irvDLn1bfjpSxtNLEnSOa8RUZTHQs703+yNX6itJucO6PcAk7tbIS1ItE6S
5+W689MRm+z9JxjRdZRdK71JrZVyAm49PbVfF6MAcG9qMK67AIjazR1t8kASjfha
KdUPCHS+2nn8uR1Ua9vidmKwQ8fH0LAQOzIiM2jTtCX/mHwPrt84AHbwRimWzIQC
B1Jt6xo/xikaXKOW+IJqAWTq2Clin9A1cLCpIq+ddaKPRAadsfWoYoEDmLGIhS2g
E56sTb3FNBBmuvAn5b2TmHrzueZfEItrBaf6/TFHbTfLEaaXz1F7lrI4y5t1cGzu
wBBUKBLWjmaihd5aA+2klzkNaUBUA7P477Kjy9Ph8MxpcT0w/X4RVGqUA/xrBsQ0
DUBzq8YpSI6r7ye56Lx+8uNDc3/REyyLW/UToSoWH+GebRwEemhHGSZOyGhGIeqG
RpDbTm0kr6P9Dl5Ange7sYpwVVXubeEFIxPU5Qf+A5P5MHjMp2vuxo+W/mXqsl2f
k5iabP+KV5598RdztrVYDS3asH9xh4goWVLvMQrILnb4TfgwaNcQmdJUu5QzyQB+
qIeah1PigUX4UZU4rvdlrZRuqW6Lnoelzps1bWijfq1ZzWgjBP3LmiUhz0/RGJzH
i927izuCedlseHGz/+QZohMgRqP8T3M7Qk8yJORwILA0z7e9xkqDi/ekHtZZ2qpP
3M1deLPveVlZsijjU1/1G7BD0+mumenaO/8UPdQQHaldjziECWBhJdtIV3g7L8nb
0h3x7K/RduQVBa/ROZFP1dw09Mbhn3PzLNbFPyl1ONt5DSi/K9qeavGIWn+GYQld
Zvuri5EZ9E8HsEjRCo73fb6cLkeWmNVpIJ3L0bmnfBBTUARIisKdssCAz4ZY8jrB
Qv7Kvy7xeADyah33ljL/RbZ1P0p2F42iCTUhzjz8C20UW2xBIzclrJbdyVZI8zPZ
zbDvCZjw51uo9+9JFaCeJbq94XKB/3MExDetVcG4RqvJq2SRLg5q3UG7CKw23p5c
v+z2TKrKREcAwRt6GeqczVZt6IdwemgpXaY3jNAt84DzYesTfBB3lt1r6GCNn7ih
jcwfqqoJ6Xnv1bH/GGWdvcOB702yzAyU5xJ+XepW1jmBOmDwvhiKkapU7gbh/za8
4ScYkwZaDJhFEjsCv0rZm6n/hjxwvZafm7iH/P3R/jRD3bd7RZA0ptFfPfGntItn
Rwh9GfQvmiJ0oEdhCqisuyh2tvcbUW+gdctWVHd+qgWIwFABaO8g43XIPR8zLHz1
eTKQBdWsEiPvnZd3kDea7euFThxb3k5zQYisTSznj3oXBfsI+OxDxXd9xbUKgkmr
TQ96YyGxteP+wLdeahjS3HytDUu+k2ibmJ4+uDRebK1uxReCMOHb3gQNU1iz8QQX
QY0n6xf1UTCqtmMAdJZCI0OLlfa7ky/TMc2aqjT1HZa8dJ4xI+7LMczzSHy4Cx7+
ojN3HLv7LE9uIiGI7aVhsu1sbf2mMxjY2INRt8Ies94zpMoLmv3yif9EQPdpVu1C
suFP1PqcRXucyiniC7S5ZFEQDPJtZi6gBfCW1cL78HDcu/7klH33JBcifbC4aNNF
RXpeWDUVMBTK7EWQEd5bTBbat5d1ZITeDpyy7/Ym/QWUect1PPv/jNklnZyCDbMc
icCY366dslu2x+b6hXUpnEF2sKoqsAeogF9uI0iSR3BVFDuHl+D2WqoLfkq3R6LB
ek4pQPMEJFCP8+9O+b2J9odDaQYxdjuaHabQoO+9FKXuXXUFXQKaePdavoEuml8G
6LUqz2GHsvIWXuIkRUXPKDgHrhsxkrc6eStQ7BR+uCxWDpH+oGBYRdrdYgqxcEv7
DhdOIATgKeLqEMgluLhxbAvXjpTKlDPCpW6E8K/3Y/S+V3L9NUnvw/1ofKd3K+gA
LP/ZIsDJuFVEe0+hLX3TGWPWwCIW7WcrSYMDTd+DzMc7naghBo6wHMb0s6eiJcO2
bSmN4KLpYJf/5P3Tf7W5D2FBBVVm7QDezid+h6pycNOGSJ6mLpI4Jb5HKBidodTN
ZlAW01aadfvtfNL8H+oJ99MrASxEgM8/r2hTjSwZr1V44L0bh0LwGLLtAHatjYHi
/TCZoZTgkblJYZqmNxlAmb3GNeutfeG2R93w0mxsHfPXVBSUyPoUMOqELY3+dtgo
jdnz7oihOPrT3yxdh/Ql+lBBeMQKWSgghHQOehh4JfwIqBGO85bfH92Ua7hmhAb/
MZS3vmGSl03RCbYQtUviGHdnyAiIiYYhxs4EIjhsRpNALtjHoTBaK6Pqq8rbSlG3
BE8TSnjGP6YqzR1uBYHHs3H9vqcK1oS5zIp3TtAnOKWV17HYNIiMxq6d4H3q5ySF
En+1hWQyWxuZP9R9D+ywhZsA5FL6r4JqUBl3PwphT6+M5tE0R3hlQ+iPbsH1SZLU
mCSbt5waM1BGqSJVgCcpSr421bGKpsbs8vjddCyKd9mIzoXDp1awhAxPy1BCRXKL
QtaGDDbXrTrWG00lMRq99ivIp5Z/qqrvTzeOwXGxGcVs2yYz1MeD9GtQVNmYhoKo
11U1XpD+8nMRtN3Av0megCa+ZtTpPRq6IQbnj81ovPGpM46TsrfwhvjbNNJ4v4yI
FYAiK1AKijwvbQ3KInesmuyiDe0PlEvvkh5bJXjH2wxni1fh7LBT8v4eIvEg+/89
XY9GMKM2BjnbodbxiPL1fYAhgKB5HN+4QiJ33LiVYwNqTHksBherojfBs7BTwfE6
F56YNLPtPCWL2v5yqVLwlXRH4nzSd2WSIATXaxNCcMKZi3yc5Jbimi2389j1AFOF
B4IbNafxd31sTn7vdymFfmY8yywWRIRlNAdC1Mms2XTvw8+DGSVB2FNRMIUFxyPc
sa2W217jbcQzUfH4D1LAJJyCCpXZ2U7vdnMOgMkmT/5GnZ4kNzSbs9bLdgJyoMiQ
NCV+2rL4TIwrrXsM6zmYakTr+lC8Kot052yP2s5rUUzgPECy1k67M6np5bQJ7MR0
b7tD8XSrDk5ThCuUu/rarHNyDa2MIpYHgEoZdgB+dxb5UOwMGxx3se0Tu/TcmPfk
1Sx8F1FJ33ZEacGFLCnmeLc5vJIiXHB9OMhFjktbBGUR7ZFR5rIUpeYGIAtxmoyF
Gjg+XQO7L2AfsACptmj4DVO++Oh/GxAAhRJzUgAaMrkC1G+Zb8CDrMB72/MTawxQ
tq4gxLlVyHlArN85k7xOMB6i7MqcNBLZgMgYzixJ1ad4GKnJt9eIVV8DF2lsMcMP
ATTUJ96VA5brRUZW72NMmNsFFpVjHr6sQ8nxtiO2GBjf5C3wvp2xWkt4AmBfdeaK
RNtd/Blo1A0Ovkr/zyTr6el0nBvDOcJAupbDpy1k/yXwzDC5KcXieKkX0+JO+vmc
NXnU/bFJ5vKUv7yVoxLcU8zrLfXJiqYHpSBQ/XdNbCPBQ+9gcKRJg4I0jzh+YarA
ST4AhJQdKlBeokiUYJKixtBHJtx530lydUY+SptgrKOf5OAbJfRrbveeh78I36jA
gXhRQuSHF9Mbqj3YIGDOJ1Pmpit8J8mZ31xRQvFRu/EvsXYDfxaZqF5E8CPXVVX6
uukNX4Pq/RFel9D3hGi1oqmF8kEvbmbTaDtBCFYZB0M7V0SV+Jtt1leXzoXY8uDf
/L+SRg75yon67AOPN53UEeYBuAsd2VVv6GfPhbleyF/O/EDgWxxgSdeUQ8H3u+4u
CXufcBLV1KXLJtQfThIv4jk6fQShL9Dl6aLM1VvaEVTmHxY7wTkrUpm8pLQFPq3S
9e9mTMDuaGGhMRgQ+dHZm8EULCS5zwfVrgnnvFtrFmp68Ffv3ksuUikkzA03KaP1
3JXs+V5Ty8tlQgE1EFPmWQGwZ/B6VrXCHVArSms8g2U/TLA2D/OoUxSA050P4dBa
Bm/SvTcYTJ4OnMO5Pwf7DYm3ur3UEDMuoxlPC30R7PTDaDDn63oyS21eZcNtpFL6
4tkzXBAKp64cRAMATPLP06JijzrDyMyPLeF+BiOHrRrs3ER69xgj9Viw/yui5Wlb
PBtgUBVXSXKqdDtyoIV8HBspP5Uwgf4KTDEnzpNRVIo4nPAJc0F84NV+/vSVBpTq
4zR8/alPH84aV6Z1g3FN8oEK488kXFE0UMzm9JFMy4CkBZuboGaGOK1tTs73GD+6
N9aJF3a0beTVIHoIwvdCfkTDhywxKpawP6A1La6cJoJP2dxMGCVbbYrEQyCyi5c3
4ZHP0miDuNp7YoWktH25LGQXOu0WGXmfzixHH32yiKnZM0xWbJNezIqVZvCnMAv1
DvKo3ZYWoG2eNI9IwLQPELTARbxRsBYI2axNC9saPNIHzAAOUExX2HEHA+pRm67e
edTYUfkTDSCM1V8+SxoLgFyGohEtcPlCfVJPyuFzjjRdN0ClZmOfuyeDKPl5EEEz
+rK8ABeQbBEToG2UJoeLL3xbcuO9GWn6xR28M5kplbs/vq5/s5Ql4N7mfk2UZiG6
6x5WLNmQVNw7zBqBSWL3Y8h4thoheBxv0gVys5TtleS+ZBUHmmuG5cYroXVzzqxp
e/rA8DBvlNo5uElWZIrEpSDpADO3mCDdr7Agk8WDSKmzLCpf7kGyOBrjgpjAxa12
Gqo4pb/WMRvbIBUouI/KEwkpq+4MI3iQ7peGDLINhPkijdQQLXmAfmWoII96rvQA
WULCkkuqp9cG6F6IcBqyHwNtVIIVti3I3G8e1K4iu5sMkL1AqT9Gqm5AKj3rpGTq
fAd3j2huew8gJUHnN0gxeQPTlm6C/YKxGCVvQxbN/1GVvWOFZLPrjXXLxBTPl+uW
ygEypp3x7Q4lgBJWyklQF+qF8FR+5+MZWn2nJd5g1bj5eaFVAD0d1Hqu1lTYeIQq
FeFIuGzae7oyf2rJC7QBMy+66xrxL5nVr9UtjE2cLzRcRnU/BNdNoAkbZro3S4kv
F9fldbffhNd1Fs0REySPatiwvzSaKUHXWjGBuxIbdzPhiGAhqueYMnOvzfAn7jBg
`protect END_PROTECTED
