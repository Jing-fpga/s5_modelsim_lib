`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pw1Mdz11NrG0Gg/Hi0UgjEmi2PUsr2hpEj2yYOMjEFEJBgabcQu1D28N4q6l379E
9TGxmRTAcgMk9mO3aJicsE2q2FIN7/w+K0tBYddv76WJMdMEh6RewDPjZhMfUpGN
VW7y1mFQJorbIFMKLYtsOf3wwqooViPzTS922izji4uGrutRzidYMza9Cj9IE702
4PEJwmYpkFswyLM14Xnq//SeCJns/+gcYoXewhwnCZf0peRqyOpXtKwmIxe8VA09
pYS1IHzYFdGU+t5MRirH9EIBYwifTWbkwdii+D8K6iW7X6+O+hPWHTi0CJ42pD7g
K4ZABeb7i47ZS1AsGFvOYCa23qZA+zKri1g4lUu3HJScLmbTguVfCXDqE3WfVJMc
HySIshOpticC4vC8woIXJD3WpItaDx+uq9KvkprsbvDDem9d9BFYkkLjZJ90q1Qi
Lgqd/TfkHZ521q+XAr/L/Da7gz3VCe4CewU/hCmhPJHxMLnJEBQ8nbO2cMwa8sii
dVsbXq9xPaYGXHJGlDosOQeX+r5Sj/Tsgcbf5wDM0J7BnftT4lJn/JyLHHWTSng+
GURSUlycjqdjooRxneYr1Wb0rXT7zGPjZH6O04KqJZ5ZqnVLAVVRjRt21LAKjkVe
myFLaD3fq6jqU1AbNl5aUIFRGmZp7E3szXKOTNZjOx6eb+Bbpdp37hCDG4vQ8RNl
crrpphS93km27eVXdwcYVqLLuvHFVRQy7rknCrsNKZ0R3xKKk/lP9KJOGelkTh8r
gUmtay6Kak3YSM9TwGvJjtKXuXFHibXiShzBK9ffuFGcGbvTTjUpmrLCT5o4i1iv
3WMZoUvDi3Z+qugYLec1X63SPhc2cU5EM3zv+Yy71vYJ0xRiIctu/dOgkxoPg4dd
5uzpWKh1hIBnC1RzVlpzDLfpJSFCGGYogCBOT5FLyJ7rSLg1CA0hbA/Ny4iLDrBq
0c6/0ubZmi7dOolKEJXWtAnLuKf/8kr0eFN55W5QDpOfcYRzbKvaZ7rVd/p6v0/q
DGBMheS3suAQnY1mvQpaY0VYzrtLnOVieVDLLU1p8jxNzjSOla6oQbqYYRaApY8T
8Ya8NGIC/yoVltUYAvZhHDNnFKONvXCiQOXFLre/p2wyTTbHWHTjZ17MKcIsKD+I
bym4WJqYrNnuhSA5xzHbz+qfO/CpMItKScqftD+9RT60DkXXVHEmp7DDJGXfi39l
wvP1zXEE7s2uhg4JN0mCV5oCU7H9jZ0lny70N7M8GSjrFSMc9pm4OAgWNBofEMVP
w67GNG/azXx88lHekL5MDwrg6J0BKmtL1j5B1eedWUb4wAR2vlaPBYFXg9PhP5+u
Zqy10aAAFbuSIWOJkpubbv8E3qMQJGpGun+UdEVe0xRj7riCI2/hoV/9x9Z7PjDP
lox5y17v6fqnvDXucPDwDdpkzwASNInvo8KgnnhzyddFz50ecm/AXHZygFTfXfip
8iU8DIaokCYVSa51cUqPYmspEqB06LZvo3Kn6S/h+WEPu/Iy/U+OKSsIQG2QHE1e
TY7zjMi5o9j3DNziY9/0XQKZ4yU3eUN77AuOFkX1BX4uaEEmkwSr2zZkmyrapS4o
duW0jyAhW3LCpNtjafs/WyrdNCaIiUKmyhoCHOhi1J8uPDa5wb7Z6VwH00YDXBAS
bl7JbEZxTQ9QlE2MbmVzhI+1kIo1iUp9i8Ar6EvKNKOaBp88JBmwvgYIiW1F+Fwz
Ip2LmdHWrxQDE0xc959Ad/DfWEmdrc1jLLDuL30XCAtWLPS2qNVcCM+Q4UWLyieS
53O8twHA8uJf6WQHwS/UevxXKtRSfvtrteCTiXpH9VXgyLVoPfAD96kQR2mbQW0Q
1f5reIK3bu09Gys5xownU9ei7kXMaEsieqXyqwJCfOA899g9q4eIOqCTntvLjM/e
Qvwvl96io7+YDM04D5SjqCVc9nHULf2tlpJnipEz5kwbVlG8UgVZiyU0PVEYFjr4
55Cuw3jqSFgKZFLZsQPu0M7XFipOlUi5VKLOQwsiYPAQPSemtGAh0/ieVLqEszhx
rYbJ2z0HjWjyIhF5WJORKl1qbq2zFC1yS3ApsT2hzPEBxdweEfnq5UA0tLxqRecO
jPWKgrCdP/e5EjlF7GAY+gTxV4R1Pd1SrgZuuSkqM+E0NvKFZCHf91j9FGwgTv8p
wEBP4DC9QkpYBFUUTjn3GbFvbzHZRgNlqFF2SUJMSzCeNG92NvH+IDrMQ1Ig9Gsz
vDMhwG4dsrG83Pw+nczCTw4iGWdgNF7rDsUqegUMqj3kJ+pXi/oaXz2/2zcEmZQx
WdRh3jzt8iJiscBymW68wkrXpeIFuUzWXooAwNh5X+DcKDrdFizTwWAW1LFHq9au
rDnpfZ2WLYzeDHS49jyZzURH1kUflNuZvRduSwYSMvM7POxzaceQu/gAYdGScmg0
Sc4fhCVIVIMaB6U2IgDojclo40jvdDzRLaJHWFd7bcj36db/KCF8OHDsIWVYilcT
mYotkNPxf1JgRGbbbvrJzJyuUenS7gWjOT43sqmNTrE5FHgTyzzZNnVfXWFHy4Iw
o/0fpnfAZpsk4jWzrEkdcpxBZiwhyMxVvMcC+tzPRz+osvr34NFwO7wrGozpTot7
2DQg+vV+Dz9Jq8y2KyTf+0x+Rxca/ddKrufezfXasJ0=
`protect END_PROTECTED
