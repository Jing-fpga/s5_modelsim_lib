`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hOVsdrLkS8iTofZr/RaO/w4+ejFQEpcAavZ6rRHcsr01O2G/y8x2CJqblwxYxXHP
ocXh/7+0zUUFfmMTZp5Cr/yf8ogSbIkJ1m8WgL8f0mN+Jy8OeLMpOvokZYCifZ+j
eoqWPBzATLWNbifFj8dmmktom/o6+acWi5Yi4Fw8zGymbrR26xic5cSwqTci6L12
bc5JGJRdORoy0lULb7nn1RVlCj5tXpvkI5KOxVCTL3IBkArK98RjRH+qcN4ejEpQ
Pp9g4NaAvxPjHzUMa/m1GwjwSTH+1lDJYSnMchw+KQQGcyWKGN/5rw4IuktC+oOd
Whnd2pNNM7uLiQD4qPd0mk5IYrOLVRbCTldd/P6cvQyfj0uUVYko6KKwpewOe33d
fJdk4ealDJDOgAEkORvRsDc16wbA1AcUT/kGh+Dwxd+l1PB/O1NvGkbKLkt3lekS
mpxjnb9bPHdwqRjez7EwJg8wCcbCPdArL9lmWNXTGmd9cyqEqX5ct0gFvCl0EcbZ
OsFPd0p26VWExR00TjCvq+i1oVe8yXd87XmbFKJIbhBbumenNF6+FpCak4Nod6Da
1WHDOOYPdihd6OvIIrqoAZ8WPI57eBMZZj0CUILFsJwfjV+JkdQO3ZTUGRGISUWC
2YDxjjsIblFcEOL36UUsA2PD+ECZl0Y/rD3Zsi0SonI0g3RgJHdJhmv+5LwNc5z5
gd3dNUELOyaSUnAQz+xpIWAExFli7Jlswkqt6q8Ivoi/sG7Uy/e3ohYxsEiDHDtm
27obBwD10w4KfqIDYDX/MyVr7aJKXkzAmCpz05vqnlLdE/kqFjgz2jXClPYwzw19
+rR3tnSfKwbrA4SO/ZEYi5ysi529BvfDyL/W4dn8q7v8iw6omTJrK5aGSAAKhpVw
9y6VC896omNrGUdHz26/UNQx8sM7Ti9/dCjlBZUWhLr5WnlS5R1PUUOa4/3Bop/r
qwG8TJx+WMOL13Qt82UEwoH1qlI6tKNXi8lOF3OkNzV1djasitzqYDqL8SuCwmKv
7nl4i2SIj/0jU4DXniZ3HgiONKA428D8zXBxjECKJ2xfRPiLQlqVmATIPLNv9e2d
JzdA0ZgX3vop4ebyqovmIfxtfIpWD3Jleh4AMDrm+GIYhIDdmt2jgKcVQN096Pu6
JwDCPxYZjAUhbhseurokIotoX6ZyiG363AEerEetrIqpo9ajtAtKuiXmMsbwKkbk
XazJRq0Bdrm2ZM8pz1OjXR4XdDeFv1A24Of2BEniXlFw89ZeJrf0z/9er7s1/4fg
bDCMaktefqN9Gq5OiGVb43J0w2YzeYs6dLD3M+GnPHivuKWN/trrCCgbAi5Gv7/x
9h4lrsmrySszKlEn874ce8ZTT01zsWwWkdpBFNcLHbPfN5S2vtWp9Dhnrk/Tr/ft
ai1XiVmOvxsuXDwBVFfGnNmY3RVEoRvYMKx2hV6DjYLvU40jam9CNm29jreboTk6
xHLgZxgh9D9rktXHTnt3O9/joxyUjNCO3vA1lphnMKJuncM7c2DWhv2Wmb3KX87t
vxbIj2mE4qsOndgYrV/fc3ResrnGL9ptw4zmGKIJtQMadEhWvKUwIBM6fWl3qDqB
jIb4NAOjJ+riQDx2+MTIuE2jflj1eAi+e2eKD4k8/L3jeVM+b6vEhFmUdb2SwFbc
kYQACpA8Vn2sah2mV+Wj2XGLaf67/VUJwJSiA0Rvqzt+BvHedD7ikMYjU1V2A+dx
n5BkOCzxOidXGprBbWo5R+Cs/cauEIePI3lbn8/JhsZiqx1fEcGRfplh1/mGub/c
Je40uhj+Yr5rgnHZZRwB0X42se1YgncWKPpSLdr6qwnQousawTQTgVEzfj0L99PS
d9Vbatu1OeReMzQPK+jOxPP4cJPz0YZ1bkAvy1zfc8AE1O3Crf8Lm6OjNDbDO7wB
z+8wiygHRDhtkyfTlWVTWDJGYbBWbSXTKWkE4hTJLKVMA9WPDtFbzDQEphwSAFLA
RGbdpB6hJ5OLr4Da5dV4kCshnDVm9YB1IABnvAHU5NKx56Hy/bUApoNyYmZYNyfW
XgxUHcBpl8bX7bVPQTFZKdyluxEOqS6n0eJlN+JVNGu4Gceo+yoRwfg2Sn1003B4
xGWENvsVQ85rrtGdZoDUmOfLqVnDEKhgbGC8a009wz6fRPXPPJtPh0331ERiid58
YPFXyvm4K5sTKe/fejcOzArR+MQqePuTwcB0cpohu3lt8U4+LVXnVN81OCcZE/dU
yqQN7r9BzfzuLkk2uwlBwAUq3mtmd9PQ+hBAgZDzk2shDCWnw/1J9cdmC0e+kZ5N
UeZkKozynUGQ6QZsSNG7mV3Bc+AfFsnpoaH6jh2yfavuo4kev96gHinBKYPbu5Hq
mwVY5ijB+c3VrOSLlgsgLFiECyPFzfEVv8Fa1M8C+wgdKVVzXKzclpyCs77uPJJQ
vKiVoFHMKjRTzYwbVhcvcTx20ciLcwBeuwBa/mMYshEIuKBizZTgrYvM8+UFYsUg
1KOn3K38PSaiaTPxbn379c3Jk7eDFjZDRgo+7JxOUXxvgsOoYufPPOyMHo4G93HQ
gcXpl1IGv+rb2uR/UB48A+ZK2xyD0ZcOIVSBEmuFadT2bukpXhIQrtWktUikpcn9
1ghh6rktqQr04LWdygqBoRu9dblr556fBoAq1JpPCqeLy+Jx9IMexj2U+aesNsRi
G4wKpddGRf2LDm+NQara8k1sz0de2nm1WjBvMLmaDaXfiYA1iH9gkhLm1rtk8FOW
YQ+LdPFiuS1y920jRm0AdhCm6xcj3AfPiU6UYklFhccgLzBFAZdf35vc+y2+jfRH
BDkrFzwoliJnbsccs8TmwgvYgFeT8U3KTxUcqxBRVp5pfcqndlG6p5oQ0D02ayUs
7AphCX5cjx4RwJ2uQsRFfK93zfJ8bDzhcaI8A7mNwFmAtyvaMmmjkp1Pi60ztVQS
whxEhHgUuL6dJQTm1uTpOTjghbQzRJesOqU6j/Wl+3phVDFeym0kMk9bdm9XgBJB
/V5bF9MnkUCxC/gIZe4vJvixKyDBv8GoCXKLCEBVBnhNkB1bNqk88BU69pyjLNt2
dddeghgYKT8/ZUl+Dd/H/4G/Fke3mqNNQAPoZDtbUYPVX07b49dtjDQZSXEu2qqw
9TlvfCelkRrAcTDTQTqm83rPdjZzZurTikA2Voxs8wtnjItSl0khC8eCO76PFr4+
V04i7nitAt8lX6bVdsI0XvjRrSp+HmUssT6FCfIxD18tonpOKwsWcgHI0Su/+eEF
wGWvnoL3xj8PYJO0P8/cpaIpuiAuhUNh6NHwvpe1TtwqUv3ntCRBfEOjdG/vm/Co
qamMWskJzwtQ+eVNGMTt9yCc5vBjQaUlkKhXYGw5lMLmS5NWEsQz2eSNSndUrd8w
fJqZ2ccEoUAPkochVvfUrwuh/MDNS6rfeep1pu9TkFJ2ummBH7o2HpuYlNyMvDNz
vKrh4ntG/meZuE79tiVYimyrRRNNunGWsLXuGJFAMtgNl3Kgx4Ow8kYEvXNFyy2i
vSYTpPgaH3Q5yBt4eUJ6lK4+4cU/okZoJHKgzYGMkye7lZBWY8n7KdO11RAGitED
GpRSj0vhWgLufN3fdi99azVGfaflOiAklBmmtCpzB5wm5SpiRgnbwmN33nsUeA3z
JZIjMLWllZfez9XpI00sNU3X3tuyRrFI3bdxVPhIxESShTgRzDG9Ax38kbpcjC3Z
4YkyKqQAgE2mWjjH8OM/GFpvVNBSJv0R3KZxkqsyyAJjK91nbcY8m5JkxtB5IqcO
gtPxtNf7VFP1wEh8TKjNfIsc/r/9XhD8e+XtU3ZlC+k2432sCj58ZlCVooNGlFYD
By9CRu5ptTYtXN7oDbKzSim9xkC6e5vsz3Kb9BW531lpP5C2GH0Q8uGC2KzRo/MR
LonPSHMOpcDwpjOGrmlnPUjdi2+QDpDUmyB56U8IJWr6YCBvGcEs5A9urvxxaIDp
3QcN3gvEdTXGV/S2H7FEbPS/L1gB5S6Pol/2JyDwGd5Hb9TJGBOVA4iKve+J/6Sf
JGw4/iBU4G+gRymy59+5xQ+fdOWCSTMtlV1hZoN2hnm39TWlZBSjiIfNkodvJztA
UicSptkV/U4NeUBVWvKlCba0BQ5gjgeol5B07m/3j1NCZ/KKVs58DN1mGOtZNLN9
4+A7AryfCKW62YWiEH+UXWNczxTtrL0gGRvDK3ht5Ua68y1kfQx9sgMVWAgsxAIg
GEtth1zBm02YuvNlibSw5cpTGO9jmqR+dG7uZK3RLfPR5GV1zzAVti+ViHRBu6NY
Z1wMNxai4ApMN07Lih9AiT70lPOqyiOQ5j137luxE4chrtKOTzYLnA7vANZ6TjnJ
ONHpKwOnUYEPVBaCtHBYhSmHEW5f6JDjkbp6nTJBT/33oJiz1/sco5SKefkMYUQo
yhKoyN4pQnE0nB9o0lNc+iaTxCvs0PdUIxb69tzMlbd7Uvhdy2WHkW3s4tANNabQ
DDIxEZ4H539tpXvcipcNRcWL53ztGnVoc59NqrBv2OJl7uhQtP6/WxX3aLbfEg45
10ZHG4LlldHwb51W5llLLzlPLQMz+lckVLLkH8m7r3wNmdCZSYpQYcSO2a4QblMv
gbADoKPa9DGRnx+KsokAA+a9umGc0q9M564NBu8gSlpQmRJRpKmqduSYykmSo18u
2zPesBOkDYtmIVH+XU3WKxWEqpgE477C9v+LA+LyBNJF5Y/p5nhbTVA7gzLd5diH
vBHnj6IBQLcSGXQoMyCJGs084487/2X3xeMBRCXPGwwNWrclnzBNvpoYDx2NyGxA
NBOBmz0j0rP1f+J4xx3XrWzFjMz0NWtSqVSxjGQ9PVjEg7vEBep50xW7uPsiIhJ/
ldas7pstzGWeblFnF66nhwo3U/0KyC7Sq7UnXR8u/ijU94UPyBeoweSe+OWCS2V1
hQu3chIhBWGCGGRlaUhqorm7PKAKj36UwRcPGbspdDkR1+qtl05llLWFeiQ+z4S4
8/oeEoGzqrcMCNgDGBFcOUIBtEJqLQ6VBbknB7e+MtaZAM+C0/L6W4v7itglBeHS
tcHqWt5ST9wx3ND+N9nCVSOaryXTR0J6danUqcZQT9AnLmQwoSwkimUXaNH63Ygy
lz+vW94G/SXBsnA7ltVsf98fxBE/O1eyVZlujtXd2VvRUmKE51PBtZ+3vp1jQcCP
/pLJmW5C8pB/tFyL7twHdY8wt7gXr/mfXkqb/jjkLK1r9IJL4SMHXr6Ow/3DGzn8
g8B2+wCewORdRvMZpCpFQOYdAcMK/42UsVxOhli/GrNbE4jCJNOg9Y4EKaJ0FxQT
j2yxLysE/tp3DHBSn+8Ae/UegGT8JgTfAgkudvKMkbAHF86V+vfIe+i714z8lr79
LkdaVylxiHDkOidK1KZrfGyo9w+KDIaprH4YHf8z8heszT8RbM5Rkh7apt5XIsh0
a+dJyfdDWhLWaPUgozyIXkpSasrGdjiqmP/frajyOXuSeG1GtpFzzWGciMnx3h5J
xR/PCMKgRJpDCLVkgkY8Hs5MAbc5WUbteRyfvD4W9bsMbPJO5QH9H5hE+tQ4Qaie
vwESCN8GCRujC04BMXKlDRdceESZGYSKNvDb82oGGCO+iXmE+gni91TTw61xxWmJ
ckMHShJV7CJWeofTh1Icc+FEhO6NMkbNaCwQEAaSsVycAw2EfnjNZxdN3+29VYu7
bc96gw/vRCzu2/uUNYgAJLCW/6IeZBNAqvPpL1CjBM2eRe5/Uujewav7wgZ6PiiA
uewG9cSv6wMD2XA6QcX7dI8lxCfnHMDc7auQ5sJ7SvrsheStxOnZnRTHjJ24DRSI
suGVTOvSheGmT+w8DjuEvhL3dMi+zePHUlAZ5sm7aRexvu7/KrzZmeIRlUZzF2nK
SjjFnfmvxwoQHZDneqMmPXnNG5hkXSysoXMXPcPRdnh17x5KGV4pMBlWUhc6XkrA
lK0SoM5LQbnk8oBSzWT28v7u7jA4vM0Y+6I2ug2VOF9T/aWQ6eHE1qzXk7BSW6km
x1uQDwjIJOHLT0tXs0D0470FeGQ417JHLEdPHvs/EVhcAS+GJyAl6Lu6PsQCxulz
TJ0Ls9MYgYPW4L6dRRDm/rd9qftyigVYTWCcv/DuumeW0OhVt4zZz3DA8hhZ5/3r
8TQOUbRHaFvKVQJer+DWew5f03jJVFSZ2Jung9BKHXPOzMECJiDD8Jt7wwhXReeI
amjqQSiqD0WIzjuUsidlvsRPtJkl37i7ICZM5APJVidwXlu06VgxsIW6Kje6+AuH
qcnN3Lgf4iyiFAIdVmTa/ArAPFel+Kyb/uu8gd4Y/Qnpw+pNUTJ9+p7qd1cwJAat
B6jrVmqjT15LBytZ881kTxCC7iABD29/bqdgMt7MxxY5wcmrfvm+mqkkGTPSmUCt
cJkFhoYd9Zog0szl3DiGcruU8wpQUSkbCHUdmar7THqA22XR1DQ+cMT9kxSJpec+
M9f9sP7NwZYcQRfSqF/SdBfvNuV3uDEy1BCmrDPP3yEwQqGoBGIuaGkKO9d0TCPr
58CyO3KjBTFnLVz7mJy5qJtWOh4y9+FBRf3m1p3GlkOSp9PbxlIfUK+osdhbw9wN
NsKA3PzApRDM7xtoaXdc4Z27nCWoELJNkj8UMkKiLrct5qoOy3QcpKoz9/yEEqHw
wGnVVwie0NWmij2wh00zxmyUmNsQORBF1Z8HhwoZk7XWVy94tdxBeWj+mxypQEMz
zPKkc1VeXvLclf2P8W4BjHR6kF3+9pKl5lRhydI/81Duo5UEc1ZmV2+m49o5rBXk
ND79z30WYwG+9bpS1AM0KtLuSQLuULiwtQFS6CjQd0U1SBETuwzHR8JlXlOxLe/A
R3W79eTBH0548XrafcMmcqyhsZ73LkxVb5KeqoezODIienbrlcSNBL4VUI9Agc/m
2Go+4VybETpiZIZtAi8Sk45JfabDIT//W/pS2tLlCGk553d5DPeHgAWoFltrUhkv
bFiFo9xjPSM5SM4YzU0yYwSusp4VaJS5vp5fOn5ucmCbF6KVVSPMpUQNdrqOQg9c
DLlWu2Uq1ouKQDCpjqYpLl8ujn2ilO7R24yEuLZ4nnzHMcSIw5gsSRYUNARLp4n8
wnMkR+NE9Eeslmd28uBcWlE1pnAoYPQCY7t6dCT3NCQoxpHwXGBdYndc0dwvcInD
sLyT7y+BJEobJf4D+k2Z5ODmGK8J/T20hbAqNMrvjUoO5flbWyGw+TEbVE5VnI6L
3+5+LZXQH+ef5/s3cUuiE4Xu3o2TI/wb82cV2kDgaBa2ANRQ/PkNmMUiXWtrJ/uQ
5FuaGd7VvGBvgZbY4hbPDjdmMP//QIIo/cYHDTOdguHB1ZX6vn2KdtlrV7NkO4uO
Vb0s8OK16jeXWJmcmW9r5kowfjc6jEFyxpGd3eREp1V3G/jaHdpMH1Y97iY7pgQu
JFPpoZyXbIJUXeet6stjIHgVYx4lEUOsNz3YIABVJ97bfhlenivu4PZ0eQrA3gxY
m838pWNo9eaACXNPWzTqf1ryAVvxL+Rh+ysYebYBcMeBSUwDk+UbiyQkcGtBNv6P
QaCFFaoU7uHi1aNb9fSQOVnrCVupM++6qE8aOSgiRnJXLBRxA3KyUvUGrT9iGqqL
tpxtUdgL5kQkm2mUgNCTjIiTkY/RPQLfN7G1I1OsBDEMqoKN6pJuZK4ZV94zo2UA
b1311npwJwB6xMNB1Hppza0qO+VddV7nUvdSXGr4TNQn7PTwEBTmhDBO63/AZ1EG
jdeIzogtjbiay+JxtZJDkIWcxIQszkrL8oZXSulYuqg1VOtkFQR8YnNXzgmJzORM
EN3Fu9wBQfE1fd6hSM0q974+MaEp1P4UCaRCh0N8f8FxFiV/g9JeYK8LCwEwQCV/
g56tVpbnAeIoJxZsaFVGtfuMJ2gxdt/LSGrsIpZ14ioh+XMM8eR9XcMmk22r7tmy
Hdt8tlb26upvVqi9r/lm0huARtFfZkoP23R+Dk3Bht4j/UZjJ0dItLqBxqmTX3SW
Asvn7Z6UT8ZPbx2C6PJ7g2Sh0eo5n+nhmMXyutVimRs5nNeZ92RJvQ6vmO8B0/QT
UI4Sw0HCacC2pTsQZzjiDu+xFrndLOQdjDtSjwSBm2tCLlhzdG38IuuFCkNYMQQR
q307QWrcVcuQXJlIpRlyN0QKWeBEb35VA+u8pl+kwGYM5j+rcHguC4dcIUQ5rElO
5u697cm0bBl35iXvy/EBwcD8mYa99Ndd6ActW7FWao4470mbgZPg98nqUsppMgYM
9dcwwTWXUL4X34+kCYTAv9AS9rVBma0vz86V2lswigA0giqWLNFkcabW7ze+g13k
NayatAgr6Hx0h72aEqSZI8lXcylux+3LZyEZD2DaM1HsHo/FSB4k54WDNlF4dsnS
8Mj6FD1SE6Dyn2EbkmdE9+zJOo/hmG0BiMXmmPS91p8HzUSgHBsqqiWhbbWxJ6A1
Hmb5eKyJiWtD+S7HsKt9D3fLGro/NZoe7YCSHSlB0U7h+YY1mN+aFObrKC66PDUg
iSSIxGCuYToHcjFkaDjrlm7J7AgLy+DYx86TWkH8PDW9jbUx5nRjZOmuIVkqnbzD
XAKx3kgfPNxSnt8bsATc4/frhNLhC32Vb81zpe/CR9i1dMSAapWxEkZXlMcNUoXs
XD/wgwVHY24tWoPPpSGlyW3neC1cJX+vkdclM+kMbOABzINYbgym9L2+unAMjGzN
Vd2G6oBZZ5fv36eIGS45jsHUATFgOB5Ohu7TRVR7OQz1aVl9c+GkkNk9/6lKa0gC
QUeqwH+ez4LMHDqv/cYl+j0h1YMoLg7YjOo1wWcIETTBMg2hTj1TjPPLJhCFnqRw
/48z2qkGmGde8F03FGzlnB0nuxb483c7/61IgZCCG56i0yd+06UA//97ZV4ubWsB
yg975zR2Q7JvO92lRLEc92VDUZFTRX0BRSth3xyS+/zIPY2OOgBLGv8eejtyL7PB
1twu2SuYR1/byeAzLGAhsIyACa3xxcG8fYQHWEnRcPL2muf9riD1N2DPXbT05zTf
Cw5bygD0vhIN2eMz/5COiDMx822WCgnq3Lo1EBkwYfhrZB4E3h5WE8t4S13uzapf
kCwS2UvMTxV6/TpYnFIqQYSSw++nxPyoLe2aMafbIEAgse4OwtMqQNiSXrf4Qcdf
j1NWEnwIRgsg99R4+eXihwk18hUuykjxPiNcC3+vpC3y7aI5O5m9OwtTZGmTsgNb
VtKxokgNRtD1nIS1pERHule8gk4B3+V9EQDgUg9VbG57otMKXHKrBGL0PDB4QmTg
L0pbTabRhX2LtK89uwWpUaHEnzj2ggQ4YM7pCscbEVd5jN6ChUbAznA+hvqTewOa
n+2Y2DW6PbZjb3jQEBgI6yv6bfiyK0pqr+ti0WsybTPDH/nylpHBjNC4yFMbcy7u
79EiS6+chTS8OKHvhlwhKvEMfz2mPXyQi2mthw35iXwZM6Qys1z2RyxpbgSKVeWQ
GxkXUI1dstH/G/NL4ADgmVzzxObOjko/vXX3xZaBqAbIxnu+2wXX4fKGG3xbKFkE
QPA1MVQ7SB4dlAHS8hcCIFYcuQ8vGI/FrXJayg/OlI1H1ECbGx41Qs3fn4910zYy
SW8FKDYjWrwxl6NJqWoYBrTuvROKqTSf88UjCFjyygxOGuw4WLqKAbnSERKVkfJg
T++MkPp5sCTXw77GWF2wQm1759D/lnAXX4G8LxkUHB05NBqFIwKHUY0PViJaa/TP
o1dd7P1HNNJKtDJUH2TEDXXpjW/j0v/KC03TbQ9C6m91pFJ/NZs5eK9cAucX1AnY
y0vZcS4Gn3FrnRp/nxrX5lKK/rlngjC8M0MJzMB/bIKwDmFLiWcx8Xjf5JS8mw8I
JiH5PMpTGuRLQFp0uSDMnm9dKlj3vhkA7lAld5X0b4fmPGbgPaPYdydM8BcbHSNv
9mDxXuo6YqywFSAllf4/8x7pUANE8HC0KPDeJw4cXfRzGUmOfCygJhvH7rWm0ctP
e6tnC78TwD3BiMCI4vocXSZPwpxHLqYW/S9IHmwSX81QosmYF2uNtdCGTw2ulZRg
0W2ahFknkNFayOrWilnNeak6eQT4ax2go3pcUzVY5A3O7z7F6ZvYc9ayfNfCfO/y
WkwveGAVX7ktCwr9QrUtAvVO4gZR8F5w/1AKr/0UyHtTagClXDnzm1dy0O7nPjR3
3VR6Vd4YSbYVB9eHpAQtxS7dLeFzQUlaZ9vFsZCDnnXlwCgi7NvfxGw4afQL2AXe
tlN62aPkuLn6xOHdMzYJESlYkk/T2LyTyJb9MCyLS8q1qU3OARcQMlb2oLwAB1Xo
7qiAd3DDd7R4TM7qW4VYrOHm4nSIpEfVNGPXRGCuGO+gTUvYe51C1RKrTonhmXmW
XyIjE7kyLxuK+9j8MIjXLThy9sAdcLKWe4WUtAuCgmOtb/0cWsv9FP2Kh/IWqN+5
UZc576k/XMOKFkbnieQ7BpKpxoYAKKsee/tB5XA0pIW9YqhQYGilz+jstbwf1f0T
MGUzw4+nZqVMOMHlt6u3rvikJ5498n3UgQrfgYzFKVloOj7B3u/tIKwB50qRG8K/
7NlBoh9Jqp9EtYZB2RtXuMV469QBtnPa2xsyG1If3CxpSrSEifSQ77YB7vqWUAW/
lxvZSRgshhJFP6yPdh8KgwAzkOj/32RqvQ8wS9SYT7zeoFyLG2gpslMEpFhV20Kq
kfH7DyD9iCZgIK4DjfNchYkj9pyjUOgVR1Mjnklp2L4jJcU1a16IpLYmG9K3rWRV
hj4KLN6pTquoiYCSopaGQPyAS3/YiKOJs1DHwG43YgYGovniCCt+fwSdEK/Tu6Kf
FZXv0DeTHQWrJcCZFfKaXkBI5w0rh0ObMKafkN9pb+Lkhf/Ga+1BpaP6qZ/nO/3m
CWVdRgVg2zBC7HPrj8E6L1/I8Ztl544E4IXZDH7DPDz5huC6NkpdPWgcdpcBpYt1
ystefmcJ3oCOh/pE0NNQwJKIzsL19LIrfuA6gZxTf2NZ0+BiWVKiORLeT9yPDJVa
14g2mTunDil1feNjZpOjm+M38uIhjW9yY5MdyjjU+ZSPirvY4SofVZI6VNt/NOuM
JBvGWrkMNSkOB7+BzqszVo4DKpYe2ye4IUCOj0Xr302zY7O6PIHFlTD+J6Fk6nQj
6pnp/V7uotYQb6uBKoFsiGOynU0BRXd78sA/04G/jYAcTtQqLPH/ZTUTaU9xMW+V
wZxNmM7XTSyO2on1t3cdr8pAvek/ZV4hnQmGytiKrxKznHr/aWI+tVbWYBvxcwnk
5mu5x1aX1OC/zfujeAyuFApoesKa+vtnHmzTj33K+szRgnAYOTgxXcp7LpfAuFpy
HW3bJLB6LcaIQFKIVRpi/tZxlo72SThBMoKCIBpv4Xry9TqkUSpeHwQw3hS/RgsN
`protect END_PROTECTED
