`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V6Tb9cTqvdwtu3T1OWfT8Ka44eeNXHgt4p8dHiDdF8SpgsZynJGKrykN50X/X/+D
oE5+GX3h6Tf5nYq7KaWHUTVbiF8GS43atNq+J3mRw41fM3/3VxoqVzu6xmab4Q3A
amxdu+T7BF20WUiJPeZiythjZz9tMiLK6aLRU1m4DnDzysEPmWKN6+Ewaru4JT5Y
ugG7z2xfa3TyaWsdqmxrfsrzcegv9tYMsk/EEKS/eMteVz33LUk/EmOqNoYvvnh8
FSsrcdXrCVezxup6IRJdyKdjfV+bO3x04K6E/tkqXOJaAlpKZxlWNoZITYYAJ2Hw
UUWSNEGFTehWDnR/NvayrKjI/Y1/P7R+2WPn7zBU+gZ0H9Fn3CxfDxL85KF0S0xL
GpXQvol9eU0xmCDEgxRDnzxeIAD2l66TRTSDxsobRjtXBsDzgCYhK6m6GJSqkEUo
nbIBw/tjQnrKZeZ+hQsb4fI7gmH+85P2MkbVDVy9Gp9ooea0tXj/F1KDTYxqg8cF
cpFrQt8IJnqwcco3m7vAgIB4wDFJH7K/gg8uMO8jtuvkxqgf3F8qBnyqLFBVvpyt
dVWq2Whzkqs+YGQ7Aj2t9HwgBrdd/ojDRt5AqWRAngoQn/zUeYU98/vdNLR0DrMZ
mNHhgYgWlq/Fkw/jg4S0bjY9iIhpNFpQBUFZGlf5Tlj6kqs3rXeN77/YOfHKpx+z
dfhpZaxEWtmDijwGfD1wMyL8vhA6ckfy6fLXRm66TF2To6EeS0pXIo29Mm2te8BD
64bxDXCp+vSNjin7iyh4M19nUcHzrO+DjlUUpy36EOQ=
`protect END_PROTECTED
