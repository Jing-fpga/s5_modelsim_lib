`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NmSA+t6eRxuq9cjv7sx9qDEuU6NLvNvSKakloG/HcsF9M70CAUqLXzac0XDeunYh
Ym1oRNJ4uqjyF8p7nHfpo+e+A7d3T9JoXjl7Ab8NySPIEsij/9CnQzhlEr3oQLSZ
7J8Sr5G3t0WsOTfLsPRBg4dvtQj19A9sQnuaj+8efja5r0PO3ulGdSP91bV4AMuC
PIddUvf8bwZsfjkil+ZsJAGecKPUNB2JCXJgPVT9LyCdEs6kEavD2uiW/77majl2
sWusaGq548w6u6XCYLw0mYwk77xvq6zYutvSi+ybXckWsAOWb4twZeactbzsrexl
bQ7UBMELh66JKFocDgdz5V4nniiASNmEFow4g4ULvMxxSB2aBDcFtzbG7otYiaEg
f+TNeoEwKYW3PKGtm5L03HlCWz/mTVD9PkS5gNSHILgK58N2dgO+bClSPIIapAyW
h6nT+MYijHBrIp5NXgZj8hWEeHrmtWHlX5TeOaoUmSbKncd20TFg278XHNoCaYOD
x/JHWU7BlLJn1ans9NFTIOjIc3begr8znNs1CqzxiDvlcENw5Y/4Ne+0yXVOvbZI
eSMvDW5om7JtbWk8VteYp8GzuxPLcSttMMVs/NwAmCBRbB2/nfruXqb6YKWSdjlj
3wqv7KxdsCrGe8YCq/w6A2Ilu0vLwH2pd4A90P9sX8r0C4AbyFV9ACM1pyTbxxHj
MHIWU48dArWEiB3j6Vj+UNVdYMEx8O3lnxg59Ne6Cbxa5cYzF2KAZLO5EQQ7I98W
`protect END_PROTECTED
