`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qm3V60xv6sbwHGM8ci3LdMrmIb+gTS5+ZnnFrSP7e/rMWCPD/hJfhPDyuO7xITn4
TNCdOhmOvEy1YBqhDxsy7AX7NDGfR9MHpwi5R5QuQcC1z5F7VaGbvt2Z0z3cWC9S
uw/My4f9Jyk4+PRixUOUaVLLbyGhDCL28Hm29G2Nmm/KcxZa6RtEnACl4aFaLoI9
5uGSOEklDCPfdMw1FdckUmWghvhSfHUf4y15jcVqxIHPHz8cpclM3FOQBoXpxJEP
bytpZaRbkRCYxBi3PnJnVOzM5VWrZkxnyNMzlBIsECesUUDCEKVNkbX8EtSf5g/p
P53NAfVZdRIIw8M0UD+jsea5DVGzZdQtebK2AEe7cvEG5fe9rG7QCPUHM1Hkkmh6
cfWQH327mMObBs15dJQ6Fkk07LhU5v2GDH2cwCq4w13dpkWSMIzdCC+8/yiCu7z0
NmHjf/j2PhHBN0+xOYlHnPBhuaKySuAX/AkhRv0mPbJjvafIWLfU7HtvRWB+ldBO
amd8ZFtIiHkOku4uEXEsMt32AjWF6PHFanTctmYN0i2uVtnBCOVE0fnJpP+fqjsk
Pr3ieWx8EbbR+vdOnQhlLgwQ6ivGrKK9ECqKlaBj4rPINm1ZrRQscB53Qtfvy1lE
KG9vvqGdLHKGn4eapdJdBIF7b9y7K5FlCl0uwwDcdNa3LtXsRrOO0RMViMazIWSC
vtJyMHjq802a+aB9CLP67m7LQ83F+Rl9M4J7EyGTEuWffzpVkN9/YpGbmlsGixPS
ArbRA49nZf6SJSnjNfrm4Edi9mTa1FCSWtfqvdUEPq8S8ESqSX77ELD+DCDNT9zR
tGtRe2+DRZd7MM23Jg6FMnXIe3YakbE0WQSLjepH5zz/xeXLntTg3pTy0UgcYg0A
eS33zmgQIUNNXaYId99sSKWVHo/CLnxsoa7+MMwwc+AFo+rTLkvuz2g15pQdbRGR
VCuP3ZgsK5uRwdfAYZHv0O/ngXZBtOFzh/IaiPAD/Z7QvxCyJq61e+lssLvOlZYh
YvTE508FAT2MSXN4uUgGRmErQD/hXIkJLqq7EBv9C/6XlxZJZaQU5ZiKzJPofWZr
15od2UlV6BxbUCs1jF8nyDsocRJPGG6le1Edy5YTmaest6+Y6bk5E5IV9nYCF47M
AswIlFr64EpVpsHrIQffyNZgcAOwnAcwAX2wPTPGGrYAENWFvWG7feWRHwaFKBmF
sx6qeBWNSpKtwa2blLTV5HZZrNMqApxM8uReF5qgsf41Lup/mMOpsU4tCPJa72bU
O63/8knh95Me1bxKG8/Igs2JKhPRSIwGEVtTNrzYfecYS0avy288WR7hk9cBOwar
hNUiF7wTrjkVCZqZlBgFPZ/Fm1QuM+kisHD9GwOztU+KaVdB86YTFhO6EMxVD5gI
1zzPtGeEiJ9bOB05nhkz2oztWQZ4X5cBL8/igPiaqRio/qFTCaSfgWe7e2m21LrW
7Z4uCAI/RMbGbdifVfh5q+A0oR6cp/TTgKbno/l8QatJC1+LxbcfCEpgrmDLyw/4
tDwkZgHgnCYUyLnKrfZyUYaunUSggrD0fc27dalCddUllfAvhvMZt4AcfSdD8+4z
7wKQbWg8zs2AvVemV6EqoLp2bdWxqvp2oepMa7jjxauWEvCXhW7WM0hsrbKCsXbz
GRYXZ9FjVuv6gaNU3bjwKwMYQMnxVsgonTiUfDf/la4mA+xnpbSZ1rGANwVYe7s8
obsIFDyAiuxWdEzVenH+F+rAZV+iPZGvvH7INebHkpzXh0kZKL3WQhbwYEfMu4g7
/jIlXYnJ4DzrU9PyZz7thx0/gUfSSAJf3/POrFiJbGi8yxDI2EEPJynfauv6DxZw
nCp76C5/+ZxTfgGCSeflkUqEKc6hg3En+wwU6bQWWgQ=
`protect END_PROTECTED
