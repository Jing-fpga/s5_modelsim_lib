`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g+pI4FNmXvsjRi9cu1dskVgtg2QGA/7jzHmQk9obZrJTLLu4iq98+2ZpOS8WzT8I
+nCsgp3s8MJTzUX9c7Cp8DvFFpkZ+IuLAsknANUTxe/5trUUU0CAipVlD1PedMln
JRfGg4BwIH7DXKMo8TfZMChLSiHEQgZvoQMLcQFeOl8RMm/w1K6zB7y104a0f4fn
h/tkmu0baZT1nacko+HGES8WvHN4CLXF054nJ8KTtCtvouHPmCnn2aeJt1EoqmW7
YUq1vJJu4vbkya2uhJM1QC9zC0JAUCCzkzfqL7AFmbocnmYrjLgKU9Y4dfP7A+KY
dJedXY54sXg/81JDQCMaQ/5GQh5jF7pd7ztoAoiq9iMFKFMlPOBENwtTXgqE4Jid
4ehg0Yxf34LlGZVTBCUHoradcUd094uG3X4e7fDigELFkzpsgXQxZGj+QMYxHkpq
VEO8u6LY/lieS7PMhX4JOY6iFdpUhx2xFsXrlSlFxYiNk7L0WAQs6xiMOkQEOuqd
UlLxfWqfVdp+wDrKoP6osg==
`protect END_PROTECTED
