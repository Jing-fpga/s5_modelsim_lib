`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
snQi0QsEvizIaMTVi9QTtaRevNCFNvTp2TCKi/utxL6c4fJZEge8Kr+NXUUgqfAO
CGfwutAoBQeR27zt+5nTxcx1FvM91RL2Iw9AoPCx8et01yj1fIWvBiAvYYwHTCH0
pD3TS/qv+mpPCfVyaTiklFHbJ1svZz1H3vtO2v/HvNQ6qV/seRqcXQ4qT6idMpdd
IoDSBFjQIOqGzXGjZvExLbP0kodDvzIPME7ZQo+hTialZwE5l1jcylu80JLA6BMX
/I5v0Zi4qzFQ03OeG05uanfyvDFnk9Ed3EwZ28o3O1IKde1tnj7UwsslqVwUa5QQ
BI6XEosZGyx++kPCHy6faQmhIme9CylJ5xD4AaMZ6tUVNJIR0cggpXgRpNhKg+tb
fF8sL2pJWqKRMTDY4l/9/YIO73oF1Ic7BG7wiIh8d9NOCFi/yWrcZwuIhcWBVWNS
zNQbk5mU7sQm1XrfD1cvZbum1SrvTC+Ngh/gSOBbZXIyyw4oybG1BDn1BPpMoITt
9Ll5TndydOnbv7tgggUPZ0Wyd7vKkzmwDp/SsMJG1ttbEYL9EEXYwX6fk9oTLBX8
JiWhxEVkBXDAtx/vfBRYsNLKw/4LQVjJEpAGPZMyVhwdqD+JRqrdc4dFc5kpvINS
M2RctAmy7wiv9UREVzJr/rns797sNu98KY5WqIywy0JWBeNe29gjZvDDSm5+uPRy
Lp+cER75Ii5rI2pJOgJ0ooFWFutdSsb/AeT+ec75sSLNHgdViKXEOLwOdg5uI/bY
F0XFNVd5p90/j9oA/hjsx4/oAfxujaHpBmu588+xqrrnRetWNZO0fya6KxK4yklj
WNzS+DaB5qRLMRKO98R86MKJ9HsYzWtel/dm47hlwLztWB13CHE6E54ba0oFyLWF
jha+JrQQ55t7/1lElAajTeI0ytw/Se7ZFh+A4HYFHJndKjQXQjaWwi7Q5/TOJH6B
9ui9mAHGMULSWc7A3PXdXaVeve3d60IIxzwYf6NdNAUAB2OrPI2Mn3gRiDsotyqy
dqMb7AAlDvencaXUvI83wAKaf8r8bpqYopzf59jqiXnkXRBEqdtH0o6Qolyppa/f
uVIIokvaqUkaC8yOAhnLgTzAiVYhkPBUJb/mufaXeOMroDnNekvlknM5jMRSqMOI
2ZNGStooftkgmSAqdHaVed5IeRl862QlJqo3TzOP8wbcvTdMP3Tj/8Nst725NdB7
8tFx6SWvDKcoLMGbUWxiCQvMfEYvQ8BseVPIK7QN9LRDJ24JnlmRdZXaV8fBbb/6
i5LgXTcpupAkvIcrBfjxTUiK4byTC3vzwGjKBdCUb/BN+GCi1GgVM+RK6BnFW2Fl
thpwmDoahmDb1g3fEU54u8R7EP8rlVe6f3Sk5RV1WhoNVuGnQ8tgHGCyRohHrzub
GYtba8ecEzmXzXjCbQRKfmrcfPfXOdyP0twciDlHrb/hgdcSWGU2h6ggDDWq9jFD
vzLbI+hWxec4f5sOTzjlLdJQ1rEQLYX5uYbjaoVNDzzaouZBZlri88s7T7X7VOym
ssS0gZm/FdhEsVFSI6Lj7I0N+wV4jKajw3e3a0bP5QsAujeis0WqvtGsFx43q+g4
u5kIG1PRYMTdUZN53xMCDaQ5pAstBrSL8YBp2JK/iJojcFz6MYrsPcD7i5kRXbf9
WQy0BRbE2Ny/lYiKt0V9/PVnr8miYHRfsF9baYWT81br/Pm6dg6BRkwAwQXZGPcR
np9BUymV1dhIvQmt/7E5mrM9uyd6qymAm3bH47CmYQtwhJVED5rqXpnapXgWUK+H
FiVfAQ5yfqXO8Qyr5kuV6bYqGdT2my3KpNeh4Y0DeIieGGNAbQXdpTJ2lM+Yvob4
IoKyjVTYfcGvpzmVtXP31I3zhQbb7kq8J/HZEqPOUzkROCByreYgjiiMeMuvMe38
CRWcFa3okbC2jxUsbtxDEoDaSJ7EBrYVCb60FHzam7aU2BgHjZHpz6ohfj0cidTa
cHfrgC0hZYWmyZ/2Jlp+xZjO7qJydQ44wjNSSGGTdkeZpizM7J3npXDxkTQoHo+u
AwVUqv5i4ZsTcWLyz57/Fg7ln/YDjLxUhSwxGZx2E/BZHqz2o9ALkWm6KRwWP7xP
RuZWK82IEWudLhE9mGrJmmliEgISn2h+DNf7pSGz91vVgrvcTxSOFcJz6/9UUWpU
eh9bL7st3DDuxjY8yPjkZlqMRX+7ZndGFtzRi5HEbNSjKD5vh8hMD3cDYNzLBdZa
xI8uZ9AWjXTREHzSx09uHaMjey1jvuNvC7IPAQ/xKdHMuvE0VkSYJbL6gIwmftcY
a8j29s5KlPn4m9szTWnjqbMahwhvbxL89grQiWrchDH2t9LO4vJFoEheAwPaBvE8
B2NHaQ3u2jn6PkYpqeA1fNgXA4xy2aF2U/8QAfdzbCuocGFXvIAQTiLrLihOGe/D
eCiipVH0gAY2EVQUUHg8giE/6yyVjZRtudu6Fm3ZBTv27s1CD6ItpUtrrazeW9Q+
16/dDRrAP1jdlq7ZagVwwVFEBOdDDRXfopnzcTfez7F7lwZ/LbNF13yLlQ/86QBY
8ckNSeuroVOM84SfhU13URelhmF/m6xxlYYBMjuHhVcT6a5BHUX4Q+pd18hIGja/
dQsJbQJMG6MSLNIHps77MLQ3ZRRdAL39Z/ND9K/KrOotj5IGQlp4U/XKrI4bjYzd
xEioll3kSD9f5DViGe/dFNCjHl3mXe4qQxo974rD0xR0RSlCY7rJyZH5DeEK3KJk
uA+PQamUtK8lrUgshpWZrvvit7XeK5upvy7o5VuXUgd8ARaGr9G6c0P09zi/4Alb
Hc7zQJ+CGJjzTdkIfOib2fFfJUHqkED2FmBuwEuhru9eJOpOysCLTFIjMbhUDYHu
pd3fyP4ys3EVUXfjZkVZngkh0OrEWGAf4rlZlfhoxVfFEUToqRfcE+EN8RpyCNL+
nHfFCC6Ycv3UiPlDyfDmykupADVeQ7gUjaDbQPEgMPYxPXwtp9eV8+r3fBfFOAVD
q5yAxUkJCSTDfCFZ7yu2e6eD25IkyombNCkBhQgF4Vs+3CcwbNT+Ros7ZI7q6m6A
3qw1HRORb4dVqSY+Kzr9YqFIvnxFDwDi4CyBvr+xDN/zW7VtVPaBWrZmLaP0ykM7
RJwTh/o55MmE5X594DtwXfBX001w9p1x5Asxx0bnwwqFnru6oSgcz6R9Rg5/NIAQ
z50wt42Xvt4FDimgnNp4h8avL0+LC2opGcdaKv9fe/0alNZrqWTrd+Pe4XRghyKC
Z4Zf/kO5PFb00cz1nYqiHCo2iDig0GqmPOx6Xy9Z2Y9mzSEQ+1gk3KeY0iVGUhrp
YLIupDyDVh+gvfvyCkX+zSe7We3O6CK77shZ3GdcBeX8T30QzC/l+TNEjWkPF87P
M40AgzThiRqKiYcj/+lUknVO7tQshwl3mPf9MV0NlwQ5rUJNnayLFXipoMPrfImF
KiF9KmtsV2CpuolpK671CJwleAmj/ENDhP8jIjHpm8xtW6j5mi492AZwtqtH9bnb
AgmRlllT28zyOozdFMUFGtY0NSqBG/Qp1BpOYuNnkuvKrwSMT4/YV+XvN8NY7I2q
dPCUHonClsS5ZCwEQcKJR/uDtOrkB+pr5Y0RDb3yPwnZK9W53RJSRFRdKs5pYv7g
V9lArfMVvB358L3MWafuEjL+2q7g2bq7WAyCDAn6M9qNFD9eEdPbhoVQuNQ8tToB
VhqN1CLbcD4llMAIOUdOmkyrcyM53Myd5W9nLslxgEuXdpCdeaB8gB4WpWZw2bdb
AGnTbIhvAX/ATsV40iSia92/0E1/DZBaTG2Bag37vm0majCs/jMi/du6nfx7OCaA
ABSbcq+ZAHeUPHKx8noE/5OCs3N4dpPR3aKAdhjdan5dvqNgatmSJkYZ7TFZZ0Tn
yMpoTAQPSciV703ULvXDnpETvk775zJimArUUvhT/tn40v0tS1xcJF405WtyD/kg
OG5uKnALNEZh/BpiXdD4KeKj8FtvbT0dKFWyt3nPofDFAzq38V3TeY3O2UbP/P7N
VU094+aqqmqNDVfoLcFn0uwN251GnMluLqm2a2p764QkP7E1misOsRBijuzV2+T/
zmMJfxQ71r2lbPgTHe73QaeCia2wC5Uy2pebHYlIe2av84A0B4OKBME0/goyd5Q1
MZ6mfLEhv0JQVO9olIFG4tFOEEcYHEMHOBLT1ySpWy0QXYNaP55Ud8f/8JK89ENY
aUukP+4tDst8hIkag67sKbutNNMmiaDM8tieBSqEIbzwI5K+/hn1OqSGJ16qsm0f
nawnEcE2KVxImpq9VYzhM/IK40BnKk1msIrjHJNGa0Z+AXZpdaZuvJBEMmqCHagj
pMitkfNqQqxVQ8XKE1lUs9qZVOkVNmb3pstSyUYwAsvFuSq7NeSHXW/PjE/oMB1R
cOv/iNwNtuu4hKliyBqmFIRD6tFAQSOiy4oKsvadjTU7rM9p5WOzThifAerA94nW
tMNXWSvCrlkvNyN0NEurQ0/vmF2T3oUOYB4gEmBrxIb4lXWrj9RbcNFFdnWm/Ke7
2x++IUnoJ2j0Jhfy6hCWm4bIyYOsUa25Th/rjAl3fx69aqBia2AdJAMOFuVYiT2S
MDLZdm9nyoCIS0ZioRkmRI1nnfGm4aBeaA255mpiXQO7q6rzZEDtOaMfp6nCU+mn
FFG6lpN42ptS24qh2t6H34Tb3dJFEQ5ALc4gUZT16WSU2AujzeIGVN1yfSGLJo9O
cuitEC69n0NG9OjSmZIFLen3hC9uvGObRhRcZaM1FmXAZxFoUQw54XKqWX2tBqWm
lb/eAqy5vNnGoIptLfJkzfFbKqXZdsY9Vg233h5JG9oXotPuxKyjiN7gP/OHsl+2
MHRcl1IZr5X0fSUmiaGdPqZxtNa2/R5NlX4o0PcHCTrU5bK4NUpRbAckeMweZbVs
gLoLh7HY4UToisP/6UPqk2rfwcWXRHspMqDKb8Y09ALBI083Ix9gCDOHYYECSGXb
nLzNOi2D7F0UBU/7D/yR+03iDul5sl1uTwB5djT/OAaB16hLFm0dtXG/qb+kh7b5
SgkSmhQnkTKPaOBpd6wxaM02udEz57UbFo5lK+pOHh6DhblunLWXOniS7zIA6v6U
DQNHDcZOr+Yl+nboyn2BDPOXb1sPGT3RTxG7atC7QauEaYm0eBYbp7jlvkrUIwWF
4mYKVBJopNL2BnuKPivGrbOpro+CaW2uwGDTIqDAVy6/GEYEKhiC5Rs+hsb3dQ94
/8doTIAzPXrlqpw7rsIxn2l/orjn5M048556faHo7C31yfVJz0q6bERJZ5RYJU7Q
`protect END_PROTECTED
