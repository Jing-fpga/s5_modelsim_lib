`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7oKttIVxya63SXVD1NfATcRuKcwzf9LnxgEl2nledPjFnIm9ttlWRyJfosbOz/1l
0d56INiHhNEzpGwy/uAXJMj327OHsfimJJJKkfdIc4QxfkjnTqZCgTKbM2QTCgZb
4GV/Oo4JpCTnJj8WplUjanqgEaMWKhmstEGSOYCB8j8TuTnFEGxyFAhQuAIsyvXW
ET919bdJIlDh/bgqyN06tvMiZtTcGz7NvgZRPwzEWMbGPiGC+1/xXa73HPgVywg1
IWLw8ztLWqrreKcn/drX5hqO2OGfN76/H/c0rgZTICcZYw8eI0tUiWIESYcVAOpG
T/vCxC3YrTQGMH41DFNTmiVcqbY18C14QvNUx7YUuFCNCN+O3K5vpL5UNnl6z8sh
ZsQW/LKQORaSVKfbIviJNAxk+0LMDySsqem7QmEMfRFU5Q8W6A4QCMhCr7FpuHaV
bWpEFYuOVgUECOl9C1Vo+tgln2m/SFAygfKlYZv2F++2e54DipkKVLhsX71VSSc6
Cm/ObBNFtklEWHnchyN8K5egGFIJhPnAz7GyZXp35ieYITET4W66qRWXnqNX1Xsv
Eb9B/uKfrY8mpOMegC08dMaVejIqIRfFXGzH10DwflDQKYf5X7s+J8qFVDoo6as0
+qmVR9Vz+cPMzPmpjuyJxTALJ4a8KwbSs9QSNQ5MxVYr8KQBQ5pZmqvPKIckCggb
PnnpCE1LRPcLrUhRm8jtV1DYV7I+k6KufshXuolWhk/xCTyM8DTvRuyUiWjZYOmo
jevmB43cf0IfoOaXBXoOegUpa5T22jw5r1V/bPqCQKrMa/DcJSDaeFtVzZGqcwFx
pjWmdefTUeSdomzLuPYAgGc9q9dWQxyNxGm0OvB23bh3SBp/Ssxgh4h8v2GtN5+K
UnBPFfC9iR6zTMX7IvlkWEgIBc+MlYzXkK6og4ENzRSDGorOxVKT06WjzCXOc1iG
KG6WlGPHQnTqrC+2ot1nwgmG/JLkDNSgFNIr2x7EKuvFhsH4dVO2deHgv6NySPXc
GDOJr2a4a+HBv4Uo6XbzBhSK7ESXZ9OcIMDCBWRzBzwOg/Mmc1wx9MNK8NXsePwi
p+iq9yYqWqNpmQ9jqPYn7EH98Pudci8youtkOSaPp/u5eZJlQ/rZf7ikb1C2h3dN
a+k20wsV3bf1kkxNHwJQz9xcy2Kn0louV25j7jCDRio3jwmFRN2bOgaprLFDGyor
vA6lVm+MtOACoSK8m5UUY54it5k5vTl13xlW2JLCsrvTboZM8F78nZAqaxexqWSM
g62kGfHJmNFHmWAxRJ/pG2Mw6wewdnU1ReD/kd0O4dYUdoxemDCDGcTnZ2QKUNc/
CEdrekp3MxElJ4PwQhYVDnbKUkM/BqLIIXcxz4J0yzQB5G/uDPfSwQ21MaoZef0R
jFa0fzfKb1g8DrZQkcj7Fo4fFdS3ysK3gfN4VpOMbytQ9ySUJzv153KmEqp5QcUI
2/pDVTgolis3xcy2axBCKvWg3Ftcrcj7p6q+9uMy08A9urPfAVJAl5XzdQPBa41C
QfddHUvzQmKRTMUdeN5+B24Smc/UEYUXfIhIKEmHJyAJgf1slWHNN/JaZqLMvOIv
f8tKrQq5T9oPIKtomHYoxgkq6m4JrnFDS0+R1tyy4BMiE5UDPsIVzn9v0XQxI+9p
hiLcul0BwuC3MV4rDCsgUkb60KiJ3vDpsHeGsdwTXdseCHlLcKbufUlrxCf807J2
pvSnoPidk1/aYdQttVzqtaBdF+sWwwVggq/J9CaCf6om79pwg2PDuJyN/oLeHXxD
YwM8Xd3+JRvLsWdZKnnlXJ8CeN4sTZo2607iufBtNICEg4DZXbyfeEjXpHp+sc1U
dn1KWwL4pI1WThjrDcrO+QfsI5w2pRBqQjei/JmopacnOqCHacXf530W3Y0pjyWQ
K61+CCNgsguiJ8dkzd+G3UuT2Y1p8FOSF8BiuqhY76RZ13w4k6xwS8blrD6HaQXN
bybaeeMhAzTJk95NcybAZtFO3hykJEWhNnRgK/TfPt0RmclGUxlatpR+2LBHzF9k
`protect END_PROTECTED
