`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+mIwmMWRvU51qPe46JHc7p4GEIC4l8Cgi8j9YU6JYEf4r2sN/tiFdXEROJRn4Ixf
aelZO6Hk6+p3qqhUTiIO7I6gp+Kd45TbvmFs3jR7SIZW2AfiJVSA5WmJ1ucN1kcq
P/+IcVTrQtcHlxoKYL+unJkljSvAz4A8B+p3cNU/8eveGQjz4bVvr8BzqcELPiYh
10/tTs5sI4YvWuE9GlAY7pE2PcmdFbw4IDwNaf1qpYPE/ep895G1glR77TVCdkNj
q24zYVOjbM7hMeopsJuQL+JWDCCuNr1b6MLigN5I105pF7QiwYDas3ZSgiPKkQb4
97bCnrBfdwd6FOJegzgi0rxMMYvLbPN87AKjJO9oIr5y4trgBFYFJzK+Pk5kB5oO
fY3Lz3EPpfwOURaR8+C0RvH201ikh2jgEDL3lMjv4y7cn1Tp6gkyocvTiaNbW+JP
coNxfx2DIlnqz2b8vbR8O261lkextwcgxe1ooEv8pkqGZmdkSPhMOyqy6Qao3LGi
RNnqeracqJXhgU0nfLsNvhL8ioDfkA1ts5r8ykEp1yXPyPwzIh/SZeFgw66wByQ/
EVqXN8q02sK+dzixiKV001nqdOqBxo3A1O185sVdIm1GRkOdwRB5CJPCLordO28Z
1IP5eHtNEW/eKKmI3ecDntjF9oMElXdYgAiaMiJwGC60kzJUFoR1tcI7fmbm7v4T
qk1D0zsBtfgnq9I8jPG9gnyhh9fEC15m6yfEinye6w7FFTGlvKZDILLt6z6w8pTI
hXARLgrl06NfcAvjrBQMP8n4thkymgDGU4fIN1x3gX8i88s/HqCgjhDXNgdGkLvO
uGmgkdRElxQ0LQcDsM3/50P125KU8AM6p/yUu2mTD4TMBeDl+spPlShqyi87SDK3
Crv4FyYzJWWFyqKP70X9a7StJ5f206ohHSeu8NBlDE6KKuy3oejGhFxGjKwweD9D
pvUhuvaBW+3HetBY/QNu5eW2SqWozZdOYJRfhSchsHG8rkLdqaWv1bME7/x8IqQ2
WYUBTIyhOrsw8dzEY2KuyionqAXyGtqwr3B0G23KbWqixTV0oK6UXbSfFoXlc0JC
+riOaZe/w6+V4uYe0W5JwJ4/ow/N7SoLEe+D1WeiIp8JzvlkG3DUG7VQxbcLEbm/
vBq21hL0EcYgj5aymOh/4RA4fYohYyaD2rhk8Xfs3di3wCeucizWX6D8HrGUQLcJ
Y6gzmMVOKEenKolMAiJrbNMGduRQpD9rGmYSMSZn7q+lfq5beMNI5ZTf+GXGetcQ
fuPFJ8cDM3KIodASjGqwfAXrEi0M6owiam8A3rOjTduc7b+Mj/TcDVBbzF7RirmA
Hn6NZ/5f5LzfKyoj/lRvBJTnFL5Ot1DPZOzrmgUQv/a/wKDq2j5yfmbjqu4RmUEc
my/qjjBsivVTqhA09CyMMVjZ5bzHLlwJwBubj+5oJiyMCCxpTNrLpt4eGp9BVb7Q
RhHaaOoZX/oiMrHPjIgK2NjH1QrY9HBM/uzvxIv3aS4GzwfWoZWQBY8JDGrYg4Le
F208gYiMpODG7dUh2CbVK8Mxb1JLxW6Rfm0mHFrCcWu5ArTp4MRPjPBQtMTygErg
C4UxVPRspNm1LwY53VVA8jjA1l7yi9jIs3c1O8drhaT5N5pnTda/Kjrmt/0BN7lT
xA6rINEPoCFfPFgtiPHxP75FI7wwNh65Tg2Fo7S9Xbi6PnJCoTjiTV3OHkw5SvZQ
KZzp5L9MGtunmIEp1b9RezORj7JiNyXZiIGs0hCCvyCm807J9JqvtSCd4oq8L9ne
jxqEXnmb0/w0ewMxn2uhGH3lmupsKGF8D8ijY6Dn5/Qs6yqtI1FvOrow2by3ZkgP
NGEaVJrwKGFTLdXEZAIeui2dAaR3TnJXxobVBRY8l1V6KJ/CRY+Fn1Uu+QcYzB9g
HB95KEX+tWb9rPpA2ewRusIrc6SdBjBnrQiT4gFvljLqeoH02EQR7kfE39dVm3ty
WK4gxozD+bUaxDsXJD/y5mgg8cLFZNGqxPrb4a6sMTMs9eILblK8QI4OvANnk5GD
i7edSC8PT6ILA2fP9phYfngSPkC89vuSKOx/r7tb22gHB4fnbVRNVQl6YmPD40nG
kuStpRzH1eODRXB97RSRZuJFVd7OeHN045ALxOXV+IqCA5XEJWHDHtnF/+WjbHiw
Frx06rEIXU0B1FPEIp3KbG0KKmLpnxNgPC7iyuRpZVwlJpzMOTx+YD2Q5FuOzaV9
dNCTyY4sm7HKlU+L+ymLB2GugxMN2jSWqA7EyFD4Z5+i4dwmSa2SYoA7beC74+Jw
HXsBxN/LkfgWx+O6u/z0ZuJrsjAlXUfsLyMm+j8ofUrvMpcnvf0T/YZ+Lk3300dF
p50ucwkd+J3SZ0YJKZL1JY4ZxojUp7WKhkblupUirG3WWwpoLIx+rwHl6oUdd7l+
23q3hLeWnPBGJzcRAs2RmleQVd9fZjRd6J13pcL5ZFlZpdu4tgdIZVGTfcw59ZR0
l/amXZlwvaZrHmA3hk4Zet64vy8WNqNIHnQIesXyZgZnNRZTnTfCXPirQ+l9cB6B
XsjEfh81RnvRl+NNNoX2f1fPralY7mVHsKLyExiiQWD3IQFz31fpI23a0T4bqqS6
D+Mrxv42ToJpzXdYqzDcJbd2ZCop5DwPLUefIHLPmiNMS2SBZe7LK066grjjXxlj
FB1N72wnsRaRfLDiE3D+5gUzq+uX0hZg/uO0rtSMA11Tu283lT/YNtcCntOECHP7
Bj3AHzsCW9Tu9FC0a8Mey1WK4vb4kdA7Jn6DdM23V5YWDk5KNQB33Nd2f6jv5sg4
g6VgfqXHOGf17dfN71RGk2U2QEHhwn0hZRUQ9WgiJ4qOpZRhGbqalBWUMAlb5bg/
Iu5iqKQ4DsJ0GI43hZsYkm91itsqrelSBzpQaQYionLsntcjHuIMON2S98klv/x6
cMhctiFg14gjnkYqupPahee8x2ByjaZ3sNkw9jDhAZSsGxzx5DndMP0CfUqho9x9
a+05WU7FjzSlKIkqz4q2e3nbv5UQOeeAjDTNjSuNwxWQpglj3KOsZx8ktLgaLJnd
MQGUHsacBgBggmi1eppS99Ei6uuYNWZdGFWZQPJlCbBzxtP6ZBEDgV+w4tJEBsd1
1c9LsuYdOd6mb2OpIAcEdSFzdi2tIF2Nv/N0Hl7qOBXVK/po8XsZH2wHyi0Gk8uY
02EYuFksTX0V5LLUbZvoLFqcubT3D+I2AwnSTYL+BQOUwBXE95BSdag75zrwvUuz
GAgfPDQTQPJTf8b+Ke92dR80IyQeAmnGS34XGhEJGOiBvLdxH93CRfuwCQXs9KZV
8j4K2ef5QffhykgcmsA3pFzfm0Cq3eqSw3Afz+79/DB1cmnj25rH6H2qyXsq34Wu
uqiIzVwJJX5OsMWl8CauY3fD5NhGk/RInQ5RLPprYpRQMe2x3J4FJFIR01D5JJT1
ndBUW9sPWZqr2V0SXiZXsqsRWhhA36uv7uZ+sRVKpuUvi+CdEMt7VACLTYdWepq3
2yykxMfuyDBrCBH6FBcf6rJ5tejYTFHe529S1kxn7v6Z4U4Dl43b79cvpymo4910
gSG3jOdG05gaZxKMpTApdPYv3onomO2yTak9L/LuI9yY7p3Ay8wRVJ6vuwxFdRUM
hIM80Y3lkpVIyFd2PbsGjz50IjVzMsnZscDkyzOf4qGH8nIvGt0D09NzdT81bbQu
BT6nBZbJoQ+mizC+xrU7YcplV1g5eK321rATB30W29NwlYQbg27mN8WTxQi5z5e1
6XRsi+CUmPG8J6Jd7crvTDcdeQb+i1/BV+M77ZFXYiObu7Qdsm3YVdxxtDPJwhvP
HXpjOhY8bMHaErAZ5QfLvIw+vv/79bxgVDKY+JxPwFmlzdFNPU8acQMl1Ms7bLf4
/MKv3dSE1uIGeZU4aa98JHu4XI6H9ZUS3Ye5YFwzt3u9ExKX3Ed6WheyqxkluG6U
1+Q78V8ilg96M4YvRAuLzlC+dqFnimWsVLg+5QMauX50ziofwHl1hCPvXQTyJs26
EXUIYd7Av/A9x4LlxND+6A==
`protect END_PROTECTED
