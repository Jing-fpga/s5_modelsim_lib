`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l2xGeT/h83xDEMf7pAziBfMlnXsGNOr1d6mHJYgjPJyWAFb9XecXtNUXKZ0+Ow2b
RdUA0V2DnOugoJMVQeGrPEr/QbatPahCGtBY4R0dUWYlz/9qLZJo8oMtOlGs46ZI
z0XqjnkBkuEtbVF7yh9fh53Vx8jWmilppLhhWOVDDXU7SOhbarU7YkAhj2Ea8z+m
36H4ZjOH7Odqh4hJJAOK12OPWeQtyeLllL0CUGjCmuydCqhELDjSBTwPuwnM80VG
crABBoElyBhBplz07viMf0xyvDx7wGwWuvBlykA1yQnoVRX9hunUfEHmz6DfD2ju
YvVhLgrn3r5S2ZNPmlpT9k5MfTrh6Eff7V3GdrhciDw+bSYwqZi9sOZW5t7E1y3E
Hn0YynRn+a6hJHjeuQiE/Am1ycMa4jZMlEzzakE8cFeZJSN3kH0ATlVD06lgN17H
6Yt0/Lz1jrFyk6vuuOgg9jElykWmJ5KpUGC2yT7X6s2RJgHer8Jgv0aueKwAnPTK
29X2c4/BFfGrYDag10d9ZH6NlEQEhYKcC8V1fiB3FcE5m+nL0EzJsXvf1n9VCTXQ
8IB7lWB7jmbRLlY0lNlNtwSdoBYHITcFn31/TSOCirrYfHbK/sTT9KAOSvu6ImGs
D11cozWDOJWZ1jWA9y5R+2jLOdXpPagx4v5Pq0YJH9sfyZ0rikKrqcYCG+I6LYLC
DFPPHF+RXg8erA2fqFX6o1GsbYYmSS86k1OZ4wB5IyzBcchLeWZZGUUi/eTO3da4
cvFd070w2xAtw6U/Yv9v9G5O8C4EOhPVkS4M+t9L64mZJhncssuji/sJtdcpRIGd
vEGVr/er+nHnJ9vsiE9jvVdaBAAyaI8a8o3BytvKgICe9F6/wxjgnr+Y422ZPfbE
TXE4bAO1B1MXAFtmuLjX2vMTL5SAjsS30HJh85xkz2onYYbH9ucR50rM9a5b5iBk
GsqArDMOcnQXf7dUkeHVEThhMh9AWZQmXl0ig7odYj48qiDDDrQzM5/joACIeUSy
sDZkIBcf7+Y5qmBbOAAKdw==
`protect END_PROTECTED
