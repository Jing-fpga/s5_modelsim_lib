`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1QkYcIlL2GIXMjQDwWqeSFJQ4F/lhVaFaJh5+L8egZrGfSse9PSRaXC3b+G5gRQg
xArEszD3ug/03uFKJK6gBQ4hpocaYS6OrZ2GOnt6q/j/6N4bgUbecMSX/MnKbDGM
G61leUwJPWuRvxJOTx1y+UQ19CMEkdMTMjUnemLKsuqP1ZtHtT3a4SYOVYZWpATz
5ZXZ3qBexGhy2B2xMLE1z+SvyPjsCm/iuItlsoPIITXu07zNUHxi1Gy/qbUFlNLo
wK75VOmiDDBOk7bVUL9FSUnFSJh/vbivBWhRufv1cOj+l7BDuxKhx4ZDspF4Gqvj
lTJZolafXuxS75+Et/g2wRMy9yQL2H4wL+AQ9FbVx3kkGx4eFJqFWcU/oyL+5rHi
Q5+VpoN8u7Wx+KDbTTpZMAHuP0BAVuC7K2OiRMStnck2ZM7OIqC0z4xHUp/m5i/U
nJaHFn5ppSjfZAZWrqr7ywEla/dUElG2XjChUZrYIsF8ixsVlN9Z5ZFi4GlcdCxb
Xt8vbfK52QvVNbyUYTGmAhUjW27F0ZdOutD6DS+1uXl/drXANbIOpVrfEnfxmCuD
SqlulmbSPHWT//aY+8usDJseIxmp+7ugcr4n33wNY0MgR2PBPUNfV7sl5fI+jAZC
r77OGw57kpCHt54iD1Aoh7lu8DV6CLYxI1M5ppxDK7ouOWXPS02DTl62DCok/bk/
a2Vrgh9B8+XMl+IX5HH5TOt0LZf8iYQg5Ru1t9C0VVAs4oT3ZxnxR1WMnTxhyltB
YQkOTYIwEyfTyU7qo6mSC2fvvP8CzJlJtaGphkDCddVlNTDiRJ4QL0dNLtSAHUhW
AxYlCSHSK5gypZWoa0EQRWDqlRzj+6t6V3ZvljFwCb5K+9B145K0p68XGD00RFJP
NG2x0gBDY/9ma8p5rTqriSTz36XcHrwyHsqiaFlB4NHUFfpEExhEvWJufHowaIXF
T5koO8IzaNMJ9x6uU5yvqgb/aMRoztgg5yXlKgCS4GaqyQBBF0OtztrH9o+W4AFq
x8+Qj/g1SO/Avfe36u0/ZzjyffIedpJwCDiCqG5qJLh1LPh0WHbovTOcAzOHzJgG
9ALvon0hA+tOMhnw/YnlpQ7StAGjiP7vhE4vDzUMI+EaEfZ4tYQ0TM00Ta3pNLDt
tCSGH3Nv6sQMSSv+frF2dbiqxY23CU2WeGARbzGr/1ctIX9G4LDtYCrsd/1GbldH
D23AdtX8/aVI+rryzUmq7DaYzInzuihlz+AQtq6wJW47ilOSABxdMa8UaB28a/5L
+YobX5yK+bSFRZEc3R336NRuciCUwpW/VlgSx+8kXmeLKxl5PQZ3ghu7oSPqGrva
VnY/DCwYGLeaBHXveFivP9s9MLuKJggv0UXRjc+O47UKMjiYKg2R7n4jb+fCT0VA
p5ca8QPNBkPfWLZenqANrWPLHA6I8yRQ7zmiTTeyZ3rkMgjT3XcgRi0l3T2vA6rB
O1RHUxL363AV0zeZ5D/C3I64Q/Wd6BKycKar+DK6/CBXu4G5IyrxFZdlq20kSK91
uGzg+Auze4h5xZp6JwRbutTRvo70R2TJSRQGp+/Q2aLrscVMrpq/A8aog9Ck5/IU
`protect END_PROTECTED
