`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ou18RyCRhi4ux0+2amuJVgUWTHbgLSj4ym9PBRUZz2BCSE9IOS8IFu1XDX/vQEHm
sWR4fl8JZPnZZn0SnHUopn6X99iDIvScVGiaDmsCogxVWfU9dsYsHMxQO8lcvpCf
lv1dIrPNFhleJODKgXw72HQHMRZPUCH4JOXTLk0oEYm+Iin97zqFRzyVW4pkO/Ib
jHidkA12ZwfZUELv0IAsXPKlZhNZbhZViNWgafRfrhq51N1rmOjBYEpFeVqmCj+F
nP/RxzH4I7ec7PT4Xki7QO5OmhZgENTo+v5LE6hx3L7iQ3TgQwoxwmzTILmJo/GY
hfK/QQpqiE5M7eCItAQ8CO76KDT4TXrpImVwcMIHNmIhJ3eFOTcNdL5dvFCh9wPW
OKgf1kyd2MUvGzTTOSA8hoa6/9NvfmFjUDG8SUbTQxRdIbwLSZAh0F26+MHlsZZG
TuQevbVxebqMHyYM26q0YRl8xRNt2AnZNItp8hU2Qn+Nlov4XmGb0gzPZEK00oaM
W7W5X0PvuihHciyztiXYbrgH5gcjj1S0dnmRZ/Dcf7ZaVHF6UQVwaTh4lnwPih09
UMMZMSoZXMWbSdVtsEfAhBdwlGwxwIdy60CgD8QQIZxmgqA0Znu5xXtAaa6z1h8l
4r7zc6RURVlB51iYeOEo+6oQHx4zmF+rJzDhTJWOPAoeEtlkFtHIyTPx23bKz23Y
4Sj/iZ+IJlQmKBGZRD35xZemPTZDdgHvTTLWkZMjzslP+BYYTJJC9C1vrFJFP44e
D2KticjL/B/iit5vPQiCpxDaPPyxaAKvoid6YRLzeAk0MdJ4pBgbi/PGW3ivDtzq
paEuB+PaVEJSdRzk6EkQVqe8AIjg8ixkgG1nFnRN9N5pCw+UajeYoZmU1FX7aJl6
zVqxHgZyXQcFV6RVR/HpXJi5J9zdr8anzLeZ9w+8XYyksgrs/kDXs77IOnULXzdD
txwkhqEBvT85PoSo/xarABjjXwzslVnEgEzRceWDAT7yRoFdMxX/yiYsmf2Uph+0
/ZZhSNc9fuH/z/RPk4ZVf1/0SvKQFnRJ4ojGeil/y07rJngBeXgxPEFLr/GN2nHv
iTyvMAXFBuWc3N8fVwOWQH7r7rYCeJThNXc1SU0Y6r5Vfq4tWflPBMpl6B+dUuEk
AYOF+cGX8V+oGWAm5JewinE8q4Uj9hcW8VSXruYMnIJBzAnmjAhqIJ7sSunOKeWw
u9lPf+oT3/+lSQQSXHZC3qtKKAisunePUjXSMPgdkAwveH95lcrQG2xbjIOrdDIe
R+D2hsR1NwyD4l7SpwIHUtuWFSd1EQzrzS/7B3G4gNxFLJkMTLZboJEwYajHw9V9
imKfRy9ShBJssk91ScslG5pob2RxoDe9SvmiR9nPIww6SSuTeztAq+NycYtSp8LU
NmEv3lgo0289EwjcZgHmZaZAvZOI4uaaQhXX4fF0rvKCJ0r4EPQWyiWJ+CKA/eq6
vHD8q4LRL3q2XQ+FBYh0I9SHwec1C5KGIdDLXws+pY4shdwimG53ewKWbjr20G1e
WYPF4PhjP4twImCHoW1P2P+dkD1cOtEP4f7OxI0aa9VBMQ7jWjfAywE9MG5PGZgO
fNPvV2X4uE4PRyxTNmxzl84mwH6v2mfuF5nmDaQxUNYYfea+OPFWYiMSJyv3cGvu
2RggVBfCpOeaiJAmuvgqcu9Ufh6xHLfdraXLj7Fbb1/fy05qTPFM0I04NWORzpFW
WrniKX56afz7rVD8kfiZys6mtlwfbEls1S1SD0l5BT37ELzW+tol+0E+1MRx5h3w
DMjLTRX6jT2pYcgY1aTY2UGU9SSde2yj4aGtSxjGaJdnjHgmagqU+k4hWCV9MwnK
H1McbPm71G4KwrK9bapNLDvav/+wBfzXE85JQGfUw2ui8WaPzTGHL1DoFnkPcuTt
pkUnNye/ooBNBnm5r8wWnDT9DPI9uDoGROktmRjsMQ28yvOK00XbV2DND82uH/QL
xcfBo/p5aehPgrXsmO2LoczpbC5HZrqP/gn/tzjwFFPJIz1o1lBgtOion0ramAQc
9+bLxIxAPTFR9you0531Xk58NHdtOpkXYhD6fXBz6zVCjcBLs/kIIBJ6GKHB4sJz
FbaLcyLnut6XV2AW/M8NBY9g6+cO3U2QmS7t2gnPBo0MFEe1CZZR6RH5FZ49qDl1
mGaGNRCbdeLKP9LdNAzXCys8TjDMvkVzUlHLArFZzPfMozUUs2jTs8/kPY475f4K
zuGygyUwX+d7wZ2Tkv3apv0r37MDqZ4+ULu7cRZZ/7nNDaFFCpXaPqGTvUKduzKY
RZ04UQ4pjyyutWwg2tL6LNiVo9aqeWyb7vAZeOInSGnJUA5eJst6VOTbLG+dGyur
A6h6m8IfacHRUZqLFBlWWm5zl+1XyfKf4xjtgDxStZ5EI7d+Fb5u7qjX9QpKgBvV
2Oi1EtN7jyx38meFldPw6OSp4+Fax/oJJ0TgJrV0N8oLB7r1I13wKmQxNltHBion
U01wZ35x+JqI6RtOQZcUfhimUtw7/j6IsY2JZihjZWB/E42g2LYBRfJ2U4Xi/rx9
3N/gKDzfPb+YTv60rbJbTvb0b/8ND9uud+L3LpRWbOSca7LK4Q0Q+oFNwkGv+GmZ
wRmEgXr7u6+zPO4FQ+jeTv5caKU3nWQRVww/C8RA4hLfSdot9lVD8D9BS4r+vk+q
FZ1gVsNRickWRvHUm/ImmfCsCNSxzcYfXK/OJDZ/JX+FZlRtrtgWWIWUEeRGJizg
PO6lOEa/hjxHGhlkem2ywiCP5sMiBuYTrXx1GqhSiOsqTeY2t6aC+B6Vq654dHHd
9EFWC/wJDLtc3WIiwkd7Vt9/EL4P25MhvEa7kiNhJN6PGC6ojAzXtOzPfZc1VRwS
gcSc+MV5MOB+1uddDgEOlsqnjlsygIVIWl8YhhflF2ryK8pgGdu923AvEmGb4bN4
lTwZf1CPkixh4vkLQ1GJnfdcS+VtS2md1d3pCpMr1eivWYgGfzswIKWr+CERCp95
FzstuOg7COXj2s1ORnjhMuoIh7x1P9VDMqt2b9LL6rzi/lgXCwwlSHMpchB2jEX1
B2D9TQ5hraaAa7de7TdQ/s6Dfcu7fploYoNe7D+/o5Hin0Q4PkdgRRugAlCOXbpa
X1j5irslvUE4zv/M8nv3tE8eSOq1/7MIJow7RWmoDxsfCP9//HrQS6Sg6z/mfz7c
N7NXRJ7E9w9V+yQu6ycFi/CzMxNvyIZnKipkUK10miafox00wwG4i6HdhAL7FANA
swO3XYb2VnteITyWJ2J33lSy/DVi/tmMbHpRNSkAayiRDCk+g8SPIZRq1w4sFFzR
Ylnh8uyF3TlK9YJqGcSHtx7hImflZSNFDwqv/bIXiIppt6EffaAqjwJ8xklfarJM
hQcqDFHtJzFiIG6Lx6Cjb4FrN9bqvLh+3NAAccZChlXhC0NVsArmK81JDBqoo94V
rKXUe5ihd3Lrl9JOxE5GtZ+VKDmXBfH616b/QF3emhRd/Tuhj4URW9E0QGFgPdWd
BGoP/vnqepcrbzcg0mVpPVIAwe/mTFhLycqggQJzm0E+b0lwzcnufmzBxj2Y8Xmm
FQUB4IlVBhtPwKRTEaOSgOOKPhDQzvxFoTmGSDTqrfJVbfXrsqztikzYbfEU63ZT
zAvJAvZC12+vuM1cKJUGrK8gwKVYd/qihFSf05QN2Whjff9UrmaSOYCo3bSao1ED
nuvEj/ugt5X4DQMk4YAnK2p4qMNdK/8obzluUGIWikGYuykZ8cM38O7chYOCybAx
fmzxJVjVwVGwdUgsrAfq1lQicwt0EsYHZcyOakQE+4MiQteXwhRKcYtPC6xGABfn
dVMAGtFbsg2at0/XjF7vq/AD7nWEDcM8OF0CnpfeBHxlkR5zZ3nUvZ/AiNajM+BH
Ych8RmkAxHApOuLidT8yi0viZztv4/ud9tlypSWwuXdtAwfSgnVI40jTSceIbiMB
EF5c7y/QZ+8d4IlU4g8+Fy2ks9vuSQD+jnQ8orJP/6guU6z7ylwHwnDq/OlZceTS
rzSOwyK47l3wdc1BDVHG5pnxN7ctRcIY4222yaTByO8xw5ZhizkLoZEVHmzAZ0b+
g9vUE4eeUdIBy+fM5zfDq8PkSTSxBc/SxMFJJAlsoZV4vRFB3+s7rxjeK2lrcATg
fRk75W0RzMzYMebeG33frm1CbBWZ4uSEpazgk+AJxhrCUj2tZ0dbM+XjlSYQMpEF
PbTGbTZsjOLgOzU4Gm66TDW+gHYE3Jtbhe23N1KDdGk=
`protect END_PROTECTED
