`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TFAWk190tzsbxqn19fe7TUYmU7qD9qbSVOYVV4u2wHNQ5E3tpgjXthidaB5WpFG4
ctImXwgi0xYi4b+KkDEuJHj473NlLfDye+KSA3eO/NxigbvDFE+Kw7DvB3A2riMJ
4Byf1V0s2cnGnU9YK40nry137mPKJb041TRxDzHoBybC7vY2PgqplFo02vr2Dght
+336R/W0M8pwBUCL9WVXIw/FrLWgaDmZAAvfIY2e0dcJbu1r6rhgIAd/ALruAWQS
1Az0PWeuZsEp4ePOlUIydPcxfLq5ZfUGCT+LnWGvXe2iTFqEhHP19E4dkh2KrDTX
gcdKOSxdxuhzmeFkza7UCZHb3dJNt97PcN5Sr82KV0p37p5ok8zTa9UL3FPcvu9f
lh/62QFHoI+3AVbpG89eE+fkBE9dRlR9N9soQ0qra/Xzgc8hg0BrwetUJzr0TDXY
km7v33Z5N707MuNqrdSg9idYSPHnMZROeLNEFmLgcaWw74gplpv6seH1kVb5v+ra
VUoTg7PQAHMfa+dlnmQ+KVAHcNbxKXwviPQ6nRbIF4uhOzL6+afpoW+gxc/8xgDu
/5SXtdvQ+OZfb2X/gDnQYzy8fs6CwPL2QYOZAZuhORgpfVmFl/JThV+K+sQHHMfL
/r9b6Lbmp93an3nqzAexUD4SdELtcMrL3JlsKL3SNBOmWbCVRzM20zAUTBY5+iJi
UlNVnA5LwJcl55N7lOby5+0lKni5hyCPCp+Vca0fl3ObvlCjLQ13AUF5aQCAZ2s4
RIlCVcESIARUoIMpV13qLiWYDEFeQWjZ7xZCiaMADJ+MR1P5VSfU5XsNCEY6TZoZ
/O6EeYknRwsMp9iNwWnDSPE8rXjzvAHff+KmB/utmvEtajrx0D7PQEtGXh/xHTGw
mS3v5B1PDqldE5qejKZRH7/HihfaTvbtwmtzRtp2ribWS17rAHKGLTzF/Vu1Mht7
sPt8bvfkFhxSv4e0NspNfdACDN9ibPVjGblJVtl+jh+ZK10UWfBVp8IV9K/EXDmm
ZnwnPkGqJBq6dNxj+YWF/YU0vrvPJTn21bXa1zyCl3/l6n8rT5ENXGnLWf/te5qD
57jw7rFwoZMtl1FRwUaCkoW86It9ReCQTdEVMiPSSv144HeSQM6JB2nrC/CnTXzc
pVx/5RhyJmjaIJRO6SZK440kjFbylpicbDEy5DB8EK41ZF+07j68SY+hxJ4KlZfN
mKsaQlWcvre9B7TzSCUezLgNHcbMTcwPBM6q1FSRSXKDZIBT5c8/jegMkdl4UbMC
OQikPNBEp38LbM6XF86pjDvrkPn5FVczKhsnrm5zFnM5DWew1L6SHgu1rn9hWhzQ
+iB15FZxyoMHS4M4+Zw7T34NoRpFZP4jT2JbllQnUh0mSfr5N6wswpEPYTVFx4Fx
HtouoY1ciAPNu3dpnVhnAEX7m4MkGNqXztrX0MSIc6XGAx9hxuc1yRPcUeuQR/R7
YO/qUyRcLWyHLXy/GkjkDX25P9MH/E0m1Et69dBDVkag93LpILtotlG5WaLy4Wew
kJsqjSlAD/xJNYzrxu30SrdpLahRcGU9VABTMaU4dicCTLuPUc31FyN/NxVO7ozk
U0Hd3FeEDpTZIyrlA1xRZO3icJ3Z1jjJ/c193qsP1H9yDx7A5x7YP7Wv4256rSLY
3pn1aG4HJl3sE7KIy2M1stKkrMrjokKqv7PXSnstq+awx/mnjx+Q3lXYqxD9wBVp
h0R2qilAFICQNJAy834CGna5buZMjfzkkI34SEsE71+e8lRNrlRwdOohZY9cMSuj
Z0lTi8r0BQv5+vxVSNcXUrD9dpI3pfrNgoIJKhei4A3+iAtRrKajD83nM4/GTAdG
xo/AAfC3VP7giyE02xrLmLWpwQndw5NfcV3wHsgVNRO+P9fKh4WaVBdBVtuzqQDo
i4kFdU/1IJpZQHsq7CsmyZRLw+2ORJYw47Kp7LXcl3tCeltWPCs4AtZsLdTj0uki
0JjTL9daer4hUYNloUZWnNIc6lFsqwvotQ7SwPfEjUE=
`protect END_PROTECTED
