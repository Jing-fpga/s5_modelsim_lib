`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LTsiIatt6TrV1WgvLGjh6p8EjPaEuDlJ3sGy+TF0apVlJNcoE0315nnmkOP8kxzP
LWyfFmxFZYdILqIFJJZEPkRg5ppsfJB84qmnJ5SvHEOEoNE/49nJiAlGQ4N84OTw
oBeGXTF+kVDYsjEJ1ZOYfM6VFaj0kC3WGINbhvGWZuXfxV3rvGkaEjpIKikELYzA
4AbRcu5rZ5VKBwOa22qoDQV1PYSH2OTxatS12yBdjfrVHzxD/m3aEZWbQ8YHzeMp
ExSTzQqkTFhBOsWrDcV0NlQelj+WkTfU/oo5iQ8klyyzEGgcv06Q7FcavU0pz+Xg
8eMmqZ9aL8bWZVzqKov38OidhGSFJ4hLMFnSkAxAisX5dTXNJPuYeM1pMJCS+xwl
XVgkVG5wBOY7W1eS56/BRxKxjWkSHtLutuY+OiRYjKgdvU1v6VbOQxS94P5N4OlQ
vOW0ZTzgCX7+xayaw6QgaVyBUqtxLEJzXTfdmqjPhx7E+TDBDrnMXZwVXfRLw71M
oI0sxRU3x5/GnYmDmhMg5kxYKJPZvxkv78EU3cnwibHVPG7wP+tc3/YReR+erFZk
2YFPuAwxn5gXloYdHqDZEfqgLzs2UyHAnaCLyx0QMPdhfELoEoV/UCfRwOWiiil7
EC/+X4gO0ePgPXP463jRLZvKwsWvTES4oZgWKegDV9h7x1/9tpvBSAR2EjfNRX7/
MXyEwptk/wrpl8w+7RE6YZ1BkTJDB/mhVMfLeBP780mq3bSpO9ObgusaOPyEpBs4
GH/d4heAH6pXYT9AOBmFf9gTR9eT+DG2H9b8K+YF+2gIdOL0LYTZpByyq36ByOXD
mxc5XBTHsNk5/NLho2pWTKUyOJ/xuRPdpWr7LDbSk7Np5bc4v0/HjD0L81R6Nk2s
hqNzmwxDk5qHY5FBZh0bdxmh/JbTNbFDE785Ux7kd+WFnxRNwCZC1JMvqH4JKkSe
sB9TswlnltlYxaJDJeSK+eVjzuXua0fhxP4t24w7O2anFTuKqXZaWDkGKc4VznEX
iHk7kyYtGqv0/xDvuAArvkYWqv/m3V8jaFdEp6L1TIdz9FL1LXLAeCg1uhqrLS7S
nVpBTW9nWr2Ni6YwRlchA1LTdQKmmtkP5nfqOpLSXwH69/IOHFFfIC56JP03LIkd
Ow+mYlqkkHRcnkUARr3T5rMJj669i1hWgngH06L/z/f7M7jMA2rrwF5sO5tGIWEm
Yy6eLIW0tDART2WQAVdJGh5TpOyVo7C1ya4V1O+8Qlg/ShO8ive4k/mD/lswYEI4
yEYQGk7T8wyBRQsyIAbkGDaPR9fK6qq17Rr4tFu66WKcglSrW4Jx+lxLeAMDGDat
gcsTir2A2xCMypwDSp/dA9blBaZ/dA+3hQxmZEMneGH81xsi8FK61+9MVKf2ezh9
hRuW9nv44iPFdJP4DSLQ+vVw4mIqsNluRI4cWfjwkKiulKg/WQ+20C71VnG87xkd
y5FMwxwCFDCoz1AHEPMDua1jC/Z8nSxy387jDdDSpSPPrSPc4L7UCkGxg2TuGG1M
pV6f1KZ9QaC6NzuQkInMcVLk9JttFgFiy/KGpM1lRHFHKa8798iUMtzocjElkuwE
MDSZepz56r1X+495cOrKYiRcqDaTH434fax4vGuAm7CyVsXR+UTK2rhfWN/SOyxh
07szwZVvmHzefXwKvDu9BlWwLqdTXL5yiVXyrI/0oEBk13QOZIXjGnmIcgKIIXEI
6dlltbTeah8xS8OxRqa9pP58MDmtl+qI4nUkjn0FWv1QYPjnJyDlYBmWTtFUhBtB
7Zaln867LZIaOR5kMhfXY6InXyjibyW+wKVlfgMWHLX4MD7rYPni4mcLKNGN3KM4
AQodyniSYcEk4KjLPxpLfFVajrCEUCAFDN9GdHbaNtc3PUevL3w3D0oh7p2PXgQl
XUwV0UwinW7QfHuKnse68HjhF0d22iKPy1YAtB6Wkk+Fq5TACT90w6Oz4Ck0Eszy
BgvN/OMjCxqK03UT1HExSZnZ9pvOYnVArPP+Q9ZLZPbAqNluiNXUhUHH49yFuD6/
`protect END_PROTECTED
