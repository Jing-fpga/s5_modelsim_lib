`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QXqOq3/Toa3YgGXXsJr4fgC+KhYyJS8hSqJSpOZhV346wz/vvokwLx9qkwgdgsp/
2l2Qqi6FqCyw2uywaNv7uN0Ms1RHqEiIyuppRfsN2rPrU8o8Kr6kIhm6FfB25ytl
86yuQhfhrj+R7O8nOV8uC4LHbH2AnLL33xnOxWykbkXNBlpPaVEgWEOlYfg0uZLf
jE3RwuKtlXSxJlRHrTNHM8J+Ga8UTZ5+H+i4h+souEiNj3MNQljO6wZxE+u/wu6k
25JWKhm9Vp5/7GU0wtNmhQIc41E48/xdGjKM56JzH5ejT+DTa4yaizdGtB0uNhDG
+rabBA8Vj/EZltvZjFj3bZcQoWqx/U1GovVox9CnpHhAbEshXzq3+8BWvScTQvBN
hu0akWhSmur+TQg/6+bmrSReqrw5RShhgUBax8mm4Gla7nvJBGoJw01UIVbn0iU0
HjZwWQu2vpufcFD6Pi9gnp/ZQJ9L5yS2wS+Xy1PN6DPEfkseUivzC6CSRbyqq9im
rBAcRiwkB8f9icTtYGRdYnvO+1qy8R05gejTkabH7F/XkO/gjUKAX+EtVTvznMnV
K1lp+SHFb+S6JRSFQl6cLeIuUvirI7tA5TOlN71dhOYsd6f50sa2wAq+EQoWzjA3
kBEM9NUe3S1yunIs7cyMSV2z+LNKfXHvzC0BSeuJMGcq2j4p1hLgWE/unO1FpMou
s0KTHg30eVA3FAqZqm0Jq1foFaJ1oG/u7UX301LiO7Qkg4EysTK4QJahwOk+CMDG
HPDNu/fgV9i6pwB8HW+4ecgIX+7ieiyFMulnwV/1IXR+m7EF5AXYOnMmrCDlBAzo
BXX1tK3qj4F1SaGm3Z1lZcN5bwP/fetYkj720oLgVFuCbL50RWvT/cx+PbTwRI1c
ZfKIkbCbeHa7E619JbAku4FKcas/aTmiSQhrVzsvuwGtpDvtLAjIEas6PXBlnnPC
5odFYa/tIHtZ/5o4IQEsfuCAcZWxjrfLtxJq1F1liU63T0O3U6MdHS3K3U3IlGRP
OqjyPYJp5oMsCLDl1sw5Dp8PDXuq8256OOTCTOtS3AKbhKiOZeODwO9qhXf8vx4t
JpLfQtH5MuH7HrtkRX1vzwbhmDqcrEOADOvOR60wq2ZctBjh3nXfC7R0oXKBSyE0
2hXOpwND+w8RtIJaVSzAbdwkpi9N0QnGVpXZOHk0IJyvi3guPmXM+SLP7bEvZcKd
uq3fuY6KTJEDmHgwBfMLg/hWHpRvnLYUq3TskG00gZUV1vTV3kTI7/Kp6qnh7oou
Aidel2Nx2VEAD6E8zkXDmA==
`protect END_PROTECTED
