`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qXAedqBFh7tM3qiGHoxDuS49TPtfAaz3TFcqC1QiJof16mtms623d6telTX0Dwcb
9N4dcpTj1FSr/yX/yW+lJSyHq++Ji13pv6I6SI4ihXsvaiNoeltacBmldZ+bDbJR
RqZx2UMC7nwCgFvE62xocGK5z8onVJHRSjgTkf0BNqgB+EO0ag5l9/fdCa76N9Pa
+mel810er1rXdSjsNbCiihuHaCeQI0f7cDWQv8JiVSTVB/SLtBTSNmXF9yaARoKJ
9zD6HyidYC2SgXbtY2HaRqqTKZh92Z9W+dGTvyeOC1LKLlMbzEuXHPEVGlmEmhWM
MwheYhsM/0Tr2T7qV2+0jcVCZNRV1nM4J4kwXUlTI3WZUr3IC2lUk8hlLRpzIRlA
s5I1bALAdboiLHbEshorv1CwunGzzoB0IkbJP2d5Rlmjd4rFA7rkuwQa4uRKl/yX
SAuMRzdUpcF3XXdzXwJmum3QMCFYZd9zlMIvmdbzyJ0VQwt/PepmpjQeW2qk1NJq
pvTJpp+wOoRTCibf0aNSV2MIaWsgijBnb44/bMz1zexpiaOnhKHlZCLY05spytDF
SXExLcTV+fYxM4O5areLAc+ABtTAmwWAHrWhDSRtnFS1crla29zoHyPiGUvGzEPo
fWfW8k/yHpZiLsms+E3o7NDmZ5rJK7YX4cI/nz2gRXU+RnZzpUAibgiCR/6g6lxv
sTwqGpm/o4fZ2Q9rqG8fU7fsx9+SE+T2IkET4H2q+UWI4OQPRJfJXSSh5HFxEssg
2muh8KtjC591rUr0360emp9TydJe2Rz94CgreE7Yl8SGUX2b9QSWweOeUdB2VM9+
VUR+LWE4LWsEIOO7LS0hlfSsHgKbzvRe/CiosmsA+Y6RfzYIYwyBmiMTq8KZAyHp
NHnLOrvmJ04BbEz/uNy7xyxW8vxwVlYYnmlxadfoq62yfZAo9nDuBxUtx44Uvc1Z
otomG8Hg4cxeiojrFUSXf2IQTBxdmCxTR3Uhy2kEgUWwDvJzwPwI0DQ22zFpcf4M
wAxhSwJmifL66JanDJTMKB8qcJiZcYsB/GN9abOdA+MnK7Re9jrTL5VbRoovTx9w
HaklG9PhqEYMPKyIOxQOUKkT5WTWX1SrCC9FgZ7jF2OzUqU8yvQOzc481A2BtGZS
trIA69AtuaXJKErv+tT+QgA3yPfLh4K/MyV6W6KypIEdwGml9Z6BFmGy+u9ljw5v
2Q2MDvfBqvg42f1PF+9hbvqnAmAy+rb53huyzvymoJjeQ+iBnAwJqBSgHqIoaLSp
4+Aw9pWMCgcRNrItEzelNN8A1i8epfmkJmKzCDChhpu/sZcxEXwceOuK+WzTI2mH
8v6CAfaNwFR+ejQe3lfM5la5m43feHLB4OSITAef88R8MKx5zKDKSIw8VLLBld9/
y253XOXry4pDVmKXjysGexNfDUidy9w+EVevkNP5Zyec/WTki4fyd3B7xAwtuyaQ
xJ/LBYMTEsqkgvrUeNe2UifvLKGeEVWEu4jNpAWnOR9On9LHMlmmXpuym8cpyT4P
Frd1q0zrUjC763vCM1V2jorN+flNss1QDhQofTG8FyxL1ZFtoVT4X/m1T8LdpSxs
0J3E3rqMFbrQStm9oWEwQFXAsvzz1dSAvGcq82Fliw8iQlcWq2KzVEOdFsQl5gyI
zXVtZnzNClzztiMjGLKxACSr8beAAVwdNc9ALmyL+0FHcmlvqo6q7GKEJ/W5tlVb
fWALccOh2PS++6yAHX8cctFUpQAMWDBAXKeP/QMjKvNQocMW1dm1lOMKko+eGfQX
n65Eu7orrSW2SJ1NetquuzbMf4H3cASCwcpyXW7xFzg/6Yd6JtBKHoXjI8CvtSs6
39EXrvqCZGbhy9G166du482rxQZ/sZ+3EyZ06BzuKHN4z8dmxVwk7Tk9eBnjznNc
RPuQRwdc8ZkCd6RYDTflLoJoD4RpNiT0hyUo4P/d+AmpBEvnJixiyw0zdn9LICi4
7W1/T5YYpVCRN9i9nbrhDuMTQe2qX/XS4N07zFSTEPfe4tIxgCYUH+mosvSzVFyv
DFH2StZ2VFjKu7S0mKg11AarzW5WDwa948vBD+FTKtksOJYBEWSMb3tUBriM7Hqm
bW/qXAtTq9HjN4JhmQsFfqCwdI1pJCW6a3/5SMa99TEspxaCwZNVwTJ17IIjC78D
HzvKsf8SkZuQa57BtWGeChvLlYOQUQaHRsd9XyvAUnNhKcoIQHn0triafcSEBqU4
kxyXghF5FrDQ7s9agOK6xKZzJAWtPNiySDVxsNhs1Ua97NOlQT7DtgXIOEU7wIla
36RDYXGiS4eszsPU7xGy5Z8YtwJMkbuodkxdSJA4K26kpx5B5ODick8aP8OUlUsU
a1ZY9aYflX2RiSy9+TbgtJN0JzSK/tK4cv6DgTR+X9cE7dmuaLDyosBvNJ1G4fZ7
6zPXs+ddbK+jbMDG4Y3QiijLcvasLt49jMiWTW6LtKMKv8RSzu5Io+CJFuqfvdkQ
L/rPDLTfqx/jK1RNfZZi90DVmtog0iDwzgqub7dHSG242GjVn+UUOEfe8CDXTrCD
`protect END_PROTECTED
