`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HFIGm7O2DjOAxXthmTk38SVVt0+wPN1JYimE4FxPV+jpPMIMgNRFkqTY0UAB681I
NqWAe4nOrVEhxZKdcKWPp3MTUxPRqhlqC9CeMrt1tJA8crcC8OiwRl/FZSt4n/CT
aVu/XXWm1rH5riFKN6ZusSo60sujWihKs/+AEgGuIAgeKVQouxduMuopawPQImWG
s/2+AurEy35zefqEp9opZAVSdtx9U6Z52ata3tyaZxfC2XlF0o8OdE1KmtfntH32
//W85yWgM3g9tZgqnRYtYXT6ij6LwCoASA/8gQO5LGXwjevLO89Y+2E/8SZ+2j1h
4cvX7V9FqtWmzYrAV5z6gEsiJ7EPtU2rtmDnqvL4qq6tnh6YKUiBJa5wGtn/bQ3p
oPGy5IFB6/rGvjLmOfddQeLyhKk42e7F0UtvOEESJEZsQ5vRiL91tvSGD9R/1kjM
3RVcfsPAC90nvDdTq2FvrPlgf2kFQj1XWc7IBPwI61M/TvEu/P4Dw2TUxRwshk2U
dICzF2hyKJWOeiY5hcDN2gAUHyaokmbz2ueXgC+CtwnYSvtf45OzoHEYVG7LSidU
u0rpxSJ9nLdR3Lv/PNldJNLsBeruUL5OKmUYG79O6EeumMSXdvqJXfGzsPAy9J36
771lcERaACcytTDHb9hFQtjFetWpwTHG1txXwRAnRVp29chORCqaQYPOrBDV1C53
811Hu0ImUaPLhraTvB3tzPW70pqel65D61WaokgEb1a8ZLNnOb6m3nVn/LAS2xxl
PS/3wP4LFb1ZI3Jc81KvuUBsfHF5l0aEeunfbjiUHnUXVhebO4MGUUedFMOyekOI
hHSKsybSw2KzOyugJ5h/mUC9VgPkYWor6T+gOqrSglxKLLvsDOeuArAuel4PYITz
memzHM0sXedUuGGz8D1oH4JY0HcGwYqrcBODRdMjKi7ga49fuXsPbp0FOyxRA+3E
9l2DGKsQkfzP2mTOGziozGtBzSr3TLty658ddxYxvINF2yGceo18R77vnHw6yB3R
PeyVam9EYcqOotx138sT1JV0V2MfzSqlb/tSs4cFEeqqhiZJhbE/uA2sjrEJNJmW
Os+o4eQ8ER/wx8oLWXTH0NyYhzu6S/DVfdkP0PhOOuMAd7l67+DoF1oX9dZeoGT/
hA6I6gSz2Ufa/XLcry97nR8TdHWjis/LTmcKwa53xJp64kseFo00FhVTH5577Gx8
okz9Ozm9NZ2T5690rlQf5GDiU7UntCf8iTd/NCJpqdRh1A1tJHUrLmZNWeoZ62h/
1BIULEfxN0BU/0TRXmxtLsH50ria7baAQNzIw960ufYEV9v2r85R4egaRUjUbEyD
mO8O1Xr4U471pn96JubQ98lmgrordQthCUld6yK/CgIaoo3WK/J5eT8yRHp5016z
oRPEb0p9emHlvJPPEJilctoT9VM0Y0tYX2s2Skoq2cwLRZMkfn2tsdLMjOVFCnSq
QskRcAyuF/E/m1aqfcsZDlkWibOcQtXk78/9Iq+z1++9orZF28S1uSJUz3ccPr2D
fY1uu9lzMI5nmd43Po00uuDrh5Eplyl0r2eHurvmRkBNdokBPmTYdukfNKTLoR4C
pc2NxLKLw/rBMQhWCXMa/3AOniXX21R6BJUURagP4q9Ea/dD79ynEHfHes7txNO8
xdXkWjSp7AOuau1yo+sX6DOo3B21iK7/2AZxnpli5IVlGUIt/2FXHpafMEwx3UtO
8Tu+gNwkFqf9ZxziLcbFV704Vm1zmQ1Y1No2SVsQsI/t3TBkh8Ht37xNWoWTqAvf
NTYZeXEks23+HbN8I6mP0/UPKrUICmJwyvabJWNZCC0zmnnudoEtbBajyvCWcvoA
B2xzDDZ2OKykSeT9Iwt0iYAUgfOUDrJaV3ydfJjorpnieM2LsidUWigMDORNb2B8
dkooMOBAy/gRd4qYNQ7HP5dmSaRgjOUV8HM8WquB+RrIBESlOVDSudYQxlnIr+GU
yIVoT7n04awAww+2UWx7emzwO8TQKAqEI/NLIxbnPUEA5X9i9HPGIeBfXoh/BGSW
cJZOaxrlZNq1Ck+dEmUT3JYi61BP8VmUYfJE/UhZLcns/4c8GVTqGSbPARZFk6l4
6Wm+NQwlx0EQqnt5jpQJV1YTwDXLt/KPQYXxtmAoTdvcqnpaMsTdIAHy7RASYns+
DiZ7dIftxuK/1iZ3VjjcG0xsq4jWjCl7YYDoxO8oeTqX+CeY6tmMiDHZwBHBLqaY
TAHcaiQMuBDZiDnKWOTEsfkS86EZWRiyqOhJOvF1DW6J5ke6zEJw7unFA7Y2/5pS
/3D51URJO4u55845b4cCtfTovhhS3IkVl2k/rIs3PQdEL7LUgbkRVOFg/MDgloy8
hPjkj7y8UoYA6EIC/x6M5rlfAa/oPkCD1LjXechlpY+d0cQ8pb9ZS0BF/J+Uvgot
p4+QUYUrhwplgLCNUSMK4HsGJVxcB3ceSFEFc2u6KE32Q1Xh0s7JN8uocEEhH+1V
zIndl8Tdrc6ULL31h+VQVEcBbrJErCaN0Tdf94OXg5M8KDGYXxEpnAzI9fqu838l
HzWsG5tOrNuOikLg/BKbp3KfMUzVCLkYkXUoY597adVul60bxTDCHBl/bndJnmqG
eKcPIMCF7zho+ZX0YzTvV+HojvaynGfiN8Fmr9mSbLS0mrF1PZv3k3SxfKqU/AIY
b4M1ZU2R9AkL9bjj08kOlxRycs7jmf3YQfbXY21pw7TcjWYCKZHml/UiMrKJTIwf
KNAa57LCikQO0vvaGcCzF9uZWwNC8jAH9NK4eQbMWdz1D8GjIgpO74Fd+isdm89I
6DamijT+kccE8RErdA2WeU88Tuf0hEowNvapEV33UHV36AE4BQjTJN9HT5fxt5UK
IdeYSkD+VkFzfq5QAarFGqsT88bzX0RZahfgYX2ghEhBAHEwc86V6dJ7Y7hTHMwV
HeS0/+p5+7Px5oNJWzOa9xoZdtr1DPWy4A+kSHNDsFBXScfTEnAkX1gBgZvH6DGM
oE6DcrbpBahsEsf0y9Rv4YMYuq747k/QZclpzUNp9nZCQnGQL+XMBfVnPXeNXgFc
MV0Bn/yivPyOeqgKC/ybTQX4RcCjhXh7fHHFuseXKRX6pNVHRWgh/6kiSpswS45F
fQd2CjwOqGRiTKSQg0Z/msvt8uJbMZFmvD8jLNmDkEBw+f/9dPKsGQ0RljyNMADH
FKsFUSMQ3eNp+u4kr2qMdcvqQ0Uv6T+Y3GXuxPNTe9ipLCStzWlwH0hwd/IucxcZ
CceACOl59lcfnLor+VPl2sCOAm1F8+kDuQqvhf/PqZXsqhvDTVtVWzavNoKLxJKz
5+JKtUuyIwcxDTWSlzQc7uR+H26D6ahoZxqvUfZwQMrC5E01EOP8drVp77OXROGl
qKaJ5ovnIoo5BOtj7tEi5/ZWDow1cbxvilxGDedzyj8JfCy7J4rHUQhcceJ2GEoM
wnROpEzbGy4AnVU+octP2Q==
`protect END_PROTECTED
