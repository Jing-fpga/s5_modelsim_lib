`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xWHKSRJfzoIei521hFomsVu5RDyqmftxtsJOBYxFtw3tmK57OpMt58Borp9OL8vm
1cL3bIFcxOS1VrSsl5K6oeiL08vywjU6v42xqVZurQIEaLey1yD9lnaKM1XE3Prz
6lNNxbx2fihEcvhVq3sR9CfEjU9jXSnjgBf/6M0mhYAHqu4ICJEO5lRAK14eN11l
czaWgiZ971YP3VoOXDzIPeCJIxOvtGuGIyBi8deBodwF5HLchfNWpo+qQhfjCC4i
CEyb4Xu26OmJf/wgP/xOlhY6fqCcO4TqzPp35XwYXuTGMT/39VwZYEpKC7kK5sZx
UIew0nvoiEdx58pq0OV3WS42tcXOS6Fn5zetB1+2+IpmagvqkeAjnKLPtNBl80pl
rHcyWbmaoagxTMgmjQiWvsrErYr8gdbpCEeLcKCMGyMEPi3XOu5y0RfcTfDdb3Ty
5xn79SLNqJgcwxEXS+t1swo5o1ssWgzjfLvFQ3qin1+YJ77Pj3j+yObtlnoq3kDm
GZsp25op4HV1SnXovgJwqXtpEY2drP0aLq4C/qJ1054b7JkSkOOS0qw+j43jfV7p
tKIA2ZGRiB3psnNaxzJL30eAGxWVAJ5PfiBOuXU6cUjwIbWRAHd2kbyJVMhn54bS
LmGEeyOZkFo7Emly0VNmbsIolxB/Z4CKQgkcrd/gjd9Ta5vk2q0q1a5/faLxoUZE
477AgkNfUfrPNuWLOpvJXYnZbm8J3uei+8TCWruhzezjDYnJhtccXvsYG5/Dw4KT
t7Ji1dUP1uBfpMYDUuZYSAzny48gMblRmrWEgxqyz1DuNSG0a9o0ognbrZsGR0+Z
Nrl9OJVwNAvAqpmR94eh/CiAUhQG3AnwD1Icc2nVecwoR1DqxhtSkc5Rdkw5RO0J
EP9KveFfcPCuvSfXgqZTEmfv9qAwL26w6uKIZAuWHsvpS8pPaiG62nHO/VBPhRbN
hvCGZl5WdIUAYqS3Q9nnnLvhp83jziDEZvcQ0qg7pXZYweZJZGYSulvxGn5a+QPR
1jn+DwNK2jFilWAhMTInN/8I4uqnoDg6kfC1+UW4DwyriHeD6u7rY4S+8+t5OiNt
SMO4axXWlYYqYhx4cZ5cjGQoMTp2BXx6qNP5936Cc6uCdud4pn1rIs7UOfsOpWlr
wHwzq8fllTEcP5DNEcJ7NtbOWZeObzC9rsvI1tMZ4bbOMbqZzlanNk0ddGOEmmN4
wNUvcD017q4euXSG+y3Ge8jHPEKxUibZzMuz/aUsgOlYG6/NqEIpR0yFvi59iqK8
us4LHjAjraMKee1PPSXOXkwxSdBKl9XFyWGBth1nUdg6BTIuv1Wx5du9ft4SlJjf
qCZYvYupzQ/NdTNUwZlmNIkjBJazquaB0RmKYP+guFKVd5kPfEn2MApwVXefig7Z
G8VX/mpFmHdIl0VyU5UKEzrxdbE4SEKsjvfpkHGglW5qpbS8RV2JNjA7wnoRNm/U
H9xgKoavblGSznS0plXdM7+Wi1IiVRdnbJmB49JeFWAVXXW3JvjzNbtZ62nYoLJX
dKPr+/Uv1ZoJ51BRnO+bMOeeUp/UfJl24RaGpZvLDqS1xwk45BE1/4lgBR+UiL4C
LQ0+G9rIi77HFwyb4cxfXcybcieNKyLPnXCozTVpwyT40MqG4ZuD0uFF6vxy87Un
iHHtHrkAb/egdUumWQEWFg+ka+syKStFXVbGE/6TdppvYMFlXCxL6sM6vqPxwZTQ
tIB+ucl/QBazYCP3grqHuZJVkvWsO4TyUNAq6encuRRP5kBAt2mD3WvDDP4Z6/3y
J0TuSd4b9q86vM9pReLNr0hwIFzmtyz13cupIF78UHeIsVbew4+nz3w2v/xYYIiO
sZfHPScCWI2EGf9D7dn8sXl9S2DPdJDRB0gNlmjF9x7ushb/mjRe+BLJEZdq+3DQ
R5/103WdKqyYC5snc4ORZll+KjEZhE+qMyL/ltRBHKrHiDl3Fmt1vLNM/6f/ZQ/v
3Q3mXt7bb0S8wyAiud03IH603JbytK/uj08KeXXygWQk6inqZOTz40LxZLy28Aio
PUjeyst2Jytv/80sRRxXkDzhx1zsNB5UTg9gos0QPfg99DCwdfNwf2ohP6S66atg
ZQdF9cqUXdH6Gn4KdM0hKaN/4iej5TAPseefU/inPrukEA9JpeuIWzNRmjVcu2PE
NsoDGtBf7K56Ep3U8NLnnh3T757xZc1f8KbaijH2QrwJNEGuDE9od9Bq9sC+iS6x
qnN9qpf3GM/BrI60NKKDYez/+Udcrzg4GanPKUbIeG/ZUsX72FpvPD6YJE6pAHQx
r5KK3yHrCu9+LeKR1aY5khD+w8uMpis0IeQDvJSyvr1SQ/9crKFiNPbp17mk6Rta
zAWPG1paJEVZXloijgNwTMU8qYuuNxS0RdT01pD3ALW4XqD38heH2+Lwb0URroif
sPhal+SIqogdRey/nYNurXTJQyNvlzzXfR8a0juPZ10YVMzY1iM2iAw/y7t/e024
o6O/bCGa6QbKeufw2pWYKQiBG5q2+eXlOd2bsD77Msds879vTEDA5JNlvcr8ReG9
IH0AcoR94rdNCxucEKe1qrL8alQAmypQNVrlc3YRkUwvRiv0oru3hihpTzTknDDk
QMx5QhuZ+cU7k2tNxlx3L1soGCpz2n1xr4sj1TPnYdfQcefrdvrfM0/sfYDxOySY
gTfs7Y7fqLopKpvJfKhYZmhCKSDCxn6YvNA4/o725QZojCaCw0oNbzpBJoG0ypaq
ip+2H8tiPRkjZrs30XaRETqoRD9Psi2WfjXCyTfh+GHuj7FraGzR05u3SzPy2kL+
/Zg5/21wVH9gg4McTXiq2lxHg5hrWaTdXC0I5YsJx0N4xAFqQaTZYrFfoIVvZAUg
+jQHpLgpIvSdSPWhJMfYiX+ZHUEvZLA0tJ57wKjy1cvBwO+C4fdiSE6Ij+yfWX0e
7tKNiqkgaMxe/mklWN53euWwf3fViNOxkfqVYlS3z2zDaWcg7jwI0QwInrM02Jg3
tL3rMaJ/qGKmKstxxpt3WKVpfjJygDvasY489i89PVwYYND2TJp+OzFEjcEYxunQ
RMKUzUn63Qq9dvte73P6iHTn2vl95VsH4br2O58Tp0s7fzDXdT5WS0NmhtRsyxne
85pjRTu0HCdQbzMyoRoW0D1BVAlpbBvzoZmDRyQ0qwbOgG0sYyYuso5M7kdu8cTl
InWJ9uSocVJwoPlrb2WRAY55L7dDGTfElNvhEHhuFlyB6iSD5bRdOJDUEyapV1Sh
VRHGlUCBmTZ8AwOaOtO5iKkEBwAmoS9+Ivir0807WCRTuAgEBSp1a8F3V/+rWk/k
tWTwq1psMJmgxJtEKYuzd2RNyd2kVmzi2tbHkCa2GcCQo7Evj2kZz2Lyh313RSbW
I7xM2qV0NjZ2Ed35a7liyXcPBxTqhWKNV8MwafBIKh3oThxit8OJCLciHDgm3ZZC
jcxhhAbSLrlxI74ulL5peuLI98GTwn017kMeY/gaKggOJF92+Nsurm5TApQhcL6I
6hgnKyyidC7ZoYdwgnbzlpQdl5WnaWoiGl6LsQcwgbjz0oOCvabu3k0Fn+Zm0Lh0
BHzOgIZ7OkDTCi3lAuHuKJ8Ga2omwIqa6+wAXmu4ojz0iPeodGubz3ZaEviWz/t1
sZRwV00z+6IWK0nLvaGkCS9JQfq1VColFFYm/R7+MB3LtzbwrgmzrOAlwYQCd3LW
HtziZCsBFN4M8OF7auFCFnrynfd+Dvgm9WsP5pa3y4iLMLr8L/caaZ4A+Mvdsa1x
nfi7TCtyfq7tXDKWaDL9UI5QHPyNWuUHx08n3bQq/Mfb6sJeKW7WL7zXruEYBuMr
YPHLFEUcbTArbxWXvY41+ePNBbiM20QwEd9qm6YU8aJy1ggnLT6QDLsPd3CrB2a1
XIil7nsnSrXhKT0DD59tloU+wqQ1WXW0pvhRl80sScKSD6N9vi5fmZl+bS5GdVAI
bacEPsq1Gn724xkSEdMWgaLwzf3VM/dfF+XTa7ZyubOlnG6QLu5Z1sIeOWRQbkCw
wAXiz+z7Y91HE3I9TmrJB8pFWYk9FJoEbKd/mle//6V5EqREsW49aQYAXX9+izKR
jv+Q3IhPDuoL67lmUnAQXtOogMnFlAz6K39XziOBoLgdhvk3eWo16eUgXSEgsvTa
XgQnVI7vOTKXf05/RPZDtVfKPZdN990v24OhzE80rNBrUJxjUOBEf8f2OU/Gm+SF
Z3aMALh/05fg+3dwMDPGCONXJX5sshCvpqMa655zfcaPsGLc7eZkfYYWDOZXzwkF
WHrY7He8LK7iiMgdSMS8zfkHX1itGkxM1YEy9kJ47qoWaZJM0evWaLUpq9XQOi4J
wfaS5V5Rx44CzL8va8sDX2EXvPPYAtj39wklEbhFOUJ+6L1zjUJIuJu/St9+mFgZ
2Z38n78nMz0WZh5lop+xj91G1ondUrkzuSce+xt0WMuwoDholTOd4hVwf4p6h9Nr
h3y8WIcMDePh4sTjcnNCw68degXfjozLHHxyWBTi0VAaZpRsTlqDh/5YG3bQvsuk
KVAV+Ke/OPZyYZB5IT3ySiwOeKTfBlcIYblLGtN6vc6pWQqZggGPeaA5sGsiGkXg
pHyVzY7wWpRFiWEYipCb6kFTm/Q2RgpUQ+lvnuV4CgCbvuofGcvD8A7l04JDgu32
SkUrS4ujyMdLKDnceXlVm581j4EvUwsrw/K4tL0sH6W0kGlREK9tCE7oxvUZ+fdc
z+exuFF3+Ax26VyD0d+wRpkAHcMCto+iWNQjkG47AWxmbl0uyiGblWOai8h2wHm3
Mkwi852AvrHvWhrBWoMDxhTvkfr9IoNssBiW44Wd8JQ4zKFW7A/0yoWUJ+XKyMtv
Z2dkzaE3PPB1PzECWZ4VbsMXu9V7WTjkBLcbizNKtsW0PDZiPyyLWCSyYH9Ctx1/
6cDw8zgSpv/sdd+Q6IanVfr8516jQWhrnEfvZH37VDqL7Gt/kaZO7HA2hjiZjGSw
6WIcgCfOvttHC9jKj0+d8wZ6qE7IBSDGyBaLq/TreFKI0Jr83D8pubQ2eRctkhu9
lC6Dj0PY7gMVtDmMy9Lpb0oBz8X1Gd4BIEVkfEQHfHmHVtK0hRis5CC7oP+Eds5U
hD7x/FRNYZ42RZ4WeBPmS2ScB952Mz5FVwDqqqttQlCpgFMhRcakeGD+veQyqkIU
N9f678UI1rrl/fcUjAeDvd44xzJc4HNBSwURYRznzy6v3gTArVBWNCWhZQ8vMkDV
q3GhnpVlANzbzN0X+SfK+7TqoPwxrLAPq/BsgmeuPTGvJG/s+zl4IAPRD6ezBc9K
FrTDkAC597dZO6MktOVWonP4XmN6NSkKkhUp7Sg+hpjPPKDZzBBqxE0wI1hsJ2vp
xAW9joyeQzYHtXtw2I0GwEKd70tyHgo231DaVaFIlY+dfwHGzx4sjPaQbvXIC5cC
AtybrFzjft8PHkNSEYaw+T5spl96BQH5mc9CiSNmQCB9CXOABVNYxHWe+fcbKwlQ
HMtiUxwyGtZYcfmAnPVlsx6rAOR4o0uq78T9AGW3OBR7cV2dord9B0tgIcxXMhnn
vwkukr5jRAUHwkXQiRPHOpbuUklv9efdkHhp6qUl7DD3EJ/Ue5FRId0/AFa1jop6
PK1frvd7qlpv+xyL5cL1zorllwGvy8XhtXmCqghyc1zqTN30r4sQd0UmJYWbCuFN
9z9078xfsrHgbE32J8fbx4aQCmYwiiv//bPRKskN6nmJIhnmyp4BByTDc0Od6mou
hcL9VIcTSARzHc1WlhIoiGp1ISwaR6lkJ8HkuwjVfXh3qNDHHCmdCg7tsPzIEYlw
+cnfi6Xb0HuRmurRxD2bLMe5gBzLBKmjSXzzHgqt9D+c45EqFBOjb/r1wj197flV
YRqnB4jaYkXvNcGvbvdOIxp+vcBKV+g6CylJ2nkVSmkk1OhHj/bL1e43u4VGDoQR
wSqNv0cU82fbtLUSafluvOSw+GiOkHIgU2H3OHqnT9Q019LxGGzvluVGcQsLptU2
Z7ziBavxfCy3QKd2GoqF79adw19g4wDxI8jkn2TYica7qMs09PJ+5mkzMqTM4Yx7
DqCYkMzm/S9vo2i9HUh/IHxlw2PwxzaYMUpnoKkJhfooFqTYsBGbyfwXM4Xx88DA
1lxZPIPZTxihzm7k1nynzPFAC1hYtZI0j+GdyIgDZf3VPStJEGXgMQHYTOrgvvbo
tV9iVln8s2gtCD+LjWjtG4TlRAm0tQpXvVLe2iTrjIcsOPN4fu4qFrFftv61FoWM
AfI/QuMfWKXlhrFCrhLJbWk1S0QiObOsXFD1lckqAuyBRJfKHJN6dPqU3tueyWln
lMdWOHEcGUyklS8LVs7CgkFoWls0oKt7zoabkdLf67RksOv0wbX6bfuLp9gb14HT
TmCQ+P2xWre42UqnJhUYKA5U0E9iWb1JPxLIFNCeKGKix+43oLB40QMR5MO+Hoin
cio/IS5QWixHOCjxIlZ5dFIDVKJ45u1M/g3yHVElgbqem8/EjTcVvS7yYLue0+dE
hXCfTB83uSPIOM0SDJsrGSn5UQwm2TxGJTggO14OICUwdISbbxxnFRput97aekcD
7H6EtDsm4h+iWmSdNE8P3KD3D+gEW5ZU4xJKKQBZCe6+ZcwEnEpmEc5hjBLkI82m
sJ3eeC4UlEhilojCfEYR9J8BMvw2Eu7Lf+JMmKr7o84Sg/jmBD5xwcuNj2Km4kMP
Ao1PaWxJJeADBmeKjq0uAhW+GzgwBPcM7gIWWkQfUynen/3wjyJCSF0JbEBfMcWf
P3VDSeo94xqdEsnhF5Fn558YrIb0AFoTMH/mf5PQeOYtKr9hhtGC/gHVVVaWvvPv
QKtbmxqiXVOuDP97RuEvmGdku/LNTcaL/JV/Qw9Ylpoh/fWj0BC7URtSZZ49d5By
WqSepyYiM8pcGixKnU1+OUAoB675M+xGsgwI425L7S3saFl23BROoF9ntdgB12Xf
QrB98oLXNXdurI1MgXMoXtzI0tAw1U6ziYRnd0L9uqy+sdyBywaEj5RS0eGFo8In
vM3ubbD0dUl+Bm/k8HE880Nnwbt5rtpLJUvsG0fXer7yDYUQsz7Cj/atgE9KLsMQ
V6CBISTaNV7CxCBsjNTT3+5xV/BRvjwkiEMrGbZpXmtckNpft4O7l6pGSU6eJaML
++uau3CvMMzwRjzOSmP3QxlmJUyICn0VcIy3L9u+zRtVOFQG7lo1I4P/NTdZX8mA
SjwbxgZ04HXZwl3pbqa5XYwR96Lz39N3cyYBUaQMrYUxr6g8s5XGbh47MqzDJJMj
IZDYadH5d8c66U1CH17WQHm5Uiqi7aQ+/2ijOa3xq5+sV9O803mfsrDOd6kpl/7a
3D6pFInd5229+Mi0f5+C0VIvmErl7SYnW+dOuhWtA5BrLfWDcS4nnVv+U1IYY4Po
Jf3eD8qRXeKcIFcIbTcrW0EMQuYzBsEM+SJKYG5NKnz6x9MTOSbTCV+YPn/y9iXv
k77nOjjONpZqvc4eutgNeLD7ZAw2Vm5exfZ7Ou5tMgTOy2zjf3KuKX4r968Qhkxu
uikjG3TXYa5ltpLmvdhIqE+AIiVfCEs//tL/8DfBX5PVYSVEV6HwjBupWh+dHUCI
bNdY6TCkWd5Vq5HB5NxZU55s0XxXTx3qBq5vKSQVREdBdJTPdeqYtqlIpUe0+d7g
ND3hBSBGX/WpscNftvgt7V8HVzLTb+sVNl25dRbgW7WdrxdcrAIQo/TIaC02L5Dn
lGRxS+MIMXPokBWgXMeWlcsI8BC+/Fwo7XHV/mjypUDltQQ9VUAHAsZd5n++myjH
vgtlGUQP6pEposIZ+IREnduT358wLPK4S8kJu3CzSl0Vf+3VgMxx/92qSOwqE/3D
0MGDelYTdSU1a6rtQNVBZIjHasVYMNZeTAcklm9233dR0qWuDqfsGddFO0XHXr0q
o9cGCkzPIuSGfWxxK9I4oC9pGK40ZTVqydZ/MrY1FwZZMykp4pakh4elrJ8gp2q0
vjzcKMTdRUAXMkJEcbxuXeNDJ8U/WKcOaChHYdvDUHS4UAwR8bRG96Jc7CCOWMnq
QSNBsblHt9NFSWQp/dxzdHPqTJ2XJLrv8DoxmP9bCko/Y9GXPduKh/yGpqiyCruo
XN/M6BRWFO2r37LMhe+T2J05P2sRybLN8loBG3K7W0g67IJrMloiCGsam/DT8fEt
hS8LSLeN3X4GpjWCKOizg1RomoFQp0CdmKPasz5CY7W2bcG1kMClLHvV9nIKtoJV
U341dskn2UjPcOEDtNNHcsFGoF6EfE0po7H+d72/5DhznpeoVc97NYrrWGVs1/6B
7bOKK36znWjaIN/29BuGFuzR46tGN2ATp+RZfIUQdfUV21RTFQGtIhEeoIMCPRN1
jsNXjElrdej0vdeZnP9q2zgrCzkTCC7o608I0dPEV1yFDrFwsMUGdxUxN3me8JJJ
NTB3DqwLLXjorRfVrcBsOwNbdytcLR7dfZ6PPImFmw8XqfXHKs0WMB7Zn79Kqf44
b9AtUP7yC5+5acH5dyPUDEbxWK7n34omilUjTMuoYvGkECfaTRf69hizh9tPo6bm
pM0NVPQqe3HpSVsBBD8xgUcFu+YEhQhIXG8Ky0jMxjC4mt0mspFHjo7hv1OCX3AJ
f2AAC7fJBmI7wrW/ZvYqePD6YIG9a2FRHFY8Ub9np2GIIJiaSBHB7oAVfmuyw1rB
Bnj2Qs7y+x/qEnwMqudW0KDZKgbxSfsCZ467yonVz8+E5Ut3yA/zqIi/fVnnhKwR
8pGXpNuC9ucMSCmPCMp8fWnRmL+q6MLVs0BOb5iiW5X5VShIfXr1+fkj11+iNfIE
W5nK6jT7x3cmwdljs4axxusZctprU7rA4daf8bSAc1bG2DSHlsiO+ligDQFaHe/U
lKE/9sbj4HfYtIuMSqwId9CjMEjG41BHL/a+O/eXSPKzem2QT06wuafV/SYApdPh
SJGVa1boScOjv3ghsqbm8ORTq6fwv9qL7k2kNhSjtcOd4VxxIQ8lNleDdPEf4iFQ
DvIAjc31a/ks83MMnZLKDOzI+s20sVBpmZApGdnRQjOXp/5moIdlAOQU5pBTuhMf
5WToLWL2UJ/ttdlGl+ddkIjdgs3YE2/beKKvAtIIGKZqjtQetj4II6unwr884BXR
d4pDyxPc4qWzjxblfIXNMHhI2iPemGZeFTP555tA2ELXAqp0ZuYXZwqST2LkihyW
t+GQDRxe879M0qOFeEQZ+c3sUeA+P29RKEf8PJiFLGidAwMNcVuJasDanOEEwfBn
UbU66BYoUn6tDX/kV9YmcKLpE0DwV+88KHeHF6Exi90DRqUVCG21XcUPZh0olIDD
T8t+xwSVeRnCDDQgCMaiRZNwTfFGO+IFw/xznilwFnNX0veyYt2FgCpZYlSHJ9bE
tzkfjCzqJL6GxIy17pz7wU7OchW82hZY1jVwpjPG8zk0a8cQfQx6Z+BJqedjvc+J
ZvTNCy2YAS2QeFvBAYD15ogbvyilFen+x5i8/cQsIEzsVvST3SkAkB9+Sw4Yca/V
W5v99YJCt0yhzT9/AhzksZpuLZnr0xpXeHZLeWDTpVHPHKlscF47r3pwidk1tlZe
plPvLF1UKGvVhbosPqATRWx/xK9ht8NxL2OZVNS7FvUVYHeZjNfFv4gL9pqh//Ac
rII2w8WFpZ1yKmzT9VGRCz5OkZN7SXag0NdhqDFToGFFaK96DdTW01h6PC+biUmZ
cvFo+lVB3yj4NnQY7+hcaHEUkb5koH7dncg+lQl90I6zElEXkvMdzMM6K/aZjSfB
D6z1ypLUz4r7mfcGcGs/XqIBZoNz9P3ZxpnMJnESfTUS2dOv7EVOS0KrIKHASDJy
N5tH2bAXA1Oq73u1si5edrOVfTg6DDfk3oxAiSnGxW/r9OFQ7R63g7v9TKmERriO
YO/LCUTPQLe0pw6RS06H08CysUAI07+Ichi452I8uTCBOOn42TqIP8P9dvbU6GzM
GYjzABxJ1mmLf35+2oAbgW1GcqGo056qecVInu6a+EbtF1uHwTyVv1yhjkAoakMD
XkXS/wRKWM1cDVzSHReCqu4aYI6vPwcfpuceEryi3bdSvKot0RgJ2U1U9WkQ1ZCA
BlyokPToRhe7qjaCYDilG6hOKpmgwaO/PuelczSyNxTJDiYSFmXyhKyhXu7dswdj
6fcT9lb7B7dOcwxmdufrn9BuZ7KXvJR8sDvQ2weVi9I84PVMvqpUuzsHgnYmVNQD
2bUVoB9VZv+3A83l0WDLmd8UuyuhNOaZu7aWUBATyEEF+UvgxxyeB0NYtwyWLwMo
3g3t8cu2oeAXZEJi0Q2qFdeDhoIlucQ3BtwMFyl3Ge1eT7VGyZKpj3F395bi6PzI
MOyiJwg5RmKaN2i5nKLq1VqJ/lb036VEUWCWP/VNGLHRDQ0GHZPYpMGqaWfc17ud
nvHqb2NAaoa48M39uN2nNjCm8F2o6ZT8N1tgthxPcvZjb0bsf7dcV5YZ3WI8/hjU
yPSDXhM9cxUSbUfnOHQ4xa51OKL5HzWNCMfxOuHH1jrc9M0fT2bYUqWrQfuQe5e5
33t4KH/5HsJSCEOh2Jt1Nw7WCtMyei/s0ykyBml36eyUTy/FHWmqV2tzymVGIQnJ
wEYaPYweLNpypZ+D/vC1o4jUjIJUYCXb7tIb4q3vzveToKDoRuDfS5m5ZNI3EciC
msVt3uAsYEAyfNXRx9XDs3ntqk/2i68fy7qDuMr2oKoOtrno7Fqrz42F4sXj+Y6f
oR138YYR+yBILeAf6vWkuDStBd6d+h7ibKZxAXMhJ+XZcJlC/igoYRmpb2cL1QDs
zmjsX19KF5muDQ+XRq5uLC1SIVsbtD4nQuQ0wC4ziKL0lVbBPIH3bdIZo0kJttF2
9mERfOI+4aTAp/t1feFRt/aXOYNdFwGq8Qm+zEjXRKwkO35ez8ptqFNtAo+s9h/O
1A4tWagWJQuypgBOdiLQuk50IyJJG0vqDYx2bCW/+s/2nb4JoLDheLuVVeytC0Zz
kxWwZaHX4rtb3JgH3mROv8cRuppwOrNz60y/UnmJubs/X9NQXwFdGz5MX9lYG71p
k8whwrU1ca6EgyG3WQbOD1w5RKn4o2jdqdsC61piYxMZAVyXw8QhYAmTwh06FZ30
EEITDsRJNEgK/RFer2eS80YPO1cD5SAvSwqhCWBg4u3uG2tCiKh/SKEYdWFGBFJY
E7MgwF/K2XiiF1IDzCpAs5f2jHZwVnFVFApvYL3EmNIo6mN0FAxWiBC0sUshbl7c
gYsXYhd/BxXvMOu97MWDaduPCLxx7GGp9iY4XxgVkSt21urh8AALOwFZHFISKVwE
0YtxU4wOcEsGjqBY8mNa7OWGLxy+BuRISTD6hynSEUPP/DBoQ+dJNJz/s9PV1ldm
grscpieBR1f829+5qAzJvve/2CLpfGrNHYUOBzcDQkwRJFFeboz/BqvW7O9+Bd4v
hnlphHes6a0Jdzf39Cdf7X/bAxn2qYAMYYQGUzYaD+F4OPt7TBRtwM5VC/vlQoOs
p+KxNbkEeBflYtouAuvUyVcW8N8/nOM8sFLXqPm4OJbbjSal3REFgUQ3hbMrGyiB
uZJxf+ppKXIfJY0HjdKwalfgqa/ctpQ+xF5CedidBCiOj1s1RSfnbGuttSpPCyNJ
TqYHClr9vz8hWZL6Aw2teaaF7DT0l/yZMiSGgeuO+zOj/oEaDVBAo4b/eHv83qI1
Ov/rtQgDhi6gJL5gTWYa5EhdUuLJWfSvirEgXY/7PYdx7ViDih32buvrNCvfnazg
OjiU3QVlQ+MbbVl5/YUCRjvLwUzYiXtLDDyY0JIkgR3PI5tMgg6ahckWcfJ6Myal
Zu0ZX0hHTuU/Shz87Cv+mpD+a/I+24T++Vf4tvMVR2A0egPdHUfUyIH7dFJ2wQ0z
ouXDg/tbzdMoLZbMUW3lW83/ALObqJwg+i1G5S3Uvp/Pp0z2UlAD4zI+DWu0smgu
cY03h4QP+KP2ZbSMtATAJoSH5EbhXQmNn/hTkV/g69Z1XJ0/qzsc2G3OtYEdHSR6
5n5DMz7+7e9gPzHpzfJCywL35MnmivQETXpjXmWgE8Il5Qq39eVhmA9wwgYXARS0
6auzFYfFeleHw9oPEW03C23mrPL/qUgg9Xr/nlJzLQeY1QeqbNTLQAE3sE1F2kPq
Bh539e7Wy+pNTWsODAnC77KVFLmkO5Rdafcj4USwk3+3rkRSUD5tbiPj/izOKuYM
BziDrLnkP1LSITlnksK+Z1WIMJ+tTGCKXvcQZVwY9nbxTD5EIpPzwNGX10DBYEnF
8HoGNjYrlKk6exo3UVPyGQYIwaAm7i4SMaQw/dZuJA1Zz6EE1hLg8JzRqGXYgxqi
8ccalNfP06SsOq/7g2gDOGebuJqhH4dgZiVBfrj+MBHGzye/50u5gvln+w0jzit3
cv9bMP+SWo40Hew73whrajHip98EfZ9+5P+6uwU/fhfHMLsbS0cbJfdo76M8zBWK
iq5VHJoHzm9SzrIKS5UN1bPNRJ3aTex817FKUY0Q6EgT/ZY+Kn9ZadyR0UW4hMSW
f5DwH2ebi1AWJJBGWr/jg6N+Vf6OqlIXB0pawuuoYEpDkkPdtJFN6DFMXIpcnqrX
Sawhj1ZMcE2/89k8qRTP7RjC9RDPYoWdgxGFTQ9TpGhr+NmKzUjQKw4VazUhUXJs
xYiWjzUUr3KFjDU5c6RP28RqlPdW4giaRrM833tTJydUVpKQaBOUrnTAAmZens7Q
2FkMjW+eJmYfIWZhkzelaPzE1w5T2QIP1C+0/d/nxjgeTMUK0Obozov/6sZfrXp3
JjjnXu7BQL4kxPiG6FiSQCets3VpgML4FiVjLK2TID5rVSi1ypGaI9W8LzYb3VKI
Y5z0p/Bs5BrhYgi98qghPt6hi+DufGS4XidlSHw/Z12ly/QUwrVe1VvaCqcCTZLv
Jf7TkORm2OxLOTm/aShB+kiUzocaspx6WW8CzWmJyT8dqJE4iA0Al+28042hS0Gd
zvhLm9zy78KTYLt+vXM5pOw77voQDwpMERkyFAjAY4PrMcXrf9Uod2tgyxprZk58
VbAnZFfn89ljtVv5yzIotT/Kha2rZwJT0voaxFjpOzWYL/3YourNCHE1GeAbP7UH
VEMCGFnWpWlMWXf1nDmy4CCe01qXCbHQGfmZc4kkDGoamC8ONQbzZvmrdHZbCZq0
ehIWPACMwMbuDKWJw9atIPhkIS7ccYqUDPn1VVNokCI3FUGh/9F7ZowT/wfl9ImA
YIE0SLp3C757AOhFcpsFBkRaCf28BgAtXkH60Alpqs5n1WOcX4L8hjKIRbco09Jc
H9v0hCwUlh2qvYdQSdNjRRsmXMXudwkoohnChsp6+fbyIbCiuIQ3Y2L0i3apczSd
LGpe+T6SFnMcv2KYIHSRWjQg2MJipmr3mwqQolaS2RTDb+OUKPZ/V4CaYSuwZkdz
wjBCyDiEKi228/m8sPd2W3yj7fj7tRxKMHE7izh+q/YOulDi/X61giQM+gjvZDV4
3GCHPigCwRnZnTYB3ZbExgP/OqB1CrTDvSDjKzMyPbTJYDd42auq/JxfAaM9BYN1
KLM8fyqktS7HtVhk+/pCwDEm/Bc514RrQ4iaE+Q6cVI4tmPt73cg3dhthMDaxgkA
lARw0ZN5axtNLvdMnCIwMyGtryMM2BrA/2TCFirnAeqM+JTW6gJOyaxlK8zLU9nE
hlzk1akNajiQnblqYZedoLXd5RGVunCV/fJ3zicZped14ifGyYWN5r3+MR/vZug6
IS4IBxrog3F/Ampe6TsYybKYiBVXAJ/iKPHzsqZCH7NAtg2A1y8OKT8lzyqn/VXn
WiiEGwmrMTCLYuMasNcB05sKGCIzCXkxV/OtE2AfhRwvzzJiuPoypuzsE9oU7psw
lpZWnAweB3y8pOkHNFCP1dAbbVbEH7+GHSREc/TV2AfXJFza8RiyEG+7ralZAzfe
2HbPODHoMt1GDM47U9tWlTy2AwhQqFT4qKDxmgrUk0GXAiRav1/OkmdjM/vRy0/I
Id414Gby9PLuenskMwzfKS8QXVZfKYivFdLBNVk8/mBxEzi1UxxrxWeI5deqKNtD
FYxMDV+3IRIzva8VaaC1P4O/x2pPXx36yyVdyuJWtIuvH5RiinJcnVEaN03/hbtk
K1JV+JIHjvrhGT1LBFH+YVdrOd0p0MHclxwK2Vr9UiasXsBiJPditXx6MYfFsXJn
06UNyL/dqp5/6wMw2/Rs3kTx67uETxlJ6k0KSpthj2xv+zeEECnqSU/7f60inekd
yWs2qFJRGNaWcg8sfAyoiAM4IUqdDMLw9xQWUb19xZqOtvrBx03V+U/3Cu82ETSm
+8ZxHwuALuupdazOLs7jE4tqIvaWHVJJY9xZa4wP3Y453c5zZbcanV+CQtFZ+V1N
sztP5EOAZ/NIoKdB9FdZ2B4YfQ8RzZv8iG+m8WVuhhFzMWvHJr1v6h/mDa2RRSlG
Njcu8xcVraqWP0sE7KyaMY9T6+35cjpF3lL8nCiuFiZ3MtvPQg0JQZwNMDR7m6GS
7bbGOBGHmwqZUoGvTDwoNHV9PCyzGSKfcwLZj8gWRkA31v3djjx9H4hZjiCkWFZS
dJygQvErdYhtvwbG6eJwYxcafTuGzX1fuqXYfuu1s7BZIUC0sUs9pXSrlMfeQkt6
s7F2tRoDw6vw+RUpS1QnvUCIOtQLEWWADqoQ2TzU/JTpjCjZPxsDk9K22404PTHy
rCExW3Ac1/YsNiA79HkOxYkn4kJKMzK6cdytDcLZ2bi1jZ/I75xDL407nZe9MS3a
iV/KbzBig49xZ+65guUzUmzIW3gP3la0NjWaA2QADWvdRlGdo/V2K9p6xN9vLhzz
jL1lYxmJR9DgiYP9QP/mJGVuosXi6q7p0lD6b/SAOYCTFeWx0x/n5bKkSxmMuROF
nYrpSpOL/ZFCLek+6ZJF1pJ6jau0e51gFneEDlKN6SaKRLIa+Jq519H+Q/erKSQy
Zl2eQqTX7UTjsZuIDIbhICVreVrzFlBNnQqNKgX8BtGCgOVH3uEXPqyuwcx0F4Ko
pulU8HKX69mLVfO3MJzMc8AkS5nMZBzTHFdvkI2OqOet1hQK937g2x8IN6ycuvig
NLIHEenQ5j7aj7vS2Qq9yfoh7KN16SCX8f7eT/ZynafWMcxK8kq6UiS5QS9d3DSR
JLfoGEqbWGhg1+xqfRn4pgTEV60nW9XxMkbTkaNvuCg8pr4fZz56RfqwTvM4oWoK
Hc4u8yuaSw3uNKns7gLjWkpUi1Ob++c2ZFRaQBpdY/8EtXvzE4javgXiXRiiU9eZ
m/hiwHUYoBPEwBZ9/c1WUKklKYSnQDelskG87aBoq3bKPJGzjExM+6D/kKsWEEil
hWN9E6/hz/OYGvIZwoOfnoOXzF0skrM9K/BUBfoW35HHkKOr9FVwfgv/x5V1FEIJ
uVRliTRic6TJRCyaKt3jJwdeWJhw78h+vE5EtQmOY6y5gi+1Zg8xqM3j8EHuIVCn
IJ++QSEm7DwoULm2ziwS9WdnwSOZ9XqObyWm5sU/3Ez+rGvhO1mD+Ku5qlhD1csF
qhOb3/2vpatBySmIJZ0PGcjMAB9eFo+db2p6aDYwOVZynW0prj8oWZCswcDrAOJA
L2Xs/IFm8f2ZK1mMhpD1ZupVremFNpgHGW46sSDlYEQSSy9BryYB8zdF89Cn4hs3
hCEUiRlGNxR0jIIGDZxwcpoHeWC5uniUcJGyYDr/Oqld5fx1/6NURZdaKQDn5abf
FCuxSYiFyR8Iy+1U6Osa9s9tGK2omLAugJyJha4JN4ws9Ov05odBGUvJLucEI96M
Yu3Ly0DjAjszQ3fqjtikoPWldUohdG+ROAJeboQSqx9WsEqFuOo11c9sG3lb6oax
OplYxzWN5B18z6aWYJAdKePBMD+UKDLx+pu+lMju+hUQqwc82XO1jQVEuvgNUDlr
nX6YStxdvHs9/S8WKwGiMbT07QaFlQSd3VMkOZb0g6Uj/x1OVoQYskiodxMcwqqT
M/lD+GQreDHH170NoOEaO8GaTcjH4IFCoaL6jqD9oCQfiIY8K+iw+rP0OLOX8Uda
2Aw9rf9aIChGttUNCXKHk/r5ObB/RFbmvCePqwnAcjjxK+LG6GiL3J04rzd80Tkb
e3E5TWMcZ661GpK5HYwBwCgQMkyNJzipgHiZ9QI9YzTVQMbCsvyEH48AkgBR/iGR
10cQzn5gInC9M28CO1U6URt3OY9aIzlehXEzrzdmEIcoD0A2WS7VctrrU26XrAJS
r1H8RL/Ja5PJAvsHFAqZ03IfgqUjGMYv1OB+Vx1nxeoNwi8RK5/yC3Rn85vRAJjN
lMI4f5KYva8Uvs36VG6+PJXP6Tn8bQ93oLTESsrXNPsWKInrsu9J2vKPZTcD553a
QGxPWITY973bDiMJwCvP0Y2bH644wGzUl/IsbF10cB7jY+sseOEXv7YNRgPVMN9+
GKq6MD4Axoy9xMZGBJjjd1VCOCXVoV4ObqPMPjIcmOGdSpnPl5Oz1/+PIB2PNxAx
qcbHnHPbfX10BsjN0XO+Jju1dP+vxuXbTSRloc/ADIcMxAb99V2as+mg8pnaa7aV
Tni9oaPouhwT0h1kh6fI4uhICDRuHyDRTnaVqGfNPlGPKqw3fQcQh2nRZREyGEzO
YLaWkblMqqkbbOi603dBP+Rf2Qy37OFRhCkg7Q7Qeg2Jal1TfbMWk4EeNXJNzhw/
I1KLwCPA09gCD/3iToh+Usfh1AoEOj0sVfSeX4Znknnd1LiIaiIZPms0CtS34kGh
TnQTclJLNd5YSGQPYKLYtZYZKSYD/5dti8TRWNLu4sVhibWLZK4pfFJOpW5k5sQT
7NcMMfR+pRYWmn4bR8GEpkQBX2uGUZ5EhLQ1FqlwVbUcOW/7q+KpX8HNK8idDGD/
g+0rdGrTsPlYCanmznPYPC/sUJVYOI7xpLMmymlgYl2IFWXYJbLG7iz1o7hRuSzi
ebzXyFTbyO5DyUaIRCeZAc+dXwHB2982YKhntoO2JRMiD1j9QuPldyw3Lki30Gx9
85En/dua5ZbiX6Shc9OGpCSKS+kjnlaBi7m6+1GLRNo4R8tDpz/crB7h7NNkZywu
HIpM6XZRa0oOCxXgasjye2dzXrOwr/RF7gJZtWPXiGi+Tdz38AdOg6hzFhiHs9ga
jY6B1Hv98nbj/WSmBoVJVcu2JOJNCDYigBJHxoIyPuhxL0uczT9vNk3QJn6yAMnd
hXHPlS6vFiK0uIQRLHX5FKKKBmDfccojfpQfCN9/Flb3FPJf4MEzHfEHqW15MavN
+zNk6i1jUYUX/l3Cm8wf6B2EwlwCQO+ykLQeURmPGdLaLJJdIyhhYDN+3qgAVebF
x8Xmt8zbMQ8A3iBpq+l0JfHjylg1uuYtGKytiRV9LMcf+efFYjnANMuKPMqaH9eF
QbJCegtJmVuvHmBTuIAFgKJZM1mqQtYP401/CrOw4anj7HFObnVic/tcerMbeSba
HU7SEUv/GtbG1XoLWORyYQFGh2n4XwNBGEvOScV0oLqJNtGn0uKl0LPcrz4eJq5I
2g218415SgSxdn5kT23ydbHZ0Hcl34LX6GaCKnJvnBMx1VEAjok6qYY6A8lbSl+D
tYAfWBl8eppRY2+a3/AnF9uykOxrVPN6nPDr9fpKTnjSPIjBhqB3BZgSMi9dQKcj
ImGW6YVUrhYuEhdQuP9wjypIno5rAHb8GmaBfZLfG5OXJOzKVJlQAy+AhwmGyysD
FnNAUd6mLCIsbGsr9/NKd5AINDhdykSLHwGvyC70kh8dBl/3xa1HC20gG2DX6vLk
cnm5fnzhgtghZiyQ/XyudGBiL5wMJUaAFuAneLXMUiY/RHyga2xLnBnrpUe80k1P
/iOExhUbtbWiBGPYWjPHCNh3f7bEoLkdKHmzpyKapbaE9Fn/0QXIL9EZ4wgM1Kv3
Gx0u2FSdwfjskomUbGRsJIV1CynNawrLwrQcALYjD8XChht/CP+lciB6GNPgDXnM
QpiaE8ViheC7mBtdqyPpfdNtY88vJvpPfl3Co7Z1k4TSz9XzGZ0VyBqieD1daG1n
iCLYPR0pAc/VXvnMGKeYAK+iWt7QM7iMpzQBU7HSSeuZGyYvY47vOPKp/HGDxk2c
ubbKWwpTTvghTfxUVQwILYBE1iyrwDWTMmD6pHzxXuBzn+grU68Y1AWgqWzudjc0
MIzZUPErngwZHB+nNsPwCtUjP0iVMLVE8IOX2N58hQqxTgK4sHdshJbaHTorLkj2
5fvUngaQX3i2WhkmkaV9efJS8rDQGz/4DIdVBevkA95PAW9tOTGCZzdAFxJaBXsQ
CiWQW6TzMf2Q2rjYxuZVljkUTvczoqBYJJ952LE8TqSFK/jqjkeUE9N8ANlBtP9w
3Mks/OmVs5VO+ZTQJFgjKBe2afKDUkHhOeqHWTPHiABdnCuN44iYGmkUIi4ijA/r
L/iVkUlrENDQzpQ6P/8o0BvCq2AVYvz8FmmxCcvhVImWDPct+LCSmclJiYVn2wOi
EwCel2LhbDIGDv6x6LgqEHSjqcyEIh7fTqofh40fsl86dN6LvK67R6V4jh1umE4R
mkpCIyQRVHefWZCgx262ZkP4Y5/4u3BbDHO1uOlTchZmahXcpMAAMg9oo89cDLlt
syNbxzAJILLXRZDqVmSumQDTZCD+z/qU+Ru4afnCyYMuPr4uEIF1zhPGatgBW44P
J8ygE/84pg0vhntDLxDxBOmbiNq7T5OQLvG3Am/pQ8rEvWgoOXCd7t51MK17n1k1
PdoqRvGnpv0xLjqNKjJ67cmgklOve2GO8ZL/BdqKSRu7yL62JZzOBSHIRYA/QK+g
5/Y0PERhUNqEPll00SxVv3ME7m1nO+ZGlDSug+xd7RMmZqJlGgMMUH1hxc9EfQDB
H7JnXOe2UyV0dujFOS3/eMgRR0qmuwKEVRhxQimSo0BF3BCnaneeiHTzuHDNKnOo
sNhfO71XYKYqSd3p0WQ+T2z6xNpIv+mYZXSbD15khC1Rfjs0coelsnjqHOOrjmBL
2AnCIQS1jHhZ/eUK+9JS9JDakwMr40InQkhAkEcE1dbRnYniJalQeOfuRfLYlQSe
IUMoSm36E4CFi28V7KuBQnTLezBZWXVm5hhhBbIoS40D9DsmBzAKYNsBOqQbQ57v
RlV46tiP/YHC8/clVIyYqsc31h4YZkMy6yRm6br6/7XBb7YMCOHbrM2qVHFJ+l65
FV63xIX1OU+Lm14/aWTIHCAAXgzBzy+r3BUX9vX1AMDwWtUTAoRhp6x8ZVyfnlVE
gxjBpquaIxFKZXGEpFtf88XXc4CyplUbFC91A9kWBIE3vP69Cou4MMee3bev3DHN
FlMVgu/drzEBtSKLsmivhwhZPOI0vcYVTLWQsDtNkXr4SA/YJmDbbDq7OIWDGTb0
EEkYRJP4ucV0yh8CFEWnu499POrnw/ReVdHpBxAjN0aUa3qz2Nzlt5+CWGU82H+H
n5VF/CqAqxK5ugPblcGe8+UXpjD1vOlYLLaeU4r5lYMOU56U+gqRuWJH7ohq8Nq4
08cb8ZKDzRDxEUJhqoaMyP8PoKlf63bwLO55DTS6fsB4364HL3g05Gl0QxSITSz+
F8BwrPeSr9QfSZ3AnFK3nHJvYCA9kcJSFDP5B8mJd9VXRvqVho5betkmZYuvxGB2
mKeP4lzzpu3FNko4lbBDGG/amDlxvZSXFeiMSwUk+u4KBg3BXwg/9bSHBJE6C4cX
P9d43EISeOX7mMo1QUJCJYWIiXLKDh2j23jyW7za2kXNzgKT2Le928C7xXh2carm
2oyyT439eozfwhCuBfWjCTXMFwm0Rwd+w8MsLhB6S6Bmg625Q5+BxHwryD+9odI3
Y1NIig2vr+V5WCf+OBxaHmI4qJl3e8zw9BeIqV26/VbfizvWmAB37/bjxuO8cqPz
h2uzgJq1K1Kl3bcJfLl+53qgM94nUgf69e44SaVZA+zIiuDqRz7Omf9/oQvkjA36
G78IamCyXuqBiMH6W4temH68ZSLzopoyMZ1oQRvF3aQ6wgh44d1usWvAwgzoEbcJ
whRcvNXhHc2p0+/wyX0KoNCeaVLmb1f5JNl8spbPFeQfIhyDaHs9bodXrZ4MOLrA
x0FBfXP57XAT/udXENy1gmKRBTfaZrzpT8wBflMBQ4g1QTurOwdGGcISk4qLyA84
kCTKkXGi5Q2CTcu5MjsfO975mafKRHplvlIyhSL6BYlYp3p93iidiX7++S+J/x9F
6id5FO8tvBcurTC6pn6DMYql9ZArjc0KZ3s2Qsc03fbJamBXxL+g4XxUkCCPfxDQ
Mwx3aLGulDjwBWN3LFjdg8f8Wze1fiEplkPRlZKBCuspWGG3M0bZ2EvKexi0B4Ye
/ZQtcQ9VIk6UHyBxzzTi03FsXUIk0gxwfNlVs+BTkqeOusdrf/DwV39eO+Ifb5vX
m5veJ9tm40OWSpYwTSCI6z3svPQcgPi0qid0qmFajhyQQRlyEkdnHItM4olDJOeP
EtM+iuznO+FimMNpggLFGaOVEzue5LmpJkvlSlY1N+j0E18VhZlCe1hnHvVsGHON
ccaZ8Gn2jImwq6UBAM9va2bE+Cy7DPSsW8g+XZVFGJ7kgRTCmQeOwLFIE8usPdsB
AXrEgyxCmkFGwqrxa3stQsrXDqH6ZUNMPyfU8+2wTlm/J8OAZl/qbkq+b/At1Tao
fLOTTFQjrAAwiFf48xUgrz66IcYP4iOhJbVb83jq4NVqmZESnMFj8YeAGTgeznPm
OZIMjZYGsHSQj3ooWpo8odgTWorlB7TM8aVMHzAl+4uvLp/t+iqpO4lJILishamt
+1Ojx/QwBBfsfAEn0AEmZK4T8t60eyJABEcaxkpYCxwHwYA5C4LQXIjaYv7Ij51L
YKIJmFPXFvpkmL7cHqOlxgtotG9+KHqIs2A1dWPY4DVEcZMNf/X0E8rcSks4KwdF
aNh2wZGJSHqtj4G6mfQ8JASSUUwb9ev70arIVTJqwtIIs1l8UDd49mTfLmXuIuxf
W2x9hzmCkVyVD0QnN3cUhCtrYqxg77QukleQkkJWJf5k8pQj+JGG7rvH86MTCKYU
aY9+ehGEblX3K1MWAWoUd9bZnJvHe5QxZTSaWn1BTMn+k0E8C2/vjpBXeclEgy7d
rk9zLQPDUunDXkdih5isSzcP4eqm5i/ypxprU1EH29ETGkIVm3eRePkOWw/115fN
UqLuwlIK4Qjt3hioLq5oIPeh5SsZamjqBm2FI+NqO5cFnQ2mRXwhZfSjTsMa5WTr
ao1rwiCAIRflP/J+S20FAMHYJ1H94AVsnQAbnEpHoFeyA93XPfga/2tprNP7vTpr
k8Q889x8VU2re/wIkMqvicTL0Nb2JAYsti9Pss5MRUSfaaB9fTo1InANeKEJoNil
s08ZZ365vxzTlA1rtmiW6zBsJxVsSUTsU4zKYt6HT4n0j4d17i8p1923v5RyxLW+
q4CRo1K72qWBM/RUPJFn/m8CFhaMcRlPM9xOOFiTw2QIA+9K1XYZy2Wvx+Hr/+Q5
YVU7PalEr5ePGVHAMcEQPViZ3DrJfW67RtLWpq3hbTjDJ/l3QPoCj+s87ct05P3n
pfSwuy7H8B/NjVadqxeHPW3D5oKytdZYDrKfEtIivT+nm7eSU1dn63Qjr6twdPWN
B5H1/8ynxqSGH/GzKRlkX9OV2G17eOhrJSrZvprQupRRYq5zHQfH+PBc2vg9IgnL
5afx1ACLznoFe/HtUpoux3QPPkiH8ds4XOrRHm+YUCEzCKJGPAVLAq1xWfk+wKqx
gtWx4L19t8ee3QlneMenpuCVk/D2gWVOu9DIjmQM+K0mqbKRO4WKt/ojtpoI9AUB
t2IvFrOVan/Q7Ryj72xHSaiI2rIoIGNR/lpZWUwmFpDqFY6/Ivn9dsdQEt5cbXTL
/br/5i4rYnFjMlXOzo7Y7nxLnnEhMnxdD3G715sAOee2UQHs5CnH5a+agSCdyOJL
Cqkp4at9Q6kPKNcBm8FvL9JOhAz0Y92+LVSzk4VhzFBMe1+u4kIo7WD1MCtpiyIK
yLk2fDOWLw58vLfRFhBozzIbD4rJ9xYRJtE0iVzGW0WQ0CdDYeauvk20MErCLq5c
CgHImbimFa8DeLvPMQ4kH9Xk8ZWosQo4/59jwrgb7Nc2U5dyQl8uO70pZmlCGugs
Uu607U+Ca9cx0R5BoglVBr72yOLycB6qgUM4LDLSFwlda07XJ97+fm9IFueH2W1w
isqkmum8bBEh5hzW59Y3B7RdUb1K2eq/Zyg5XyIjhQ0vy9jnm47uqX+/iZhiRuca
SDHcM/on+0u4tMZ5fbO9aEDMGg4Dz4Lpr6c7NJlav7kJTKYlCl4U/dWad9R/QY/e
Xzffg6VPqfZ1xqWydOeUKtES8QIqApzPWFmk1Goc9W2O5mlpr4ZmlSOo+J2tU3v6
tFkQrYUmmKIYQIRtYeYUmsveaILCINHAuBlbQ3s+pzU8Ab0vqQy/Pk+CtgFFKX35
XINvzOL4vANzvr2CB8mrP7wCzmOKu8OvIE2/LEVNRS6Gs+xRFCdNrErN7UtzJ3lZ
q6MsF7McATmHY5LVsRvnw8uBmFXjRVL43Ossj+NB+N8yXm8FIl2EPGTie8ADxZqk
0sFeWnC/xPIajHFIG8e59SJ2IQFObGQrySGbbvEzF/T38Xx6mTQHN3pb47pUvj8K
Rd9+sc9VahDulrO3+IgLC6srLxc0p3DImI1T1XOd/EwjzmPUOIHBdMyVEzOJdGTU
XCEadJfYcHMNHeI7evVVpEvMHOjKOPOIeBcZQKGpE4HGBUzosaawOWtRZdFyGaJw
XQDEZ35XU+Hc2YnnlDBCq/VTuXvOC8b1OMusTENB52i87tVinnQX+qxONpV5rQc7
po6dCqG0f30JNv+i4b2YseGBy+ks++b3lu1/nyvcjSiiXrQoH46n8dQwOcHI8XMi
JO6EWsvu3G/fRiyx8YbxpV8G0RFGt4KaN4RQ1Xv0QqUfOfB5p+5LtsacRqPv0ww1
yqUt5uXXq7TkU77HZnvM2y0/diQEk6NXZKKxtHHtuEqOfjAOczcA2kRDp4XnkR/E
XbD9TmOpadT2oUGdOy0/yGA4QRTQTLcmohEHBIQcHdDBB9P2M/DgVzr9tG5BSGzI
cnb+LxqOdUY8hgRORNvcRqGrZ2iQc/JzbdL6/lHk6it5qfJjVO16EEjlG1vM4oB+
r9oO4XA3yfzrOYY7YHX0XLhFm/o5XjfAjAN3SXMTzESsEE6D8PCnsXV/3Tu0fpCy
yAfxdxwvl/vUDB6MxCkbmaRzYpcyfneLhhveEodOmHbI6p6lVCHasHSy627AulFJ
FrPTKYLxCyFrMZoRQvtWvFMTLPyyDdt5Rkii2/tl/G98qS/O2T4n8CUjPBuKAanq
VfwZV3HeBdJsseJYL0Zk37hZVl2bjzkijs7DalPcUcQLAvYg1jH71nS2G337JKOr
N6X5OHQYpVWDUg27vq0bm4+Bn4ye35cMaJiPjoq86mm4iXKoTUT8JuKjMj7gkfQS
vOV/ivrPbPYxg3FL5Xpsx1ANsrmo1jeQO1yB53CaexeG64aBTAewutwbGw2/e5Io
HTl28ZYmya7Y51UCt4+mj3McqqiEU+JCLhsCQyUpkqwx1CLxVdTsUjHrAr+AU+DL
rx0FBaxv3XaK+deob21/1SoWn2Mwza5ulrJn4Z0hpiZQwhkdHfNGk/SQPbhEQ3xo
jYKunMjkrvHt3LmaiA8PUJiwVkvziF+VrpSu0yBfDCFjXYc/tx9vHO2/NDj7gtfA
rMQdYz2ogFViqeftYpGG1XKh+OSgdxxFvBm5B+GfWyOLjp5dxN3JFCcb/dT2iH6G
AWOSQcTOE9yCkFzgeDOR8JbN5FVHigW13B8VLY+wIVsRNppHMYBic7PDevQ/GvO4
CbKK6MXdJXKFLk7Gd5NHgkXYqjy7T5fi+rDb4M4hIa4=
`protect END_PROTECTED
