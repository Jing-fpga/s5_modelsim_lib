`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2kMu7t/mQoKB4f7iyQmy1XhjyomG9yhi8oy16UbMWR396HMXHOHBZE6jXTPBHFe7
W7z4GHlOrTDrjxwQyI+M9ElBzy9SyeyLnK44dGuMSg1z27hbFL4fHK//mrcUg57T
3DuPJHpVoQV0JtCYCRH+/88bK07nJc5TSdRT9wRaTMsTtkh65PxBzXKJNesDDxJq
OsF+Irm1Wcn9Y3/bDFuAtL0jeqUY/NK7CfQR2cwQ+Ae4oYADzAYtVAbdBm75cy8K
DptWaUTklpwldGqT5suQ+Q==
`protect END_PROTECTED
