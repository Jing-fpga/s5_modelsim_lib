`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m7WY6hTjq9iLhCyBqxDm2XFRrjn9AuISv50MNOaBONDFSfECbiX1KvUeBOOEfIZw
ODyMtdda4Xpy/5epQLtVQKEt5AATRvhJS30iQL7IDK3LsDw8R+V5QuMVl0riXxHK
Xmo9vhgoM5nyj336K8JL3bcMMxNVR0EdW9+GR2ebzyF1+oLTsI0CmjgYAqujaSkO
PE8TDrvD1A2eyl9Q/O8biLaFHqDFN9vWhHlWvQftAdxr+rRfQxcJ2BzpF9ST2xtw
16EZhgTBL/xdbC1ONFzH15vzJkO89gqLe7UItoLHTz5hQRu2336yxMryVOI5qggN
le2vCuXbqzVP641H+T8CAzDH+4wufTWrBLUXJ2+yn+ewpAje/GWC2cECnD1vDfHS
aIuuRm2RlKfVhyxx6vcyXH/7T3JMoeBohvvDV+pYTmJXX4RX6Sih/+FN1S2vLs7L
`protect END_PROTECTED
