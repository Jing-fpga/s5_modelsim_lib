`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OHfoeB9mQohtkyqnGewRsHnwn+55Q4DZFcE0qHv0PgRpyjfZtmv4XrxaXhE3gZoe
gwKm5p3ZImwdGZFxdtk84j+HUUPeIh5gEDdxp9dEJk0ppXEXpnuKS8F5DZ3zAdMk
W2/VH5tC3Sxv4Oc53iBnUnC/4p1C2wCNeVC3fwm8YgnSvRoJ6rjwbLiNMYDS5YKD
6wkq4n0QthaqpNviIpp8qqknt5QcH1nsu3Devf4wAeRCNzKUlCokqkpOto97m086
NI6I5pGsl+eihnia+/qHFFHJi+fX3pF/GI1PqxnpHkCXHo3g3cKptJGq/KInWIwC
Ww3OVWrDI2E7fp0PVj2mpzVf28FgbqU5E4Vw/ixNqn1i8NFBHt6FiGD1Kn/FTmji
caLfFcrggUrEtu+UoFfgV9hhW0V7I/hDKAnPLfxUYwGXHfj1oLu4vs5dzYYkv7lx
tmCsCw2go7ubNIWXweYFEqWBwz27/snvLGF+Wu0TfoeFBJYV+hU6qJDZTuLy62n9
mAoHqcPsL9MsjlnWKn7Tx1nxLEm4cPH4TY+VUFMWk+0D6PwGaLKPSl9yC9nJTUae
UKJnt0EMOvG6rO7W+vGbPQqjv/+UhxdkV1Q7KJI0oWkorONDDE3ESgDS/5yDvmMI
aHjy9JfzyC9YUVv8UCvtPR7p9xc6B8Ry5sO0pdj/hS+54+djUKa1PQpobjIvrb/1
1HaWuAY8BpYa+Xjop1Du3VD5BEIffPjU8OYxx42grsOpGQ9S+snvtNRO9eQQHkO+
vjn+DYCmVjSCDWNe1U8yBKlmRMaRBgVNiagC3paZt/JfFjUxAeOH5BtxpZfVuTfk
xZLjY2ZFF1P/qm3g13D8Z86ggiIJvDmq+2DuL/mwiA87JGp+Fqp4285+FKC4hwBC
KJkeTsxsLKQ++wYdEP5GOGZqppf0+tjBiMG0diXVqpyLOTQvfatTt41CyogDw+ax
JjA66XfMMKR6GNTooxtEYtJnm3r7Q2K3i5nTNc5bA1NMdOygwMRLA2WSUYFpxJqk
aluIVx3m8pEwV4mVI1krjtBktQyRPhMbd6vY3xRTaej+YooHlUP6IJvlL+R+T+ss
1AdQdVyZautAfNna9hbhAvrJOenM/RivsBWtuhHSjxxa37q7n8yK4TE4AHZ5dmDT
8p2wyVk+XlNDvMB2KMahvslZHMKYeiEvzU8MXV5MOoTfyiZEZlP6YglBLq0dEsRB
ZHoAmQvMXzYI8yTZxGTQ0QJONYvmzrhCmbMXsd7cMeN0J2hnPd/Sj18PpZ7yWmYw
HsxvQrtlPRN2R1k96qSp127X1gRxTfEGsr3e/jfTHvfitZ0RAeemy2zCztyC2852
OpkPx6pz23t4XOc5l0Ttwg==
`protect END_PROTECTED
