`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZyByD6OnRco+0ahfvcPy3c7yUGwqLibNtYVG0SQPbe13Wa0SVXWU1S65hZIwnPD+
I+YpAc0Y5/O4dT47+SxLH3DqRWQY7xnzF90kdzxD5oD0CwMu4xwF2OIOH5et9PQv
tQ7xuSK7PFjJcodhLy5hs1u3Lgs2CtzLpcXxnforo832XyyBNFGPLY2uQVfelccv
I234/Y8trsOgHO46xQwc8xt6pDT1URuQHHbAb53Bz87f4GV8iMpGH5ZJvaxJ6E89
/nTY22mRftvLB4ei6v3ROpQbEkvpOtjPYA6RN7tP8NcNTZvfWSH5DIkqri9WUCqw
xE5aHHwovWdvjuacUC5UW739Aj88RkA16OJRSjj12nBfU0Fx8NCLBAu0wnl0+Gv2
y4nzvQgbC24AQt8mU2MJUbdZhw59orXXIu27yThCz3yn0J42vkswo+UPe4BJbNWo
uQocFFV96GnF4/zwg5btWImAIOIxlg8UZp21fkGuADgp0hcGCcTaR5O3nHxeg1Kq
V//YvB/0adnYyZaB+D2eHa36byFBL//EBEHnqOWtNbkTERKA9SfWVYr7CV0EDMIL
5qX1dBb4I7G0odQT2fmQJiSPat4FiWSKDpO2CdeR/GgTJpO7fPhV27UWP1EQI403
C98TThsBMzJEAdyo438YJQ==
`protect END_PROTECTED
