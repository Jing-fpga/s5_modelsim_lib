`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fRMv7TpYIhohXvF0pWvFxVZD6rVhqDOJuhgeo21d+K80KIpp7YzxP11SQGMJipLN
jzDjSP3IWwDMkIUg7PHIxXQHc+QVcd9uRR3sGg9+pTO722w920ySRGQuWoPyq+IQ
Zs7cbRprv8bf2pAAfn/IStGIhj+sgIaxrX9W4qDCsA3CXR9lu2BbUzc9VjWaN8RC
zV38yUS5WKEd2QfGSRb0wwZOukTnYK/B9NDoYr+2LhmC6rCvLZzO7E6w/FnMa9vc
+VXIy+fK2C0Y6aHjkMnVsT+vFOFNyAfoSWHKwxTB2tCWS3uExQSrCrYkcvDFn+FO
TL11SH57Qyw4oRK1NPi2fiqZArOWXG7yDJrZu4yylJitI1u+s+1CrskR7is998wH
pMSLGIZ8jSgAYSQAFn8hnERExNpfZDacdrccUSbWfZB3Mb5oVmc/CNyNdNddQROU
RviTd1Z5JyrErFP/IAPrAk2F8lA7i58SyVvBtPQyZvq/4cBbmRKQnHkjz0Bl4Xd6
C+QWOuc6QiXVfs2NKiUJgtvrURZ1E30XSR6PhLdS+cKQ51k4FosRxY95hbGA499s
2GLTjlp1H52BLu55UtIH/KU2wWmxebQllyhVAqYu+QUNXTRSO1iLPsyDeyuR4kFE
ixuKO/uQ5p+kEKFQdv/NSwy/jnEsOD61eSwHRe9R3viJBGLnctyWOHHH9p4WarMT
CVJJSLBCvdSzv2jZgK7RWojybntXNUaU5NWkTpMHl33tdBqdFnBIWl8KUApOGja3
uzqbL0TLlLmV8PgfXFJL4qLlb8LzLyr2kRVF4ji9EuWUBnh5dXmLE/cJpU0hX+dm
N6H3vJ8yxcBSS2L2O2p4EPdFEKd/WspU9tCIlftZ9WWFKxpTTFw3OdSn6UmypEDS
BeUQnhAH4C5IPpN5/sCxg4Mtp8QU04IyW5FDesH5mzt0zM3mpHPcRceNHWPBGraZ
f7rWYu/qxNDZHomYnIXwWKmPAHyT29yFGRvaiJOqIsR4eWSJ8s4z0rxZX+rXfiyE
bJopEofrWGBb2+u/BBh/nxkNDGiNwP2626NuaiyIyD/1hjDRQN4aZ2c+cQLGtPyo
A+uNygcpGNnuxhGNzj7lUTjWODNnrldEelgTV5TowZCQOUE1gkRV2fkZvivCNRHJ
4IJlVemg3UwzAvqyIyzZPheGK5a5te9L3c0aNXy7LN6Zz3BMxHr0nASobjKQsTm7
mfAVX29aU2ohUAnpTLG4X7RlqQJIWATqATd9bKfSWsWHlSEEQw7nJvDY/Mv6kJxw
LRjY44l0MJwS4ae3q50HBVmEX6Y+tVff2TjtwExSglzkMnKHWf+Gdvkbpvj8LPtG
TvzUz0sG9S2TehlI7FOYke89WoWEpywxVdgymqNiSVNQR9StzHtlFpAqqhCTB5Gg
D2sGW/gigufxZthoz8ubl0GjU+/cRs6G1ZUM2UJh++Rq+A+qLnP3odJd0zaRAr5Q
sedM0MGnxF1Fnt2GHV1i/8qpXAutY99JWnUOdp+J5vn/YSyuFknfgHH8f5TUiOWF
yF+0cUbOSQ02+sQM/zoAlbmUtvo6OEwclEHjmj40AyXqRaLE0Mmc6bQXEDUbVqbs
gw45XVKJxTAw2WpuPjZjCzK2UNpIoUo4Z11MOZYuQjTY8z7bcd5UZpgKSAty8Btj
cyajQs0ze3QoYPLfdaPMWEWJkDhVRmOq7SmIgbNG3JDslRm6HLxz8NL2v8tzuJQi
xywdK5JER232Zm/DPsFQIkwcDFU5cbF8hPQSVb+K4amImSjCZEWV2PFNeFueBXmD
vep1zTqOVEZx9/v532IdwXHqnrLfGIp3fBu+Gn+1Z7uM2r8feQ+7m1AsrwFLpSAi
f2+rTyMWlV7Qxrcoqv0XavT/NKghGaL2HQNQmLmwv2CsmE/87+a26sVjBm42ffvC
pLhb9WQEjk84avuACA8MEwW3HQv3tk0UejP4zQBuecTOxlf/3iCQp39um508BQXB
NfbTXdI4F9OVe0vcmSUlDxKpD9nsMtlhLqtSIm5KdDVYzGnl7FlKDxTbtby7fcVL
EE0aLYBVkHB5uCIf/BGNB6Lur9GhxDY+J/eEa42pRNBkW1lcZjCjQ/BJ/V/COAjB
gbUmse/EXiA6DmBZhKN0ZLAUy0QzThJ2vrqxyJQWMrRWbVMD1aYKll9TqY9wcoPQ
pXjDrxOloKXrozpmq20MFmz99L9LJ/uP5pS+25mSNEATBPP/cRvD5WRHfYwrWxSm
nTMlcBTNvJvjGPRfx9Vfd9kuqdavnYP+1OblcpF4X1HgyyyesDDDzZLrF2EsBx6Y
adxyuTt0lCpg/AV+Tkl6K3bvvsvrhLaisNaa7cm/mDGRWOL/jLZ1eFABjzjj9Wpi
fMVC7lpXMKwfUCl4fpI9uRo7N7hujKy2lg8x1DMqykheBg7kp4pkSzdEFS8x70NX
MVmzeOBkoE6PAl+ZIyV6yPqoyeDX9tEKbxUOuOHFY3LO7cfbJ3ILkpduEoXFNarK
jFAGORNGkxwQXzLCjhjcaB6kcloFdYsrCp+GvlyNWq/amw6nh+rt3BiAQIV+VeQK
LPFj1eRrn5jmqDZgTeXq8LU9CRRX7zvTzKeDUYIhiVnxJphVFYJur45U2JDSznpC
pwmwLZ3c/wnogVYB3QmrMeOdqKnaBH4wAv37Q1tIww6oUkdKk1YnRulT2dTzFRE1
PM8TnjcP8Qud2rijK0ZJvX5S2/lekAidrsAy1ZoGzX9FI+vng8CsEwz+XOtk++iB
tGWublOYfMBXggblbTpIqSVakrZIH465L1OKjc36VrC5DO7+lFgY+Dx0LLEe0XtA
0f9Pa6ylza5OAJDbWGDc+8g00WAoW7Y2PJFm5+ZaarYlgrkR4TZdrGbRPhM87tWy
shlIKNKXdIlmGYzKQQXg0moLMLBsEge0bNO2/kuXn7HVmcfU87E4i9uDJ7j5pC6I
SdEnw+rXtpzNag3HdwWEdfnw2JXb+I/rahQvaa/HjFuJq9+Xioxq/Dpdc305cr06
76DLTXq08OGfLVJJrBXFJUACmQFpeFUMoHn1v3h7WhNrG1mQObBDr9lV8GPdeV7I
Dw09iXeVzMu1+mu3sPrHp4D9YmfBH7pcwQmfNCMXhHf0t4EM4OMByKadeY6suGKV
Pm4/KyhoaH3xxt6bmX2Zg7WyZ2jNmu220bs9IPQT0gV7QCVlnhpxXuJ8VGkeAvyl
8ZTb5xfi2LdULuBPOpdD7ROLmDlP++GWbmHSiMauVyPncqKKyoDhlEbbzy42nIkv
fbpFmQO5xBCPRderHtffAqMJpCYnT/uu7fajddopQSrbt9VEibUNWBTWEbd91Rb+
4oqJtGYZo0UFqnD6grayY28xdfesaZRg8PCHPDtsefuLXEX2X4go0HwSAPaSQAKF
Dh2FNFfFOKH0G4gpoxAnudF/WAi7oLC+b+Zwil9IXT8wpw+zb2PhOOwqWpFtHQCn
izXDPc4dBlt2f4s7rtY0a+dJg3nkoXqQE05sMzGh/rg7TqPuqLyrBpMV7z01JzEw
VljNIgiJa4taMT2CdVPHURX2MBGNUos++BXWaPdjCtlP/JdJXsXT9xI7cTMxSBHS
MmrJW/gC/yig9zerQ9tYSi5+SWbgNoVMf20Im4SdBqQKki9NH6v4zsqh7EEkfwLR
ZjsMUcA3GO7FSY4bGVuOhZXJEfJpSXbwiveZTGwdDPL9RSzvGGFeDGmLVT3DkzZ2
bMAKlhUdIfWF6lNbnbYOJDAeG2th7ybjVLPmYhdOFSH5d8Rh66uKoF2roM4jy8pW
vzC6Oo7fte1SUspGaCzwcy88Ja+B9V54TZRO9tCrPD8BU8E8yT2JqAceCVaP3yd+
FJ0CTt9+kfWYamI/JlcBnWXojX/p5SieocoBRfz/BeVZDQfFrSiNKjVzbrsfpr5l
a5NvRsg83dHa6kZviOBTJKET++ZXfws9D0+BsQqvKZjzaShSJ/I6ONuu7XrxlcDo
EWJM9c9mV59Y7Ii4TW4HPJgKaytjH00SwjeaMgvQho1YGhC5ARbxX5MacNba79BE
i/QtvtLhzJcovrMgU+bLsdgvd6/XCWVKtWkyh82JPBY3pSnoVII+6cubQJHQaKAN
01AjwZxk3o2+tHKnM+ZEl+Xw7vJNP4AgQidvEQxcShyaJLxPWds445URggbBhvcX
FmGN5XXWIhtlnFKrsKKPj2tlQR025Amlxk9VZfuK6rnsp6d8qckV3twvwGfkrcPR
07eew9hTY/E+jNqbfgiEVt+c5gtjmhjT4A9bSJwiog8iWq4chwBjPnKrsLazfd6h
oWsFlVMhIhsvaGm+bEpVAQCI91jA0vNi9rXHgWNgNme7mi5fycAOB5UPTLCSjB6c
Z8I1gJ8SXkZ9JLeJmBc5PamtnKx+rnYwM//skCZxCJtGCDIi1ddczcTeJX+If/nP
IssJZEAHIj6eFsL9wmOfEiWjVVm7mj9ZWnMpemyRFoS6MIUQ1G4vxBWbrN//GEdc
4gTGXRXtKC2jPHvcDXMh71Ab4rPncLi+jpCL+etGBMHZAJexZofL3BOZ9FlQVbAj
fOyuHAAJ3jKEarB0Q0tKk3rdydHe2RfsXfhVS8cBGbC2qufPKnFP19kHEVyXkBUq
+31PpviP6/p5Xum/dGasugKLc23eDHZu63t1tj7M+U2aGiiXySVfHixi0IbXEes/
mLdWrtPD2dCB3aQoyT17fOufdQW333L8IRz5RxI4nB0TWNBLeEjFfEOscUBOOiTs
oBVOb0tIuWWpFMII+xZpsaajHXe5cNQZ4sDGJlS5L2lor21ukYU5EFaUbS+jF97l
J2oOEdVnFG3uZwXNObsy4eVnfbh1ekY9nTR/WqbeovIAvweAEwiHbnWBB5LLmwM9
UJkIDjWfi1AhcppTA9HFKq370EVgKPzOeX+S90FlVFgu6nhWYS5P4dfajrsHKfEW
DQOuAnrEd1bLGCcdqOWituxLbH79Kv9nsnoHI95bL46+7nykXfcf+/zogGTZHV15
RwXPDeImXhHoZ8B7aUmnhDVXdlqJLjY3xFOkrVNIIaSWqnN+xDevlnsd+N8FfUQe
REKWy64i/ChiXG8jc3OyQtZuJk5gX/jsPAQ8TEjJpOhi0B3Ob2PxsTId0JXqwS20
ukhWNf2KoJ8y/HAP+5BL3cvOMN4vtCIKTkUiCBoOBwrGFVF1Qw8XO/hvscr7PHLo
2QvZ/7XOFAKRPzkDQsHFURMCay7rCQzmaZtdnnLrdSq0QAgkMFni5sGGDvSCycQT
xiO31XJKyn7H+cmTDwVD8P0SdH6Vy3/LUx6fB0hGW2KW8Xqu2s7cz8lNYcvfA57s
EAcHhfaOZtMVGllZE26v4HrLLPLgmswGBOE9HUmE5n0UObW2S3NLXirtk6PPjs8k
8Jn2hOApXhLEax6QLu3cERicKwBZbVwWWSJN48v2iQyutyy8J0BoNiOgxC/fynsR
lN8jpqVro1Nav0t9Z7Q+w2Uo6QapAmb1VQYxC3U96JfZyGyO3Krc7HxtahOs3Uze
grpZxvGBLHwGuv/1J04afd3UY0D9MZcDrEzFcq/ljCyqqTuf3QSygpYsy2T+hOyh
ScGe3HbneK2UNAast588uSakJTAzQnJSDNOhDCgfQfpER0/HCzf4vei3V+3QiKys
k9gxYNpFS+0yK0Ezc0HBxk1Z8Uf3fxqDiC0fs638QBc2fSd9WhqDkM6R+NhkdGNo
ufoJwspsXGp5nMUxDXtpYBuE/5FKXrkoziGAoMkreKqS0PGLQR4sOcNYou17a4gr
/+XqfVcR4GQB7CA4JPsld3I4YJVoXcFsNdEYZpyWNUmSRzvxLqO1dNliuGLyDq06
RlNURCmtzxPFbduFC/ygwavc3UYKDkf+B2MJAkMUP3rzUf7ixU3YHtY60UuincbR
kbmc+4qQCf6Q6RyI09ZsArwf/v5ttL+nnBUlhNjQ8wXzEi/kcst+ayoKsbr8Gq1l
GQYXA9H/Hmxa4tCzKLFEmQ0rdV9ciV7f1bofbAoTUsTDJORIyyVLrSNnRhxJDiXm
GRSqn2YTnxdq9zsoyM8WVFiPg1hI72Af70IdgkqZg2M1NP28j8cJgn+P0WgmkWXn
YJu5mlW0p3slhI1QWzJ2vShYyyi1/TGxZguenhRWIZA4P175icWrr+Lv/QhBwzDl
vQCaUKrrqu8rB61QFJjwCeDKWZT7rYaOrxhn0Be7cAl4Z6yK6sczbNj/JYdmPztR
03YCc9DwuMHgWqSF3kauIv8QqQuaa5QX1TMwh2XGAnILwrivbxuCb3cmDFWhK8lh
vkdpB2H77Li54iKMH9ygKjftqTZ/09bTV5WdxS3jjUfjC3lYoifoVsJ9D2fey4vJ
x+/YyQfP8O0eb3UZ8lilDAlI5cE1/PYkcOEqoCRQQZImX5oeUDsOVWvH1/h+bIAd
7N0hIhn2IyQIQyno9Ly1upIBzybnlXjahUlleeYtlOI1pnJoTTk3K8ECG4YMkdrJ
T2hcJVzmxDDQbaFEH/ZmtJJglhLQp4VJj8TR9BnBqUANT5+MQJ2GtjcTYpsHKLzi
Kv2wWdmegJ1qYB1bNGl+aSwbhYOzodEy9C/joQh2N+eLLAmaljIq7bB4L1S4Rg3L
Y4/ilW7AffhYpuJ4vvasWyK3vECW9I6XYKmVjeQrQFdFjO5gS/ClsyJ5cJNFanIk
MbH5+TvTwOzm59RmlK42jaIag/3zchn1LpYkO6wYwdaKgDbWNGbf4GPVSiq/sbb4
i9/6rcH8nY56VL3cCkV0QPcVTstY5KpJ1GBdqS5NzLW6X4PAz9uyKI1o2y525X3l
LgHN0kQaW1Vk6gST+hi+kPcu7Mr/KJhHzl3L9gC3xHC1NN5ceH1G7xQUoWi2bkeU
LQnbgnYZ/lXpcQwKbgykhP1h410ewFrupbN2TwzhWKNR942cJ9FcF80ChcOgaiaX
/ur6+ct4SRXeN9/aRbad6YZUu7cRbBY5HtCVMbUbenKCT85z8EHnh5JSNGbj7StB
RZmaPO8uJDmmJV3dvpEshbL5cqy1GtkN3/LG45c0H9CybzyQWGCJiPvVqqJHzEaH
wChrkpD/p5hHa4NPDGJ0aSpUTTTR4qlnOVkJZ4wTaJ3b/9TaK/kkjCUC8Zjuh2Tr
J/ogwMO0zrbaBezKvuQOtUkoWipuSCPJy+/NhiDQwLEbHdji/gwCmgt+k32p+LdX
YTobsHEDxHkw3QhosWTzp7/qdvubmfb0w7fGuQqR+zRPZH1Nympf8wnfOfgPxYbe
Xgmu5frMFxVjvI9HTlm2JfEVk8KxC1hdh0YQb4aLuLK31vKKcIIHPcYa9AgoWN7Z
DU7ZtYHULrqo+j52NKk3sz+3I7yXpIN/9VrKT83RUBbIrlOW99yGBs8B+KTfSn+t
s4t95iBHARSE6F4dEuAG3kjx2iQniOjZCRUcSFLVJXiMVcZ3p7M8t5EejGtU9EMy
15e6mcn4sKkuhtQ/mzkIjc+j8ISAYAQX26hF4Nf3X+rxUyV9KZZ5oxtedwiCLIii
0ObHDq2G7Pm5XEbthVLLVrdiY+ZbEWcwxgCdvuIWI3TZ5Ln/AARXkokZUSPl9ofT
T7EIkN82Uj1d9LP8LAhwda5D6S8Tq56on7UfvIsLyMZaZvY86FA6RohQFkOoh3f3
i0IQoaBEYJsdMOlRTXS3l0Lzx8VKv5/BtffIXllfQwJ7cPImxNsu4oYT8lvohruD
1PUWYGGPcvick6c1afbCkmSJZwIkMfzC4e90IG+Dyd4HtI+BQWPmbb76FbZ0anwI
vnLlegFH+GIn8PLkIrKpCVmnfsxg08+wFFFMokaE0srAZEEY9t2vANPO86tL6MkT
enBfjK9BvKQM+tn4hRlV3F8ChE8TJYII3Oslv7IA+4G4AxtsSEqWgx9Ltmpj3hgE
SMg4J4BuI6+C2x2O1dH1oNyZsfxqUX/zEjSnisHcjtsgl5q8BLcTJIdBVzzYxk2v
FiXiGy3yk1KPkjzfk56M80azVfzUnPmXYdQi6gDbPammrqa/DmYVzYkuDKghdqPj
59sbC2T3PPwhhcvh/U94BRKNHxzuADM6IsOZhuHZciAQ/OcLTC+hvNQ10gby0qjT
FiiLL7OZWwrbmtlIpqUHJ+8Zs3OVQDeMYxWtKmMmH2bB/iddi2cvP7TCmxW7SHGp
IAgPIMNCRFzk7NGua6qzRNXeN0WhyILcrRF7GWAtWQ7O0E20mDWCXE4zhEveWWAs
VB+9Iwu+UqVsFjmP2FOlLZkHArQAMvuqUXvmp5P8rpsjN157eYF1b7VtrDXg/loG
e+4UhabEsG7Cx9UN8K9qYZTUkePFLFjjupE+n3ugEjaQQDxOu/ZarmLKRCeXXgIq
6WbMvgYjNCp7E3J/VC4rl1bF//UrBxkEX2GTojTAcjJVDEaR2SmtDKiKvTGzw4fQ
ccJ5GTNqkVe4/sGmxtTxPRnzslesJ08BiMt7WKuM3oE/8JdqOwPtrk2QyxoQR4rx
Ec0va9CIK8RgK6/bgtF+utPqPQsytyAlvmQ/0ZgElnlY3oF12pO3o9wzGgyKiKcg
IDQnyCs95BGiZJUcBi5gkQ4W1VhJOK/wXzNSVdw1Nv/vVdjvTJhfqfkSW+SeDPQ7
e8oD7xU6B0snE544AYtscBopXI0sXnFKLcBFD98sbTLdjpJxoEknlRZ34BYUswef
hgxXyyywRRqd9N9AO6aAjK98XAYYV3xuptZIi6f53PeVGVsdvhVG8g+nHFh6JBhp
dFiKEvhERbYrlaQxBNR/Rw==
`protect END_PROTECTED
