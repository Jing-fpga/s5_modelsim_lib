`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pbJEy6UV3ML3ehiGieXrJHgLKrB5PoXvGX17phUzJOH5xWMhSmfG3x1m9h0lroEL
azwSfMYLW+iUNVV5f2bPqpE42z52XBy+/STpnGIou4DKsdwYMgonyxYFdFkd/D0i
5jjhcHINygyhPd0p5LetPbfVJtFLAGeHB31FPAA7r7CGiq0MB7B9IdB30Anx+MJ1
KQ/03anPrrSBU8PX2qS+JA==
`protect END_PROTECTED
