`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
68T4q+xRVvKS78061YH37sr0XubEWK5ABfPnHXGi8XGGfZ3g28Vl4Ej9f2gGLUtY
7j1LmTWqRUbc0rIG0utRjez78JrxKWhzDNrhm0cpT54xNu/+GhDXCNwQBb8ev4cQ
y3iLKRI7+XoW2YEwyhXLhxQaoIQqcP2VPD3BUy4m3tLC12k2lro4rQU1X6YeRR9B
+vBkXHln0nqG+HtjUaCLvYCjs/kW3vpoafD8cX1uTCHUKcmH89NnOjKsrlAfjiEy
jxxQypT/aEwpkU9nUsj9wimQ/htTxL0bjPEkjiaYU+a6JzIVW6V2J5I15BqRNdSB
osOk3GY69IZ3CEC/Wzd2hMf01ItJneMiX3RqVzCQS2WWdi3UpF3kb2n/nxAJ75vF
RXcIOerWPGhmBMVYKQxe/AESkfyyyvfuqrvAAe+G1c88cJpYgmcJI9EYjI3oET9s
ocxs++jbDi3tHq+c60GSKaPLwVsvMQH6D97MfOlNwq71APm83YooY2O7rvOh4PH8
sHQsZ1Yqdo0/48pRIj6EFmSSym1WRE/AHRxcnTNa5/qFKcGKL0wmzCLep+/CKrNu
nbcoDQp6V7Uu7DlKgCoY/UWVueZ/m9kxKw3D7HWXF5odHEtAsgtsBssOQYxyhXFC
oz1SF/wZ5Jj6LVKDKE0Qqsop8jVRSYKbVPOZ01VPbKAz6O0pavZXlHOVJ2sQ34+9
P0zCBQ8Tb5V/xfbIpXBeQ81jizgQ4CauS17ooD11gIVQsMVlEtVlFvPfgfQz75nC
IGtNBms1b1if2ogTKuqpHIR2NlFDc20CpqjaQKnMwEyDxNY8CSWbSjVUQQsoTHNw
I5jMNTp5XhyBMMyAjGQv2TmWNcvNZFlec7+az/vBX7Dj3HRHx4fCA5kF2/Lvovtf
oXy4B9WO7BScCqcAoyU43y5/1zwa0lKakl2qp/iOUwugh432shU50P2+Vpj5XYK1
6pklOSR9pOtmI8iDwSffTEerawlWpHME0CHFUyHLh5CHovtHvCZ8vebq/pXqcbkU
uicKuxLmP4/H9nNW15Ix6YREiakGrYSkOvE8xxMHVNUZYaeYPiSHbbkd5LlJywlv
zO2UOv947a5dl3QpR59qkB3nVZL86TmQCCNeQAcM72woyVFD6u5ia9HsAxeXUxvp
4cB5EQ/bCYkmtvRjXkNGUZ0cPrbBTj+Oox0smPpXRGSsXrmdJ1s9IsMovOEKUbNP
U7eDjK20tNKPwgVjlJJPxeDMEN69UIpHLsrD1gVAODq6fvmTY4XK7ZqFg8OjyBaK
BdRch0l5kgGx00o2RwKBBZWM3+PwlTavEqr6HyoxhNw=
`protect END_PROTECTED
