`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VsKUpS/lxwpBA+vzpy2PzTj4k2xizDudp+E9FEmEycBd80rD56gyO00qFsOKvpOO
qWBrij2xKRCZWWbuzMONXDCK3m6eiVOqk6usnTzxLdSYm5hR7Mu+nkntzYQhfStA
DezMyzMGn9k8QE7w/lPVhl6i3azEo5Wx9s4c98gQxwE52ZuzChGBV7vVzFtJ5v74
63xpuOuz+QjqahWSyE2fJzrnaID/+iKXQ6hhz1QisY41qmxKTkipG0UR9huOTIJz
POzyU96Glm5ypXqxLTWRJbBAHYpvFW60Rz7nPHKS46TXx3px3hhYLVnd7VZMGstb
gzRT0vMzaLNZSipvvAT/gd60gfJI+jQi1HBT3y5m0+rkSlKkHGHXx5ns3RQdd6Hi
ayWx3rCQCNiDayUMYuAAsiwg0lCevH2i7kpCKFgHB01qXDYatC2IthNh6cMOCxFL
ht+jOygHoMu3NX2veL+Gag/+Iu6nLAjdXX4HXe40R1of4NNUqWVSitrYWIfyCK1I
vsHR0vN2uzAcu5IX4A3AncTdGjvnsyBSxsjfVReLEK+mpBLKxaH0OiObyKW/ms2o
Nn1IQGnje1fsJlvHEXlHq5rwj8t8ieE7+vUZ72w0m1KE3WlHAsfRjCUL84YXQgJZ
slaYaRDVE6feB33BR9hz+FhohCk+XpjEU9/kEONT4xWCdGDdzE/HK+0ARhozcHY1
b3eak/+nSrjjueWxkZHxNtkvbcvWKHZogNb/rkp16fXTyPGPdLgLuGG0lBrLLRYl
V+++lvmWchYs6NoArKxR8df2xaOSOeKAHz+cmvTPHrrCMuDrpEMpLSmc1O+qGc9d
FU39k+OdCm8ka1rcdxQaA4LGOvJiYBUXiJcjYLbfni5uYuZxabH3FuWtapy/5L9K
w1/6LxQIxdLpkqv8M3Ex/Dzh1yHBWeWTlc3kta/bf85Wgsozzd5f6AFglMtBX9xz
GiGpmmfVyyaCS0wkwjRTNy0LB7BtAIVW9FamUAWqomoEVtyYcbU2T0ULM7j4TcTS
aBqrH4S0zMUbQH8OrvVaJU+8DYdhsNd4pqJWunYGsS6kLJeC2XsgIsx3OMH1gjEr
NUf4737/NkFU1Ljf94+FT/YvMSdSHxgQb0oVpxp0TPFF2zrT3SjDp7Z5RjCOJnus
wAQMlU6JMdgle7xexi313TWtufw/1ri58m7jmJniAi7bZey1qymZ8wRP3uC1zz1u
UeaFtXd7bc42vOMBsRDNIuMtuGaKqxi7CqWjjqU120nNtX0icQxpWelOCW7OEQta
qBCHVAZft8FoV7XFITks/OVKfeb+7lc4suFJIrdtDthCnQVh5/JCfAxN67ZTk+pe
TLGwUsiLtgWKrYHNDoOBPdTtLQJKxFC8kjw7jj2VZULdvzuQhmXVDJYVBGV5xm8x
kd90Kh99HLsJKd2PxaGlN1aXrleKEB6kLCowqQk3TXzGjSAo+n9+BDY/aMk0CAJ3
bK4C8UYY15UHbZjiYTzUH7+MTV2SVsna2W61imWpeu0HOsa42+/q3cAnDTjpjWZu
oF42uhAjfWguyS+RtpOYZp17fpvGTZ3ayRxB4St5nkK4LD4JV9QFZTXS1mep9JXg
G3SOQ/jJlC5LtBgrBam+CWQ1sTqkVJSK84P2bKd5e8HhJxG+lGUQnChov3LP+Pku
Q08Ncq2ceVRY4Ni9Zlr4o0TqSKd6D6xIalxIqNWtsJfSJPLfRJjv5e2O4R1dJ3HU
/dLzMIPdOpKDyEfceuB3dPIBe9vdXzZyZVbUU+mbt18oPOue3/GVAGgXK6L0zDTR
1KxvNek1geSrU0pUlODLbEzUpcHQcovx8MpM1jb2kq+HDZUKCHIpLteQTQ9LHrOp
F4lpZ3FeN9lLb5DhJ7V4O+pIqe6TY4+UKH3Fpe5WHU/RF+hyFI+fh1eGIUoA92sk
eHAAzrV3tnZZz4Rs2tjPGhmEhAp8OuxhflT4DqixgTyw3/9EX5QEzFTFWAcMyRqe
+dc9XlxJjsBCZui9dPczsEvY78Ac69HgkdImzZ1mVhMHUNQvmplTBbg4dUDzalPU
GJ8QzPv4b0GFStQZNSja2Y9bCZgNpPo0Du8dVXEOwV0mjFr2OTtW+tHckN2csOth
s9ruluDx4tU7GPzd2i12SbsfpxU3SORZRBtF1JLzcrz42bYHzVq1IC0i6I4znVDp
Oqi+C/1qicY41pmJW2DQeY3KTw+NQtxsqojIfkkrRJxqBHdkXj2fGrhg7YkdyQXi
94BnIhHBktNZqy6bC1JdYF2wfO/1FD6GcEnLPig+2GhwWkJoen20zM6EYn9jsKYX
xImd6CCbONDHyPTLP39zYKvVChI2bq6fG6ryppXCNJr5wF/7n1JX6jHgyQ/a06u1
r7zrqH4mCC5Im7soJx2qDiUO6GP6sofo/pi1mpecbURP7MR5L0uP9kKt0L2wTd4r
jp9SIqXKhNj5cVyng2qTXbK143oBO+sBdld7c+a2NfUpCV/k+VDa4mvqT8ONbbAy
1lNVL6+CBOWpAoG+KLq5/dbIbU8eqo0GYLLlMWCvB8pP3bOiSK5RDpaWd8ME/WkF
uluQq9RuVaBm+OmdZyqZE8799gvTjpkW4/ag1wgVuxgyMi59hpgrGrjovHi8wYpa
5X1Aa4FtHcIDgbgvDkaUGILnKrSXErBpq/6et79Wwt5/f/W2mDmveLdWmj8Gl9ht
`protect END_PROTECTED
