`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gcAnRxliR73mVG97uSIOjjH6O2STmh4XVC1jlLwVmBIz8TSctAAcnKxaQA+9mLPS
kOsTNdiMYS0alReSzaiL3p3o6TodW1BR55BhCSHMu2LYxI+FigVLVQHW36KH0DMT
UZFxfsmCCMNDP4zGNEBmDI2HCkCDN7W06uOGbPnTIdtIyTP+pS8Nw5SXyfTyZL20
L2bvQCH8/MfMPHX9cS4FmdOrTV1LGAoWsdudUZZcUNxmLvseRpDoB/d/9zpA3mtj
Rcv9r2RNwWUCRqizl5uBRV0EbJGBD/yLv73yAt7x5Bxo50mSGKWzDy4OJPrHk8n0
XT7QrQqCuB/BtvigzIN/MwGqBqr0TI5yg7RlD0dc8Tmw3foFWfpp7Mzl9K6MzLzE
e6PfE3wviOOlnRAefnyyTL1cmgv5HDS/ns+TJo1RyUcJT10jkcw80OzKMXG/GWGu
R/hINolgqbdfRi9sqT2IiOQSVRD1nSR1PLTBVlhRgd+8CkqstHNqwY1L6oX2sFAZ
nW7X2UH5ewRzD15qU4fu7BG/MdQ/o/+0mqb9TDLNEqyOLOmXy4pW9I74TIAmqCZV
RHcNzcwZqiPOsS/xNw93lhPrH9Lzc6OZwhsnJ18uBNdDgwTX3TegT54Sz92UKg7G
z8GD/wTuC16O1IsExFnz0xU8J5pM3yg4mr4zXC+q2FZsb/PG0Qrs2oheOjDRYd/f
XuULBx1iCCBt4Vvq0+HwU+Y4tyo8TSUZP4vtLLbweKkxfEH0UjJ0RMGL7zD1qIxJ
8SSTYxvvAwGVVo+bsTKRB5J4V7nL/Y8z3Av8q35SuEVi5DEW0Luw7I7IUbhA3uGP
8W42hzGEmZSiJITscH3SOLwSccSuBwOpNS2LhocTaEFDHx2LyvWh8ToBP/AvSCcT
i945ldXlIImqw6NYqLS1U9+FCjSfEIDNn5GiCScbLdTKWIq+TyH0S/TzLqv3Kg5T
hkFP3RcezonW7oPWU3y0UeFT98EL2FJfIPlktOq2WxQZJOA1282vp+NRezNZDcyS
REOIWPP2SxkxKFCCZXalO6hgsIRkPCXYDCFQ1gSFgllroLhsk9nua8i3yOcutIsj
gdhVZR70J7+g2CMnXcFwdw1QYKWmb3lrAmzQOARxOWK7Yrn+zbDYEEre+IUcwqgI
baS+tFEBOp5iTPAfAf6cxbdzs/eT11QHBMmNBGLI8eXGhOFkV001L6hiYGU1VrIH
xeG19yxXCDhknil0ckTldW4lPJvbmrh8AYG6YigFS144g0WmFS9Q6lMlVjjkF0RG
Re1+VrFDpx0Cchd06EMBtTHpIcC9kpXyWiQKlMM4uCprwfpwmdBmFY0ngvRb/8Yw
j19s5F8nEeDT2m/0kF9/LLj52vJCSz1Yb0yfTEFMczwkEiliKzXKqGYxPxs/pMh4
aN0/g9r6YJlfIqJdKoS0vRQOqxEB/jUhDfvvGrcqm3zu8wWDF9xXvWGY2oTzSqko
Ksj4N8h9OnfADiAVIVH7/UIANDSNi2t+bwNuJ7Gpie4dYoWBtqELN6dD/hdmdjDw
0YBx/im6qXfLKhHCYgSEUZrBkXBqf9nlnAX6tMQ13u+KXLeFnK9AxgElpvXRA9bd
KU0u9t4dp8JLerpL93IwUpalYtY4g7yDX09DDnx/iJAuBXolP+Wn73VFz58fJDvn
5f8pnWRrOKCwXSLunaker5cu4PEHY/EiqEAltSPPdmHRiFqPnP+/qhknmvdgK2qM
8aYLrL+lzC1Tx++Fq7j+H3figPd8IiSfFAq2QgEAzPFZBU5X2aKKRMGbOJ9nwoDd
y/HjWQAzXcpCO6W2n1SoA1JAXKVMN1atDPjbROaWiZXEK90a93A7BuDRq+SN2Oh9
gLf/glA0SuUSXt09Tt7ddfGzn3wlJTNE/EZxc2r7CQo1MlS0MC47fIzw3FhnFUfm
d/4czn5QyAsthBLtt81v3ygAhBPcRJCcNISLJrSNDfLuypnzRrVor8sC4134uNel
yGDLwkt3MceeXCtDTdrqB+sfqAH3LkkKb06zvEzlgZM5XmLhpzBdEpDkibHrVrlf
PGl6ACZE8ijcIIep7fIya0ryoC6SRBxZWuB0iQ1miwpq6i2ghdRCeo7qrJ668bOT
Kokzhq/FH9kOtN+1Xs6FB1guPcGX6HoKFwbLpySVvc3jQvs17Foh2MqBJUuf5oM3
6/LKyrlYeZCVd1ll5zyZLPNAZInm/ClC9kabIGMr7G4ELcQIR9YNgY6qQMPTXySk
Y5mOc0oA9BMnBfUj8l0QVJlPcKdl5XUwqpnrwQRYsR5R9s4wBD491MAPfu9wBxud
jDRB4aZ4aXnLgCDSmdgagqVaYNWAi9kXKf2cLUjZtQVDguPBwBJIEDch3gAo8OaI
ZDoy4XjAD7vWqUIdS4bU1EJzMeFNGKcTikkjPQ8h7SJ8sd+5kXHcz73bHhZXE5kl
fFSWRXRUR71paDakuQVX423urx+P7cUk1ZRpcWZNtTCDTsvk6BAnlcJ6irfnkLwu
MCtfu0e/BtkP3ReXJ24jBXlitDb5IxqMDE27uOv3k1C3tAf57WgDhYn6ymKzzSIc
veChD7I8Y0uH52Qwmmz7rygS/wie8qUo55mRuPE1sP1jsVLqWc9MQSUo73QTLF37
Sn3iUgKVlCEXPS8c0fuNvAUffGniDvIWK5QNurB69uMzyBRc5/rfhHDp5vkOYNTE
/sMeOLpfpwk1v/ETjfo+bItwd1RBkQmuh0fG6iIeZKeFP/NoYn++Im1laZ13tnYJ
LFL0E2MpKQoq0KIaJcFFsh3OLLi1eBFLIMxGvzbuUFxv++3lG86LlenqJGXEgXDG
jn99nx5uoS0akk3AcBRY0TJT4wjTl+35JkHXJrnqsGE=
`protect END_PROTECTED
