`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mS+QT1QUuEY1gfjdEEN3TvtheKIZlYI+mQCQZ7Pd6I7cWYr//fc2nYG9mL6z1FDo
wago7NiVJBNU/T6s/MBB/PZLChludZlASiiq5bctc2Fwkza1w0P+446kvg7CeGQe
TP7KwkQ8RJZ4ftTGc1vBqSU0k8bvEf/e47laS0PuHGnb+041DYrv43tXUkchNbnH
KCaCgr2SdXozMvR2fcrZfpwYZLJjSl+iaNghqAUVKyTPmhnfNJPCOGeTX8WPg7Sh
ren8hSAzAYwGQBZqs3wdp5O8E1PkO+OO2buhr4Tkp0B3aGDIwaOlXbsfXtPo/ann
Gu9j7YcSGMDAQXD55FrD+RGyP4rZLpOtRAT/ADl++fFpTWp1reqFYTKmptIZ7+C6
Bd4PkWKZJ7GNJZAdbLulaEJNzjOXzWksxAqee+9vBZhydpUfuY5UfsZcM9plC+/y
3a2dLfuB5JBuRmGIN2RVsQlqeKTa+BNOmLtG2GhW2mqpEMZNnGOGj/dXFfnRvCdR
Hjh792hbnESUXGYdnZTWQ5BMMemzBlIZ2KSzl5aFmv6B9CLOTE1WTftwP5R+r8Kv
xFwOFAZ80R7zyue82Fvga/+VXa9SEL2LcR2Opi+/jm0rQyHNlI1eVBREinpFuSMQ
IXKV1QsgbtF2crRxAPheEkue3j0vFi/Fjst8TjUsZUsKUVa2bG1RRwYTPEF+y/LW
5qu83vfuFPafL/8BmCPLIiCKZOZrYr9DoYvYfmjeSWLK2rjRB7Sg3yy0JmDH8Xyu
XZ3FAdWteCnxgaU0yu9XOUuEFKmEi8oj2c1SlDWB3CoZSB9JHPjEK59909DENo+G
StudS78c9J8ILVNOPxylFe02pyERWjR2MKbgus9lGsmXwsy1tzGQVnN9JTM5SDUc
DSnoFZCNGbmhgsSRdg9BWRQerGqr2KCyOm1islqqSGQ=
`protect END_PROTECTED
