`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2gCoSPmBypT+ME1el9AHMPQ2MCPSJ5rieHia5TkvJjNEj165Or/gR0+tveIXdb3e
YdDUDVtKS79GE4GU1Eb6Rfh9VGLf7ucAOmvpPDN/xepyEPQ381nwSP1fb7xL7kVw
J82KdlhfaB/6QKD1AAw6dJGdPkpk1WFgmNZgDV+i4bxM5gFh3IATWLpZDgy+i05A
KYBAgzkxU8qldpUKMAsLsaaEllUsI709dRbzCWP3kcSduWzEe5c7pqTqN3zW63dY
U7Gdj+jt4dMvXGct73b3TnnaA5M7kzxn4cI9kX8U7PJEepS2S0MIJd35mwWa4m34
JbNgcK0U8PVQaOAFKxGOUnNa+c+DFU13f7yL2J3Eat6E3RYQxlQeqqDyAcYAVjzy
ALJw0wH9alUdDYvY2iIhpODkQRm7RpfsmVheGkmBTV4Wp2SbMxaA6ZeW5URWy7Qj
QVLj96IUYIfdqZ7t7rkudhKIMLqE1Mux6LM0koJNaYFDc572NPQCdt7Ky1UN4aOU
j6YVEQtfCnrAuj2TS/XHCZS96QMlXHEnPHNYBOIVg+5pHY4YwYsUdRVlNvz0sEyj
pBZ8bLFYhHhT5WGdAXZywhtWt3r5nKA4xZZ33wOhoi7BoPpxb0dYtF+UMU1N0uxI
bzkOJ92/mA9j+YJVMxF3XJOYjBBLBh1ILtoEY8JsgcQVcMmBKX9M4+27foj7sVSS
ToCPwCh4IYZNwvWJCb+pDwXCaUbVchJ5137KFpn0GubjOAT9VUjrFaHOxLbor0G2
kWopkP/NrTiptTy5ujDXcaseQt4m9hhaDN/jJkEfLjqDHN22EwAXxpcmYDD7Vn58
koo/TXbRsFD8qqd8FSJk3shxrtR9B8iy1+KILCHMbDv0vxgjXHp4v/DdzDbX2nxO
ZZZO1aT84x7ePAC9g5e7SksDNYaS+gNcZJkFzF4yrrPsjxS248eUmIt5YxF3nPUw
TnYKkT/1axQwrDytdsDWJJb2cZOo0pbBb6kfQx0k6mdIfnuJgFyeSN+3cYG6aq3E
Gepyl7HAp/5Hl9hd5JRTKH/T6dX3+TQ5Afj54jJTry/2XzN4R7dXeL4xMuiUsQ5K
mALaU8Su8qO59UqMgL+hOaUHVM0Fnldm0VpuBLBSuqJBIt8MTABVUGflKIyY+Aua
igPwhJuAMEY7w7/2OxcZAd8oXOvhNsTkmrZudppk88PpDqDfmNNk741+sLvyZsQD
UnrhB9zm8oQoQikUub8DkCgc5oc062VKa+ekgP9jazgf2BV5dARE+aJ6VYLuC9rK
8JuYF+7XiXajMfqN+lZyFz34Wv/+fKCb1EAezXM+wDomU+3IZuu7KX5vTHQlT3Bm
T1VZiwYkz4FK6eDELARhFiPfg1DQGKDCF5fR5IuOnSOU1LNl+aMhTIiGS7uqXgLg
/aN5NAGzca6N6KyK/TMAg03MrSEX//q9qyUOTjTeYPtyIDBqtnsvqInV/3+tsmrp
LpKTCaddZeEt4tLYy3nDAw==
`protect END_PROTECTED
