`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e53E2UfOICijveHa8rNjrMuVYzqpF6oceswpuSV7I0s17/lEHfq8YMlhqBs09WLa
/lc7kQm9RDWV/IDwZNMGW5gq8ERCHvN1uvQDKF/gCZmfnOMuJy3C7AOV/RxQALdV
+Zm8Rh0MpZWQaefbfrKHroPRZthn1/skTi+PLaOqFkzxLxB6n/c1gIazPTvvaLxF
jD9haL9AvtFMFLIwX7dHwvdrXdaasusFPaUxqENrhgt0mL1FuGazqTaRMInqPCZn
4dxbpabwEm1R0ynUXrfSbnxSlu8ici6bD+xVZZHRUqLY/v8wg3E7nwHrcbNawTYS
rTjZrapcg3K+SSKxabhUspu62vMOk1kAV/e0bhYh+VVqD2MaiTu8AMPYEYtrMPP6
fBYh9ZSQi1LmzkhVcQn7Xwg8kGfcfkMnCm6rOrNddiUYcneyrngFF0vw07D1YLUG
P5vdY8WnScE7TITQRcJsKMQz1RzdZ/skoTDI7SShSmxbzLVDeeu91uV1CVTGaX1f
5h0vhktS7Pwxgi2IN83//Ps8tkZjaBePLmCQEJ01++H2M58Fd3W9PDHs2lkS9yXb
wPEFONewdHiJ+h5lZ/oaFADH2awwnYrBiKcADUWVoPZfXCeCgva4EUAN68YDYFIT
fFaaxonYJKPzCXkARPchNOmOTeYWOCYN4v6TLfcnewZG0ihJRVc+k6uYyc6/O3T6
yUzFEKakViGvPUbHARTl1f6mF3YFVmBAxFOVrst2QRLenZuiDukRE1/dKaQllMQE
fN8nn+K47AXU5EJonWfT+YXzyjXXY7OUAgPj7kHdYzxzSP0v5dqjOpUGxPc+9IIO
XxGsnrHtWI/H5lydNTIY7xpbp4MAemR4esN2eueIHpQ/SH5EiIOyp19RCPs95HP/
Ll1dMEiOQ5o6k0VjrhzptLdRF7J3bFCy+OkIZlDP9lckgRlh0qiCixwI14vSp2r4
0+mIMnT6djuRtgZ4WBhg6yptnj/dwtn6iqNBTDgq93YU++MvszBnjaoPOw6f/mfx
P8+FxDVZ2mSogY7ONcJGIGnHVtIoisG4njOdK4w4DskpFP9FZl/0soERRtO4f/mT
FckUj4n0bx2WU+mMrtE74qs6AFqEmhDy7IaoqAVRz6Vvz6MiUyFljEMeEhCombTG
WFDJJikPRQuZJkZvP6jwUWGf0IW86roUevjjGHUk9sVEz3XzgMmelSII9nfnIJEG
BiaezInuerPFovmKAqyC24nGJO/l5Z0VRK3xiHptuje5lnz5vxnFU/Q/VB6zh/HW
GsQIBMrnKFhhQ2l/861KVhwaKjQula1lUgHdieESKBlaRjI6sfbMe0Pf69qOx8e6
Fyhr/vUKgh/xQxl8+wf9+if2fmXP3B/BOaFMYQQ2fuV/AsbVkJNXIvKtic8dX7sr
Osslb8iX0KaRBbM1Rf4hAwk6MG+CNM9VzOVvokokWNZkYFF49s+8qLPH526PSg4c
sn9wDHfd7IsGxAt9Mu7woY+6SLv55Oq4ol4kI67uJ2eyWMaSsAFR+ZJKblP/MnUh
iauOikd1jwMzrJEu2bcTPfqMXfbvfvo8JkB48S0iWsSc6fuY5Ve0fFZGi20Q0D3E
4kuu0JH8iwOt3e3Eo18p3UFfAfAM/3IHoLcn9gP76td4vAiIgz8cda68kl3qPX4/
xHuu/pDYdp3nWgXZDqzuiJ6q2+vDvxi0SFrCU8uBUu0EYEtALDG0dXVZhFSTrKlU
vtzu6PdGwW53FeoLVDZXdIYczhWVha6XTjFNAAo04zkClQr69YsVD3ajSmZzQwuz
PTy3RLQTQK2gPRac5Uq+o+YBP4pRwrVgXcGLAv/0LUW1URpkEj4EVh+TcN6o4TOQ
OWihtB9v85BSlFgamFPE6aznKJdszsVjAg/aZvUhMcP625O4EV22hlcK5T0CWrk7
uS1wAf+AQk9d3qqOwQy7QviXw2HDAMpHLNnsFAfHHYP5de80m4WS5U+lQP22EI83
nZy9mwACF/ix5MkUFcduey5+I3L+XGkR83ZjzuAuTRsWEFaacqFlgKN15cp2YtfG
lsotRAKsVSA0NaKdB/f9cCGijsS0ZZQMnxhDXm5DCNFOUTURpP1dSeff26nQEcbX
5AgZZQg/9BVVJea6VC70fYrt8cAxPCGFb1dl5/1bj/4pkSEJM2FG2pRmqne/oxc6
uzQAWcIUf7dzMfVzsdEPPP/GrT/GvavEUxrT8WUTv+Gz31p/GIF4+YkbH6wNjI4y
OEVImkp21oK3V2h+37feEtteqwSTB8UW/5/4OT9NaKQ3xs5trSokU6hoCYA8o0e1
MtETj4rHW+J0E+nfifX9Gn4My2jXlcKR0LiDA0Itdfoj+8fCzd/pM7YY6ZBiLw5H
djWC2B06jzjvh4jVp2SHR34mO/QtOSB+M1z6ar+1jCr/FhQlEiK8ozFVGnou3aVu
WlvuTDmp1HkQXbCTm3AVHVXtTkQhzSI8yctdT8IJ7pIvlT99dujA/BnTKpKm3wHj
J7Sles+ot+mCSvW5hedk+TDGvYrGeplSydtp3N30PKefMa9Sp0HF5DhESr19tsMx
cPQnxVospKlGVwZzCzEvhOOLx1+fNY5B6etcOURhryKJ8zCqxkosITkZrvJoBfVj
LsCmJ/iL1oHsg4fy7aBcRRTlFQjFRp6w12LjWUlxwQK2rPxrqV9hDvzQlW8oB2lE
KeFXDslxcj6k2FEhAYuhqMCt6ysxuOVxeAaiCayvyfHZtJUWllLz4QkqMlMxw9ag
KBctBZZptsNr9Q8rVzIpxEQLfCgjKO8jPylKDae3ngZDdRqkt7Uw1osnVXYWDcLu
+pCuqnnSfhwkK7keOury9CleoBznyambl5WPjcHGf7NDYM9XpQ8PrIPkm2wYWoZx
MpXxTC9u+hiPT4ZyhLKCeE+wiN8oJckJkgcl4O89h8xaiTuXAd6PqlaxCPVL/aLt
lbFgIrFWFncZ87FsVEaGEjCLNsJ54AthYXIl5M8i4hryZBJYUvYe6gEMHwC3vDZC
M1zmvHQqK7V9i6txQuYmGdJk8THHNoKScDFCYgovSlodQ761KvBHsTUlyb0Hpm7k
98TCNl+DIUvUnNYUNXYtasZnhMsxLqg89K0zJko4rBf+OCalte0M1x8co1kbCYrb
nM2OwwoErvdCrSmGkB5mjWVhqPZ/ENXvzE5CTVxCSqfznV881ygTumeW/RdmR2Y/
V7Tb6KofkIolRQCPj0Kh9nRcB6Rh8CIT+cgIP79c/0SHFnrL5JLiQCQkYJjbpOI2
d7TFYAzWn/jCndkXPY0vfXmv7xFxbHyhCHyyAdc86CSdjJZId4g8iHIo00WV34Cc
BIeDFxlvRWxR9dLABVoWBabVB++sssS2RoNK8slgQY2p/A1SsGYD/Or6xhbMNrve
Od6FxcCgMIT1+DyusA1fd9HitirIUY9cWMa3fmCSHFOufqIQLO6/KNvQ8u/abymf
rWnuVAxfAoUaIL9+Av5ff6kRSy4TZwtTLYdQWxc9o7Ty+ytsUFptwWKWV/3f7Lzb
xHXyuN+BGTjdGup6g5y+useotqWNLdbh2E79tpsgszyijLmhSkv2YY1vQIPcHxqn
z9oh0dkVzn2JlJocral25q32dPYIozDPOdevOKCl0QFv24qtNeWQ1TbTJE9FBD53
l0NRV72ouw1/BXvHycNE77Gt+yYcL8vaBQWnh0jmoyaRmoBQudoinK6BE+0V/UbT
uF62oguODrFUWI+QQl2lH3oi5yWmJ2yNtbqOGdxi69591gjfD8fDIZ5eA3wh9uD2
LggWCoTZhpvvgWeyQ8MNWRdK965u/7O+gwL/ZGHbrM8wT0HEvs6gwW6oBpNVKTlG
Fx7KY6ModJkvy2tgARzB57ZDBHJ/27+ITxx62SnDuSuMGwk1vGvlE/E6+zMOlaMX
ZhoyrPH5PYXng/NU0x/wcKdTR4z2zE15zTLoYZ1yHZ3L0syJ99JKDXigpTU1onBw
wb94u93deuZcBElAk1SpKDscXesb3zZtEXx/rxGQRZV+GdoRzqdXyhlkOWXaeJR4
32KtWrREyjyRJCxDdE2JyNcQMBgJCdHr3Ht7P6QCefVGG4DfPLltTKqxZxlALU0t
/twKjeYlveo24z3NO9AOTDRPKjLPQwv3PR9GQcZAfH8lRlXJN9hNuBzHBPHB8NYr
vtsBXsU6mZoVzg6c26dUqmeIXRl1RJLf6wx0ygAJcx0kNMVLPFEszUjZG+4HVTVt
9l7nz3lTykbefL/hCZLdfqsgVFKfAK6B2WlyPv9rS5XmSNMGVrsu2hlBEunQUq8h
q9+mmvHvi/nnSZCPumXkx+465J99CsOOqnG4Gg/0iKb7GcfrCgVgqdFpxCu1aPR8
QVSh0D2O1Mbtsz5vPVFt3/syF4xmrXKPvbBG7qccSvBCkFVlvQeh7gkVvuUFQtky
hzMXU0+5sOSmVPnukafFruPYJMAFtrwqwIMTF75M92z/HpsCB7GFyl2gqSUrtrpg
npD31wkA9NvfdUcu3HB+qMGiZQF48j/f6g6OnKpnrjMW2QTnqPb5bwgi6MYk5w6B
G5myfABmd2OXHhsKNx5BIQboGsbUbmtFuburCCqlQoK474yGDi+6CSnHutOB6H0J
NNxRcsbMTLuIRLmRwKg0CCxs4dxQ2c/ZAoC4kWZHOYDfhjGR3x4eIjl1g+WQpezd
MlO4uAZrBa+UjmjQb6553DhjStc6HZXj73Zw5BJ4dCOBpcnRUJ6ZSPyA8vqD9dqG
LLCOLh49Rn1vQUZfj8Q4yxl4bux5CAnLSJyJEEZ8YGp3X5EY3uEJzfE76gnvuXsa
Uq5LuDlWg9n6SH3c4UmjC2nINsDGHHSAw/hlUmdplVXbrXIf8FAPN1gsF3XNjdgT
woWKhD/DQiulwLJDR0ZEYxNgb2etMW4SAVudvNFL7APp88PEkE29bbfW4ar/PiMa
jK9nOH/X5yrUfxZsXYuX8PJAmRBWoRwHc6RXArVrmvLBqe16/Q8jmLQfWOvJZuYK
z4ndHVlahmC5z5PqRbVykrsphmowJEaRdrZmdV4swNw8ti82SWuBb3RK+prj8P3F
dtTIO/2JGy0u6bTh9XQ6HKQQy5uxSWfNXWEx8orZA2jC4AMrn1rvgryWHr4cC9Eg
TGahn+oD/u8yOjM23mX+efCh1F1NAkAWjBwMeI4szRNaM4KMmvTM1p/G98ScqMUD
mwPbQK6Bn/AMy4ZNtu6350LSRY+xETkqyPB1Vlrz8IrfRnIZopDTMfNIPPck4p+l
bUWPtIVvQgZH5jLqP0hSyXw8ma1ru/MFmPY+m/SS/XPSn1D6hscZnLPvviwZPbq2
ysGPcRMi8+tJnOWoueyv15uIkiYhDMdgjryN/oeg8vlaNWord2HRfmf9gbqTLV+R
EIxzH93gTe/QvkgX9y52RKeCkfgnZu76vtr8Erl5w5Mz+rfLPMDqd0q3kIwPVA8L
FVGEK1wFwsI5YRXBVm3n86IUmc79pUbepqNXExiFGdElv4DuzpuSf1cmYsT/Ec4h
o2hM7Yonma70ykkUbm7ASY1PqCT5gmXNqaO7+NpPzJYmw936PA40jtK4zfq0rApq
U9FgFWUNfUUOwFn+WZqmhJVEdZYIgVM1/xONPH10+y5zqC3CQEOj68h8wXO1n+l2
0NJXhKmu0ssBOtxBRUlikumUxeFqYoR3efC3gUKCdap/MBuqUN1x4hAuYbSMU+Rc
4gNjo9wcvYOQX85D/kGywMqCYmQKFbCwjre6UZ4kd75Stfpne9mPxt1WbDOCBCSr
Mweu2XTjK5uJCDFC2nMqVwQxOEX+JPyN05G0WoK83zUtWmn5aCtcKAkx7AX/lYeS
V2NVj0gbLU84UO6wIKdRWbplB06B6vfoSoOJYyGHo4DIF4lIPhbxadii2Hk/cxqS
npyOTLg09nCBMhBmPnGmGDa2RGfWObiAW2gPVlEIIXXmAQWqR564I2MunK6KpqiZ
KgcuQRdl4eBhIiRJwgBpMoOs0SPmbmgRtgLXXYjKOjkd4yj2h4YDIcn2GiV8P7xF
qqn3P4XZ6yKYIqgvtPXOdc+WOPKitAalSu8S0e7HGoOjj0lixm6GnM6YNMfD7dXi
KYjt+b6ZRzye2ydir8Q9mveiLDq0R30p9COwN3dxkJYYQfhAfZSbztSXtvSxdsq4
4J8AVyUnu19SZzM1qXqvfS+9GdXDc/8kJJtptgr192M8RZSb4K2g1N5tzwGFuCSw
6JErmgIWHM7WXdqf18MMWheEigw8S0ZIGy6ApAXRlx+53bCcZQi7Umz4vcsIfrut
VjkYqpPaPZoTVz6lKj7s4H9j2F57ch7XZuluANuEcUsqEnuVqQZ4OxhX6Yzo3057
veUMjf6LH9NTn41Kf0vIKjiBJ2I9mIiGQyTKn2FRbeghsbJ6jnOpxMw+IURsqQIS
fwoBQV+BCfXHPChGEz1YwRA+4uhmRsclR3oaT1KPSPPb7JJbWgjk3Rb4knIuLl01
Tk2ZGxTvnn7ILK0EOi8L2bdWuOcreCKrly/qok/8rP0TAoFKnvJoTFcCK54RRKtu
f5rx2dsN9Rl0RWKP47cbXXvpXdIZ2hjsZl+ppHGJydiBmbpszvQRrut2GHsxsJhx
uZdeUC4gP6nXmkqU3f/5NneXxQdkItSrdGVh2EBRiskt4P67w1sF5asCzhF0pa9J
DLQuNaW0fdEQAoQfoSchBuL2yPs6huQ8b1mkAgzPlj7DO87MKPkYcfjkdPA8L3/L
nRFrG6XiFwX2rD2PKgJeqaTpUxSBiWmSNRPmGwrqxcpnM6Rl2uriFZZUCIEAxLh8
9KiUFg+7glniBqHwXVYPvZXVKJpkboCMkbmVO+OmPh5e5B+oG5vANh1xY1IySptW
yuHOhMZS3S6apL9seySLyyBzTohsnscSvMf05aeD7HknxQoHjM94rnca+SdHTY4H
T3LGQ7/SS8hnXCUgGq3XkwBejjTQu1TIk+ggS+Y+nZWiSoNPIJZmnFWdLPHw2aR6
2tHof7BHJO8hKeqYt3D6p4I97tPfzDe2QTcI3EyagEu3FTxw9myQT13BhHwbt2tH
8mD7/3HDYMEnEnflWzg8djzG3cVJTtfl68116SkZp6udNlm44b1Y9O6VS6d24XlQ
1s1w3kk0z2RbLAeYoDlPvbSKOoPBibYzQq8hAAyDacVtGnjfYZRqjoHUIb9Vi9jn
kwcVbRKj2bMcaiJ48/q4O/AjOTE2DGQ6rjPzBa2j1VSYwl1EwZnmBnAypytiLZs9
qi/fSDWYha53k1HsH2mRhpnd//lCEfsqL6qJCgbPiSS8m/RJm3Iosyt+foE712KA
SJ69hRzmzgcq/d8bGd6UcNvFdq/GO/rXHd2AMMJIMaphEGrnMThKuaUHGC0Z/SOi
cb+vFNaAJr6EicUoNla1FxT3OE/7ZLmtNpDFWEAHy8Vok3vOlJh28XmInbvVpN7s
ZQvt9C34C8++hlTFhNSmKxyjLhGb5uIRa3FZDi7ocmkw0u6xGhrXdus/JUSnOyfL
uwlydGcs1Wy8pzfE59DhL58iL+C8C507W838iVyfIyZ2uHGJQOFZ7t/3TH3hlBhD
+SY1FkD8JkAfzs3Vj2R4wbAp6r+qZ7ScEmSM3boSEmMuS8kDCDokHzHMms3doLCR
Eixr+4X9qZpEOCQjOHnpZSAqwlg24jFSouCG2XPclQds5ZL1vNabOnROkXUO3pP8
jTcnikUXnjp3og4acbjYcZFoj0SS3N6coLsc7ui2Ls3pejOQgJlZOsZKBxWR1UTl
ujqRMFV6E9eSbUaDWZjY+4SRLCYmEKm+h3s31ke4d2GpTiaXRDsYSlLrwoy7rlCv
PGXg/ML5N7vUJQ/Zn+79nEiD4aYTnJxV5P/2xQ19at5hmsnpxDDlVdMngJWe3JXn
bJZ/14up3niiqAwK0lGUmx9gu7HCWxa9hlsivhTuGJNnhkUgsA60p4/gUiVjZQAl
U+0tWIfLCo/kG1QPyRF83JdFzuY+n0VKSO6XXrdAQ3vSP7ykh7sJ1jXdcyENWu94
m+hO3+2JdezZHtYHOwbHdxHUANGnJjpBjgk/KG1Il9tg2+xbyFM8cTVxxqlyxie6
sBisOSEyRe8gWiW4h4dCex4dMe7QBEish5okkHBRnGGvSKNn1xu/2YGlNo9x89tl
aTq6xi0f/jx0U6Dx8VPu2vwRLtQpfNaWhNtOucx7nssi/taj4RIKTvzJKzis374/
+odn+7bBadbaDTq4HcTurpFi2Nft7bcCfeFRjK99WGepCmu4E1RdORTgGFGKvuF7
KxHgO/W0a4/yu5S79EZl4lM4tCI7WUCCHtT22tEJI18En28HeBJrtlsklI/2Albf
J7SbkBd+Fsjg6kvXIzPQCWLjmRnuyU9j6acHTt7wPvylltWEglPgQUnmJYhVTMGq
3DtxAUGPRyERe8c6m8m9a3F7x3VP9b1JWlME+5tpcQYf2V2XfZ9zrlLKdlBd5Htg
8j84A2ceQmDCLnZNAYHYTbuAp6mSNFaRDN2ZUGV2lXW9MKIkswDv6SNxv0pwcCrx
vwEY17BtJGYyHl4Pzn9YCoMHD9IuNWo7oECZ4wMpTb3UW63ywyWyMQigp6sbfJno
ZcPKnyW56R47dKuFGtBywH6VFDkY74ywDxXc2A9Rbh0AkFvEIIoAOVWrSVhy6nG5
Gh9IMyXRV7zuOQoXtKeokcO/vYiK0XysVhgvic8c8lmgXnkZ5BDGVSyGTobJ+G3/
It20Yl8QScbkN1tElyeV3gg3FX95EjrNiy2s/7PV1wFnAMqeX1/m0Wggs+m0P9A3
Iijz9WLWT2brF9U93KUWmXeRF0h11U7/qisUModuaA67y1VHjtEG98CiVksk8MTh
BXpyEFmQVjjzVEgeQECWxqK4zs4zTCbrxPA7+OVupUNggBpkvC0xLAY7l2D7uoFP
5gxE+HdlZGazBpETrJh2gVdlnGdGA/Mbgo3SGxp6rNkv8386/Fk0yRUf6lHx5MF5
UsDBS3O2ETmcnvd/gRGJza9hiul0SkqFUwF5ZeL3UMxv+92X+Bw8LbRmbeqd5S4Z
30/8njCovDb4SFfoZgyyxZXerCkCRIzTlbYlyZE7P4Y24r7ZKzQpi7Pxdf6XJQGu
N9viA9DkhOCgkWfgpJH5NMGhAkJJeL1Rf4HDi5COHk67qZzNgf5CpyRwHVAl5Ofd
1o9oshQRNq/0BCQKT3WYwpTel0gHU1pQWAZA9yHp94k+M/Jul2qI+NnegQ5Edxg8
MpMb9ZHiE2/VC92f2HXQsqIywrN0wJewAZ8/3H4xm+0q7bc3iU4F5gsRpVpfj6Hf
0y9Twr+O7z7epEUPjczFgCXTMmfZBeeJe0FPEK1Yf0rzJfRrdzeeTPBbetG6Ck0W
rOeO7I4VMWlB6skcANoFeCXG8GQT3//YX4HYMwuClgSJhSP0gWZsADP188LmiUMB
2mFgLdkUHVSlC+TnlX/INjMfEvN+J4uKreg6ZogN1nXNb7J6rCbsVIkEHPB0i2vB
bHLcO7b5ydsGoHaMM0SUZlx0mboMbbkJVtVTvBtoyfOAjM34DqHisjqIzff526zE
TRO8ChiGNA1zYlVDK8jieHrtB/SL1oDCVL0uJQimtP/wyOyBP8uVfYsF4Ud5JaY5
iJgXOVIjJdcHTZFWNVpEYyt2arSNS+OphvEZKG+Rnj2luZpUJMYR9KK7bOnqtqV5
mH9drAPO0KsFuJFCMMQdF26waAGLz/8U7gmWSXgoNk5sbc8V2VNmdiUX+pyY7wWj
bTMTpQu7W3kW8quJgsBpkYba6wjCLzVGkKhOyl7llV4Ym77GSokJnkJ0eLSFedaJ
fp7bKWrFwylL+oA/3PM2o+JxH0ctAcqxelL0diYc1yJoYlJYeyUEOQa71cymxypq
R4eI9/7EHh96SxldLvbK4HGgfCgH0OK8CdrAJoVPMiQS3QUx5X53OBqpnWImDznQ
uKh8uS/nFX+GXDNAuC9DYSE2YwhO738ExlMyUsee0hJ6ie8AXBhlBbIj1nl/kUsz
PE4XdfNVTtEMPrqSdPCfq17KpyZw81loCKpalrQHrFpPFmK3z6aTMOmRJG42Q9cG
j6VOVHJ+b8ALxhs4mZk62udkMN44aUMJL79lNoLc7Fp3fVT5CdAL4f2ZE6yjXbOx
Ra/uI8ZsTVQy3Zzn6RINYPIjqyIAroWx3QIPN3Y24yQhzz8tSMGbsT0ZVZzZaaS/
fzRfIdS2cwewN3W1XfX+JSomEDuyMINZF49zzWHAEDbNRaHtTNh/njVMnzJUK+U4
gkTqzQd8g8x1hHHQJK76kLzMfUH8D13ftbKcjAt7YmZ7rGNBBkIhitnL38z39uMW
BRkcX0FWpxV/ohCgyUGKACzPHK4y4KJX6TV30+J2a7n+ganQ8LjY/e/FXwWVdFlj
7gl957Cw8pMYm/GvePFdoKSbae6mz9UlAPiuQPuHn9vaVZ5j7ztN1OX3Yzpf+u1k
9GaZxK85wefOQH6e1bC1I6crMTP4jyaEbqIcQp1J/eW7YYYRkz58kDu3WsbBYXBJ
9pCq/b6BXXXyAfVT+sCptewGWLXVzlp2mdHh0bDH3sWNG2a2ts07H8K1QC+OuUn2
80evISsQo2BrjLNpaUHJnYwbgNI6jPWY1+QbX9DCZv/6dRa3/QuWmCCaigus5Ms1
xRVHrrc/aa5AubhcQejJON9S1mBEPgt0U8HRO9/8nHsGdnbUVBblWdwikSLG2n0F
zWts7S0ZX7F1fYnQDDjQOlv0Ru+38OEImK0HLoJvuCBh03EASnmesMLxDpTgoKc6
idloM4W5OHdXpphsBnUUj0NmPoI8mzRtnoK4Z1hBfUc6zgKG+b1vjdHNiIPcHFnE
IDlR0HfE2StAB6BiSlkXyXmoFu/KClpBPCDWmf3SncgUqWKVzyiJ6B+Qnc5sDdaT
Gn7bZsrb8oS3Y6fpswect3gHS13vYT8AXNmgQcxRHgHclblWFGRY22d5ELBvQlmy
S9v11/HUJJc/x3dCXr7EZv6v16NBBPLU6epc4dVrHsS/eLDjbJHWCnVzdOj1knEK
2tQEt3WmtdZTfnSAbLazGwpbPcep64aSsnphkNSjH/9dIgpknZkWGCPcV/b+cUVn
aM65flFmTI6Wu5hdvNqI5Ggb4wpUa25qEqQ9Rnv1Rgqv2Be47L2u6j03NAbAMZeN
PL1LaVipYMeJNrlWOvyFN+LIhrcWlcWicNKH1NNM5g8rA0Xi199w8vVf8xV6nDYM
5iDis/dCJoZndGDCv3lWAopp0bNc5OquDNLxBFGJQxqCexiCqbL7nTSaEPRDNVkv
rCMNmtW2jz7X3yceXxSPO+tTnmMFe024j2kRuN4nCxmjCc1ZuyBtqhOPpQdYc9rj
pbsvJj3tLPwK39upR4Si6Wee2zSBhudaI303pY3nPiyHRZIqJueG3ze9WL7j6o0a
xPWff7GrQsHc+ZviBBq1WLY2aG6FnOh5nWhqV1HdmwQVIiN/CdZjnyJ1S4sQ2VkQ
B4NHE/G5QKP7wXFu47jb03DgKLuOe+4FwXPTv/yaIxtrCU7Ghef7hQq5AROv4d6y
nzXmvqXL/gnTyX2eT93JofYa6zEjpbUXmZAbnWK1Dk7aSQEmaAcOYfymJ/Np8NSV
WelS4sFdvoIf/9uS5EB4a/THQ9ma6g1jOCksEOLMST577N0rQGvlrT+0o4n5HlyC
yIUK3n2jjk/CzuM48gghc1J20U4FIOzEDFenOj73YmTh/P0u/yJGfPliY7x4Taef
/ZvetZNRZfgrbS8o5u2oeTm2hoIXBaykg82f6X2WWGmt/Fyc4MQtp3tR0NBuBwNu
ZoXVA/TOUwSOYwc7jxH7ZLlDUvuK1F7qqugko4sjodLMeB9etClHSEooyHy7R2Ez
dVvknRfBdnVb1xevlH0w5CEqoKwAplFHG4aDCn216BOhM/dzXO8k3Gm76d/ByChY
ECNHH/uHx1CUNYaRPSuKyse2EcAfTpgrABN3clVrYqCaESdyT5Yx3ll2P+qwKgBa
PIHi8MrIR+LA+CoCPJvIzwbnjV1TQ95wecu+jt2+i3JZ1WzMSDb8y+WX9wi700Az
KIeaGd1oUGIvfYKNfXzIxXKQgSWNgFznn+oi3Ho820iMZUloCL5365OcFGFGhsBb
sV7vl8wwz9m0UAvmh2E9YCOODEfpTwgx970eyNrkdvVO+381ibZn4dA9rwfbhXGb
XJ6hfk7E+nlIEIWEUT2dPfSVl7d4cNVmDgG2zJYsEPVSAVNNWFPHDaC34eNiOKya
/HWrWmjRc64MBq4r+zs9sDBRqCOistNfQZ4+JfB0wEHq6j5bPeI7SX187u6YAjIP
T1Ppbc4XR55ebpCcWHigFbuIRtpjiKsaXU6OVlYAIdvCwm4CUzw1OF/CuA3XcU15
zKhsXe41dnSjofMbtIWx9drn4Ui1vSnr4DWjmqAkKsuujpmnwE1LXKRFK0a//l92
HyPE2hqhuTGp21I94sp5yRNKE8CKqvnskACKTHCF67PF4BlmH/BmLy62kaOx8oiQ
lJrr8O4wjSw4Fne7e3/2ksAsRyHkh4UlpLVHBJTEZMsAFfNss2EDDcqEFiwiL9MN
Yc5zTrxflBew2Ez43dG3sz4fPW8ozqdUSumEHs0QKboSsEmsmcoyp+UF0E+3p7/3
k55nZ0gW7q3nr3zFDNMgHklad+4Muo0tUyfg5zQQQ/Nhof+dXUJp04B3lYnD2O02
mEpXKS59gUzB+rwVlK0XPw==
`protect END_PROTECTED
