`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WleTx+Zxi3Yq7NxABaO8y7pUIUKHZKVpoyRg6MUM3Hk2n4rL/qdk+EwYoSY6bmjs
nYEG2HBXN25dTG7JW0caNa1vW8l1ZsWKTI64BU56Ws6eqVjulmHAD3VxnoBTJBU/
oBgvdqSGzCMJGzRGZwoOJvHXKVn/NP+yndbbhhLqiihCKbss7Q7t2PZOb62UPzmI
8zC58KYBS6IkgnK0mYV7zCd2FSdx4JBvN4a8kTSYwVtn47GN7lPrilR7tQlt67b3
xXpAQfMqq53/F6kGX5t6+o5t74OpCezmqYhKi4FeAIjBDXtEf4fPGv7afyrn03Dd
hDT86hcP4wvXg/2zamYsiYBxeQDCpTfgvDshvlCj9RXe5V5JaYOVQXRVY3AGhokE
XVw+LpJmWL8ahE4ZjAwapzYP4h7vdjdUsfaAj2XS6UQRaWzkMtEQ+54QgQmj9zL3
PM0f5codgeWsHdmyB2DeoMir8zn5UStpY5fjd8ujqaPd2Ni4gu3Ukr5BgBqv7PKi
ITbSl1P/ivx4E4y/4zWHevSJXFEv5qprUtGoJn9RDizvsA4RvIKi6m5Cn7Y/Rox/
dRRPh7zTXsik87xRktWOwjDEBTsSZ/cK5IQU8oVCUhcCMKKFy/2q6+6+YbHjxyYu
X19YPFscchJngpZtIrtE8A==
`protect END_PROTECTED
