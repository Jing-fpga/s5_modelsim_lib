`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WgXfZ4ZYxQFreirbYvLe0MfvfwUWiTBLohbJRlVPOGWdzwflV23RAIENNJtXBI0M
SpCrE8hR1hWHP1ZX3iAPfdFxGJHLM5DUKdZNSUuNBd/+ymw7ZBdl1Gbaka96O4Kt
NN8BwQrwe85P/SjrLef8okWQPMaAMpVLjJwZfCH115fWerfFmI6Awmt9fKXc8k8a
gJHLCuUu+5BSO0BLClsbjcltfGX2O1UBGYs/ip5W6LskaYOKP2Rb8KTUdTlsCd76
zgY72lyGq83bTMj23RHLcJi1+wvHJWZ0WIPlhCTXb7W5Lp9OegaKc7CanQ+8WvNb
djKanM0f/NAKn5R0OU+rlzzDKDsNEMCLGkdYZUNqvcZiETPDQG3mpmMUiWQuRJ7v
gfaM3TDX+TwVBnbdBDAFl4mgcCCga3i2/OGppthojCEpyvzoOt5V+pVdfdQcP++9
ryHuNtciwWaYbAHuUemwuluNSo/GI7jZiF4bKrvXijg/FfIACz3uz/kvVCt8WeMW
5DEBKjsU1/pUnZuziPJWUxLbDSyhdQBaSth6+aWeXOOM4YBb0Lc/A3BOhCq/BlLj
VRnTQcDsV3kNfmkBBChePfQDhHhcg2KcGYarpi91hNGg3mKaubp0E+YKlhUm+zAH
sywhsidpx1lL8biHsw/ankhs+itJCfwPT8UK/4xGYk80PUsQUqv3XU0gqT0riRMz
2h8cqP/zhyzlvjGAK/9l7YYpE9GYSdpx6l3kFzwlNO73QNg4GpRQkYyCDeQZgA7d
J/gDpDGNMNeFkdH8y5smIdu0j7+1lq1W0bqZjYkFz6ncxaKUyf38pPu6rKsQQkVg
jlagyX0VtPfMBX000b5EqPGgiYMAvB9nSoMd1T1dH3m/0jTlGxVkl/rBOe7bAIRb
DVgqBXIGg5sGC/AgONbQ2fKUlgex98qqfjAsyhvl4C5VUlu6LbblVJ1S2s+f1X7u
DPFof4syehEGcTnjLuXqBcjpYnJazSu3DveO00lW/DN6SKQE7uBaqkEpVGQubDi/
NuLR7U2IsOvdzdu1awKslm3pfUteeSNc5dc8qVLTIVMt/I6z86zX2x+z2Hn0ScrP
qpTV01TGRC0JXjukHIOtG8jn5zcENHBqKxT1+jj9HhYGOW74P2/HZSauHAeL5+eq
UDfri/41DHi4VNUdPI4kh0G7ipA91fP/lI8uIsm3p2NZ1KZTCRxbh7YkbCdiuepK
BQFQgjt4BLkjtDhcE+PEyw5q7VrWl+8ELpXkC07zzi2V9jctq5C/mNYF4y0jj9qO
nHCwK2WOW6poTi1GEKvvQpsHTaA3JQafLT1uH/775kaYw0So3NvrLIOHpyqdq8pT
YzJSwZkspQ+ugRf8BXhu2Kuf25oDVtCtLZVKlUQ/EbSxKnUdXWS/NoysUz3GA0Ks
0oi1s+C7zxPoXgEwidRTHJWCOhCDRFvrwEdl/enHBS12ciex0rO9TmkCtYDvZ1nS
40z9EJ1BjXHLODlUvXGdqVDxMCqYwbniCQCriLT7T8CTyUYcwvyVEtgee3dYdOeB
EgSqd2koZp2SHLkX+pBVUYcFR/zS+ijpe/8MW1v+BvKKGAacGLHj4Zz9gPD4BDVO
hRidn8yDk3pxeLPNekypc/sVZBr5SkbJfLYZGzzTDE8y47Ovz+aINlQzTc8HN9fO
pp1hklQUdj9gPTg4Bg7EJe3zJtBSiJqvvo1XEdwPSTQ1veU/OUvYwZWMR3+7fKTr
G4wLid90oQo4GZaD/mJFjJdNY+cJNrqNqcYzGSLV1y4wnTmF69ACFbcBMIdNaT2e
SgT7NtG2jqc/rHyaMxNCTypN0Xq6ayUZWWGqX4kHxKUrKA4zLoJnbZecgml6Hqi8
E4U+fP6vRk1UZtGiWaG8wF/xqVI3ZcvDsgyZwX9325R3rxX35tX6wPAUw77FJQX0
I81lA99PkS3CEVR1+DqgZzbJ10cvBdFhdDdu2eMoREPOQ6niSPs09uqpnwNpT+ER
StuQKYVCS1/BXRbbed39i6uWlpQYjeZQ/OhlDNXniiJPp15zZNIZgSmHm/XUUmpT
lMqrMA3Jhk4j2JZk23jKmKj5s/+vTgcAeCGdnYmZnqvDjmUrkKHyozs/BDTJGjGj
fVbAufeP//4HVFVyiF1awernTovz485B94BndF/e/pgzwPxn4m/oDMYBiGsMBo0e
kWkulKYhIUdbyLAsfF8zpitOH+lesU1ytgzxlZRLnhPZPX4q1IA/wp6fJGXWWV2N
E43ya1zkrC2aSp7rPsRNac3w5YQ2eanhQsqaRpOnbRw20fLHDCbwumxeiH0irECY
Rn2EdVC1PEtucCPuEXpDujZb18ScC3OJLrezFfYi7tNcBCllUdiX7lSvVSOJ3PEA
tbFeevZGNu3+fTGU9+8Z5BqiM9xu+VyXeX5J8Lsu+Ibg9wNo2qrcaAXjEx0W8/A7
wrHKWdkKmmMxP39YE0wqL6NPN4A5JT89KuoUNOXOdEPgBP8TO9XORx4l7URstbgG
Ap8rEj0tJk4QxgRMsIYtal9AoT3P/BFrxD24hE6X9FEwNCUhZ7seCfW9xXT6Vv+Z
0HHY272jXAzPS9TpkqkENpIm5CQihwGxzp80/A4vdBU=
`protect END_PROTECTED
