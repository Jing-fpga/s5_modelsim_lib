`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
swMmWryLH1iUBEkiEZJJkXpuB87YiRVu0/nUB0+d95i0BsFF4BxZdrODYRY6++e8
KpopdMdPG/E4cSOC8r6CAVBIGng6ki1hQz5tKZBPuNOsb7UXOBA0CD6I8QIJjTZp
MsZeeAYsn/8I6aytcukmtoJ35dUWgIuFCVOW5F4NScvfPKlH73JMKPzp6e6u6Qnr
W2ICLDHS4P2XcjdVG14hcbFyjyRdgaCT8q7EuCcU8si7oL2kurmu5DF+Mg4MlHWC
+g5i8qKRUebWf2c15xVU3J1zcDyV+md8rTRK7N/xZ5yEoWUcaVdEj7s575Y35TSF
87ZhxP93+3hmnYXkPkz4DhAuqxoycpE8sq3ugXWtmsKlCLkhRJdi3d1c08A4i7/L
TIg4SmCd4LLwAnfUoIg9jmSAbdlXf7XsOm60BGNSHNfOaXaNy6t2uJhgVX8+xu5H
VkJ6PGfk6+LC2lTbmS2Fufegx5Av5CTK2MI9iTETcz0ncnt1LFLJDB8hbR+jYAW8
FLLNWhxKaDHzXWqwp3WK/2h6QmiM/A8brfibWiqc3BebHWCxdK8huyZAyzPAmDdx
BEKfsfidbcL9apYchx3QLhoImBpJscxxD3AXMpS56+I47hrmHK0MOVkIUKHjl0Y+
rd09NRFSmPwrybwEwqYJimuUKWiy2wIzLXUN3Bfyeibs2bHMeo8ztJRTUWTAgXHx
NnxgS4mx8CgPddjHn8nG0EZyZmoCLUlOZU0NU1wDObk=
`protect END_PROTECTED
