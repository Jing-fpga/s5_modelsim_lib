`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j6dxKHzu0+CJaFaKj/ycQEoAnJDNaOslQSki716VfJAwbFQQOzlLfIIaDKtfkNwF
TpPnNJRDJTrid7FURpRT8wID+PRUhEKXoqSW8pzJTAgkOUU8HlrNk3meSu0uG/fD
69/2FjfGhP5pnIBRFgV75aqD2hnTZSjRHqPopch0tOWrLqEz2CrBZ8+1PHae4riS
ggieJyo0qJkojonkVU3Ly/t1kgqt60W/xPShj+SwIW4cHgXRe8qy9gqugYSPv3Q4
hS8j9v4rj5i02uO+wyPstqtNzny/FGy+pNyB0D+ukQb2qf451kpjfYDBjs5ZB7re
j4COyLFkNZ/WhMudoIfOL80h3J+6dBNllS09ey5JJ60gwXHbfp44BhoXx9LteSqu
y+Ztmz9ccWM4/f24qKsMk2B2KhPBn0KLZhQU62VegEYk8vbybmg0nNGOmCFfqDnj
Eaf4cAFk36I4tl1PZupmBiW28WhR5gUDx8uJ1H13/l1MsZGSKggWF/XK7zpuw+hD
vR2LWG0G5u3Z5gxL/E1p+KizPlq0Gq+RoL3eH06S0Wx5OAvbsq3fJzFK9zEbl8Mx
WEnRlpMMrjm2hcSsTurp97N0kz3YoCUgzkdu97AyYvUoWkc91X2OXj95aFBwe62H
inisWTEaPlLYlw9h0OvbZnIRPpF47ucTAbH6+551ecRC3I1kApQ5spGpXMBuPBA8
Do1cpLPtxPLRW2ujCrjbavS38gTqq+lUDHj6YvqImCBTH1jicQNJs7eNBwpwvEq1
db6ZxJBr1NeO6k6K0yKW0nmGkcfxvy5QeF8wjkOmV2XafruNDIoK9uUoIgmIl6YG
xQWKhcyhIUEmhMDNiMWv+8ZYXOwowCVLA0TsSXAhJSHM/Yc/krp19mh+iVLeG1dZ
/CBQ0SP4Ks32EfMnxKrUjuUbNFjMSZszCbHjRP5By8wkhbSJxYV9KkXUTdx5sWmb
1Ui4qcYOi3MhwxvzCazghXTRYJg/IxljiNgYpTJckDPWc2IyjpD+CPjPZ8I6VNkk
qAlDvS2IEfRDxyZ1BDen7RL5ZohULlZYB0rfmCvyOy1Eyvkw6zk6lNQQwrGpLpCY
5MYhd+1a5bEb4aQ566It5ENKQ1nMatQPfH8Ba1whNA4sa6czgPx5Bh+l+FEJUnA8
1oUEp6Nxi9MPl1Mq6dc2KJm4SQkElQQEP2YOe7o01FEnErBjS6GF6YSuTptgeVJX
YV1MKv/Rl6u6zI2XUtuso5hTtkZ6tmeuRzvW0dz6BVf/NYkf/DRVC4z/2bOqLfRN
uoG4+vpFSVBos67nMaQH2htGC4shTwAfI4xEjUC1aUHZUlrrsBFR0mLt9E8wbEQc
TGrRbO38qFZencjfOCWYxDbVUtKOuO51gPpxwOpw12/iRws1jwTbbuDELNBTvibe
qP1h5j9SGpGbLfOj63r1b7LIOqC81a4ouyfuV7DuDG8swtGJohPZ2XeFJ118ay8F
Ue2h4NralVQu6Lhxj3AeyC3FxgFvsLoArG9MhyLuSbLmSmYyXTwLzLakZA5MaJ8N
1NqPNUtD2tmcvWgKpacHPAYDL0xNZ3N2p/nXSePS5DTE8FO7vEgkN+/PYLkiLOV1
SQa0u4PRI/LvaHmnUnR8HQ==
`protect END_PROTECTED
