`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JaESQCfLnl5nNK3raVe2dDrgjSXzJvsqjyeYPmfBaaq9chU+oy8NX6OT97KntogM
mzEMnvKivFOI5s2gLHmYAk3uJZU6ZaEUGxYJdNHHVjGVfOGL2dpQ0LILFR80JOyy
xUlForLdbyn1erMpAN5e8B6zu5z+k9AHrl5GayMygw+dW3WJtHcxLxYdVxSBwWBE
zGtj/dyyEbXXXxZnMM6NpAHzB7fjPadjvsgSvHIiyOClHfF5aUmxcYDGHzl0+eQT
f+avQvhtmBNehAuxFVHNiXPT99esuhumO9HAigckEq/jpXFI3US3L0fQ3a3dC4fX
AWYZkwcnqMKwKpWydfXKZy2rFk6AjzQrDjyzkR5ld2wksH9YHOoyB88tGmrKaofK
Jw+qc7yIcxoJm3v2KpUIvb5LZva3e37oWzzLxyCyyeXOLcdv4rp/gv8P7xRriqZ1
91VnFKnIdhFE9m9kOV5N3bYftC82n8O9fK9sSqvgXpb7Zpr6lVVWMFWHu7BnDQ4L
PD/wt6RIJnnHIbUhHlJL01R/R/i9FHVhl1dxP8qFUoByQHZHjNjIySAk4ujeTZXI
`protect END_PROTECTED
