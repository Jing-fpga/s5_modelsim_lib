`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EUpN20B1asnYYwHazMvsTFWVDGUk4YFVVfGzbAsYcTefP382dKi7WiBly4+V2GKc
sGOEeYJ3ziuL01pG2hgUbNsPr1t82AabFec1oSKnTTsLQdBUssM25iDCnufO5Kdi
rJJPmKXactiL960ms+/j/k8HE7hEl9ZPsHZoyZAZVhF1NuFPS4o5rDiAC3W63dBE
oDioXwOJ69r4Grivgvkpm0RNCqMk6dJarBFL1FngWWRxCBDWYrhJTiQcwdmsfhfz
DuGycuh8Qtt6w4Koh0lAofsO4KoZ1U862FQRnCZrUVlFK2HpKU4YCrgk99tZoZ7r
ALebqO3jXXpmIJMwTIrwvLRqRBDV2GvNZ1kP46ogII4Qdr6RPkti/v5jeq3jo41C
/edW7awk/N+4zxYMnPPbEnMhnoPitQhhoTgMVMA6UMxXhGcx36ukAdwMNFGOeP5Y
qlVJYjGCo1g26hWyqpLSsgquxmNjoihnJK3J4/ZrVzHBvBQ7Q5Vkgs8azDmTX4pi
unDTaMtnV2f/jr/4WX1zDTaEX/Hrp2vaIv85I17zGoWd9Q0nzowdMswT2cOcHPC8
GmbCUgFnTczbPPmMep96A662Eugfm4Ase1ogsxAQFQsPcauyP8P90/vjGq5Hk/GY
HdIUqzQ7IAhhQpnC3rSws7XWV6L2rA53xgeB50/bjimefrNH0iMWOMwQ5kZqaYOX
SEp+HD6yAH90gMM38vZ7SfyZElBglIposhBkU8OLXCLavR45+QUraAV/eLQYMPQT
L/hs7fCRAcC8sKT7b6yx8m+pCbXK908glSulCimOj1xVI2DLW0qA8HWZYl8l+nDn
oz824FHPHeIVASYHzR+ypnqk6rQCjU5FKfDdqfG2aZtlFpvt9MOSUp74Qedq6to1
xgxUf30JMKmd8AUf4kbeVfrvXI8NqlKk2r+k/7MQounkEKRcovS22b5ILZ8fFmFU
MnI12iHfgqhkrSVeKNPe6iJcnIo04+C8Zpuu0MH8D+oPI7zPsFRP0LIshFO2bM2l
Qj7Rz3JIM19nuFNyzT9SyvFQcMBW2dL3+XRCFs28dBCFIlW7GxA9xXZUvrbd7Zvr
LtS0CYTwr6OQwpd1w/XE0Aqr9pyGy0w44lTHScz2Od5Ed/857sKx0ek77qjnLJjQ
7sOvHvFEdqUBXBDHb65fAM0VVYh33KxdRC66fqmCZQ0ZlKs9gQSb7m1mGtTejdB4
LuprQJKA5XEpjs/1cbaoftd7o6pkYiKPDk2jifMKcu1aTbnajcKZvSQT4yJUJh6z
c7AS2QguGO6hV5CfOxbfSBwBBmww6W0BOnVIwhJ9mR31wxG8CF0WE2aV/Hhm6Pp0
s5LJKn6gk0yuFbcsBH48lY8JdmU/Ex5cS5RuWZdRhPduKqY4tQuOwW5SDpsh19Xl
0XM5ufBi64PTk+XpRNnjdAtJZwou1sjM8taICeVSqhrmBdRmlFEP1fueBIMIWr3c
YzZ9e4bu9do2zkw/SmR4uaHLgq0cKbUVwJXjtciRcIusKKW6Vb5kv0/LoC8m6xPk
AFBFLvZXCKRrwzK+PibZ9+hY3+ckFrdt5O0B4wei+FG1av94M0yYj5rKiOYovTi3
0Vy1+pL91pT0VlSlRA4N/ijxp6Pz822xW6jil5t4NTc=
`protect END_PROTECTED
