`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vGPufV6MkI0ULMBAHRgX3UpiqC4q6wZPDLiWElzABnbQCo7NYhzXjSGHiDpD38TQ
KucvDEvQCjfE3lD5xBnj0zOh+JHHuJrReVwO59l5BK31T4w78kT/uJAvwXPcNRJc
TrO+ZIbXsmYFkudfjAZGmXI4PGwWFzGTI8+uIWoLlfVOUbXP0YLvVAAN+81NI9z1
R17Udh7OeQjhXl9BONz1jLYnBZtrxtaPW+6eWxIgQ3qcWRrMat66GI6jrBHd2KKy
qdqIMk5+5ztVQFRxWBCUkhZe0ky/G2axAq4/WTJEQOAD1fuFg2lSRvJSvUugUgpD
tGQcLXMTuFCDL9ua/cS7NIN+RJ/qj170Ojk1e75CWj4OeCm9BQC5vQd+65Jt2o16
3N6u9Iu/rmy6aHgNbGcwfNwOIh4eGAvvq9DYnIxmmYtFTfhYI+X1JKnyJs3sJCqW
FYUayAqJHfYcRgKlEKBfnhnegX2X78Lflgh90Qnwe7TDmjc0Ha1H+3R8OcfaEYZM
6PT1L8FENzPlrwhDE1Z/hplm06ee6nKz56WYQ2p4z9+hp6QkHaAJM6X8uvid+3J1
xPtUJnqxOfToJcuAnvTKC0lbmOJIAG49c1YFA8bB/0Mx/hFwsDp57A86/F9ZGx1I
tMY5eqBb9KwTacU7NWh+F9eNXL07vscTDuy9FNQql+WWKB9dY9GG+ACMMaZ7Xz7G
Sxo2HkgQh3kRVBZesVy1n0eBRS6RZdrek2jKbFZ8TKmoLJmCcvALdom/TY31+9E5
+E7IvWdcpHpdIWhkq8HSGuvTMcAYwHXrY/eTvHBH+9VSewmLdVyoLxOAqNsfK1En
SS/Qjzu60mb87oVt2XM4dq3rY3ZbwS4oh8+3rIcfINI1z+K3xu198lHUQerB2ke2
1kLEz8TRRKAj6Y5oTectJR79IVc1vvZcSN2fkPb8+uzXnfloZWdvbe5hy8SJ7UG+
nJS7qqyqodTixlIxaH4h0XSAF7O6Ip2oYzdb5IXayE56OWvKUcrHGAp7QUp6x3+5
SCihXBGkqnJ7Qr+JYfCkd7zJRUaa1hmEK/Enz9BE3QYimd5mxRBT1BgRz697cplE
iJG7nkZTu3xrrDDy8aGF5rMULVGJ6lV7qeK76Kt73ehovC0NelT18q6xehS1wkv1
ufSY9aG2CfiUcqPGeioVhkw4L4SUzU/bshGhCZYAnDKzebo1cKbYc+hIEiKqo4Dm
bzjo+846JDYRrC4Ac/cK8Ghvd8aYBpk2pG1iy4cnN3JOgBe1HsQhaoT729HBxfz4
43IBCY6zWGZ2KrSWWVnj56Jz841MfkD9FuSGC8NxiNmZzKg7wZleDnmq4TBKfx6Q
LGJfyVZz0flc7jq527Nk8/d8OtA/m3IitWinK+8VwVBkp3HadTmY/7DV59ThLosL
SGI7grvEIWp+YODEpIQo/MCuyAw0nvsscq9QULxfARu9zBIn/ooPGB3U5DmBvrsw
s4Pz5jOlYziwGCn6mQ4nV0yMIoI9TUh5OGMgDxdDc18FRP7is11d7vMOsBOHSd/W
jTv4wcxQG826ksIjwJcGzsF19q4iq11NMpIH/txZ0EAuQUFbRPVz9Vgppj3dYqFi
Mqy7+Dj9vbnxpStUVKgjsj5mw4fFfX+aPm69poA+SFB0uQwbysbh6/Cr1z7RSHq6
JflS0f7YOo3MgNr6zoL78pGx0rt9sSe5YAa/52/GIBv1sXbq4siZI3QJW7lGtrOU
yKbpxtN7+ieBR/4PRHhxzYq7ffXpIQBWoWogKr8ZTacrGn3+VVSSKBozeBT0PDMj
SK8s17gsxdSz/4vSoc3+2RXsofzR0+1jewuzHzv3YWKb/RPsXshrzHVyOHzz3cch
b/cK8UgJZzdBI9F2Ii7a7VWFQoglCSG212MbihKxJo+MGuaKFUPf7wHuNNrK8hqv
8nQ08ZyZfKthpq2KBQPxm37/fNYkzjYv13LSkerCnRM+dxc4P2i86oMbVaeArmDD
SXnbQAgX4fK+l3gwK/hQUA==
`protect END_PROTECTED
