`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XJ3w7ZsSy4KFeJ0dAr2VEERDPKe56zPcxDxnPHTYdBptw9lXHRwutPOXb5ivi5ye
jigpC8xxggeLjq+emuNKaV0BzJnBUW80jxsZZRh45/IteCQKRp90GX43DNK5QVZe
ceusCiwt3VdKK3dsTQ2btFuDypH8++OU7L5NFGmahakAmJ1OrRCJB0wIvV21QyF0
UViieocYFk3C785epvIrYBWYfJeY3zUubW4Id38q+TrirRdlcxaYkyKU3L0snYBu
Itq5gXJozY4X5o8j9+e2ThD8Zilp8ihOyNgqM1PWtvLeDpo3fw1ng3FPhIbGQ32w
99ll8Im+/b6GdpanWxC85Rr1sqTAn/k6Fc6DWeNAUavenX/tEampY+LqqQ3Z5wSw
dWqcr+oyQG75EBxgzIjA3ghq7/+IXzTH6YIBHH+7TmyfP+/5OSe+kle9raSzR6Wc
MoGyjppcXGskeQ6EXazQCQo2JgDxfxTax0QLQVocJtb1ulleXoLn61GyV/7t/Nr4
Jhy7crFGmVFmB+p2lwAhChzxaJys0S68ahi3bkNjEWeNbEGwwABp8JN3a2gVlJzi
a5nOrn7b3tPRCFuMgt8E0PtiGV4NRsVN3jgL8j5lhbn3oItKzQX+ZxK42yxZGmo+
JxLBjzkgVss315Z9aRsWJcRqEZdtA7uU9UeLrK7tU5f+pzefooZRHVWQ5tP0Fhtt
fa0GZftf8iW///qGRzwqcpVRp8fQQQ4HM6VFLzigZ3jxTf/iJ6BhYiqcflGrSXm/
TC+sxXj9ceahnEQpChu434TTUO933Of7DaHwB/6vrpQ5YB1acG8DCl18dc7gy+50
NNzLb6ypz755J1oUoAlBX4/8j98Nh1iqGoiMXTytJ9AudocLKVCwxPY4kCcdv9Yz
KkD+0O9xBGprabVn3FBm/IWX+eZ8ui+vBQfgA2x9S7A9yphMxI4LaIu1cVeyc/OA
pCkKN4faP9DFkFyIV+YvQC23lAUisISIbOm7pLx5xybK65PlZyvOKYZ1aM6zQ7Dj
EVBlZ/Trcfo4cGwKN4or3BJRM8lBaSRRKPgZTf4FonirnNu36J4L5f9YdzjMtdsh
3Nt28cVPRHWLHOXLOUj6g3xhjdk1MPzQr+7jqzXh4Ex3W8SeQCnRLxefDB68U58x
mefDjQKH68bFfkSxJvsryM2uNtzPHBf/52fWCuVRIHN+nOmOuXIkwY5i8b+0PRLG
PAA4UDgRG4tf29OO5WxPz9750DSG4nnYpDGcZzXfkzXRbelbCKFqcv2SOGlPyOzG
WiaXIbjXeEiZ29n9c4L4Gw==
`protect END_PROTECTED
