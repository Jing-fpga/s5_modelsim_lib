`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8vF+8/B+HhPNM8vz+1JA29++TRam3DWWaXq3d5q6ssLUFpd2YuZcoQ+Cmvnx0yaF
2Ett+rQK3IdQFmddUJRoQiTQjRnF9sOJujaIXAK/3JZYBylAwL2KN/DnAaVFJxjg
QjcQ2Mmpqh2gf3RSJBORlUb9ClOMyXk4cnXHrL13+0QIs+YwSTSsyCQizpQes0+P
PqzOhAtNBbsjCG2p0Ao84rngimTX3t9YIqYMi/sKP5HoU4RYI3S30gb3Za3znCh4
WpHq62jHm0kbrxlQzmJQTMJs3j3ipY/cvZ6MyeNzkf6ClL8epR3KfX56W5zHFuj4
IW2F6Yfkm/hEM+fT1LEv9AX5TAUSleW4UlDcgFek1h18OVYji5ZUe7OvNqqeIhcd
uYafl8Cu8qps02s4NRTsGmoPg5tamJp7pXaYlV18LtdG91bQp1Ef1eVE2feHOsgq
/cfx9luSDeEfUNj4CqVjEM0jYv35Kw+1ncw/+BQ9wNiytqMwrLtjyE3OikFPbMLF
ayteK8VylHNOMTbeiWuSpDijRpKn12Wfc2BM+Orof41QtRPmCmEwVcDv+C9orWor
WlJE5Kwfx22xIuHnB2bwAtescrsgDsQq5KpBvRKddekM9ImFSlbkCoYm+9UcVvOh
k2F4Yd3kE3/xPC2GtixcVVOp6l/TZV49aDwOoPJU5xNm+JS8OL12z45pN1x4WpUP
DfRW/mbY2tiUgjofVEuwzsq0cJmEstnxrAEW9hRzImgCWqfXiFFrprnZpvaGoea/
idA3NHeizqXdCddUVf7kDe1JhNkZQGKVeERPQCjxPCeFCoY7Ky/6mU942KO3zReI
dBuR6kltR/nPdFWOYTby43RM42SS8DwkYwtD1HFngg7MTfP1LzYYBrF9aa1nNllR
9pUeKiuMzelhRUmcGug9bJi0OniZuEMj4CnbKiyAT1UQttO2UIblj3U8Y/7m8BtZ
HWe0VI0i9IacjrTyti6Dd9Mh9FaB5Xp3o2u0m5mlnTjqysq7IoZurkmrCYw7LKXS
yjyg27T6XREufPyOhtv9t5YbjTt0/g8ns4MWWJRIvoBI1gEd9n49CpcJwHlG4yaO
Dk1oN9XKCP8nskJPu2KeMiZLwkoDo3BUprs/rem53g4Cp6Fdy05BUZKWYqFuKRWB
dOYnXTx6pBEPJUVlGeVaUYVpcHAREwrU+kTqzsm/8UN3mx8S/Fdsc/La/et/8SxT
va9QAjpxYI/Nrwu04XQNAW3dF1mdQs/YiPcb1STC5RuNlRu5ezV3yX/exLDHXslh
Nde4ZN9UCxHek2uY1fh29WhqMXnU/kgndq07SL9Bnol8WUGNjOYiFXxStWFRvXly
hB58C0+3M9j3aI+8OE1QR6AF28mIZddSbxSQeBhZqsoY/ledG8B8d8zXkd55hTC8
cobCqVIIBVgWfdvVNz0X1vCgqSSEUiiCyxp32JgSjQbdIDsFLk0sWfu/8gZZWZ8P
MmsOwm++6MPYj/uvQIdRxd9pYvAS+XsiC2D0fkc0Qv+hkHnJ0sBihmeaQLPgj4aF
iqOy+ppkSIdP33SwqIZAanxkGPP+86LPtiNjCMb/lxHuMnGj2V1qMfI9B7azUhaj
nQCT1d/vHK4kUVs7UKj8s1Tk49YehYF+IAUqaRVNXhuzOMwiRaVxJLTnEf+5R3aO
/via3cZaKOeVkEAj/pBHp1JGVuYHh2EI438rtZDlQU5Ofzj2FvJa5UVNoLE7vI0K
DXC4xZVrTk6TjE9pbABf/Pw7bUx04gXlJGqfcDSRQs1UPyPSAUoFcIpcMr53nMa5
oubEgegEsLK0ZyvMuNGgwV5mgI+KGXJTKn5C/0XAXy1PXqGgNFT8twWKpVGQTc9E
QyHpR/Dgk+HBnjDkw6SpxaFA7AWpXVDX9zbHlTJIqX78pcE/nAF41O5HxWuHBTnZ
vbSZlIZS+lhWJL6TYKbDtd37JtUUMYlhQG9hiepNBWhegFbVXEthBddh+WC1f6tH
ulAnq+0Mb03YChNdL83PWFt9Y5cPu433g6mplnLko7lZkcw3Z3SJzWpQt1i4WSHT
X1EKq2jIfZq4ROaXjvthe/aj7+LIklAc9sA6dvTcM6il4g/8vPEVHVLTzQxo3+Ni
huJxktHbT7USlYTPu2AfZDBm7+jLkmouvB5By7R6hvHZIitQNgMmQ3brvUmPWUe1
rcrQNsfpupSvZVpvYSQyozzlMCb3C7j/spRxgeDagEIMCOVto9+bZ8q3TLNatNqt
HjoDSGMjuw+RQM7Lrr4GcJqwAXGpJj0IseBGqNML35fQzqZB2cXR4ECrrzhoYnzc
OIdI63UasfPjvgZr9kuTTaEu2cRsK5wTbqAqtqu+LOqFrhGES5waHDMiUVSklMlU
Kk7+ojMQ/WWFWEL+lC4Filkl/UbVBNpjJZaKK2y6P29PC2inqFRpCwE7iq2KVHOr
IaYXo/m9W6/Sndr48joseunF4wp5oBDqKRlUsxJ08jKplJc9Q7OTLrgZL4513/n/
hsnUiBZWXz1I9tdJQ+IN/4QM+ms6WoURmYSxYaehHZ2QbyPJG7MWC8jBMrKbHy9C
Fv+YMPD2VbHgqUy+uN//Tg1wMj5y60BDtH1hwbjb14H1c2wAj+6ZjL5igClY7VUj
N4eOYTmSedL7v1O96G1tHpxIVGjJAhr/NztlF8HHnY+7fdWI5xQhE4B6exxEbbH3
BAHUNQBxYauDx0DUkN9jSQ==
`protect END_PROTECTED
