`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v0nAyPkFPxLFXazL0DkazCJlVW865MFlOvpxJE7ivK2wPPrkMeBeN9PQgF7JrKDI
99wsd0QKkz2FGlZkQmsOnlXOx00coaMLGvYCBLUKR3IW9flFmdn5GHH4AbIW3/MQ
oLAX2UjiR9yYG/9NpyaZB/JYV2ELBS0Q30zR/NkDHhTRUOqhGdfvH+O2JguV4kl+
zsh4XCh6MywHwJ4DdEnfNPO9XUc1lSvHw2IUk6fExTYi8q59+P2vD0Vu6Jdh8eXV
u2Um+yLV+QNXIdEpJHyNN6xd8GAeR0Heq5GAgpoLuqriRHTTgqpRW2qDUfpaQoOp
IaX/WG/B/If9QoZsq7mwWS5Pn8QeFpQ1gRQIwtI2qxiVBGbRbx1IKqXS4T5PVMa8
1EVUqvLh/YMKZYJlO3Mmkh0DJhV/VIixdSStMvLeKRoc5rHkOEFRruG5iHF3qXv1
IBLiqhi6Wdi0sMMo8lYOGiLTmnuPVaK8RjqlkvYfXhlizKBQKLxYnPs80d45ZHMq
PplKdTiJQxfGzq3ZJujo07dKkOCFlLisEVqywcrvUYEmW43oxnKrvWr8K4SJRw+C
I44YrbFUvoPXrYcFZ6suB0CtUjAnPuCmkx1wiE2oPGlFwFLdRTG8skM1Q6HzT4DE
UGlny+028YiHTnNnsjNpY7yBHC8Z89N7K5OrJfFYYDwHanIZmh53IAM5zFRgY+Kj
n87DY7heOEVD0nDLYaNLBISaJF3I62Kgzsc+R0pXzQ84a6FWTTxLh0sZ9rECAtM/
xuyN0Mpn9/u6mJ2xm/7nu285xRrrSh1YsQsn3iXU4bXHIsrPIXMbfhfyARYtmBgw
H7GrWakdXlJYhpLjhL1H8M4In0YoE8vYKp+lOYENa2hDyoa9uWrJF7xeDY1v4UpC
CaVsM3vlDwsTI0djELmMUvOp7+VESBoJcK1wrGKb4BxrLkaT1EdlLJnaSCSk7tPr
BViIh+j2FHQJgF7h4z30MHLZGW5OhGt3Zg5ZPdOBQBQ=
`protect END_PROTECTED
