`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MA7DVKXeCeDL9k5PI52d5vg5lghp0maVUKWsqQdpEvKwY7AzNFFJOKCJaABgq1eJ
4K1vC5t/ByXR3nJpbiuyO47+3YEzJhq767iXjCpnUhiRlDebhkn9wgcZgzScR5x9
3bAq/GJxiKQVz3Ui2h64pAwO+9rtVuupHjBvfJcsTzjpQsOShbqX+t/6kTQomdrr
XDlNR4KWyPwKKZCbDDuYbGgD2J72A0Gkyp6+KHx0WlqKKD9ufsV3nMmrxTiQFUml
hzHUMcJPpP97nRZ0hudTQqIZDZETDkMDFYA98UKl4b6UdpxhX30d+fyjruBjR0bZ
rP+PKcIdMmEAf8fz/01ujH51RV+eKOlx3wGXh4Zz8z20cGvnOj/xX6x+JdSQ7g+A
kK6GcRzsT5dVTOL3v28zA02G/KHjDZTX9P3q9d+V9fElwWWB2hv4IE2y2HKGsSyb
EvlTj13pfI1sbO/XJ1S4tc0aWAK1Ti0av7wqUU01HRmWoSWZm8NBbcIjc/D0XyAq
0nUiiWskpAPTkk0I22t5/H+yVvqTDCsIcdES2VDSIXBH6/9LqYl7AVUQqzg9Hq3c
MkhFRxXwSYwwflzhDJP0Vne1fcyo05Hk0nP+mKEuEVinzOQtVfZn4a0EnNJCfKi0
MX2dTJf8V0gv3qlXwbSIsGM23Mzl7l0W4MxYnGsihxT/FdoUlc2X8Sc4Qego2Lfr
dQGqhIyCV04yXekIskbzN/iREKwtW7GAb1Xlydec7YVxascl6nszKZ+7adjFwAs9
W6dZu2zNIPRFDf1V7pPLFgyijEy9ZMJAJAeqMC76iVa2SYbiAmUOPZY29ihKrc3X
NfiguXi/5yE0Mo42XtQp25HU1JFEA2dNil1gAK5pkbF5DVU4I4AlWaJ0QpiOZxnR
+LDZOVnVG13LJxAlXd3BmGGEpY8y25qNBSpRVSksBgLMH2jiiLVvw1bu3BzeRlCf
qqqELg4zKCAgM+JDsYDMuIiESB66HJN9hS1dIa8mfUOwVsdJdOezHCccKpaqtgvC
P+uCcX1+dZnjE+kgwwb5DZpH3FrFjA88REvSfQAiuNAZ3VWL/HXw/fOO3mrf2qA0
`protect END_PROTECTED
