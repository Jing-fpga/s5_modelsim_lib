`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u8WtIbWh7j9txbufc3pjjfnzNhPMsRJEbvgq7PajuFxuz1eAnqj93EH2fQ8OiDZ2
ZT4/DiODvmCwNEYqugrkLcajyzfXC0NOvxquAhnSbtXuNA1Tb5XCAqJs167+1NU8
luXLor0Zur3QLzj/oZsCoPD/DhbvUIvW8O612s5APmOW67ilJzb3rUCjY0q37dJQ
dZOtofjcZkIIRPivQTgB0sgy7uBJEwyL20MmttnYJLkYdPclhCYNo3QTXfgoLlYF
LT5TswGPsjHsnArVSBgRoGRrhbxe3WMvt/59qNHKmEtSXSVx4HH0hu2bM2njWZXv
JVJrh/ti+fG2zsoU4c5SElOfnm4FoYYbkjrppcR7d7rHvMVM3Ddt3o7tsbLsiKPg
6/sVELldIAzxIV/tOwOw+3vooqvmV7Jn/zSeFsdEQiidLTKn4V7H/hFqYkFb7HQl
aaUDkkjLfw01Ou2G3M0dJbTc8mTFYgW04LeNQubLBajc6bEF+uneSYJ4ieJunoLt
JaWmMUfHP3F8JIeT9cmzFbkl/Sy0QU0eP8suREJyGqAxScSy0WYLaiL3YN/G9nyH
A+nqu3t5DtRfA/0ktiw+FkRseo+1Pol8hLvTe9shFS0vcT5NPU+6XUAbvtFyrKC8
7x9u7p+IFojLFjr7/I4HaKBBd6pf1dw04cr8Wlve5bWRnxA1ZvDL2B5CF3lg+kxq
K6HmIncDkwI6u0uxU126+KcV157xhluoptAmlorJHVICRFVV+BaswlmGcdLekcjL
uVWHGyWSo/X67Xn7CQz0htpzUblyXR5szBKnkmE4q+enOUgxlBT5rXkPsADFzry+
DCQFVWLB5QHEC1cUmR3GhhzGr5Xd43MtMlbv4ZWEwLpScV6aCg9A0tPm/ldGllNx
avD8zPj41KgkQMIR1lqQVr0qeMh36aYuUNnNvWUumzUwnys7Y0h4VWABHUiSVfGN
kdEuYHXpYWZgHWq3jpHAbkbjwgkAhjhgPPTQeE1udZrWoP6nWI05MH9luc6Lu2R5
gylce8yZoXo+KEfo4EkS4xE0WsPhs9NI93KamSHobWdNC4X5/WLolDhosA38QF+M
8pJl9B2z1mD1QcXaUan8xoThLx2lBQNTBr6HenRIL2ht/tmjT565z/rx0LEL2n4K
vXp+ip4KYBrUddVfwVoMS1AIxdhvp5NAvHRy8elzujI9zQQF/kbEIS9foF+qxbbc
GXDHP4bk7vrQA3rCQ2QJnY+QDzdq2FnJasnpcSABuEqbfd4p1MfM0Ap7UzntIwV5
QkJYrVBAslVMPEfckymMk0HRpZQOs6H3yEPUJ9MkeJzzm5DlbnhgezfuS7phS25F
EIezpXn/pCHd3Ed9rk6fo+A6yADyEGIyImmjKZeAOXdGScKUmBZ67FmT6fwIC8Ax
MpGT7cSRADmkEs7KA/sXq3iruQ+/h5oqWeqxxRXmnZ9pommrFmJ+7GuIzQ/chNfy
8MI+wEzTQhhvV0y1/xPDtDcW066odLjQLFELTjYPMrq29ojDabGie3sh9/WW/Y3v
SKiFI6WLkmL4KCah6wBs4CFJ91eL9oMdhwbj1Jp2FI7Pa6uND4oyKPGFVUw34vmr
bLVLlecfNVdLRZzG7i+F7Uca2K7b1SvvSPPD9A8zeGmvFwPR2jnJ1jQRKU0TQj/F
VHUFdlt49OfBizdjAJYZYY1+gDU6F9EFoRU2/E6zV2Nm3XVrZYjo5+uAp7N35+MS
ArXCWyLROy9YraQGmzp4eRJUVju+P2Pp/iW/wAuwyPEss9i5sTfOzoKS1dK5zHHp
/a2HeOUaUL4e0NOe2yVlyEOdqk1C65ds2DH2bsp94PUDj2OjJnQzDGFOA7WvlZxg
YhhsBvrq4gpaiOJ87wNrO9OYjUb+k5RwiYmEXlC4vKphe6MYya5q/49P/MONktN/
C0LHHIOrUesC6tsp5NNzdtAcQlqP+7yB4mzbw71F5mrTDHb+5JF9cHa/bLy53UfA
4+hKyoT5skHU+QVK4bRI3IjOzWUGlGh6I9CK0vx95L2/PLghXUfdGCPeQJFBl4cu
We3Mb2FcqFRKVPmuDyr5r5Lt1TmQzEdP6Aa8ezy/98KTTh/aBpQmKxF+46wX0IFV
pqwYvmRb/Dq+kKaE7ct8JXN8nEucIuU/j/vz33dUNVdolplkx56gSOSwQJQU8rA9
vgDA06WAJk5E5RFWrLnZueNllsc2q6vxrde77efWW1EuaDfJ1Wb9ItoJnTznQ2jB
5elFjQIQtYTesWSe8ROxjqHhmFgUsEthGm2e4PJIOD4QwYdSv/5uzqhUgMN5YLlu
62gTUhavnE4OAC4YghxlP67xlCFAIM4yPYZyVs7ZvHB1pKzK6rAYB5Shovg9qHNj
dEjboe3SLGdJt+8PkYk8YjsUiijIpZiyNjgblaY0jcB4xGDYKeuRvibL7U9QDxu4
R+zD55BxUfQzMvj704UQsaud1r7TDwoJOG2iympKg3F/sn4hEQu7t3sjk9ml1om7
Iyb8Z1g1IBWxjhl17TGjlzd2Whkz23bz2U1A0NIRc5dGuYbCQ5+x4tY8Vr5i62gU
0wZSBFw4BMAc821IrXZ8m8UxBkr/vTsui1V6DEPkGSn09uF5h3I5JDD2tFMb0+eB
WPGfBiFwnSD1ZvSA2FTdso3Kt+uTqzh05fYvXVKar5i9jbQaASV748vTDjIqOJky
wffs+lr1xPXGqPTe2JIQxGxe4ev90OPZQ3SudBmhLCA0h1WeuB8pRXCPU7DPxhA9
Xn6x6Qk+DudEoZd44I59/Aeds9TiZDxQktbXJQp8fpgrQk4DO+AMN6nklKQIIrV3
Rtg015ebdQMfSZksBVyMBsn3P4KD4/H0+U6010wfh9hcFVfF8ATf8M2ukVnPc3bC
nKTA9HdKN7ZU7YM/Jfxa+RkZujxe7vb4dNSVJ+H8XLfm5KWVIqyHwPkeGuzOZsO1
SRN8FeR3bB15ecuyZntl44mL1jsq8NAyfIzbT9SIcAAzi9XkG9bfkkITeZQQTLzf
E269CdhwBSVVmVAAvJndb3UgjLatFSauypX0qi4dmywJKF+TaT5pvudIrggCKX/9
0F0xydETDzi8B3K0oMxp/JXofTnn2hrqxVkPnd9uO6j19D4kseKDLQtsJ6A+Oicr
9tbQxj3hLUbnWVNszwHPK2lO/+HEhSiJH8yo1bNr1Bp+3D647tE3jePZVVcjWa8K
vwXINxo3Yt290adQU2l9hCIyraPh0UII/WzTyqSazDMxOURoqtdsFSGcRlqTSVDW
0oA0Bm0gQXT94wzCcTDRgCChn2yMDcx2x4/3GhibC32Ug0GFDUqjitC5XrsgtXfb
PPt8/p39ZOhhir/8J5zpfG+HdbL1NdMupMg+lDxg2rCCFmRZ0HsUmANROF2x7crL
osz3/H4hkz9q/ckVm+KcYoXoJ91o1mZ65oLQrq5v6tRE5E9lBsyYdDUjgUJZD2AP
noejmto/sDrBVSiGCbqsxJfpTxnH19UqckgwHYH+rQlYe4HepYBXnv/gTnLhpuvr
X+/dMNXNt+nbLX4JnqgnDg/PDQIZzwUTj2aJ3jqNQUhxN9VCtGkb0b5Gvt+4PMZk
CSLBmyLHPIzgx6KZhXoZUMHw6+ySsJ+Z6WlXdv0pbs8JSqcx+PlNFdUtlB+EwcPj
Sh5b+qEzu8bLd3cq6OiePevEPWPRmhYRTD5B/Dw8DbtORzF3O6+zR03uM/5ubs0g
zIAY4uGbgjVAEMqBX+OCm0BUSUU3kCq5byHW+5elqLQamFnmN+C/N0I/9PZRdnfo
LtdmRHicJB5m0sFQVyIp6ayoYacnQZXcVxfmEZvfWbmjglGUejFg1TDk90JAuFjp
ctGz+CkWuzEA4Q4/oKw9Q2Foy0bvu4/yg67e5D/U+6vDSu5QbISu8Bd+zfZ80C7t
GgLFogQ1j3coVIQrSUnMpt3akJcTEFsTqVY9bOp8BdVp09JIB/9ndXXFyAx7XOaD
MB0sG1qW5wdPqTs/IhaNTrcMLb27Wn+akYFMu6eT9T5Ux6mNqGRfxwaZUvavne9Q
bT/hs3+nYKAjmVpWXf6M2wgY0hvnOTmszSj7jeRiSYhUjR4Qg2/4IFM1/iSBcZsi
yO8CNbQZedwv1mJ+zqjGiy+syvXYVN/R6SbCk16AS8P+dj+JgciR85aqoLxcng8q
f9WYcORQiQFn9233JCIqXb4awatsT8+H2sxCGlBXXEgMXibefdy29fKCraePo5xx
/2uRQga6yhyey8AtW5/9pXjRD+ODoMyhS1ZGwD+1RQiGQ8Qvrz4cGlJnlsNdm5rn
U+bH6N7Nn06ieHc4EVRbGYPBeKr1zcpRpEA+IaXTejBKHOICixaLSFl2oRzBgCYA
YJkR1wO6UKRzA/pNLhONT44LNFy2+GrUtZ27XRT3tyQqfYAypzJKkHuvZMZacSlU
6est26Euvq8cwJ3QkpXVKUAHkvfmhNUo6oWhrfsMbetd4hmLYB4huYYOWfDf/sXv
Dj/ZOeRHjB0yQjaS2cET1ggV69ydRotpkTIrcY2LJ3GXmvHWYEi6PHRhipNfKrVH
3Xt9kOaNdQFxRjCjDTKLrIssUN9DwpWzKr4kpir1hTLbazoonu7oS+n/Q7jHBOVB
tVxl/hMZAb41dagDZDHVDkDz/ZymoeCH8gl0IzfYPdRADMwcVyVSYy3hUrQUfN32
tcs9SX8N2tQu+z6zrf8VZi6BI+Pv3vE5Jqrmq8tchAm/Z4qaPCeIRkySHurahjLk
5RUXE3V+bIuSFXTDyYJpvGUICFNr+uPBL/TqlmBDW6FVNCN2hYmRbLRvj5mpaSY5
xJyN/7DanYdHpL2/LSwOHxmir3WjhX+G7YKasDX8Fgk68UfRs0t1+lIdQ6yBIEbk
Lv9T+J72l86bNJGCSXQvA/8ozwJmmtb3SyZrGetzOO03ij5Kfb0NZn4usXL5DrbV
JTVqkT7/20lIqLrs13IwyVq12iO7hCwBi7elWcCsmdzKHfbYBRVFHL9JFUV5yTU1
uy+Ss+rM6WLodAb4tW4BSJ4KHMvf+oilh0d2xRvrJrbi3fhs9RyTvBXStt+mASd7
LXWNPyHm20JNhG40HZC74JbrzH8WNcsIPtMjUMG08Qq48SLUCmXqAIHu2mIt4htq
Dt1Fj2z1iKNwCw7OsS4pjHQ/l0Ea/lcUseJMn4qbXe3MY2mVutdgoHepBrj6G9Wk
MSyXR7R3mfVxihBA+LO9YO5GhXHN8nJXRCbRRbCD69E2hcI9gnA8Fj+449npw4PZ
gnyKkKyUcOzCYP0gwdllVKCSJSS59SWSpJhR9tq+GSeWkhlLu4JV0fDDOpy7btSd
4hz15/qBS8t20ILzmOR/OOndQVqHska1yxUhzqEY1QjObWZYTPdEAsaEELYp9hdV
HkJAL0dOwQuXK6xdOi9ueYRFD8M2w7CEqJh6zizSvCWBMm1O5IJLrenAqQ2Md2jT
8/iH+ZlfM/l7AxJNUdSwQmVDWxMrRW88Ma60pUaLEftE0/uKBPhTtMEPgxv4kw3N
lZ/bsmqEcuIjHm7RNnvydF61cyNKFlxHIH8HfLr19E6QtIceEGJh+UOahfabqHPH
rjsatK7tWdYtmTPHuF4oYP2yj+eQA+Qr1oIBNj5jQFjQdo2/oS8YHWdbpD/LQP3z
hn02cSCA1KTxOaSt6vZUkB/ABTNmXlj3iJCVVmKnF+hsvhy4QvKIrNw1ZRfc65y3
SvDNY+saYRq4XyZXjysTzp018zAow9R3Ck5JSQA4qaITQkXWqdUF01L+GrIoFPs0
JGRXoB+ffuQYOJuGr6mknYw00sd4Htg5U+AIruEzxQUezGhY5NNWTTNYfC+M6eyh
jByDVAsr3nTEtidiBjpMWvaZ85O5RXMLeuUmeZg7POztxAROwXeUyFqi69jk7F3j
ZunHY5HypX2MqpxgIgTjKYPjF0CIt6cl2e8PrCowr7u3v0h/+6vD7pC2Tn3wIFTC
U3vRMZN1C81Hc9NYayUQs2jvxFNwUaNrfXDvqTpB+m7HoPa5weuaxij9t5ouvtN+
bMk/ldX+T2aVoSbRGTfhWTsFxD3dDzfcdeTSMSWv+0XpnkWiC4uTZMvbIfDIuQQn
qV0tIagfsSg4yA+n6yOheIikbHBpX65Tx6FtUW/UVF6s56SgCFviWNXAhvTyLVBf
BrMwHka0rxeOcBBqA6YRAvq7/sd/RsXGNjsLVumk+TK5BcPSBD+VqfnJdPWUM8Li
Vm4Nhum/AtMdzZOJRpY2o9Z38T9q0gBP5FIhm6VqyHACHyG+imVclAti2qUYWErr
xuR5Zd8qfqr3ohqaxQ5e7ZEuQmKW4rtafpR4tu4Q2oFLhQkPPX4N86P7HUzDtMIu
Ln2dlzohybfXrvz/MAzeVFs5u1siS079bFMixpkceHjTEm/AemxquCX8Z9Vb5iF/
FGERLhT6HGBhrf8RSNvuLzuvZVMtkohw4gfdOkZavxm/0ZhsD/WlTWpJ9EWPZUZG
5w7KHMG+qZs/lRr2oanqw0Pt24G9ySlSXUPT44CU1n7tTqCyX2EIq+4sPlttU/Lv
22LNyeT2E3WvQBUDEz6QnPzcZPYYP0gw/UAizlhtPXVquJB8XeH51hJlaQSRam0N
SrCFH5/QSs28kD7z56l1cy5KSwrGoGoZj6lgUHQhNp/6R6fo9wyjd3N5XRlzQdGz
J5f/KOQJ9UlkJgfLKlO6LGCPc8EG0N4Qw1SfKhA94sWEMDuPR5Ebmc5wS+s/Gl4t
V/2ZXXzr8/hrGMzBNuGXyLY8rAZTMonZ8ObWp+stpXi815n2uWh47dFVRYJOcusP
2w8CLkLZag6Mg/isWsENT/SNMpcPJRXh+lbBtTgEnPrJXV+mNQzsc1jjxBOPp9G5
cC1pM9UO/Leu2N2fL4LuvvJxlTEebqoAhF11mAx7Gq4001MYNElHDfnZa+9+IR/8
dh4mgUX2pCl7glXvvCg2VxLcbdXn/vXBlIX9OEqjipIFQo8IYosmldxqnXSKl8yY
tb4EQGGwFM4xZlkIyr6RhbyVmls/3x3ZfM2Ue3NFbUpRU5IRj3W6B5hK/otLk/jI
cPAN4rwcB3yomEVm4VjSF5YW+VJNTl5WQhGx/F/OadYXkSJCxbhmBMJr02E95tF2
lVZkS4c3KoCDPsEiwbzwgpvKiJF+tn23M0uRhoUw9VpYM/w5E0U4qguqEiDdyQ51
v/b9Rs8nDA6h4LP7SNJmAA1bm8wi2KUZBZX2iWM5FB26pEmNi0GL4rUHWjVbOGPt
RE57FUlt0lUmeaN3dQ+e5HplOYaIh5LmLMVL9FMS/qe7Uh250ycIek2ULXXS/R9c
WPgOEL5+70Ftoe7y/AZr/40pRty5LP9MT7THLCp2U74Bu007oOLJs+t5joyXCjqo
jvbihnTdvQ7DxHlMtBnrdD1BAiIyVyLWhrl5Ejqx57XOJqOpzATEn/cmuxzho7Oa
mM1w5oMWblu1Tioeki18S4naDRAemmbq65K99qhlBtYadx0Kg0PkxusdZtcs5+wb
4Odhsxopkh4YIuGxzh3ly8XP4RX0e8HH8k6cDHlKKku6gXFbsKImlKAqxgbXfvhf
26GgCq8JsoF6VhU1IuxfvbowkX8EBxwAbLHQ4KtN0GPBno/SfJsiPccaqmklI+G0
c1oz6ljt4999XQ6XW6+5B0kOghOR08Z6vVtqd7JH/MG4LaZjIqjdYUbgSPWQd5w4
hkZHw+p+pyz0xVtyDzDt4dNiSQVtSJiLcO3P9BUsdHHwHyPvJtEgFIGBcxxCxItG
hRXr5RhWq3aKdM6+mhT6uQqyaTRs3J4MnU6qiCPPaZ8FkvQuO+/sIFgb6Gvpmdn4
So73ZUap6AL31NVyBfov8p3E5Gun7XKyO4xamUpDtUgbbb8F4XuInXSMVsxxGIco
+tj+vb+EsLZftij30AtMVs5VYKFMoOn8G8NmmaR3zDYk4LIKeC907a+++V4dV3lV
RosskgLxfEHAkvUkJV5hHwTGEF23ZQkU8TZZSrp3l3a1Q/80J1WebZWJ16tDgrfd
1s9mwfRB67rwD6kqcx4bJci/wL7NPjg037hXVi1ntyOrbUeOv1xPANyJULA6UFxT
ZyzJvPzGsIXRa5IOF377e9GKsZ0BvDJ+Rngoo6q0TFv5oqfsrRT8ewwAgAQFjUMd
3+gIm6SYDjF8IZpibzR3wl0de3ZK8BWmwgiuS9v7YoFZuz9JN0pGwXXAMC4RuKoa
wT/rpoUqdfAsnlfL+7p/e0uNjxgdphvGGakbqTFUooVjM1JW3lHAqUktDippoV/i
zrXAs3B5jXvG72IKNdaYlv3RaWa8grs8VFHKs6a6V2gkwmOpQ3/SHJu615OpqhDN
RbKj2pELDJpwAsTZDy4IguXcdcYBpY9I0GjyztLf+80BEm7sfceCjUQ2gyskS6Wj
fwHF60+lVdgDwnYkCuEl8PQ4l5XiMwfJVqm5/RDXGGwBMMaJE4wi53PoCCV1kMhY
A2gJMlGCRwcTqQrR01lTAzQGFEe7VKbVwoLHXTdZ5kms7rxWcbVnU6j1qKnJrIEf
vPCUK/MTOlFIZmGG7uuBjimBLcCB5/irIUNnM2iUn3KXRWqBewFdq0dtDSy2gyjk
L18mLJMVsbwXzKQ/x4bFN1FCW4QETelJ3ojqwPT1Rgrmkh/Pwr0LWHxW7mMOOTuF
USDPpfj3fRgTIEywtcE9AljQX7LlwRDTYPV+LspFAnm3J4kZJFtAnn7G+rZpUhsG
jn6ByhWu7ts5z8SArIukHvkt/MsTCYt8AJoN72A18SWCD9Jj9cFwmZHyp9CTq/lw
yjneD7bwI2jvtmbzHhCK5MoqAQmSkDylizbvtm7PjexeE9BPjUo7eX+c+bvXBJjY
JshtZpPcfgnC2bNGHOlwC2pDnOaShHXwKLJZcnvtOsWbUZUfxf2RBUhaLgZv2NjA
+0I3j/adFV+y+qnluXNaYWpLxItDajtrV+/G0F69y3lA3s6ZdOMnc6oyQZDCpZ3H
HtS95UqKzk5Ygccq2zj4ZT+gOBsokGbuB0AdfP0IeMAZnFPUfhnm8M5EQrSz2Q6O
IZ5dZvuyTZOgP6G5ouKzYG5LzGDTSuDEgOep/IS3UsnOzNv7rz0DWs43BosPZVFr
407eZVFLFsObjue7YuNkwHbNCNLWgmULpFmMuIENCtrd5E2O9E+NdT6waSZBXPNH
R/I6ymQC3y0c1XY/qg+dvdQtfTcMUe4aTF1CtUrFU9uV3eJiNl/EkYsLl/RhNmpN
JM3LcNBxDN91ItbZ6rZTvaS4XofQpZQk0m0+FUV+rJnedRTkQW8BluV8b05buMU6
OHgPtcnSGyaco60Lgi/Fg0xsiy2ER3cKMVqOt8jQVPPvJ9pvelnnJW5PvAvcZD+m
tFs0uyWFJXo7bXjZbVW8rPmZTNTjO9IdhBPRG4WmNpXF/EX41bo3xPoZ9VeVc+dC
njTLwgp5OmUibeBxQ49c2R/Wbwq6CLx/PWREnlC7p6nRxZqkJH/LLv7ovx1hrfZC
`protect END_PROTECTED
