`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yax0aqylCW33SBWl8nGoy+U8E0c90grIBrPVxsOC5hMtF8Y7MiJ7wTRRDJE10PTx
wNCCsPf/vYQYs/rgsMjFOXNgvcecLhNwRm5sgP3ZER731sf2FqSaGUwAWAL02VCc
2VW1fplZafdaV7gTi45H4acfFc6baImY9eWnCJGd7JRG/ykgdTUMSVGsSH6XFjRt
s6EWf8rHmP7cVsWyjmZv/rIx6aZdFSX8PSa4hz28t+jF/Yr/eMteecmVBbwSt5HS
FvUdoPv4yhERXTinRXfvVKJs+xjo9rFQfeP7dkdp6VhYOhjwEfPbET8vbLwEKUBa
XE4HEbONNqgToxprOceUXoI1WCjX/9kwf7WCCXa/SSv7JfBFrKwGy8GqXPc3xPhe
lczQwt7c5txcRLg4/qjgTAZOf9tsu1vHdQObk/0Mmj74VXcSEskKtzeNDjV9862m
MmgLOPd6znSho5Nt0lrrsurdeZOQY22LUfVasFjPInt59s9dHiqHGM/CcI0b+fmQ
O2BKfJ30lCRkiryTP7x7dJAJ+bp/aVSn1yw4f8p552LwfFC6yyo1j6fN91Ve5qIv
ItrCBpA8clKFlHPBQln+Q9VlvieyYPd6KW3AIevZtn9fN0koU6MeWjMP2r0MdQ+9
juvh0oNCZXLkZULyFqDp9t9VLVvSu4mh1gPhIXIvKpKX83UghG4BlOF2gvLeUJIC
Gl0rzBh1Fjt1ReaGN9OXNow2WYMUnYWmZeQLT+V6Xv9pELZhl+ZaYZDSS8YN+irH
nteg2vkvSbmBNeuQHXIPMiQI+xbrL7TGnWHozA4etF8ePuBNt3Vtx4D7tHloslBt
Z/+LrLF58wDBnppu0iB8JuzYik34e7sHuz2Z1d3ZaQoGE4wARRQVF6QxQ7krxuoq
/1Hn9E+nf6jPfqEsAht+Ags/wLhJoCt+hDnAF1YsJZLBuH80CfIckAkq71luHOVR
l0XJickDlAiriiwPVMyPyMZrs/b51IXfPSHHNWh2zn/cdwu3D7HcOw5XOvJ2Lmmb
LyvRYe5a22hNwTHk3wfsBmP5RGckRPyT0/ko/2X+nEqa6KLIgnD+D1ZLqUONP0xZ
7oJCDgY1oM1heEWuj7DoLeldPU/L7eadpk/CNqEQn9pOE/fIqiPEspwYuW1vj60h
LIML57JgEkSAFIQiIRxWsWaRRzF6/0+v12b8nWUEGD5J3H1YdgFQerXYGR2i/ITX
py09QvRK6fe/UxRct+8DBlj1Tg1jrEEatPIv7FYuywPqT95gPyRz59dyhFShyDTx
jtHVSGT5JrHeXDghRb+XvhEnGOlPSisd9NS6r8IP1Sv7rs93eSGtgEeBvvAqqpBy
xLAXPmn+kntVSW5bxOpbfXNKUWxNJWrWcVcjd739y2mv9orV2H86VgHv/iffcPvK
Onq8LD11jy/qw5x+EyxznX96vp2/biHewc21NM6wNMPf9bR1rfB6Tu9H/9CUG0RT
+6j1iQU/8UTjF7zXadnV+O8KjwE70EP4gQ3mvs5gNilT/5n7nE3Xbt8mNl+BRk3k
n2pQOZXmY7UfNmqD/UwmDemwN67p/tqqhcKUjiFZ65XW7haio7lpXpCE9DkN8Ez1
Vwa4E6B+Ga02QZywECUCJR0CLYjKpjFkpAsdsiqlkuT4JE1BH7OXU8UgF7qZDUar
9vR+T6Wu51SbvwdTRcXnZo4rFrugwJ+GiMkt9sHiX04DESv33qKrL+NYBG6EKsV2
iJs/mcpze1NreF9FfUGdFLeDAuPsRw7RkOraMd9g7pMZdty88YX+evJkySH6ndcD
ygIAkduzZ9ih+ZdzkwdOr0Z6nIxDDAftmWObLXydDhRbrgGw/x6wuQBYfSkVq+rm
0nF6Y8+3nz0MarArbsTwmEht4ECl8MSh+rkqrKmSRgxcgFnWnOeYzoiq6A/Dgb5Q
i9hH+E5snAChVFPQgZMgPy1o0qh+j3R+43XWb9WFbseAjZa8rizpIrKpXZ8rIXJs
BabfgBX9ny3aiAbCqxcw2VDawvYNmokD5hP5J8aDWAEe0GOr7no11h9VW1s4GRIh
WGv2kD1TMGCanTr0p4EEqpltLPpV/kxOsgt8a9LyVivN79KbrVyXyGVA6db8pnnG
8Vd5BaTGMekMlVQ5Ee+ALDfuWCEogfE680Mcp3ilJMMROjWknPjNOlxwaCaXDobf
f+lt8bV4Oj28H/Kk7vUBjK/KwMXKKtXGy7O2J85B+4+sM1dLLfaxI2tqBzLlpub+
NLTUKTerUZGv4E6cSsKXF1AYU0iOI6ZZrZrqWt0W+sPFNXlolUA3ORcmIC/NTETb
vhfk/Lc/L5KkLHLp8kC9qXyEZUVgG1dMxa6TjHDzNMNFZzOueGnGWa0oof3iXyRy
eqN97CTXKZD3wgYfRQtyED8ge2wOLKdRfgJNjZBaKhizF5OglG62ycFi49C3xvlu
MfS3yD9fpMx8q+HIsfvQd8lIoVHFqaRTKTAzq/KGzjFMxNtHt1toQMz2UMyF7XKG
wU/1CN3uPn9X+hqeHz4fgigb9hd5QVhLWGZBJSWdm7UjhUdvnEqDThHFe4/H1sKl
gbUkicBByyMO8QOKWUe8ku9nMS1+5ibQWb7djzqHGh7JnzbVz1UhVBJ63JhCfv7w
3jPxPcx4snEjtAlgNv/XjznSI9EHXPdHIbhpQm0ZdyQcZ+MsykOcFaqkbUk7/ZBo
ZbXKPlUUDZhA4V4PKSdma6OgL8FFPcpMmTkjir3TIKDGdRtaq1AlSjVglBXWvp5J
Me+cKpOaLTrqfDYMrP4fSTjWfRIzhsdRT9dUjdo42jjrDtZJDmUh1C3uIgPbL568
vfHUqGRTvojDWZ+qRMmH950QgfZXX0n7MoNWcGmPsy0zuy89wmi8K5J7SjP7NjlU
eqI/qbQwCZMMFKpgIOVUOPI2eCpyMHQD4NB6JwKjl1f44dGGEe2h1ydJN5xaYdBd
iek7zrimGBOhJx81VtITASTEGxvpDhSet6QQ6JsrDkmPIx97nCD+StcoGn3HW3x2
JtCXWjEB/3IuDod8fyTVmEPw1oCaY1CLZhsQ84YTx4BeYwa/ZcOSEj8yHZE9fjUh
5IXmh9zFSMSTiF4uyHWCR+LXM9ZPplfTifg8xMuk+znZkgbtkPexER8YJ5fREa9j
nELED7p0XL+C66l38ybxTfey/gica700pnV8OVour7Rpn59oHNy1TcY8qoHcyhNQ
/5uJAGJM+SW+pcBhPX+tXdvZuE2etKtsc/YogXxjAZmJq077cAiCkvMSXoM4eQOl
OYwACJgzSuPyOOtokDfyPMe4lJVBlZvcvZWOTJomRbQr+IQEWA9vE0MT7QwO0uzS
ZmAquqnDwknJWQbzi5Um35fC0Rh1hY9Jed4rfe0iF1TbLvCUwR0e2v7nxRmAMWqY
2jM63TcGen9dAxg2Y1wyqa0Dh+RP3rFjT07pn7qWqnscbLYRszMcXy7niLF2nEEt
wWlDrR8pZWT0e4s2YwCxZ0vbAjTBJNJtRtxHAVWTOB0b44civYPGuIVJDapjiq0N
gK8bvE/8hm+gubDROimCzS/4qJ/glWvAydWhf2KyW3hz3ccWB8tlmFXYjsTcGidt
icGtWbISksyl9VnsmWqEb4184c2JwTVkBpjjHHUjmIxUSIiPbjqq+uqU6Nus85Sp
W1vpSqlur1a2eOCISp64u0x3uwJn94HJYv8VlKKS6JS6rne9t7nf7O9Z+ZhCQMR1
GgzKjXrdK9En0T+l3Og731mJL2sbc17NfgCt1gSFGrVRxX4Z24fiXFpYMX+D/hJn
NPGEi6lgAkzxFJCMUjHVwtAOCg8g0il/ssLQXwgYChbsahIC6DaqE1B3z8SqmEsZ
Mp842hMDiCn9ApVph97oR3pS7vcV6gGLJQR+0nXAyzJUQF2IdvKCI+e/UsweCTWS
ahV1HA8sob2VOtv5VP6dOmXct+vR/QCld9jr4yZz2Kdw6d0l6O4zu2dWjGH19RvF
8TxaJgM6BAHVPWwDkgiBHA1SQldfBiICk0FGFdU6er/EM+OSTDSkkdS01R+omPZM
nMH3xiB43Rvce9wXNbyE6DTAHytVu2B/H3nqS1iATeIoV06Jq5pucPbv0/H98riQ
6qwgQzqJvlDbRdA+3sWdafAsqpopCigDqzTeDBnwr1POvrdh6rid5KP9bRq2LfjD
P/AbE76Oms+M2WThk2ylnlzdxQbFAf1p8/8gEt6UYg2myaM59UXYRf9EpyGPo6+6
ay+odrzUOAks9XMaXew3os6geC0hX0GCC2616spqt8wq0r81mkcpTh+HBQwpZsfE
JyQc8WieM0pHNyhpmNpg6xzR26dOmmkQRAOytnrAD9sbrZzSbT1hpYfkIYrpvvxF
fb1V+T7poUAmvpZdMt7GaqAwZE+LWFrzPUhSynJ2gpfft/gXOB3v70i/rkIRfog/
evz20JtFj4mZTKsrGqRmQqYMhrfJgOW120QB1tk4oadx3XP9I9S4c6/Q1IqnQkRy
gjDUdNcEFdF7R2BL362MVaXlWZUZKZH5Q8Am9RoTG29+Kf6KWUu7jC6Zdtut/MR8
oFapHFR4P6Zu8DIGxPkbh/5XuFU8WshTCVmuCzzPjU2+e3XsHaQ1lJFmqbxWtzCe
OttHMZfwD8nb/ytFayNSJab1KC3BARhSGNYAnTq6QuJU4asGuMNUObBhUDFORPUI
yI0Ukv7cW1rsbAJcLhCyZ+V4qzrofEcIJ7KqKp3xIF/hT6iD0GP9PULNy7PnaVCb
M+Q6RBlMznZ2y4sQLOr6+g+TJvVgo7eQJ8Ow97xcdYWs6MIOneXYT12QNhQrhRTN
VrJyObAZredRIX2Fo00EqGqI3AvvxJpqVR6NkdNBWhEfkw38/OQ/20tWwt108hOy
Ix3NSLJKHgXYE+zijnqvXPEgX05snHsXBJtwbBMJZ2Tv/J4J5WZpaqI159eP+9wG
BBQbNC4SsDLQjbH2Ov3yH3E+FLzRFAvJuzsDuFKwik+QNA7xhu+z1VdF449Q7Dem
LxA9Bz7blPTDKTO/2aidHBUxNberc9PvjJDkM7T/0H3YyKCmsLSuiCcauBH228yO
XaICTjMZ2nS/a+LR5y/f//YI27/E2AJAbZrzQ0zNIKW2dnODS9Q8T0fU3CsLuBVX
LH9pa8Eic7UtN+XUg0sY4ztBbkBVHqbgEp3DsR+F6P5VLSQUoRAyydAkA7PmsNSU
lEZzjcIv0iYhMO0szhQxRo7rfdEKmfVj5CCYrEIBDhupWjSkUMI8REKV7Mpg/xiO
pdxkKQpwJxu+uwbP5WBZhvWIZMrtTU3RTmECmvexPvVpZiWobeuK4xYteJHKP56b
0ONN+dJ32SsBnJX/mSM0HEEuolIvDybDRU5CkbDB1waTSfzwp5FZBetaAPIsfnIL
Tx0o26TrTy/dU9z0CzzUK3iVL4Tjboq7GI4Z/Eb7Dd4EUThndfu3GEE/9/jCl6Mc
2E1uCk4CsRgJrvWvWLm9MQ==
`protect END_PROTECTED
