`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7r7s8G1rzMxxj5Ktq5fPJWgqhVuOL1eC7GBSW7l3Iqqi2gURlFj0vf8m9+NLTUTz
64LF5g04hLDEFB2i9Jq+9E1jaFVcIyGSsX8l4zx23T26nQqGD3ObHHTotEdxWz0u
FrhIW7qXxIEHTjIAWr4u5w0NjeyPecb+7BxRiVAtt1jLOZyzHnW78I+AC/9TJZes
Ia7xRKgeMEsdpRtjSnuIUGeiszwbkMdFNpv+V+VJgOAOTGaQE0gjhF1a3wg8YhPc
OLW7ew4+BNxu6dhSptO8Czfg1LOUlEL2/qPzhGsZJQqLT9S8gr2OaCWGGsBfaT7P
TiUrjxmRawDFamY6EWLBrhfvrsXvgMIgPYnXVpPjnYhLnzhgzsf2xZ9ESPbjPgXz
BxTYIGa9hKBWSO8FXnt/MPq7nahNpjSZXZrC3In1XzWK0ITL74AXl7dP0hJ3pR0j
vA02JXT6WvsPgsml8MltYQ==
`protect END_PROTECTED
