`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ME3bTGckXpCpQGbHWeqP9isjlQK5/61W0MvOR+dHxwS0fv7lC0bViHxuQ4h/Aqwm
m5q+VKgeVQDy8tmeiOwZVYVj0SKCxd3ReLZJPnrZoy3/0gCsnPTpWfaIwCePKgi2
AUqpFCeUAXlP3MnegVGq0MoCalCk8nUR7vN2UHxcg7m6ByfUXp8nru4FgD/SWUOK
iR+hUPXXAl9VaWshd16qJkFD7BH01RQMjusTwPGY9mWcy8ZFT2pMaR2lC3SuW7zw
W2eZgnGHaj6s/Czox9r5rjbqgWJLptQnWAG3xntir8m7/YVnmbufuxk5p/v9ob2z
3qMNSXvMkI/Y+JKiGSNbaPdNdn4GqWWD7itDn8igKL6CYFzpUfi1HnkwbZyJ4j/q
CxVuLXYzJ8/plP/DyaC2nuj89EQk2xj0Sd664WI5xl2o0TAVJfe1WDbBTQkWMIWg
HqFbpzwabZvN006eerDCxw+UxvJNOBYd8YvZ9HULgy4NHI6GyLIsmEVfSL0oqRKP
9FEFR06jrHk0gGROBwMpoQ==
`protect END_PROTECTED
