`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mT+juGg3poH3g/O4++/+O72/jaf59mYcmzkxb3dYJ1gaf43MqWiHLY94i6QnOuxg
sjnwVAyeXGgIMNcl43YYc31c8Kv7xwrc35t/YRPOO4dqNXi5iDKRlroCguk2ojAd
cdAGXiZNe5omZ2gmywxOvys+BI0dWaTqzPfh3JTKSu5mt7/suCGc6emH2+MEifKB
nSsSZvEEa0vCGgB3UAjLg0pNR+qhhuXAWokjRfK7MC676+HunRL1LZxVa27i1tcn
C5Sx2Af2Y5WlgDaNAyQQX5p0Ks5axsk2QIZrr5fGUy9HizJ1J+8ECmz+i1nV5Jeh
Eem8K+W+om5/6mAmjpqbL70h62fGZSqyFoJbkd/sOoN/dAKr0VWPRbU6WcXxQ6q2
GMSuacMgvi2ron4RwBifmkJUbCZ4CngGDl00DW+X5PWe705cRu7A5GHRpoN/VO9B
3pngJdz1IpKkBW5VbrTTj6cF9L9zD1fqtDQleQTulpxEESDhpeeB+LeAdxYqtv0E
oAQfsfMWQ6cgELapfRqokO/NYM4xcac/4y7edbP7xRPpjxh0gS1IXitK7jtjufBU
dn922O9o6qB7B2m1eV97Ct7g3NGWDksEmFvG8+mwMe9chhnn4ClCvPxE0cmyMeFt
DNd5FGJhxOpQ0UXByq5DskxemqsZos/JcMJGAvLB+vPA0qy/yGMBopYd++NIaN6u
6QzHdPkvAyYab/HGWTioet9mq1s6c4flUNRMpo9BHmNRExOnRW5vEGujmtod3rLP
iRdFZdk38sjCFnCAujuOaQ9J+1Lv/sd0QndhoIS0Vtmt8MqLi/zAguE8Ovg9TKbP
0d2wJtxcO1sLDaWwy86+kgwAcFr8lNm0mtx6NgGj71+RUhRczI7VrYKgffaJmIM3
99qaSF9dJhJ2UMI9B9zerTmvUItsy8Rh+rOh/VbDT0QCWUbi55OU8nqUpi4ihlCm
dbveT4dVWF4ITsJhiOsOv2iCT8OiMkXr3fE2VQLkbxHGnp70cTTyD0tQ9a2n4JvO
XckJItxQ6K0Nghcou25oDaxH506GzsDBEoJoG7SGwgJcU9LXcZST9W56ZKVUCOPX
81oQKlKZBV/bW3pGpu5F/3SN42wm1WJhMyLge0GEK1qx74By+uVpruR/rJIUGZgY
v5kfrKnHZoRM1RaIyFIih5BukK7umEMQ6rmlfOWP5bzGlUNdpv9tdUszFAFu1i9g
pVLNT4EjF79mFYZDQq4ysnMA7my9qTF7AWhWxAR1aUMLnkL60t0Bq8X2Ed/vbhSp
TaY7Ca+GUt0d/Xj4M/77FIjat3Ij9ggR8Z3WJBiNLtZXrLUpZNLh9aqTRIgW5Iog
JC5oHOlxs4Kocx4WS1DsEUhwn4qB51iEZeiRYWs0BiVl8sFtYmaZhTy15B+zI7x+
NuT5bhCQEIoCTak1/OP6HtoX81GgW/wSwZ+Wrwx6Jrdcplib5LUtp2VUXv4N0nf0
xZl4kwap9ifcoqedvKxHXpS0rJFutmNvnPY+1PH6uWxAKjoRxN50U+CQUTePb5cc
Y+7FD/T7siKDL4oM58CWz0G//4JnAy/2nqZ2r2m4kfoaC8N3JYDDkRghyhCAaqrc
7rr27dIp3pRaqqhgDiYXCKDBaggQt0dY6JOJgrzmgbYnEM9gAi0GwoHoIN2kQNzy
ih3J67nIcuMnuLE10YGRV1cB1NhoCTGXNE5BzgrjAG/B3M14x1dzvzA7kENeReZ7
4HU4uCdXVTN3aGnWMkMc9BILogQXSWpAmbdwSW+gP0fiV/VG3fJemwhAg4WfLaYG
k5HucpHaDLhzV+C1nZhiZA==
`protect END_PROTECTED
