`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bJV2zQjxkKWnrTGa6kvdlU8QiQabnZ41WVTKKzKQw1iVit3gwcQrUfIyLdN0Jk7P
fUIQ8VHS/WM0eYWCOk9HaleePg7JkHqXF36VgkF/dZ2Pc2uedjpqpmTfXjYC54gU
gEwCOZezB9f2HNAACOzJ35dWWdxNDBpOMhqU0dy+Q57SFvhLqHAtRM3oSu45gIRt
rqA9asLhxdfmBAOQq5WsrIexjtsGwTSXv8ibk6Zt/uGh416Ug1pPnXm4Zyy9ecx7
CtPfVbOtBsalgaT37l2yfjjqUwp4QLT6MwYOApJcDj99x6FRLGsv0RiWmNfRfG1K
qg0eUF7MZ9V5PQvWzscuzGjBqqHkqpZVd7P9OjO2EXK4qSA2gi8aYTo05dESLsNE
/0efUadS2cRHbT5NwnaDtOzIQrKxKoyGVLOTLprJ0v5VysPMVP/A8vqXPGCjCHhF
/cgjnzDWaXREMNoprwPrv0GuIa7PpCWOn5cd7KTl+lA1mJ6QnF/qnlqcQk5Lx7LB
bwqkOVzXSdWvF0BgwbXJzJGixfBagbjyPNuQ/1pJQB8RFh+xw3VkKZQpq/7ILFxW
rhcVm2XUyR8evdqjw/Rt34cKUl9RTz2v113CPgEVPAdT65sEADUTKk6UYF3fw3vn
mCitR7vAnvG/yMA1LfH2Q1ITRi0o/CSiQPvZpbKdAxlncDSdesvPdu7BzENE1cul
iHRR1AGJeJMakkeq0Ku+QgGG9zzh7sntsM9YJbd6vJn8mjVQmimteRk5h8KYht9m
G28bmPZCger+lUUsH6mOD8vpU3rznMzOgyV4CzxZenLzs6LdGDahaqfJy6imVaRi
LSibDJCEr2DCEq+cW0xsmk40WarzADByPRduaXv3Z2gCwX5SieurJDn7bRgn/Lo6
wDHLWfVPoPy5ze+o6bjyfBlGo21E02TL0Bz0URJ/okt9YAnl1gs1BlJnvjMKTFQI
hGHh5K5UskYVA3VDW92LnkeLw3inDkoYUleTP4o9d79XEUHFgMwHkVIGk0mj8exO
f/5yemuYBgnHIaM++rPCYorIbu+lcPiJKqyovOt0H8IZOcra7h7RC+8TS/EAKsYj
/6HxpWSBavolxD/196P52g==
`protect END_PROTECTED
