`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6C7c6J9BIdqciYyGGW7DQBrlcYpbpRgbMiJGI0kLGQuhRVNPN7liZnsJ8ZXPydAy
CESzQHmua30TvVoisQ5A8hd6y5B5/YL55IKu2PGDP0JNjNmUeGEThEGlatupMp3O
NKgLHzPECZw0DajUU+RRyAvlQEoRjLNPDJg0NE84i0BRvUcyceF3t4OPREgTD0HG
ncC5gsyowQo4bM63wrhww56kRGFPgMKX2BKJ+iMxAQ3SeRRmYXfoADoJfoDEkP6P
pvJ28it9YQAhCqTdZZwOMqKIQnKM8ZXQ719VQJfcTrmNJmb4KNMme8jr+i1/8BBF
188BM2DT+7sfogciLdU2TpQiPUJX2rXctcDvBgOwAxMry91AlnsEOf+dukI2aQ1D
oYRu0V5dSHWjYUdV2Ps2Of9me/Yk1t3h2SsKfKj41uC3b3c+V9zx8pq11MfPSRmX
VMYbQ+C4l5mN4l/aJK1wpuE/gGuvBbLlz4Ee6EvXDwBHEh4yqdwZEbF6fYSnrtby
DHR3MpYHc4lDb3Yy7TGeiR/4d91fQD4oqLfUFqkzuwHa2nWEVQOYkrc5WRs9w1x4
ZNu8zOCBDjIOiHsZKVc0PGAaCZPgVv/o+rzAFIt92vLPKqjH2cLVRwE2w7ZOZdh8
y4s4G36pDL9dT4XtvCXDyejOLFfo0glI0KHWMzPUuFKpM+GIQH3n37lrUyqkEoEd
OqahN754ZwuFKrGLn46bDg25AlWBS8qOMgGxJpXz6AqguQSu4xPTWsXzSwBsgJ7w
mt0yMcAoV/SzCS8ztZlqAUI8zMwRGpPg5m71xdXMBsP5Xr4DBP1L/r6CHPkxGCLQ
j6xtw3Ec5uc6uKiRCVzhvg==
`protect END_PROTECTED
