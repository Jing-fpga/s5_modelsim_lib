`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
51unKENPHLrrtFkAHROxLYGxou5FhH8h8DxMgRy3upJa0KBWvJhj87EQSZvua/rf
oijYEDr/+GkXqfEjmbsjl2M+MAHD2st33wMwiSzjGF5RIVNx0RfZC4Mppc9tYFjw
vBeVP2jv6TCrAZ9M7Szq8TQpkkfSmE/sLwuKpL31H9sNNVCJ3S1C9fWXmedAfShM
5Rtjzo2U1YKAp/DJvxavq28gHck840/65woszrYMEMOfVb0craIvqA/5wxKOEzT9
JMtO8IXXIScpGAJ4B96lZ7cGmvqcHAG8S7brp0U4dN4SIaifYCkoT48ltRetURzq
3MPVpa6YFvfn+jUafaQpFJROsyWwzN/byL53bHn8kML1OYt154avizK+H/FvQQhu
AcH+Iv8mTPt3mjoJtWD4thuZansJadBzrJjYL2lcfSC7AXaezNlr+Kx0sxk1VjbO
h/wEjm2vQ9ytHdPafvJxaHRGdMwIQaPA3jtAG9Wmr0cY+gGpLDDHE9ZMdfkhs+Ch
4pLWNYh0TzmPEypF9y+aRnJsKYm4hC6KYJTzq6kQzXmS+071F4xNq3vUCnQFxob2
LYj1iXkFXK6X9VXsRTXcHXfXh1d1AJg83nNZOBv3W3qVUOAFuVp9b3sZ+f+yw/fD
ca/mh8WH5hdT/T2GOJYZq2Qu9OXOuTBYQqrjVN5J1jbAYovboda0cgj+jFsxvzU3
RHuzUn7UtVCbFH6w2bWz2C4Tqsa27ImWvlgKoVzMCmGhDBwl8WEoQi2Cqj9r9iEu
h35OeIqW0EzO5BoZGkzHZA==
`protect END_PROTECTED
