`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EoGhCksCtOjdhdUVMjRkgcqlA6WXOa94qzrtwbCsMmdkvXrfT0taQbfr1QeLOQ13
fovf6puQlP42kFdRpd1EsP8mqC46Xo9vH3l1gLiGaC7EXP1bh2937KVPvktNLyCU
+aGYTWrKJRrM9isQOf1VNvtaGXE+v3btZ0uV52JaSc0alW7q16TiqqrnPezUfn94
s3kVd/EWpxxazPPDDa8hEdaYuHSZLCDQ0cLwT++pmP+b4XeHBW9Y1RX1JCR00itM
c9aR7MaeofJb8qEW5LH1EPVGlhkfXxNPW6akQk4+2zwSHEBekSFt9pX3h2GCelFV
7TCCk4vmmkVBEdaJlFPKvvfu1LdjuJRwDipBDHkcW5xPmk3N9OytGmV4bRVMqNor
UvEpCEDF0U2rvzLowBfd2JyLML4LhRIBabFPIBYHT5ZhsCEGJBT2jw3RUmR0UREE
c/Ot8MSVqsybIMQ5cmIT9K2STCCNu+odbsAN2Spw2S029taprzjlL2O66fuHlNtF
QpOTidGnqQcCpC07pmyYJ/7lkt/lc75J0lr9ZC+RKjCxdZRk+pfGjeLnreRuejwe
MU8OvM7Sddief6zzu1Vm/DnSIZeShaRPKA7cqXwHWnpNyrQGNieTfGRtyV+GMiOy
xSksDmNqIgv6LzySbcSJDjhHciTRT05ppzVdyiZr9fkqt3is9P7OhKezMRmQVTbh
pEuxxGqw96UzHgpEVTxwWijGcwjNfkM1JqCQ6fBELCCS+p5zW93Da6qCY0V7fRPW
ZZ5zY0zDM1obU8OLzZscWSYabfpqZxoEIbeTCAJDGlZb/BG1fECU4PTMYi/l1lkV
OR0jDXygkc6EOONSvqNyEdokvV7TSkLfPAeBVpQ3Smg14OQ2o0hleB7oblft9+ex
PP9cdER1rRPvjpz6J0Dz66HnLmSQS7UkwpAbov8Bc0xmBor/9MEfqhFWAa9y059w
ULEWZhWniwG9m5/DxQ48QsSzQDnG2rI6VFIjJ39RuHbwPPLDBXy/t4iwZEU6tSXO
i5B+8Ld2HLOHgEfvfGr/F6xPp4cC77xfYeBtsvgLvB4XyXmEJ7+2KizMLvLB723c
`protect END_PROTECTED
