`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+xbjVZH5+o0wMyzzmouWx9VHytfOXwCe51Z3Pl3iHdNILwcV12KctC/jBtYOSSLA
aNZXcN116QNCB1UxmlphMZJAlXYWzLATtkIgGK91r5+J8wh1jaN9ih7ZTm/GTyal
UAqKkBR5B2WD+rzlXCxS0x4j/8RORiSwoCBQn6T2U9JYzagxE9E7pQFEGE6gdId7
2EzVaNWNYJk8eMGeGUWILr+gjSyvNR0lyDmO2nQ2EaxAKwk8o5KUsVPD5kTcHYTi
yJFDsNt14WtjTzXImlZMjrMhcDD9Oi9jBQMQVaa37wG1ifchb8V/371Pd45A+spy
PMWXJa5uj4e4LwZXywvsBfjRK89MNBcVuPdTEsrR2W+bPoOmc1NBcG68RUf8clJw
gVaXQMdC2rhRPVq97NfKyaI6toDT9SqRVPOmcQJd/df/WF2cAxNPd1QxmIxxfGDS
L8GGN1I6p88NJ2IieZ9ClvSEjp1uwkRY8SUtwyDtR0HGP7rD9JCalV0smw5lA51u
TDqAiK5mXWTaKViqFOE5hsj90dqrCFQjcHWoLCfNQC0wj3NO0+24O8RquVnf1zDo
2P19QRIgun8LZfKAAvHJu30nk6hTvkmtglH6lclUKkVTQKtELKnU8FTado/H4PMB
nCiBqj1ybBIM/NPnm665BB0ZRsRcfC7sESa9TR9LTpHHmKHWfkcEQCoGwcP5nfg8
k83Jy23MQIbTOMk5Bo05xSt/McRU/BmcMk8fSwi0S7lyxhdbX7hFZ18LptKZnHqA
O7VmRuzO2OW8kax3OIe8ZDGXjC0yW2FUXQY5IRt6vFpZ/gRk0CjwiR3+lKCBh+ea
1Z6QVZ4yaT/pPuO0O74xfnJEz35jutZj7XO2NvoD9MDY78z0aLOEbytg5QmyDlre
p7qwkZEZ1ELUGeAG4wosGkmdN+7krEhE3NM1eYl+pmgUrT9Z+wgM4lItYyDDTsO5
`protect END_PROTECTED
