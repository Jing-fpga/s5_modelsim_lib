`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/fY96MbH1naIz4fuAtVNXGjEBUm3rd0Pd04dhLacXfTCHxrVz+yLN9IcLI+xB0Ut
NQGYVqFRI1XdRjl0homKSmO79pkhV2mEL4gEs1+7CLOlTkWvqcZBkfjYRLo8T+It
t+gsAwgJ9W1+LmZOJtVGl+VUsveXL11tr0FvpxHdX534JQO06PpvFxS6/MBJX1xp
k3wE/99S/uo0KTYjf4wgZUzfRyBiwSW0YRgGaL8LVSBP1JI+W5ALXFD/gNSh5nv4
pPmaaFojtW5H8QS3liFzJr/p9LjxhlhwSriC4lxswEELMxiw5h0dkvN+uTxjTyUa
DNN65pmAhoIak931CDCtMoo/HKMNYumUx9Wr6SOf2il0KKY23hHs70mzL9lGF0iO
eA9FuoI+4ASrPLJZHR9YGyRuhTwynI8HrYL6X9Hyd43qRi+KWNvB0oqER+Au/snB
5hxQ4UOrip0WU8JxPug580f4baNAF9tto0Vq3EulnL802EZrX9xTvvPpcs8nOxfU
R5xl+aM9gtAbJOLuu8ZdrFSPazt0N9ocRpLo7aZ3wVSyM4tNWzLtGfyGvYuYPQuA
9vPoQngDNQYWPHVBEonNwIiFo1EEP3LXJhSmu9GDVjhU0gWPvS7e5NdlQd3/ulL7
vv8NnOy5H9Wprp/mSL7wiPnTyJl1hVzGCp1eVsyBJfD19qNR2mEeQyXSkQD2m7nc
3Qy9RalIEajKb3bX1ICSxigsuvLCb33dex0qXyAnyvjLEJZZV8xw8zpXYPMKN6u7
BIGe85ihpbe0ehKq89rAg5+4WRPWZaovWepIQDHL06jfQVsoJ1JZKr2VUEqgEPcV
tMM/d5C/uT3jyitScZyayQ==
`protect END_PROTECTED
