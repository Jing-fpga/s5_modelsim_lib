`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jnIE4JUUYOwViYvHpu0GQqZeQXLvqTIng/dODrK5S/thEQdGeZ/pFSKeWBDM6fcb
E/Y7qBHfXgHUk6hfm2lFeHVIBrDoCVP6mzaoZe0+e/ZN24qiLa2kBqNionz3NbAr
G+VmUsgFh2SJKulHDazt0o3y6zS4TJzJ017tnMWpkoMnOYtSxcDc0RUPQO3L0Egg
ig18bX5QVciJFvuoLKeAhhGtAri7wWEallT+X2llHxQsLOHEgVuyr/JsS7VY/k6b
sOEbzQVTHfbUX3PpvlW80YSBgMmd4hcb787q94ivl4UKJP4RrpPYXVlUxF93iDI2
fbh4FJoH7sPmzzdxP8p9vYoHEdDTuHDyaZEIrpD7Inc9Wi5rqhLrYsxxuEuTJR7+
soU6+lI7k0IgkZJw38Z5ksmS58Aji9/VLKlU7QgvMgj0Rham+LaLHZR8vKhDMa+B
98px6T2eSxEVo/lnsN/bqA0qP1iiwU+0ZN+CD0Paj8wvqeq85bF2i0gIf/3QVXBZ
LN7g0EQGrPExLMweNKH3uD7W4aewzmoiN6hllbjlSI6z9PlFNy1cvAQ3Mq5d0Kn5
8ViLqEq+98brMwfORxvBsk2j6d2xLr2j4fB05LmxQ3YjzFR6CHggThs8kWclgBJL
fWBlK68eWrbPvuERxTQ4UQEqg8OA0OphnYVoxVPTOxlYAjMWFtZERnbORRd1NnVo
gxEpx3cuUDFtF5xqsZeVJ1n/0X2TlwBRU7k2RP5gcx2jibEnLAwFqDd2FuRjtZpM
kk91SKHINQqG2+k/SADZRsSCJZvAbvNmPkqApnEA2ZtLilfmZZQZha5UwFfTB4LX
TseQOGH0GFmilNhv/U3R6EpD0+XD3xF3H22mRArM9kWtILnkZeOubfq5s//Gc3sP
C4Orfiq0g9bhj8IRUGXDOKpBEr9J71cJ+Hdgb3QlQkowuRAAiCbmDIKMghgRonHa
`protect END_PROTECTED
