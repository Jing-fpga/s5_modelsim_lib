`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GcQ6gf+dIrUMPfhWf9TardpFdyN7+/TaqNhRWvqzAfcwbE7FNkNfPCr3ESKhLR+L
sf2OSgJuHijAqFHoR2fSv/JDxrrZTYkIl9Aym4ST3o56wSUEEAGG42K1ePhfVdKN
OY9BFoHH1acVtZOIHZyADtLcp0WiBbxWHndocYCqw/t2gy45AJICSdrCIAuzs+5s
ljsWbX0JskaV8EGQ9DEh8QHKfVgX/faYSaHCLFgOW4iJxUVyJwSrxc3wHGG0+lye
wpELCg85yNJ7UmOymC9OcAua0hOaszXMpjk6bQc74/blnij4JhJyjRQTJFSR/mQt
Z1aqMga8LMPCagO4O88j6kXDeWteRZKVYMGRgKL+Qz3lvFnnNPPRGHVRdsQuzvET
+QOBSH8Qdu5inKTC/YffQTh7mtLUSyLu58U1hXPnoTX0KmaNrClCUmMdWw6KJ4Hz
`protect END_PROTECTED
