`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L5tb+QIMIUn30H3ynQ58Rx/G/dqFPZ/OaSDs9GWW3JUOgt7wI5CdsStfNAHJ4y4w
aQ13bQNtuj2k+VpyzD8Kx64JX+Tt1D/w2V8gXkAn6QAjH1nGTTuVZmf1FgB7Dxyy
LunOxjWR8oWGc8B/dgJJ/G0j3TNN/SLOoMjrdMKAP0s0GGxdsxydh4kx8SAhbSD7
DfvE9/GxXXgfO+M6JftXPale+Hw1TgP36/yWms08MEYHcLkb/nkZzcIqiTtedEP2
HN1aEoWkF4zhZgn6OjMDe3l3/khquelQumujaTVu2GJKYbFfxkGu5yTfaXafXG+F
jx20BV+H/orTJ48+cnHNrzzMwqPy/5OlrQUfmKTBSdyWfoll9AQ3sXnd96n/2IWJ
kSYrnNN/+PruYpuyMfYcdTAmif+O+rqbMvxEXdXFCwG8p2VTb3yRYZmXHkc4a7vL
WtgcEe0ElKFKyUTSis1JTEFTZZbFtkVEae6KlW1INpja8ABEqXB0f7YOSbWOxZdr
fFFL247RQkdduwJLditQ+gqKMqAKHV2Iih4/jChRpEhtiXHNGjDNWNQdMGdy3L83
hvj/UilZQezfKVoZOaqNuTOkDIjmy8nxc21ZonKK8ZHJglpZ4BrNY/VEqXHspcl0
kqeZwUeEC7ev1RILuREKw1b85SCb3PbeC6/vcJMavsgzO/GUxfgayhdQtYm/tKVa
Dv7V3rzFtaRhR+4jBYGSYigDEDYMHh3dlGQc4FJuAobAU4XoljeYpv4R2f+OMR2t
GZu5iforsUkd1aEbCHP75kGa2XVU2Igz2/1U4c9iELA4yjNer3d4U5d+3zM/14G9
Nzfq3ki22maOSCXglrQEvhna4VJL16DQ/nXDTDJaLNAWhSarqpVZSuCmRTaiXGMa
PCSTV49j1rPv3gWbuyqKA4eOQAPoa210EkGQ8A7jY57MmwnnmmHzGyNYukWW+FH0
`protect END_PROTECTED
