`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UY+h81OMTu3jXA/59a9m4Nz0h0oLjN+j0k5AvVsllZNVbtUkCheK9NckTuvHbxFi
Wu7U8sRgdSndZB8tyQxHvldiZAZkS15HOijxhjDNHoiTOqbgXssv0E2QSFyGvAe2
vqtABUY8YnLKmVT4zbp1mJ33zTrEa5vY01xzbug0154P2RczFhRvsETmgVW7XdvL
HuvpP39csbfOO5qhzoCV2/dlJ3fDxWFt+gDpDezApmme629GsZDzr27U6oKtNTVK
pDEUgI/5mUCXHiQx7G1mUDoxlgCc0f6rAV6tXbafu7ykNYB/U10VnbEr94wz3XbN
FE2tjhlZFyrpgnGMCgvuLF3hCiQwU5Oa47jxtXv9biKQa/M3PjCJa8EV9+lpktyc
3hJjsGaqmTsMoiBiy5NmZ5L9kWP06CsXgIfQL1AtYMpguIV6aGKZPkQN4kgh6aio
zi5vNRdgkj3MxNbCfG7SVwUlLYFVkvy4iA88xnl6iLtsZ/z3Ovex5jGHCWwx4/lo
8H/CCX+LKWVjQBrgc7KL5k5vpkFsvQC0Wo6c/d/CrZCFK1FBkNu0A1Ibf+tn1+Ui
IbJULVfAfAxMKWsAW2QRu4EzkXhQqQ/97JH9Va9C1+h4A50BdwCpMXawRxF2+vwg
/P8to1V+5geJHD3qJhRQe881FKcUERw9kDrTvQO4IBSx4pNIvq3RDYf6KXXfuUOI
Tna04BtRFPs0HRfEmrvq5IUUYjt96KcX5ZOsCOBAKXNUdyBhKToCU4xj+2NkMyjF
ya8HqqASljBZ/+1ksFTxXTqDuGLh8m8M47fRZyIHQv+2R6sjH/Wg8kMrFUP1NPlh
idWWK6ydo+yqWNrlHhuSAbXHazJhqU+C4ShmDir0rXeokF5OTxCih9ROUdhRLrtV
BFJSdZ2hKtH8BT71BuoXqt/Q9OZx+1lpZR3GVJvS2AAv6lc9je/Xit/SrxLrahRI
GGf2NWWiZIijnYhM6Boq7zs1DbzeU2hG0oSeOBdkvVBHkHt0ZM2Vg7mid82gYi3U
62vKkEYiWLBQVtFuOM0mX0hES18cCIN70eTupNTD5QJQcrnr0YOKcrrVPljopNhU
4gKeEzdI9Sr6eZdrsIGh8Djnr0ZEq9t6Q/vdVRw9u1wGTlct/0PkEZ+QZW4uYNny
9ioeFwNssMhHrsbc1YbqMd+Jd8EY2gF/oBYyFq/beWZbgYgpPgKB3Xvf/ZBAlC6E
nGnBCm/EOIM7bbJTb8mH7Uxs99FCgUvmBU5LwjkOWG7CIdz3/6304h84lBuho9aW
LfonScyogOZolxl5NnGV2QlAtXrAkKwWMsj+Ha9iy7yNk6laeUjg+LMdy3055/sl
m2wkmxyZxyDhYSQqJTosT6avwLWou8Iaz9qPXUeESrUM4jbddw3WLPsPBK4IfMiq
VS/H1C/2UBLlq9ji9iSgdkUqDDHnefDZ5pNU+aaSsNQFOGrr9iW7Q9KkeAQcsmgy
GquQqzX89PX9coBbv0IEVNOvF951VehI1ZGf9g2FXxrdwh9UasI/ylEYMw6C1yjb
hyHJoOvzDhKLcO8dTV+8nOyO+62zzeibH674W0t6xQOFae+Wb7mlzW015jX1wK0D
5wO2f6D0AYybjMJ2tQVffVjhVtZtkj2Q/AL1AcyRF48HmeiWCrtsgRYYErruNFtB
nTgPIRKNEDowa3TDtuKGnRilEWStZDJ173H3GPvIyyeQdvyg/10BUNr6yOOYkWUx
r40/f7xDrkQkIGc6oehCVpdLnnydldeB6Mp5Xq6Xld27pZLZZcCHJoMpcYS8jvSv
slOMZS2aQRnjiNBtd1JG4wK8bjF5sCq4TawHSOzjsupj6STvxPxcvaNX0r0Btbd4
FltCB9ibD1g5wIGCXD+XcQBq6r2eoKu4u/hrNYFdq8RtznWvI+iBAD5KBNLxgvDd
GiXvCgUBDjT7qlrRRROT6p2Iq8z/aisxKj/qo90h4yxMM8Ax/QIU+XeKsbfGtHXd
Lqav5mByw1LN6RUXcU1TzM9tB91fL1zDPkw5rWtPqvEvbMfKA0fTZMC4P/QseTmG
9FzkhrogASF/miY5qu/twTOUkRMNvndYLAtPDDotwNJCs8FOWxzwHkJQT5MOk2hP
wd8l83xrPi31UEa2zad3BT7tcU33KXSmNNbFQyNO/JGP+2tSJ1Rl8AsHGrRhp1j4
jCpCRttWPLP3EXAxSH2Zk3bnn8ho2iaRwk9PdW/dWFEbjSrjdEU5uNTruOnO9Olf
YfTpUjJoWovnRLsFFQNZQTQmjw8WNCrhV/IrUMQQ0JGqf1zoN6K9obji0jpP3u0X
fbgjZCxBnr489pnr0t+nOaOMco2hWbzFPeEX2zGWoDmMuzE1fcZZuAM6frOuGF3q
HkWe7aN4kcJpSn5jATrWaV/Jo0YUgzguU17W1sgcpEWBujLsniCciqqUSOrI+nGg
GDW+CXJVUkjVC7T4+rZKUg==
`protect END_PROTECTED
