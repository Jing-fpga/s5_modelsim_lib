`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MGXSKg+JNI+dT36n7HAUmeMSj9njkLbE2dcNLiFjR0N2ojmceJ+G1BjKeyfs+io3
R1I2K4192tMmskymRp1AtSl/cWV9Ti+xHBtWB2eEqQgaVqaAVK6avuiRkj6U9yWU
Gk9xzfiM1ii0R+Ok+XysH3jrdgC8Ah34SRXWoGQA3VUXUnzDRZkdW7lpL84i6IYo
4THd53E7XmYjVTCQmUqoqKS1XjdvTkCvEeo3LYjReJjS2NsldSp6DVqiHGYsAmqO
c7+iip9LraA6X+HcbCbADwWMzlPX8qpmxLo4GpZRNNZ0UgMNw8MkQir4wK2LnWYI
hhWM6mZLR5kNjC9Fv+k53AnvrbZ22oPn4ArpoUgze1R74O3GLKhZLuOjW49Teanp
x3EzlK3tMn7A2huFbkjKJ5//HdFDB80oUzvVaX9zgt6p0v5xC9r6Fq4NB45R8Eol
U3Dbx/5yBvznka/EKzgqvwPgGx6AgfdgslrIlC3KwmVxsakzxjukbsTjJzP8w8kK
1XPJon5nrVgn6Gaw+aDtDTu4B1wzmFB4WNSsa66oP21cGZ8aj5wlUsWbwgza9Hif
0q8f2byPg7hxaqMUHdX4mhFj7uq4TN7mFu9i2tkh480t1S4n18PsW7IA8wzNPbAi
qIeO1fqiOWunGYEbyNv9P6klQX2dBruI6d/HKVSlucjNMOB/e62NzyhqDeigjLF+
`protect END_PROTECTED
