`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H66AUoR/zf7WefaZdnTM8dE3aY4DkQMYOjDbGKc7cD6Jd5b+iQDVxdRDagRV1A/X
r+ZtaCshC93LSHI1aOgc5WSAECOT7by3ZuVv/440Fw9QCEoiIODWWa46RWG+wbsJ
5BxB6k+v5uLjJIeeTCco1DrJJqpc28Mqz4Qhvur4WS3kdlucQGgGPDG/riPFEBuY
b/HoFZNL5t5txAednQhz3h7pafk2K7Cl4GQVnFDPDHUqp9EhNnTMrABE6WvZ3LFr
mBuOs4vt5EY3g5mJhA61KbCRYbt/LBekk93l4wlKu6DHQbZdCVSNn1XUQcYRLxp2
zLC3ppF+aOj9aueIL9+0TzIeLUa6UzkdYx2dohLBkP22Dl+RGUmpqzwboRmn9jBY
qHhif/hxtm0SJ7Fjf0eHXAJmBX6u2B6Gn6pYiwCQsCE+vyn7nowK6G7XqBF/lb5E
yNJvUQTIG5jl2vTM2V70AOyLcxJ6rs0H5DtV6IMPmcAlQ/fN7ofnYLaX/D8O7xCt
0yzNefDqqHuzxJjgJ0XL6Q==
`protect END_PROTECTED
