`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L8xDv6RQsj79+0axa1N5OHyz6onV1UC4LgzuLCARNuDj2uXhB+9MVevgfKdpQaSv
vY3yeZECpWmlaHtas0KZjRyFHzJ50ajVkyfx+/eZSfwOvH3O/o7ZrJ5mveeFt23Y
JuFnY1CEcqLx3eqX1bZNbu/td0JV/e7A4VmLbFO4LSIm/A9ndzm54qU2zgdXJXbU
VxnQKvn9u6Bn2Bp1dIVJCmJbRn5c08srpA+y7rEZUhxC5SIFAZC+M2JFQEvzWbh0
TK98V16ayXpTtNX1ecgsrQAZf4Z0BqQzBNYXvNtmbIe6LSaKDCXF1YokzKo2ZpN7
DqhX4fqdRqcJZ7pHvhQsHxkO4BUbpS84cmnE7KKkQXkSKGl3qwS9OkMJaGvaUInJ
WTVMB4fwtx73MksqV2H6/kPvHyQqnMtufG8gVLMLuruv6xDYua78cEB1wxDKlZOb
oUVtfSwkpWEyuBlC+gR3SfOg3Fcnblr1Xj5dQEAbK8S+tAZpKrQGj8itRB40n/1q
BLhwDuQSPhYGa4u587NIJF5vgzkDENVGrmfXQKmtxEBfi5jhVKpDeYcL4nsazA7f
BcFQ6EQgIOCI6umstZRylsbfOgRu/8Ie/s3RNKIdKKnV0mtUAMYe2urKBEgQZskK
gnN3gH2VoovsjCpFWOXhQlrO9GeJPZcNzksffyR8iE+pNkvO4BAvtLGist+D1pR7
t0ztNEnf/8Wfa6I7WUxZTycZGy/qZA81vPpQ3TvPPXwmvy2bcl5p9PzKltqvqfip
Ahv8PuO15Rfp6lPeJ8Ejv6ctxUu88POlCy/7JCfZyBe9h/KfTB2qncqYWd3Zm72L
`protect END_PROTECTED
