`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O9Vvb2XKwXB/74QmRiofZj8ldXv8NxBA8fPMeYaQa2kFoJisofv/6c8I+nSiwRDI
0KyobfVQjgb5IGJgJ7LR+CZg5CtweZdKgcQMKTQhx5U9utCOZ6Z/113SkI+Ouu6N
NtxNXkgHTj0UZz8ywmJtbl8uPzdII9m/ml5phNHeTEhcm1VzijFWauOSvamP0spB
s3CL4n2+cykru/NIgAkdMhCpohG8fA/15zu2pwYAXvu6xagYtfrMcXRztsFPmGxj
fbyajHsWfCrBU47PqnPF4MHPVQWLoLYqQq8dojIYaNuE3q/1YoWhWEN1pRR5GtIb
JT11acxzcj2RptUGrbyO2buTcSqldXfWPpDtX1WklP+mYOCA1GMwcCL2Swuz87GF
evJjFXhc+J5cx0fOHm+xeHx7olyyOwjBo1zFvC85Jn617QoRvXaZDIlpEljkP2qX
IXMbCgbeUy8/CRTAIfWl/YSkS4rU0n/gaKjuxlmzt1y7QD5iDWqsYNW3JUs5aS5R
ZkaSLok7Zq8qKkU3uYrfXYHVjK2e1PsLHhxOm9dsroZvm1Wj+HTzz4yfnUZIUpYY
3x5n/qC3GI0D78mcZEoWEqC/GOpwpHEX+DqMNVBdN4pWGbMXkrcbjvRJjK7+KOQn
dw1PDers1RGbLCwTtiuMf9YcK8GTBkr6n/2DUxAbmxbgYIPgFe09sN25AVPG6KJl
/20l83k6d1GjTvHRBn98XrgrKoD208ZcziH5tFziYEt8XBoU+FT2ZW6Diio8IM0Z
DamIWeyqcxdonw0xou1+jL4A6tqFpmU8axoLgo91vP6PA56II4uGGgzUOPJI57Re
moIz07f3Dofb2VVxRspepJasXI3vfBoNNocz9G2hB+IQhycSlx1gmEaQGTRMJjIx
qogPxZ6JY2a/fr1Tb97tPj1o1K+nFZDN0WZ406qFXIXC9qneN956m/vUcNkPm7Qv
+wLSAL87fg/fL1Sqs2XxXqkL2NJPMQ1GgyWRpxW83Tu/duxsTPYb20EvK1Kejk22
j85P+rXILf8j2qjA/qT7uoFoGOruYhFKMRvHo0z5CpwQoLb544BcBqJAy/K+UrNF
EX1MoLLLguWeVKB+Z6hCIIlckfdHLDOzmPXNy3RQLY77oBY9LrG8AbdNR7+ujJeR
RrXNAhHWUmlziOdzjs1nTD+Nc88BP3IqspoAODwtH9fVHjkwUEsjtbtxHJHwzUln
/H2V31J2+IRnGVwQiSPJSgdtq2mhYuFHabUStQsvvCBqdeg5AG/dDLBiwtP54wVq
lXsqxKVL2+IOYJMyozTQF7BEADRJkli5Jxgz88g3/9W5YOLOdbW+Sgkl5R1XTd2F
JfEmjD6N/aAss/E9YSG0qBm+MaQu35xrbJOSVCUn/RuB2ETBaAirQR8Xb/gW2vd2
WLMmemtjePSIvDTBu7yxHSU/yo2TcRndvMv5FJ55AyVjzAjraIg+pC7du4EUP1rC
+uhquywizznJvf8SPgMbYTl/3sarbPQKgYFIbmYisOzVglpQF9SKRg1XMrAEWEbS
PZKtY0sTD182LJvbV+B+iYPF9legWlA+Pifzw5+J3PDUIBw1UUj6OetbRhjAiVjZ
1GqSpOSrOWxHK+qEeZNLf/loxrG/B0nc1RSV2mJ8GstR3cUZEN9zIEQVylelgMy1
MP9QplcuffuEzDHsRlqVmW/W3b7eXb2r+BU8eUi9AWWrpSFJFDv2eaoqGK/j8R3a
vbu9ZRywJkIpa7Ng6d/r/eEnhNgfSvgMjb3afBhqPHP/df0hd5WRBAUij1lI5wQx
NxpibHBLfTh42ftbJqATgM4wco2tU0SnVqPY6voGoSucLiYuhIFqG+dIvTZtod2f
e1My1Cqh1ivRD0dKPVz3VkbLndkvPsUrgo9Gh4nQJ0X11sNuWIdy98db2zs0eOKk
3AZWBxBmuHGb+oqEMkB/zac19aTW4s4Y6OXQiKnAr7M=
`protect END_PROTECTED
