`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LzMLkrec2hq3hq4s1GtrZuYN9660An5EJl8Cy7GwV4ExM0dXVRO0X2sn3nRyRihm
Euhz2zNV5sN2e/c5uQGDnMmGc4UgOY7Ebq8KhrFPk8036C5aB+AXwgeySmf5soJn
WecwNY70G8Uo2rTvsVpfxH+IpWbD7DdlGPYm7YKTBupo3ZZjz1yOdIPOWPQZEQ9W
AgMWxubdygG+7Xp7p0BRsj/Ud2RofL25tvJrH+x5Azey0vTDrj1cHXkFTaTa9Ub+
yIG5nrv+lVfk6dRtCR2cEakJWxTAYTbH7bTfog2rb9vo6RhHK76Y3J/CCU/uPv3a
R0cQsrxBQGY7z69i25l8dVViObCsIh2TmhCb+f6wK812CTUFiv95f8wE2p3VIr+0
3/onTIbLKWzRaJZuVkGnD4MJ9sPmJlocIeUmxI4G2tE9RRXRrhwMSxYF3/Q0jcMn
s4bY47cn+/C/S7c/0CAeB3AaydqRph+V5UoV5elAjvWhO4x/npbsewrmrkthPEhD
koZHrkDhTFeubKep5/P+ZWqLzpod3YJEPvsRbsKli+swY9fT3hILoovD58V69Hvi
+Nrc+XyM5FG8G3pX7wrMSWKvN89dPSk4LK4a2JK1sG0BpJFZLmkQ+wu28v6YgpHD
Ac0TfdBsz7AEZDTT4m1bDn/pAoJshtLUNoW4xCGz06EuCIUubmUHPaB56T1eZaeh
SyxMwsWkzvZ9VV1c9zx+6h0p1QJmO08kwcJblHpOSQZfsBqM3JOqyVn1beABCSKf
y2EAirpEVXmZBVvFnz6H9H0vIFiMXWdReR6O10GyFgzrOakLpuFEv8R51W0SQbbc
vtTcmsexDXJ0PtYwFmumthxTg1dma4+WSllJf6WbYh6PYu/AYsBAsIYiqTVp17K+
dryq5o1gB3abtOphxKIiB7Vd9+GwcO8SqV8uO08rfhsMc1bbMpfeBr5ynTXrgvQw
cfaqNSCt5FjlRJjBk5un20R7o1VL+UV443m2Q10u0UDXvmgy7syn/g5GNdSbpizF
PyHgaUJUHdScENprHcZybRMV2m+o7kLQmIplOfct/BdbSbVs17SV772tW8a2NStv
8ze6Ac4mPb0N+wOPnq8qTrHd8QzJeAb70NVbuy1PosIgHhFnC14vFEU8nhhw6R9j
Yad9hS14+wL5tgU9Mo4DdLuBSHmWr01aTHhB4fg3oWV75iVwUCTvY4Qpz3hNgmqX
uh7+Rv22xElVzHDJy7Loj6uxQ8XTkZKqsuezKW76Gsw+PArSt2ET0ZPlrlIdBi9u
lxGKLnv+d1z8c4PgGuwLrE8FlgRrknxU+BnCISM7gKqo8US6/xH5RHIX0LYtF8ca
LuFCS/slT4/uyurxZ6JcIUstKV3yuWDyW2gxg6Rjaz9ajsSN2nCIv8umzTTOxgCu
LOqYdv95j92e7YNF4YTBQq5dn2I5GWrgeQP3ax1wPDrK1s6067qKlfl8Ci2wx/aB
4NmNH0a4tunmmJ/QYIInmg0rlA3/2hIsMLH5UfZKkdQL9i67oCXso0FUIzeLy7SG
`protect END_PROTECTED
