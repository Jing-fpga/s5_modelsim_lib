`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ld/frViYop1cK98ap4EQIfvThYoTzFquxOIVxpkqez3rCp1u0pTKOjbDx1Axa8DP
mAeJxQ28DLfZFhBhA1uZLTPEEqHfEyrO2sQxGsBe9FgCths3Qww6OFUafcC0JD5d
yNNzfM2ZmuOmr1DqTBVxZxKWV1Yz8Y1X7ho6b/nbLkrK2XATJd+wgsyVQlx1R/mr
UMpsVrTZyNP+PIH2eWG5+s0D1hwWIfFRC4XwPxcoU8ur38gMNk9ijBHKL3DV6dpY
PqDzS+kJ6nov0m4d6UnSgoHZ40znXhpq+uWqmxfKbGahWFVK7HMMvW5xX8jSDYD3
9mZEyzUP+mA+yuTRpYejNibxb2bS2z/pe1gfPDOZmqmSl5/gNvDbK1pEq9p/Xk28
+OT3GTOs8yx7hTKWp0wocVgAAYD3BwnDDkU6VJ3tzWcPTVc6G4AuBgrQJ31V6N+n
mjJsqNn6HgehC4Te0ZrCLTditO9cmFSXrjOucAMyOV4pd8TaD2W8tREnrmNZAQDK
qdDOhJ5pajYyaZyplAiGqtA026uFEmuzKBDTihkA9IN4u9lmNhZHNYsi8dj02Ug6
HgE6GSWrP/9WQIWSNoQLaKRKphwQY9lsl4hy/2FVgj4KDWSlb0spcTR1SGHFv3tt
0aYY6C9TgzNsIQJycSQhdxXUAU5XsBgDt9qOnslG7ZwNVvfCmuiOrMFCulFs/Fjp
T1ERxjHe82Xu/kC8JTEj0HrFPCoTFX5XkwVXI6htda3k81T/6R7khILGdsPRaUwn
/eagQYtmxOaUCraQey+7lmlaSFMPyFzjCGd8iTA9krsX0Ib3b4AorxACUZMi0Jmf
esyHmWryZ0U8ShEzhXxTGDdi4k+vS9ygHcO7/6San/I/nVMQMI8ZD/L8vbIvu9Aj
eh9WYPdktSuz8Rmf3FNEl6iU2gdHIsVwECiU3oIvjmwoS5murVOMnK5BgSDiplEk
4db5s/FQ3gKxEzfCZ8YIgHdETtkHqD95GY9+sN7At8o9jkqEMYHOSwa/4sAub2B7
1PBywDOKDYv808hI7OdsFxvJwKX2Q9Wo4AGblRGpuxQvy6cO37RtzAQ/3MbmWq5t
CeOWxXpkDyi+q6npLlpug3a+XTWTHUNPOzf4nHB+HezCQIfbF4TBzPnDue55EMm2
3UkpVL61reqdCBz8kKZmhu3m+2QhDjhTMNeOZi7d1MOwBS2xNgioTX3ebFoXwpGn
DqZV8Zffl+PHpSy1WFl43iOdnw8Er/D542bf8zZ2bI/8NxHDdH8EeZidQ2U/NxW3
`protect END_PROTECTED
