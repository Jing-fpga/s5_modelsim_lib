`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q5ne3f/snlWCvUQPtc+iZaiU0GkuDQGOgpdxgg0gyO45cYTHoETsD9SQZooy0nv2
ADHAZXJWeLlH3nmNqzze0qanN9rL8q+HPHokTIKxnmuQk2INPbDWEG5qlxrAJFJO
3GyRsI/0pGwDfbIJZacVi/ZEg98tp1/J/cx53FkLg+qdUVbd0Z4rBrIxEynsMzaZ
g/n/M/oFf2Q2QfeetYi36RLkcM9HE80t3xgm3He7UGQWMGi1ISxFcAEOGvc6wRnk
d56fr4mndTgGkTXXpgj7AlqqvWi9j2hEgvpLg8c8dt5Yql+4JQSIqDm//PSeiRDM
ELXBZXnDG+XsIKBKyGe1T9zriRG3lWXTykq3ITsT61XtcMAqgYa14TiAipwnhyEz
6ixXe4dAWq2bSY6Bm0R4fTjbkKDgRjQ/6ZWTEhVN7Oolay0c0C+X8aTqH1ytc1/M
aRKBkHfXQrcMHL80LXT1vOmkBWEOXddac0CaJreZRUe9o3o2viOKmlo5vXmJylpC
m3Tfsmtk0nt2o47D0+l1S+W7M9enGmCqFfMiTeJ1KYUHtiOowDSJ5WaIygGuhU/A
40+a5elc9/aWSDEE4W85qb8BXkAUTtj+Bj5BpZwMwlBG4iRHfI1w822yOaDISOai
PDKp3lRoaKG/CUW0FrjensYbqY1Ro3ed2YBe2qlBEOkyAxBrTnDWWzc/0P/52a3S
6mSITAOxfc4y4hNNynf1IPk1U5l+zFDCiN2dsjTR1YWebCX9KA0RFENDw0zszzu+
eol3vQtuujJTm8LUAcZ/g7l9OgVm3y9fN8uOeyBpntzN1XOFEFbNQ1CMATjCfbkZ
7qvHBhNkgYn0ts91Jo8Ut4r/vMykEQEDtSsPzPu2FQDs3EqzXR+x6MAa4jXnO27K
Ubc0w/RZXnl3gF0P2/5ysCXTsxlf040wY8WUe4r0hmD6AdR9rWS0487YqC7dOBGj
Mlx1dcABYPHa0TgBrfscsA80NWURuulgrcBdxSMvT/wCWaHnpiCVcIhLLkD9qmHM
uAeDHE68zyxD7nCwpwm8GoRVHLS/J10Xri3b3nVaVVwvq2yddsmlNskyKoactPvD
afDmzN1tF9JQld6Ez6+Fiawnwc99o9EbtdX1HqCsiInGMiu9h/1KD3VwIi9DYHo8
nnt3Fld7KOsrJ27tZ+GIhyyKJblZdv62THAHtm8pj8odbGCC5YzCZbkfqkApNMCe
C7okoYoD8uLmbvhpJX2GWtyWUVlh3uNh5dDDl5NMLgox2MC2uIa9Z6DEJYoL46Ut
9gKOH3fGZzxZIeBVkzllCxydFfj3N1x5/dvxn51RPvjbTDHS1cFvJBvsWwj226H+
fmL9cCa1CPI1N1XKTChnpSEzKRoFqsGF6Bdw9sF2aU1pJtMDrJXqvRsgNg1uM9BH
7Nkuy3Yvpb/vnMQPtUA5WodGs0DDQXqpriR5dYlHXkTQafpTOgGMRTXb0sNZNzMP
kcq5+mXcLFh9rePT4yeI0D6xO5ttyQNAiM2PHxnGgcc=
`protect END_PROTECTED
