`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BQE7Tyns7lE7gLwpym1Wtvc2tOM9DAjaPGx53cPRZrNWvg0RGmkZNh9nte9MuE9k
Rs8BnSte0gf+6OqlQWj2HaUKqLcdDNJUP6Jp7FSh9KiysOvmL11moGiLBWykC1h7
HvemePZn8BwuqYZWWcL7MRWzwbeRkXQ6+Ep2PitYdq3CZZsm/HLBgi50zxmyaa54
v+Y5p/YTq6kBZHxTpufTCJ3/7H+dLxyBRAdL8B6ABe7NIiAghB9eDabHMzmQOK8C
CupXwsmXCWg424Gnjhf7IbSaG7ZXEJVbonVCdzb98AlUvGqthFX7U608crFxYOze
VkEllZD2LEkHtH03uJIzfLE07zRjjA8IRA/j7NnHBT7cy1fLRA8YvIx4tCU3ku58
NClB/U+z1JalziaEtGXoaxp/Q0WBm4KbFcoeNZaznNSIV4m1XKzS/JDPoMQp6UO3
zRZPYtcdKlzfwJaDGHeOh8Anwm/Gr+VYpKKj+XSup4dqXRgKEcjmEbTOChuPIwk5
zji4m1A8ux2LdbpetUC94mqzVAJ8rb0TqD72A08Ee3gZinlXwDkN3XAR/E+GQ0qR
fOi+Zj1G9ZK29VusEiUDsBQYN8Yv5PemIjnFwEoOqDwXMo3RS0xqswiRW8J67kfD
sljbYY3gZnmMGAN+ptzaV/IdMK8TPSVsBAfCTnmjYma+olkxh2jhAFH16HMD3bzf
mw/79Ts5O2uY5gdFCV7FcY6h8GS37CFbw9G63KT61DFjl0cF+b7T8S6wdAhDQe3b
4/R73Mbvayhvw4WoQDXSfypCPjPLryVtalkbkc1CyiITbxuXBuN1bSM2sPH+wC4E
clnmhM5OOBKG0vZZcm1+BF0r1P0zTapEdJP3KxJ4eOpCmzUv3jTqRoaySx1emsWb
w8oBRsi1DHXtEralHanU8U4qbthXS57Vs3wZzqJmkj0OV0kMEnwjWk7iGVBAoBAV
K4W4NP86DNIr3nX0HuhY9d7tRzmSt6jkQpToOVXHm4XCDoJvDd30lgKA0QaHyl4c
FezWxM3GLDKuJuYxiuoN5ohiZv54Uu1rn3DWpM3nEw9L2sY4mOX0mjjVICoPVe/x
AfG5pD1xnXsfzbz9t41rLoZK7/a2uMymTFEhIWRdrG/QY4wBcJtKBJdEyke7wSwA
`protect END_PROTECTED
