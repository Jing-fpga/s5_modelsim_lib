`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f/Kp/IWyaj8z72/8QxzBdjVGflWQiGLbE8Y2OHhMZ5sAHb6dvOwnrxpL+fFI48Gk
tLKd6MSY7mdmogZHlPDeIGoXSmnv7L8Odh2hvQWnwCcy6AmR9Canix6eK7D+A9F7
xBeneWdJONlCI73WVklygjL5H3P6n/dKxnodOBvYEkSMIP5P5Mpj4ZnKCWGCcFy3
TB5mJ43Qvl3Q3UXZDwR2glg/LXToOd4dHJITtyL/uPN5fSkvNzPueOnBUbUKZhfJ
S1KNLwkS8a+qguo4CJCnxdJe5NBYJt1qMi4GCmFQvv97BG84aWWnmL2pDLCOQOS3
VpZvr9+lbeWysAVJefq61XdHDttOla/8qx11rUdrgAhElmoVpQaaUCL9JGpw3xu3
DHXhgyn0ygjcc731SodFsAjk1L/F6j0Zur+rQhgyIPOXagcNdKnIMDhgz2T86fdj
rNaUnn+y6GLkd5YH6tSVcCgOeQBbeMioIQId5JhS+SERcGYzIlWtOXSfNi7Pr8hN
NrrMdAwfJhzEnx+N8AFrqk9vHUBLP9XvWZdR1cxt75gUIyfpqQ5FctSIwosBnwWm
5pg4zrf3Mh4m77kqVht/990gXnfj1A9U19xi0CdtTi4a3hCZl9Q/vvZreoye2JlO
AmGSJLu6Wt3H30H9Aw3BraHroUoiMFv+LqhUtPLI9xzqrpltTW+Cb2wo6qDJb88c
UWoinagT7KAiw7Q9z/fSlzpMN2k/OohdXAc+tb2U86U6bQaiWuZj/Tw80LAMTivB
GLXwtKMgKOYT3/ccW7zfsc0NH7U0rhSL9ZbH9suFO05Y1V0uEzyJ9gJL2WcmUeka
2BuV8bpPeBTepxJx3vvUIXnaQ5CPyRdMX9BeI+IB8j/NJz8jrne6yQ2RI4xX0Vko
hm91rtnFZkdo7UhDVMiKkhFNFZE6arzXaEaEFts7Y93lbFVCAC4yQw8pDSGb7GUV
+c00+XKIoOOByhaVuIMykSdGlS6gvidvIpLIsk9ZCv72Vseap6wckSPCoJ9JX5Ui
6soqmrqelIniN14lfMcIGRz/Ami+VYSwkw3tTPSCSTHPfaJrYVNDmmD4ETSczURu
j2YMm7yB65sGXrd9/GnmaJ7BMUgfboedx8JdF9CnlU3AXCeNidLn8ixljuGgI+HH
t9mV/2OsQG0g4KldRkypagK0wIixDYZgUn/7WsxNvaBNWmBVxlcJtQwWudMljGO7
0OEKlwIn1gycOKem3ic54w==
`protect END_PROTECTED
