`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GGt6v65Av1CtLTyJim7JGwOdalryibxm4XseSkhY8Xv4H3wx4U9FL95vR0FG020A
seMDUzr5MXAYzadlOU87EscavU+ilucGT7jXPvO3o+gB6wdOlTwcrc7RwaXpqtr5
zYYm6UlSx9zrq+7ED3YsKlvtXhGDugPT95+mIM8KLV+5a7TV+wDik0I73vGmuCrS
IGg2pauwxpqlOxUYnrci4FgzXcWQ/HpCKCXejTvzy7BZXepoNR6FkcaaYcaf5noW
BXJltnSEcExpQ/eVsJKRe9Vzpgdh7FKyff6LUilfslWGriKuk3qd1oFM5FLrBMaA
iGrBKzLCg6qR/b3LLAuUB+ogLobYU3ySVtlqpuBRuO5TURgQSWuBIVrvFsYObeOZ
NNe27A3ECYrkM3M65Rttu8QuzKc9YywQpENMv0M0C12wQklXYfgXkSER0PnYmAN2
fhbJNiYK/CX6v7AX2iFXgJrdAppGZdwzJhy2YDlLccARmIXnhFLOpLC+fuhCdXyy
zWYyksc5T7IonqPGwC/lPMCtz5wyqhP6VhylgV5Bl4P7ddRBAZfLM/daAVP+WLYo
W2pyJ6tVJdzz1ncJApidK3jOrTNLEyrWHF9Qz08D+VtuxaByYjR/EnS6lw9i6ZQY
psNb+16oNdPLCUQ7zE8586bmM2bQebCG3RZzElnVko/+kWKTZVYbzlJ40MlWaRxF
i8CbHpmkfo/GUvIkhJZrFd7G0eGiDKtoOPvcd6gIy3wjW7PkxltUxL1x1ej8wnqg
pT10+c0mM12UOZYUHlAlYbiaZXnHeVAiFtKY1dm04JBH+q21BfKfBY+9IytvtT3d
nsgf9CGcDmme2WMQc937ig==
`protect END_PROTECTED
