`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0FxAICeFusvFdNpxUIxLzTfpAnukXlgWEgcCxwOpJpKnBPBUaSBazr+gcSLwh803
F7ozP32CSdIU56nlgpVdom2LMK/U834yglbTJHuoKekhPx8lM42+MsXrIo9Xz580
LPbg3zt0a+6d6ywY/JuNXqube7Iho+RRB3qNUga0exvazTuuj0TfVb7btBjIdWiH
F6FmOOiW17xj30J/7exNI41TUWBCn9ytQF1oTlVI9h3NPrdvutASfF1BZbHUoVTR
Mh51ZGBcfWofs3h9YEzkFG7+a+m215ykPIaRVtVG5syPj07k4Y1VpZ82PMUVaBzx
JQopxrZ/wOa+1V58rwj+XMiuyTQFygNbXouqTjd+7+MK0nQSeypSKPcAJoJtmA79
NZavasDU/JLtS52go3kThSzVwAU1038DcumtnnZa6YXkUGIyo/5evEGvcHlMW2lR
eMDgKK9ShWIhG75l5KSm8l/ZZIFP9uyorwuaEuaK3suTDfzRS9alJaQYo2SEHvla
XVyh4trq7DNmqoHyPAZzwMfzFw84WidbYW+7pm5WurS8wvKeTJZGCS/Y7EhPBVhG
9FHIxE5ISCsgzgqtQzTW2zEZBtjMZ61FmdfmqCQO3dj0FQjqRHLdNcELyw64++03
9u0UNWOdFeA3bF9RqQ9GG3lQmb8L3ZClNK/I0gAcvkBaM0e+MrfmSUEd3HI9CTNJ
saZKyc4At3o9wnzwXbQFQdarwnK+HvbZ8Xc3rArse7gujLJjalLc7OhFBKpwy4bz
HwWx/fwGUZcRnwG6L89yeb7qfHhxXIQpJliMW5Z8NLhkndxxcRLss4QA3+lvVsaX
+cQl0UeNq1neNQAln+5XdMu45CpIRRmFcBjZYBwpzLlFPH+u9HDySjimdbDfUf5h
nbIJuys9VNCzEDM+PT1LFveZ106TYlDAjb0t0lNkI8SUc1FQqbvOkU5Us+IGoDnU
99jtk+eaHncuQq+NrKPLvYqWhEtfKfeX6VfxutWmJO8=
`protect END_PROTECTED
