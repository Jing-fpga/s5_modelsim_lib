`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ouRAJLiB0B8vUVld9HR4bEMmM/WNw6elTj8LecdT+0PqD3Mv380ES9xBa6o41nG
ZcN7zuMlBQtbwm+h+BYB4nF1BmkyNZdty6ygRnO9MsljzxHkywQsSspQh3HfDpd+
NuuVJTAySzigc2yKhcjcCVT+Q6BHIL6fbRmXcTQaySklcGnV2CnkWiikwCrWnUZP
/cePAQxSbgkS6/m3L3fHhs927wGkVoU+bJwuxk0TzDk9Tluu1HuA4oYLjR2JCAiU
vCRdSpyDtUAYLXiGrbx0ahxb4Wg8SFe4x8rPZ+qyQlOnAdivEXTovw/BB+RubsL+
Ld4AbdfqOswRzp4fDJBc9hXZPmyVR0/4yBF/4O+85Ln+ttSgvimcaqtJ+wF6DK2n
ziUlosNAsiBYunnKE8fhM4p119pTre3OqFYiyxgjOqcrDxtp1pb3Vg7K+j6z+2+j
CpwsRzrzWQaUc0nc5MCMgaQ0oJbRFCeQHY6oplB9zniSV7A/axgt3II6bXriK8bp
cPKn3I3eNHCgYouo71jDECQ0IIVq+MTQI7WaOv6DtES2WZnHE2dpEF4NxxV919pI
aSKv0EmQanViZ3C73IVwXMpSjQh/Lt5VZa7qWcgBFnaNOvCeKhlqB9hgI0lm/IPF
oxDf8jHFFhhIz+WCoCYqhlAOT2CCEG4boXAsGiqnutq0ScrEjJDNDrd+HXnYiaXy
yFo3zk0lFfDv7S8tu41Ef80YmWchUIb4yjLz9eaiaZYedNTv0VDibhRdoVNf3Q+q
/vavK1TxrcQAFx/SsbsoYF5U7eLT9QyEJa0xn6sWK7DfUifCiCRGKlPblYqIxyvs
jzM/ze18YyebhJfdD0hJG7mkptHLEeZmLDYgOuTTAUd0RDxmCl4OiniWkYPcFzwG
Fgv3mC6cpWaAIjQKKjwLXNJjLsNMA6tYyNANeYt+yZFOLdMfttFaOel+bm74I6Ck
Gttcapl/xoWuXDjzAlopbvOzBWVJCfyRP5fdRE02no1UjJ3vAzpNdh3qOSgSjADq
RsoFl16I7tWbzXqa2bihf9J46rhOaurITBWfPf5WGoxVElQgqaZtMAuedfJhD3Wp
vedLFQtRfF5aZsyvr6I57Pe+1ajNqUEO09TP0kl3j97sFScev5y/EcGUE37wr7LE
1Q1+0rugUDN/opwW6NXzzp+RrK+cw/qAGDWZzxrV2ndy+eR7pESoqa8RxFZR+tIL
+ml+3Mu7/ziBo/+I76hJhhcYN7U17SKTUwQm2J09Z09PuPZG5e1LNJKGxVPm8iu0
X+LLYfZEYKRMlhYw8MKhXe5cGOKcad2v5xXMdQGxVLI5AA1WkjDaJDVTpMC9uza+
6VbFTzh53lmqUqd7B5V2lASrxFPtOY/TXeyhoCpkjFA5U1/r9bnkE6u4kHXSofi+
CkPigD1lkyjNUmkoWbsgKlthW/FXMlgLHrWdhUWR7lAZl59NpY95ENZYUw5KnOps
g2x1Pwsd+//T1KolDuL16u/+JYOg2R/jwILgTyycFvkbN48FhEqCB14qRqqluGGY
XLcH9jBl0DIB1WtU+0R+MGMOQCdVaEIsxxCXD551S/QneLCKIVe6Ymm/7/lpUQjs
DMP7RqIMyM9GKOGr/mlOAMMFNH/nFamojBURaeIuCVfAimoXzPVbyyTeI2EnIFFd
YE7TagVi55JoHKI59nFdt6x1CJZZ635Q5NpK+LsrNyS32zDg8Ec6OvTyrnlNDzL1
Xdq7Bj9UJww+3jKXNZACirPW/gFNYOVKx4JkQdkfg9b+/w85HuOPRjGN+sZ8FbE9
wOIj5B9kIEAaVnWKdn6YQBr6W0/Q3e5ePSOkybV0R1XxhRC4OCliHXUEkvpiT6do
Z76ElvGD/KE4oUFG4suRsI+9kXsBc4iDyR1/seFty0PhwmchgCWoEc52/3WF3fr4
vf2cDSOL1lZPhTBv8oUEa6HU8OaTTwzV5UUJbaxNEmUX5FatfputA14Qwf53QlWD
ShO1uCw7U6jth3U7M/NcrnICyDCkeUOU2rrQ2G1rCS9b7DxZvBPo6MtjfCSwN2bR
QE6YDqYfJbyhc5gajevGv1ba+AqaKtPKTqaggh3EQK071UoPSjh46j1p5+eUQdRF
8xv4PXRqAtJVNRpLZAGN1VhxQJu4ETuyrcxXbGiBBUMjH9/YVljz+0sqaPc+n8Iw
pi1VN1jFgtvAouAg92AYE/e3GzFMqGnzbHqwShn5Q0ZdMxgpC6OglcHrYm3khi8Q
C6MvF4NYlM619/nckxS9nB0/zaLw/jos4I60bRlFsKoSKSJfu0DITGofRApiX9jK
JbBq3fkHmwza/SdEFkH6VzciF8ZBzgum5+eSSLfPPj0rdUwBJ1QxXgVXqkREFsIp
HNv3fki+tYFqkaeQcOivJIXBY+EIQ7tQSZtoCFISvbxAlsVngww5eLa4nLV3tL2U
zQYCDBhIxtcqf3iw/K9/M+cziu6EpG7rmOnxaU1OFxJUUMl6goDKrJJVbvX+n768
2NkV16MrAKKXi6dN/L7sL95ngW+Hhib0cYmIuAipREiD6wHrVHmcjI1b7Nn6LtxU
bnQSEuU9vsuUTeYimQEDdkt09H9T1bKjw8LinkFkGFd4ssx/9i1rC3f6DWq1RKop
UEpjZVtZvHn5EWKFD+HRoe+wB5GaHlOXwlFcf2AwtlGeQLCLqmeAcKOUUvfv2KjX
Oi0i3hNlabjhlcs2LfR9f/JflRrkzS3UezcY8FeA7eceYxjm+RnT/47weBVjzcr+
fJ4RIK25pEmucNxQp1S1PbpKmzHZ9RM00F/vdvcYirbS4HpShRq8WJze0y25vhYe
8uRPpuO2O78wRvZDQQ6jYa/irquloozBhR8vwj6I3+NRMC0YwoDwczryA3ePHjor
q/lpoGxsplIhv8amWdLPrgCiRl2B7TX+YvXNoz9ANd9aykcUnfMiqL+775uRs16U
va1QX8Yh7Ummd0iE+u1cu78lUaa9vrjk9S1e/YvDREM=
`protect END_PROTECTED
