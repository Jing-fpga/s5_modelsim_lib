`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7WVKaYmDKG5ji+ufSn0jemMcbjpEKxc+jqrYLfdpqaBAaWPFsteLN50MKyDC4Nm9
+oA8WbF+yFBxXz7Id9XQj45wLgT+8N4NzKPOcy29UDmkBn29cl2+LsGIkAamsHNY
9cZb7nGWT+K3Mjacb+VFzPk+f5hj/InFjNZOUGkhYIxPxW5NiFZcmimycQsOMsrT
vtsE9JL3Sb5LPqcE9atZcAj235wi93DhXi224kSGmdZi3IKddj+b9JKhu3e6Dg8j
Tq9VsUTB9MtrJ+kMCb+/BX5RxQnmxLZRM6hRL3bK9Kvwd/L+j299VaEaHcn9f2HI
q/ScccIwI5bxLjXr6az1kc6egzRh64E0uS5tByZckxEgKwU6fIizL5OY/Rhz4x3S
bgMUl/dmcG01BDhrT2wflJZYXHemG+FZ3k2Kgn/wz9/qzyiI41582tJh94mFO05d
Y272Dd4b44G81mfZxo71vKmfNQT9QBepwz7p+lyDB/V2DsHezEoZIh5zYdDi8386
HAwplKhpqHq6AHWszf0JQafI+5jos+5ISbGFm5Yy2dOX/nKdVjHyvhUsATTYtOpV
EQ2aR5/wS+yvK7zGzZyqwMPFlf6PWEgFTUWPVIDg+8f+2FwkJ0eBBcKq+79bYR1d
9wM4k+mDnpkeNLdi5KqHm2EHMXdm6Ymd6Z2CSYqKjY035jBFGDhPxNZiK+VHyxhU
T7R+anpoPGhvSogP2+sfG/9Nk2qvLTqZ1a2byPESQKG9FHjGzBihgJF3boIKKTbt
E5nzHY9gBosSJmnnAYtL6X1m7/WJViqdjDzm5VK1LU7D/1aoyJQx9ksIjTX7jSAZ
0cJDqlbKUTu8JvNfwFZFDGL2aFb4WdOICOrz+PphWiOnt0mAhq+tK4jPwcCJkBT9
Fr61xcQ7lHNqIrIcyGjb4zozWk8pDZWVVN4Wde6FxhtapvWtbk9UTNDtKYGfIHal
EkLRkR+V3YvpDYnkkv38xVnTkJEgE0fVGbNhSWUr7AEVZhcZhBwa2dfokkQIr1k5
swHENzWtd0K7mJj44xrgN++qkHo8qtUAwKOKKdBUpaevsK2RleXIEKAa7n8jKXBa
JILjrh+P/tFXdIbG2HELf6mW2T4JFWqftDd0ChlYn5r2qmuyg2cYTrqvXnvrbDaw
Vj5igZ1JW6Te/s8SUEceMrC3GH6Zc1dT/LkY1O518v4CneFjrJzI2laRP6YVCEUS
+v4Upz40ShxECROgOv2ijHSwN1af+NhZDR2wr2IWVxJLaQnklaxlB3QE6fRkUtFc
PkLjuGwSGO+8ONChu+H+Ymqy5zcXqsnUmedS36/rdWiFDhbKsblg0A8UpiIyOlrD
Pj0+Ggotzna4LuCBu5ZHKxNUjFM9uMes8kx6R1nkJP4fAlGUwCKbvrYZE2QTc3aW
fFF+MUaLvh2OJhkQOlS0ar1239ODLRdIqWfiHxy6ZgmKNLt2JJtZkr610cBDvX4F
DGMCpNMqPVaLLFRoOOVZOQRwIUNDBCZadUGv9ikAUR87wAZrkTxFp08Z8LFUfF55
NoljV/9OrvrUgEFmY1+TP5XF+81iY+hdbmwqbyWq/qx6IgpAKAdBpxhdehbPLjAZ
B3F6hLt0CkJ+hfAeBZji+ChJbZhYe2nMbvGYYJ1PTu6CUrmLMES6d8gv9NZOjf/4
G2e/DjygV33zrYsByr4UjUrFn5nMRIC4TJGQy+gnBv2NX3jpiznzFlahH/Sg5lgg
hVyFGH7gVxdMq9GBeD3JChhp7xWJ/BDEDhh0PXqN7DvgDQFnNbr5QU6VhK57MAVq
pwMBJTwbSWDpGh5socrWj5eEamOxw9JbcSrTw2M3Aleg79urZ3slvVhLdcJE6HCq
9E0kDWp4CWOHRMzLCLce12BguF12EwGf3rHucyj6X6RSMJ6AwiMEERp4Y55N0nfI
q0WOb70H31Xgm9VxA31PY98t5KKfPMUOzkqrBuLZmKnF2rFr8zyDD1NBM7DIE0yU
sf4KHVBRXurlnsp6wDs9F6WsdnIxHyC0XMUvsYWLJsdtnFOWIgIe2m6hgMja4ifq
p2vIhkRiW9lQ2Fqv+LnSWcrQH5LXQNiCazKU//9plWalB9uYTcRmaL8t/kaKwi3A
4Udlmr2iGs3BY5iZCCcl7csWVVQCRAErjQe8f5T5wq1STCx+y+bzFiX1kkq+lUgi
OSJ2NP9NYiKaLA2CKJrie6+SkrbYXjzxJuUF4a1f4Eri7c9ml1nEd4WGTCSYD00B
o3rz1ziufo7rbTBDkOcFR7Y+NqBzDN5x+UsPqc0oYK3VoH0XWNvN2bKCrEiqxO7+
FsoDmePu9Rjs10U1ypjcU1AfSwqdJiHY1cPqrenJN5mwrupEZ9vtriO2JRnMzQ4j
RUFK5FoO4K6z3C8YJ1QsMAFu3+zcxR1LWPA1w90fX3eQt/Hv449axlEIE+iFBfyL
RNgiPBdpi+ah74LTlB3veL3sXIdsFO8dYSyyGs29qOkebGy1YDvuRQzDKUWLVZaU
tDT8IqHBYDn+S3SlZfh32GytlACqCC/6K0ru+lKkgXOaPWqelyIOGfJMiIpx6U9q
XyPuwhmesYo2hB3bMhlgEPZPrS8JRPgFPHz8nh11AUKkyhu3WioibIbum35upO0y
vUec2jXSSINlD/MBqmljRBJSIJwWEldesN4/1wj2SGoUHv9z6/D/un8PxQLWLEGp
OB46XXg2meKObTPejO0CbdaQL+eMoX5CTjiT72h8O3oyb+u8OmAbJYjOohlYqrdu
FovZQXJGvmyyVOvVAOOcdfZUYIW9x/narLpovTQ2TzqUA/WHvPpcBdjdo9xBn44f
hrK74zdU73GD9qkc2KPEKpEMqkUWomPDNnrSGblAOUsQcgQ/xPCQz4XxcxngUffe
gAlkS73+QSvfhVTm4+SDzgKv9KooSfUVAbdWzTYHoJ0l1+0Kxvnio4ANvYQ1U3fi
laiTXHNpouc8oyUnzsFMohyQp7EpP+pZHzeiETEJnePHT4go4OnDCMjaHBFU1Kgj
KYu+fSk79rDWRn4d5wZnjESHW4vOdBaS71Xjn2XXg9GSYmxV9hlWEi2lEoAeA+lC
ReRyoCYJFudVCuU/Svu8B1ayvbBcZymVMRL/ls9b7yZgtRBQZa3//2Sg/hP9RxJV
eVY6Q6rtrFYNFdPKbYe1+Bsk1z3k5ySoUNylzzz2znoPRyxb0aXbswjLTeHhPxkF
QzceDmTwHY4Mur36iHmHXGG7VsAfPnDPEdBMqLhCVAtEpm75ICIdiLTZoRpeGWNw
DvRFHpfitMq6XI3e2u69SU8yqT8dAkCbLx1vy9cDqV24kZoUc97Ci++YmiPnmId1
hqe39gns7YrfB+rEVDGZjwglyWbx+O5xHasm20/wGK1titVUABL+JYkIS5CJe1qd
foeO2UGMvY9b6tRjo+tNwN9yO8uiNAFLsu+c7U0vI4VngV34dZRVuhf2Box/YxvX
BB1HiGEqU9SYaMV6PaRVSO9Eh8/LeEjYCGCyWpLQAvgQZ5QhKAgvHOixX44Mq43l
kolAkdHlKgkouO33CJZpFVFcoqA4jETsulMgTD7Jiux3cSeUAfpu2qTNEmkruV21
/fyNuX768Ll8XI4+Fmhs0d2AqRr8qMOMmkYFfNPOy04NWVgQBuyIM6H8/M2apqhf
2v1j2JLTMed12u3RpGUdiwRjzlLuY4e90bdsYOE2R/y0ZpZ3Hv4yHH1tYErrgF6Q
DgtYsJvkBd3Dj68C8BKZ82OwEtSAtqEiW7u6/E2tZbDGd059+G9xqCKeP2Vw/xaD
8JyXinMDT0Xu5PM0xi1U9nyV7YbEtzpAPgISFK5SMjHoxWTn4wYQJDbJwfWZHGNN
on0VhuZM9togYE+bs38LpeUMhoJ0UQ7opD3ZrKer92+J++c9m57uy6CrT3dXl0S4
Caubs1vA0bBeaQmGwXovjgiHOs0A3P0sFiwyuST5RxqVeilGWuzWoBrKgztAk7J/
2uqLb+MAE4NcEUMql0P3JGq9ESu0ul0QQ4GNDGgIjT5CP1upE0AYc9ryp4uXy/73
QqIRiGIyB/4MPlDg1CW2Shhav3P8aQcLdBXtCh3jdM65ct1L9YNgRLGQQh/OBbuM
TCEaD1WWqsPb4WZLTW9lRHa3x6220Wdl4Xl+DbBXXxgmHdzUNObuizh2iMzLkQ/+
Uz31LkHmsRFlZHOGLIArT3Wcjs9zBvoGWNFnQ9Rs948ZDhB17myyqCp+2vjSS5Bp
YLo6xLoypFPyRB1d20NFhOLrI2xYIh4p/8NSb1kDMWvxs+syyao6NLzo1oNTHELp
8aQSU98flHhu9n1s9EjV4fiJongZ+ypCYGA7Svwp+5L9s4qYPzKATvpAdw89NBKt
TozwMfnE+4oBvK80pIBxv1Jvh8lNhmMuKCnRGT6GY8xpLYk5uuaYVQym+4T0/DOo
bQCtcbBnpOeJfrJ3GIGG90dHtw9hS38ijT1RzhHNbuEd/jAo+7WQetLTuijLnVAl
EHMUwW0xmeoP7tppnL9oQWriU6ocT0mvhXfO6k9DBY781Sgp3+24Sjcr4dIICL8n
EwwxMv6yZIZXinPQM7ziE+nZFBjUGD0T3IfRjppnZbhoFS57rLVIDVoPJDIkmnv2
m2panSqTBm9zS/HqSlaOPbXPy5txAjioqTA27s7CLDWSUTpqIHYm7BOq7TDoJefl
oVBU37duIF+pP+qDI3GGIwVmcQlVQtaG0+nE04l1F3ZHWWOpCtC4vP/WTYs4nL/l
fXE+FrStqQPYluyp8iXYpadGWW3m/1BjFBUGgt8EyYDWGLjlX1pLwWbO8lP1MGvI
8O7d+x+1LmqI8hcTBhxjqCQjSvdNpeo2WJQ3+3LxT2kkOweqNAV5F5hbohec0KUD
HcmjZvkhS53T9ISMHrPiiYFA86Lj3KWGsWQx6lDHnSemiDyXkbcKxg3Ks4f9pYPc
Wah25tp2kUOOcklAY7Cg7RwueSEO8BSflS38yU0aVXR8YiYnXmfgo+jlMZ8KORsw
mghvF7MXK4ucNrQrnjA8k3ckhQRF5kWRi032c6yFwr2VaANobCAEQAkgg8meTN/0
BErZo5mJzAak9LqguBqfuu+P+APUnd5L+mDG67kVKVV5vTNVz/gmBIiyUr5O1yLQ
GsQxhbHC9lj+mUVfI/B+kZ6TpftJFcgcrtJV5TIcnP47JE+r8asZLzom953wn7l8
xbyN6WOrJNbUomhyTk15YL9PD+DtO0FAPPBppNawsWCMBgx8MxrzuZCuX8KjnOL7
obgmrYLz661YbvsOJ3JEek1rOdev3scKtBzpX38ikZdnVhEUj6W+Uw1/OE5dRI86
mLoLPrX6ARyiGbOFtnxwHFeDzxVhIFMvtE7dMItkbjEeuODc0u8PrUMfwbF5mwoL
YY1a9sgX580FKw664C6IJQD+P8a1ViZ95OOVoDdmF/lIcqYElvwltkJhSQxYujBX
UzhToFKNmfwYjmVz2+WdoPr2EQwz+uiefW2cc5J0Z0M9VqI3GAxMmXW0O3JD91vf
ETtc9mUjPm2C/Tvmdnku0OhnqOjFtQsM5VWRLWz/JKxKI5AuNWjCAxH7UTcOyQJo
oexAwr5wvNTEAJgjp5ELiRfh4BsN0v7SswDvGmUwfY3QSweETSSz+zNSS2mAAaxK
52EOiDmi7j7e4OzW99LeQnJbO1l7s01deHf8rDxMYTqe9fAp95aVJPOjSB4YkBKy
8K/ZdYzYLj+8R8OMnO6J347eh52PjjGLgqh65d8U4ls2FysolVkFQjMa/hKjGAPu
+0K1gq0y8WJQ/6acNdH+Fyqd0Qxuq6L8M99VzYGZn1zbsBtM3JmdvuzLlOcIFksb
mn3tVJbo4QsbfbHdh7gt2E+SX9iszTU7qoOTLBJPelgGKne5NsmKqebSZEwn/BaE
5DFnvqT61DjQQk0qSZL8ppW7Gl5AwyYoFD8isIDlUVZgVElrLveSYzps3g95ogzR
USF2EITDESe/SThN6lFlLCVqZlBcaMelnHe7z+SdHaFvn+uHPUtzyjNMlApNzyqG
rrx0oUaYZWZZ/B5pcWrn5fFvt/fOyCmsP2IpdvralZ6nnJWZIBNd0e7ujXDJ9Sag
I1vnaOzWmJneaD/4JWI6zf7a2ML9zKi793rxpK1tKpt7v9JwtGFkCjknvtPDmNqy
1O1cxsVIZZwWhW8veKss9+4YHjsLyPVZ2u5pWdhy/xE4rNvjK0x9uc6xCxmxHvyl
yzd8OQcMfuvNT7auRMRn+2WOai//9MQavmSeZVmJ8cgoRzlzk2MTb2zfE8qlSNKb
cJOzNx9JxdTx+uSFmJc2sRqCW1+ODnYA7PnTxX8+uRLltydNQW+WINKr81NTAmbh
0ksJSZL2q5ijI8I7BVdsr3rqYwosXgN/CWPwyU/Cm6raWl30NDCpHrpFEj92ULIf
8an1/MrM7+com0c2hBKj0s5UOuZdZ2lcz0FbW+bMzvD5CT0PRlFLcZ+jlyMB37U/
iE3ySJS3DhIiansr5utzFWP+nAyWlA9I/1qXS7SfKEwIhXj5ElNk4C03H3LJhP93
yqtRHDYMQOuPvtODVuZUVLeYPojDHcms9v4Uu58/RZ7qMZo99n5E4tDPQkVerj6E
bITDibmJub6JQuWt0oanGziTbzunehB2hofDwC+Mgm7Z0gjvxZu/HSHxG9WGbZRk
Twm10M/i9ptOvm/6wznbmbCKnGn4gaYybIi8YXUL8hmKkYRxx+22ZqFO5nl7Qsur
DeXOOMU3FReDliqP2mMyMF50zPNZE8smawZsDX7SuvlSFCixXDa9bJgUQ0qB71QO
a+QG3DEyOfN+9alUK+5CJX5jaQApeKmeGv0enoR/fY1z3TYV7u2GjoT8B2tUsFvN
lhuPLtflWntzH2z5v6qYJ67RQQp+vrClCelvR3kfTmDnqVWt1YSgJ8rXZJpK/trv
a83qtG6A06pJV/k6Ena1muxFKytO/oYTL+MrJO2Y0KhwnCAoCKLyaWoKVP/29qtT
aFJIl36fLT11sUMmIHvtOe7aqAsSB/sLCWKlh69wMzny2MLNjWkIAdO5+xw0j6au
umK8qO0DYNOL269JZMajXaPkhi+G0t6XReOenfpT0+L7IWdas7S+B8sNOQAni/Wh
yYl6x7yKYEKuIPcGnqiYEr0nMd897mwFy1QNjJoi2azikkdGBok14VjFsBuguOGL
1fm2TK83QgJVW67m14oGoVrvZalsfA32dAOOH6LJdiOM9NJA1NMjpvSzDBLqxmds
uOEPm3139wiyfydqY6PpcH6uaKWyl9ph4NmD8t0igcTgg/ZcFwx7bVYF5sM1klMY
QUh3JjuAL4RiVk6SRsHrhEDmvVeV91PckDLC67siq5Z77dxzdAKNhQSSiwV4wPhM
c5n5gH8ZQ6r2b1dFgDR5onf6oI0PstRUCGATs2Hz/zF/LgiiQh9D4iNfuuYzgVU8
A5A9lFm1jfUkpZranRAL9JVpFgln2ajpdFzgg1bSH1iCeVe4ALLXcJsszaQbJvB/
BrQg+ndDkFDWCjjydjhq4/lLq9CTbtjKkeuRGXg6oMknTZKnk+Ll4pAXmiZcuJTj
zOJYLBx89stuz8/JU/3EE80iQ+4hM+evuVWdY5lCbwuBx4sD3SPq0C0U3OR9Ipoj
XHLGqYGV++SdaTQFmejU1mPc2HGlpf1wyu54ROg5CqbBNMoSN1apQrS7UQlDPypd
k5ZtQmkW7XEYt31N5KBYiQOgEnVWENU865W5LeIry/1t9zvWrgxT8NqCqwYEKC9h
jjiSL2gJaN0udlnRhwxBVWmXLuTf8BtJ5GJo4uG4WKJM3DpM+AjST7lHt4nOjAcw
9PefdaF2KnP6+sKVon71ALovV5k56SJurxDyVMQ3/Ddkws4Q//XMJSE9R+dPxsry
Yycvd3IydohJXfyfkEsyBtBLaq+dqWAaS1M+P03fFCtYiX2J/t+9e7SYSqxp1V80
QwKGIDjm0NFgiJC1Go9OkKFmAZiGHwoYXLeyxW3My0NPgeX4cf/zFiUQoP0oC4gB
cy1tMgbPzPMWSh6tSrhHiQWZp2SRhfKJslLuNdEcqC4lFgeVvw7JJIKVv4s6VDa7
mFCForfBh81q3amtpOCOEXBlzGPV2D+oVtDjHz5SG26Gw5F4SJUciGHUaWeRXxoF
`protect END_PROTECTED
