`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cpIb4BCENSYRg705LFIznlJFv75OkVEgSvOk+kiaVsXo4daMyJMbudUpluRtyX73
skUJfqkmCqCMPoWtoFNV3pMsPwa3ysRAEXi5psGtElh5VhufqMi9Zkm4nOAK+VYF
eEYT0OH/PDUi1mCKyEy7Aql/puDyWImNrmKDUAsji12vQCtS927D+Zfvk4op53VA
RM7N3olcE3X3wwO8uVsLEeegnNfiF721x3x5S4yOAF2MNzJbJYHbZs7Y54+GLb3P
4irddmPeUGipy8aH85IxQxF0sGadQxcW22WIsR8JReq3BQzoMeYVIQP0JoLdGIVu
Scpkyu90zBonJQE449K6tvIfjbNbDDuz+MXQm99Gx44X4m1FAO5SP5XDeLi9UacH
Mm3eBa+2EHHXGbLVogNWKd23vduxkj5yOFeQ9JqC0q/WNwYryVR1A03k5Drfi8FH
a0wdxen4PsWw21eQq+GTPW8op1yUeu3mUsYfOV5LY8CH3DO2UaLCJVwXlzcskebf
I/q8Oj4TOdKMgv/7L0ZsB1MmmxGuygTeldNoWmFaox+DbhqmlciBC6JAjLxjqjMD
LC7VAaJ7JIV0GmJ2SFYI6FAAROtG4NYk/atEv48TPU04DBgsyouG88YS7Sh9AoB5
Y1fUeMavXcBY77cA2KySq0LC+xVnbGLs+196up4GMhYborcIpcpaJ+9xIepLOsYU
LO/4tuicGmSw+zQgm/iL67NqzKQSg2K+SlKNKhhDeDi2GisDY2eo3L485FGBy+qz
hoP+ns7BGvD+OkRpSTnH8ZqlnnnYtwAkIEIh2SArZ4+q2jZzJa9hPrY8kVeCjBZn
ZrHFQJeP9yyRSo0I4X1r4nZ28ZFv88qmAIiorFjgLoJZnBahAx2m2htJSUB9/g4a
+dLsNwCNZtC8jkePX17y3N5E51A9iIdBrNdzixA2KFKk9aGU77yLZHRlAuQEc2Hl
W2Yba1D5B8y9uAXLzB6Q0eSQ2Kno3/p22BUL70jgq/sa//f497XmKSy7G44mvet4
x0CERUbyJT13YW3mRqtAJYrA1frtb0SkcTpUM91OtAxdkIZvsBkwO0Q7hiuWAnVY
MSzU1ON69Yy8Mt5+qg1r2csr/9q/d27KzQvFFeQm4X2PGADzg2gHnwdOwNyOCWXg
IU5aMmUzbEu3m2zmwmSMRWT//0WnOQouxwk6qrTLEsv7NwBUk0GkM3snXjbRH2vY
zTid7GMJrE6wMcAFiZe1lr7qq/fH42fmbhVQwn6YxdQDlt5coaTOl9vVJLxAvQD9
ZNd8CvbLZ2A4oLxeeE3hzBYYekAdAQs5n9XrxC9b5ibkOqSqRDBAFEFuyi2x5NYv
bcSL1F7v4i9qVrvckrunkb2A0tjzd9lCZasY543EfiYad71tnEE95Rz9WQNt19OC
RRh+FzE5ws2Zzbj4ppxR5VPfy0i11JUOymq5QQBoV8w3Xgg7dZAIS7G/QpQy1ILj
e8rRyTMF7Etg2lB1WmAKgy4vRGnn83HTHM3t5Kduv7MSH4h+Gn80qRjKW2I/OByf
IGKSoifjW2HzjZpbgZnkuLnqxxkXXZ4H0P521JWzWOzTj8jGE9Xc4Yc4tsxhcWyC
Vm6SttLDqpl1hFm1ag5DCs3szmfb+0zdlEiL/gRQgbpMXN6dEL9wAw3q5gyO7gZY
En9sC1uW0tcmvngSRee+Vq+T4QeWLJYngSB59UcsXNQC0UnGhWN0VjL6vzfex8Ye
PaxnQyMXzCCvzPYgDhNF0g==
`protect END_PROTECTED
