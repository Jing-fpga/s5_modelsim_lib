`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9G/QjTJat1B+3J84HLDDqCfZUEISN7boYqGfYGsMYkGuPeYXe6SfD4BVu+gS3+TK
7kr1/2hYw15HG38j2KtsDY6gep8OjxpQJs90C37u0wnjK5pGe7ThvhgdKLqGM5s3
kKjpPB2Ouei9zL4GsPtKpvo7BnWL1hAY0MKAemwe9IYKkjpdS3oQtv1xySJeObqO
6j6gtIH+Q8j374EObJFGDWq+zds1n+MRatP1C2K/pVWIPdQFrlt+A0hye43bFkuS
WeyqPgfXkijSswZAwJM7FQ/xI22rh0Fo7m4z6Xbsk7XudVAscznQ6ELf8LGc9x5Z
re1ftEXk03FyiKiULeAAtTXMz2E/6Zdls3HJ7pR6gfB/19EuxqmMSiaSKC2UGF5x
dJZi5X/YgeXUAx0FD9QE6oZkRaCxIcDezFzTxPL/Ph5qPJXLRYpbIBBfxn4E0f66
vBhbkIoJWAAdqRdypHcM+cvRV27RnwH+T42lr7JDYBvvZMMTdy1yqwT7tDV1scJT
3b+Nd3BR+VeSyYO1sGIVz9xmDKcGoU6TFgysX2HOB/xfgC0qk/XbiiGn9KvIUVoD
SRGHUyqO0iA1Kq1WnOF8vIVk8I//127v692yyXSt9mv40XcXeP0nfdfK5fMKEady
HcWJzjE7U7tOwPSsega83h5a2l/JkmV70JCWcKhVjlFVTQD8NYnwz2bUSafcohpQ
WXj9a2Vd44G/WYDKse1bL3ffPXjBOrEVCwFw+m5ilwjEDaVVSmTjitHR7ViMekmR
CaZJhcee6bAcnUoP4Qsgr67jtNemY8GTncnyP4VH2hPTc7nj3W/gz1DL//ypY5/a
Nuk+ZxfDGU73DPGg1LmjkGmUVK76rOpbcuJA6s+hyM//54N7Jbp00nJJD8Tvawz5
KZB1VXY9nTzvYcZjQOiDdIEG8q0YEEdNiUp9mWhcROgibiICUUcc3dRQyosNMsjb
QRKYcY2Cvs1JlmCsIAx11L9LK75SERH1zJfrS0trGJDHqRQeHm6tJuF11RDnjuHy
xRtlEjNlXXWgTOnhKTSqR8b8n0FbUQn5sQCt76c0TVaXgCnAaSFyngYCl3+bYG/J
eEFjbjAD1mJRF22cUR3ksBk7eZWJE1tTkdpHqe9mO/bFELo/lOLy8WKi5gp6N2oR
pzm4MWU/wbzcs3BW6l/sLA==
`protect END_PROTECTED
