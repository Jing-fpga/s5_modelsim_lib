`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c1fYcEqI5nrXUECCBa+h3/eXsYBkpOgCoyNdpfKYwYWEVMXmcpu2mmuxd+KHL9LS
MCeorlPhlmV2c/nXiEErkOMJ9fLUB2+gEe88er7MaLsiCan+B8PdiYHyjQSImBuW
HmCDnxqrMA4jX24eFg786w2Z/3Gpc6kHvft8hNIJ7nRzUdqZXWjriPJO4mZnfGlZ
N9NDxEOthB+26grTjZynT+SuJ85RbMn0OQs6yWQiIskSBArfotf0Lq+n7mi+7U81
60T8Oq9zOwvqy23WG3/C2dpwVY35UZF35woXWAXykrZxlVN2eeUEVHdsm6ShleBN
20YVmkmzNf6YFqNeFauNDJR5ya2Nu8cVp7niHLancLTK8OZ00DxlnGO6bx5Us6YY
bQW/AAruyVdI0dg1jtHyp0ICAzc9HRrCL4mhLkidTSWEAGbobm6Llvovp9LOv8V1
tVHYqmokn+yu20naVhA6gDI1aODw3Ur9DskrvoLs9FKiqWjlNLxeyVdX//CQTvWn
fj4rofxbU3pPVOWTU74oMNCOnZAUzxtaXXb7TeOhhctysl8tWKyVBZE+Lva/F5Qf
BQFUZTMkoqNv8jLOcydGaufud8t8Km7Us5EV3BPzuyWVvCeJ3GijwxGhOCdoBpTV
5HwcyVUYcbhdph8uUeUBTzUwTYk03wZBywU2+TtGyIsPNWAvHSmPnmz83VqWLJ5w
dCmlCSowDcGf8xhoTbH5wnlxvYuLsLEpiiNs1+WkawF0GumDOcHUEWjWCDh531Pj
o8Ig6kxzPedqj0L/nJiEBiNJUnj4CiR9AWd+CpNihF0JcUQYNhVshQbAxWAyi1ul
UOB+Eppu7t2IbPzKWAXEDEkp9ZxoEpaT3tmw/sO3aAG7GAVzOGMiqyx54MywRfpH
sywTIvLQVfdgjZ7610rJcbzInUuNnp0BQXMRtkY6/8pcBmEdKsLy4DsivJJ53as7
RDTptA8o4WfMHp/I1F7JsKfFQ4TrQNV9BS1/qg4ZRRAruZBF/wnpLQTsNt9qk1jx
GQpkT1CNlLR3uKFH24T2zJACAEzku5lGj5plrQmROM3MfflGe/a+2ehaA08aeneA
Zx+7qmxqYArYRjd/VGyXaPgfv6iN7Z8b3gnknhFN0/47F0ZKlnDdRCgXOIJfclbn
ZUBAxYksvWHerjdZ18ukRHoPSNfuC+3JdeUDV0hfgKDvfIP3R+qcTc65h+tWwi15
D0cMrV7FAX8kUghuO00jRH/irAUvyJIIwiqWMhNnqcxqhnzvLq2fXWmHLI5l24CQ
zkrfm4NOtO1TlH7O7hxpM1VhHFiG9f4VIejNTJMLh15Ns2meFYMMvSLR62WtBSJm
uGVJb/Cvq8DseC/lERUGrqH+K8zj1R8oEpWn+W1/IgI/iRrO6wWo5Qs8n1NbKu/b
yWZMTliJdriB/Gxxe8SHO2PXu0bowYJeCj+F3DlhIznyf5wVnIYfLyytlagJXjyO
2QUConF2nw/crmY5L8OvvPxdgoOaM/SHQX74MYStc7MSIQrFqxnr/wE7WONG4nNn
bbVwysYs+s+pbch3hDZcF7j3fRyvx5safs68iNO+2MpAnIk1TvWgljVEHBISVusv
I39SRS2lBV9Z2bBmddCB/89tZxIfW0JlKYho14Uwz9/P3DLH3XonfhsADIqNG+de
EJb/qYFRMid+xqYdG1IK6FcoDR1Biy8GAUEMZI5wyS/egA+1czjyH7x7MR1muTdM
Ibs0ZZ0XZWhuLjZ5F+NY1RDSO9CAsGgcIj3SX1mCJqP2GewZIdvkLONWEpBfDsd6
9Dd1ywld2M51iDpd0u3dBnKb4pSHgjsJSIYzrNhreniU1fTRk5JYL/BiJczvewLj
ZxHVbTJIAQi6zD6ulN4xWLiWhSYQIYIed0+XTR2/Ny2tJWi/SM1NNTq1EQmCPvYW
GKLyk1igxk+SfpCDZ8EV03asf0IWidf8ugJeUHwzSQ8rb5pyZ1iAYKv5PWWw6yQp
YEaDeSd7MYbBf4FvgC9HcGFIxTUXDC0b4W21e8fsrOWRZ+5xoiKPy36Ow4eSzBWB
gmaox8IA4eraXT8KYi3z4Cl5+uNdgF6ZM9vjD0ZphHuO54Up5jDK+ldJC43gkTMH
r3iKcktnbKzkC9jv9yO3l5oekMN9v/YFG/ZscN1kOP/hE7uuXOLM1uXmdIh/M/OF
jXVY2UL63E0HkFi6AiJmJwyEcvjQJEZ5oP65f9ntqrQaavv1y9vvyxMXcuNiO6hf
K5UnwF0HpqT94Vik2fusnhCHCMTF9QmTS7Ho81Xv6UHcg37ccWNgiFm3zYzn2PtK
XLNSLsAvLBZgThertpYhLtAqKdM/tQl/toEs4KwBBd+eAb79yJBaOCq5Lk3FxXxq
eAx7220LWLE7ChmEN06dUDkGgRRLnDC7QSultLy1NCJqS3ZAskQMinpZfZg3FzBf
Je1QmNYgEgJdlt7BbJEe4+NLTC7VLOkQVxSW6GnyStX8GrGqGHL7G6kTVkcnjKdo
RIf/3v4rDlsUjkzsKTUPuzQw/SJUizANkBCpUiT3bc8oW81BjUm3mAhDDKA72W1j
4Xb9mzTLRWxXpcwU2vJdig4NBMWh+z7zZ+d4sJNhItwPvnD1t2VP05u/NEi051jR
T5zfFq83Sq5bysglSWX1ArQ34chNMggd5OVnDVVI3LAmSOXRAZw7myq+poZeQGRE
XAIcsHxkz3iODIOhQPIPAMkAM7sc6fzwc/0E9cQcP6CiIDdKpjlM/byYQWtPjOQB
Me5uwd6U89Cg86kOR2kTMg9DqkQgevjVoitP3V/boa5SMLoKLGPD21xS53Br2WFu
Dair168JLd80fa7M58pYiPWnTzB1B9ZnvF2IyWF2le+qZYjamzOgMtWmgIgGG3QV
s47EaG7nXNplR+m8Wv5lqCwMGJA4OjgDEh6DZGsXx/0FO23RlQYtZszS/kWUzY7v
0lm/FuBtgYnVoCiHmgojhykCw+AP2yzxWap5eupZk27n9Pk367V8k5tCY4whdUxU
U/4Fu2Qg0hKTMsXU9tRII5SCZWhgVPaZLgQ50OjXrXh1cJbGrR4GqeQPUOHRgsw3
Jc7DShZinoGmYsof+rLQBfPPA8E8lqSCbvuf9dY+JSNATjiEX8UHD/0BtZLS4xWw
xzuanwqMkaHTCGsswhHI/UKoODGRDB3YfvI3Vp4ZTbPYnFAKvpHoMJpLX4smV2mu
54BJoGJ0BGfZOTEcRiTaH8ZjSU5hqpo37B7h1dHbWyv1QnfQTMLAYdvmNJxgYt2h
QXOGvA4G8odd8I9zQCx307XLGEJIWxs0KoHF3D1RO+Gw/9gMXcRtsMJeehvgN9ml
HjaYmTwzzb9/jmxUWPLs9XMzsYEMr4+I/wfetitOLU1tUwqCi3XqkfON6KNrYva1
lBKkEY+vrJ+jG+N5bKrNPqGhPiAMcj641lEa9Ma6Vg+8SjJAgtInXDToeR17kAiv
KxGW3L+sz/pEV1LuixckMjWo6fMLzxp8a51AJvFFXXSZP5/DtcuO/NB4vCwsrtSA
VhSWG4fEkbH9wTnL/aCEkAU3oPHqtWzXdxw5j/PAxOe01cz581ZnL6L19azQwcOT
YZafqKUyog5uTcRFPcAxYmKfhD4it93tDY6zQurFBX03P2ngBYcn9MOgxNnmSw3s
XRkXlNzZSvspo2itFW4uRMWPjQ6nl/Gb0/4Z3k6RmmxLUNPhKnmYNUruk1OBR72Y
IsrdeQ09PKbUpr7hhULjGnb0nmkZHhmjRkfyBPNWyB6BLYsGS05e1YaiXbBZ8bht
APbKmm4iDv1Vo4HYyevoIxc7+xyE9CLPk8R5JpHXFDpi+/4TNEF0BinH8a0G3+k8
uVuFfLgylvzUYvKLOAWF+REPr4Jk6vaoTZUtmJuIYMs5QSxFtgcZpou5bsYviRZ9
4YocN0PKlmD5opLgRyvr8yu1t0TIJ92r6yvX1/g/cNJsj/lT5Ktciv709SjMDKu7
+lFRomEoydVFTIVF2PdORCIUBydyrkKIA4HyXc7FUsd2Hc8U4JzFyRHFRlcbk1X2
jWeC583BZ27xUvB6mr6hnCdKq4XlSgb4Un/R74WRCWQYemPPB8Tn/JAH6NCGrwDY
Xds85CMNAnrReaYJJjy6JA3Jc/ts3GPGuGejEx1TOBIK4Sc+PG25x6dZv14roiFK
tTiZ65Ft0GO/B9rUJ+eaHFMR8PjxUhwW5UvGRShrWKIc9TayeXPVzscCB2ziFK3w
0ibRLWkUSDK2LoKSoxAApf4qtTz/1clbIzrYoO/zxnfeYDXhwKFeE0oDKplEihP5
hkTZXPUxLSOua139/ZxDJ0WhW3VHS2cFFeZOuomjedmhnSusH9uW7glMCi3fyZbV
AMjmtsWKSUUEkeBZQ+M/NlIKw8gCX/5xf5plJcd1Cf1cWZdb+HsFeJ6am4kXvwWk
fd9iJ1bp9V2se2iR9l9341vhNxJYpvFq2TnBWn4CNvujtljSJ5iPUM3KnO2ZQKWg
FO0oYZ0NvczmtxVpDk4kuwquaAsjcWqdqJRRUJB0j4O6K/4DksQKBiHbGF4lx614
WxligeMFoBE4Fgt4s7GYehvf5W8x69dnYa/LiBW/c0KwvNEHDM2Mc0/N8bbIMYKF
n8wB2VdBl1SSLGB/Gftrp+y8XkkMVSrRvZaYwDj+Sj76nM3wxfTTOu+fHGFohE3a
IhoKCakGQATuEL6Njo41JoY02spo2zCvlZFr2lqUHoWkYYqq9hjznfNXjQIzNPJO
4DZipP1VT016iLAvUMdN3h0bNRM40CYWo/AeCO+rbixbJz1/nnRCsyhdc1371OxP
Ic8ZcrIjAqMD/22gZED62nd/l+cLQTSFl/CNz7m2QCDyKAMo6WMohc5oh6xngCWo
oUqXwluDidLuwxKj2KtlWQ8rjuRg4LVsZI2SeH5yORCzGJv2R5ckdOxiFlVFfeK0
4IZ8gLwsvkWfUEAIvsrRlYNiKFPlBx5YWvwBp8Olegp9uWh2n/NoZMaaArQNu6vF
C/PEMhNH4LmlCPr2p9GrAQ8vXj5te6zdEet1vpg142awBoA+xmvhqYsjljUTew1o
8BX/+rIp2B4rxw1wYzAVvXut/SgNZbeZ/LAlI/sUt9XCKT5qJfHLP4FW3tKGWTVR
EkXkRxSgJ/eFRGOe4S9K2p/Oma7wKtFObS32sBSIxdxSSfE/whh0ohiEqyWclIiI
D0r78nrDYi0ok/QqVH6s8oL3LtGih1pd0qS2bs/toEC2DokgYkVpM5onUyvGwwDz
FbeMW1NfTgzq8+tTd6A5U50VVCmdPLhqSZTV8mt+6X2nQcnR8e/y0OxRLoGPTLvx
AmzmRBxMe3LgrW/xZ0HkAYmbuAGv4uaztgAA8yyCbjkwMDZjjfThtnTendHxA6T+
ceSOPm3k8QdetHiUD3ha0X7ECcy/IbdbGfBP/puVTfNdqJI4et/XgX0oGE6ytQ2L
JBu98Uq68TvWpgXk+djj85kgQI06brZTjy9HXhg+S+h522BPpIHAAiMRD5aplqkr
tUJOWxL/ZCBhf652PVeiS7MW1wnJMLT0P8mXrmSRqqkeQpRZGhXTMHFXVLo2jBTw
X5XmMxD/d6ps17P6dp2Y+M7M9KP7tYV8PtvEoavqtsDHrJQOSSzOoDagnqAXUInQ
FXTB/4+9z+i5tO8UTQqMeLTSmUgtt4TvLdcy55RPV3E/CQGB6cXg5Zc5o87xY0EG
QbPK0ZUWoicw8NuYGAqjfLNL2U4YF1FwE8Kb8H7Nk9iAU8VGBWp3Qf5nTKL6e4Gs
BQG13uTiVhVzIkGFzOF7mcKVAYklczs4CgUU2vIjwYI53K7zcEsYzTG9AhQdt0AY
wc/lk7Vaiz2CmcLW6KvEMpgsoMSCJQnIDyznz2ecGvZLr6eiaGGT55pcpgl8tTfX
F860y4HOKne4XnYIJoxroRi4RupCp1ZeP3bt/joP/Y13CVgTbxzS9v9z8hqp+GiO
7E3CXuveyFfeh7rOmyH5Xwtzsy1VVkUt/F1dy8e73FATVYLrXvMc7pLnZLuN5p5k
Rvt2SrjHLgDoxf2pJDhnttGXU3Yz5BPYAf+JiFZDpCQv5FN3nVEbii11VvMZ1Cgz
naHh0RBFxLx3UkrHcdiAA+UoSgxlLkXNiWggSrAvYnKfTKgSMuK/pdAQPsZLTZbX
f+OQmaETjFDXDVZH3FlJlant+vQtvV6Rug3rFDu/ZhILhz0ziUHt3Cp5W3LYEG/w
hhSl7kay9cgl+r/sUyCMFVe2o9WmpupwaKhuPvg18XF85tC1y7ClnkeXsFvNChjf
nm9rXvS6E5FMVZmK8vfgspmXK23wHMwgN03MNUvhtR62aqa/RTyfvcxcf81DM8gd
QBe0NL2ETLz+MKsF3o3aGOry9OWqrgW870N53z4RY+n4B6HgLmQyWX6I0DERHAju
7S5W5/wpJJwtKPLCcmeM4hts0G9WRZe6sQeCl5iQULK7oVD3BLWbOlMvuHIat3kz
q/RVgNDLqIcRBy7s95oxE/Lxs7gwV3ZM0hmwSnGA4Ee3wXGtSWDWDy63YgNSjK11
tgyIKTy3WN0sugFE0KsH9HSWkwFMu19XpQeYrqgWH7RlhyQZ04YGe8+dBXShNsSQ
8TAZEYkwRq1Iafi9Hrqx8Hu9gqhFcv622ggxHy/vHI4b3vzOVHxz6U95iD9GNV7X
lDGvKDPr/lY6TnfyTKt0xeml9suBeLhvCkW78igFwp56A5T+EV+kiyQpZcbpNfiq
jVFWEqQ9qzmbjgpD6OYaKMX9+vKbcmnMyBuIXhJE9iqy2m0hBk/sQDKqOiHEOjWG
W3Y5bdmXk1jmMaHFpD7Pd45V96a7J//Mn6kxetmLEOnSws4lPtwO8cBGpFc/5x/O
6VKNPdtBplIQmlRTRFVvXCtI+/XCvVoh0pSA0M2y14ANKQ+eBFTvgxG/3kQaIchg
mLa8OfxpD/36MeSpupjXrtCdO1x4Cn2QwSoLSfUADxYPY5Iyw4V/Yc/LnmQkjlWI
XxA1g2u9OUp8BTbAXibHxg8CbSyMtb0RRNh5TGibniswKkZ4tTll+yFrhzdUDSl+
mE+vztHmUMYnYHt1SZ5hj0eht5jT/CQsGfJmwHiuRXHQ2apxewcMVf7yTltUFONr
s6HpOLfeqENLLDU7roi32J3L94fgWF/BvYbRJud546r/Pjy1b54aBRDt1PwSuuWR
JmkZUvUenaBD3pG2SJB4ofyINGAT5Kh6UJ+dDAVjHbjN82q8SW37hV4I6//buHE7
+pUhM3y8XElJZX6CqEn71yPl/1pKtsK/RmdBvaqoO2s=
`protect END_PROTECTED
