`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7RFCCYKfAEZAKrzpzc2bgVVjLI6ImybHUKUi65Gcm/mPt1rLJjksQuID7boO1290
sSYz/OJG/glXx5KWP7w/y9ZBXZqL8aAxhEs+7UL0+fktcjXyDyem87ajOMfopI71
ZLQW5V80UNUnH71HYlg71lXmCQwoLc/kWgUy7tThimn4laccuVAnY8Z3/F8ETvmj
LlAmEpXmdioMgsSByXMlNIz++toDs5XL4pA+P2deQx9OOlQHk/yqJpUo1DkENweS
amKDIOJeEt0ysWY36Dj2S5O9webDLSJfjX+49ZTK+uACYWHLfHBhL49fnBtUgpmZ
wBsrRFlFY3asYMOHFdmk26x3fCHYkYOADu7vVBUUZ18zCwDHVC4l02ZnJ1SlouAP
T1IjF6Roa7km2rYrIjXn3+M2ek+Q747s5QNwAUjkqmsZHk7vnoJZ05AtLQin76w9
3Ne/L6i+BzkVvgHdqO5dQ5FTAFFrNJMwTvcLlqm/ooG7pP+8nd3DQgstZuvP2Ggq
hQjb99yf5prsp3nQwkX6+mUnUnvszcDlK/os7Tx7LLA1sOwSoelS/cvzd2bi8NyH
ND9GfTm4jxzUeEyDzjeSJvRBa1gtzGKJqxDcKwStJjFAQDHQ/+wW8VqUmYo+r+Dv
91MtwS+0Q6EE0L1qebu+qjJeMtVgjK9VkcAIhFmDCQ4XJcAH5UnRwSgKXAko5gRg
wsjPElUf9RiRRX8hyVezq1GPjTKvEE5b8xlpcV133Oy7vFh8FwgoT7+FLJBdXKf+
0RqoyyDDD7XoJezevTc6fWqb/xWZ5LJb+ibGTLPpGpMlgY6n75u57JYuFcHa+ati
JqjfJvWdiBvIBNFh3Tdbyjp72KE2D6OHR6XIc2kxHumQHavKoMpqpqaH7libYeza
FR70E4CIEz0aal4PevCALQNNRgToHotbX4ny4MlcfgIaiRdBD2Rt2WwK6F5NzrMX
JqQpagltpeCXQgkDxyMT3TaKhtTm2pN9l8y0bVvRa0zdItyTA3dPM7UTZvV3kNy3
2u+/wxcp50c5hck0pEGOCeMRD2Ci6JrqqUiaLgBJAOPxFf9Thxt/uLUIEn4aYWWN
fyahBzFQzbeoLB/pbT1XXQMYYpsZwjW99+SDAUpKbjFG98cu8+K7U+8Kw+WQr8gP
M/WdJdY1wcMxsWBwFcJkwn6yScSYAAFyueyX0F0km/v2KQ0jYS27PuEC8j0gcnTu
cVZzA9h9JefZeQ0MSn356sWDsITBj+02fqI8uUsipPgk7rn+uVbdjYTZIcmdBS3U
vg4tnt+tklF3mlzrfUMi9ziAQIyP0hnS2DuvniBXInc1vegMqtAjhnZIaaHRUq0+
eyymiw6fgwTmDJ5Rfejaj76rZl8tbtpWy255fhetLvXxLb2E98BNtNnMIeUImJKX
TOfy8VtmjOi0DsWU88Ny+fZ88LbWKhb4qg6z0rUFqlgDbOkPrcCSutLqoqt0gq7y
EE6hBVBgiugHyWl/2f8UucFWadZK8SA+1bgWPV+AQ0SMss3HzvQ+zFsmjTRdL7qc
A1jqCHuG5qYJZURvLn8P6XFsis3h6vsIOQ/94led0bK1Tz6PleWzFVs5Mu2wpDCa
QbBfk6ANIvn420EmzamBxHK75lqr5h0P8ZzawnOOyyj9uV0UOWgKfc2hLkDmcSlD
1iviXbMKjDOwCNMmQ7t6liiblD4obyGG8erHhO+0yBwAsgEjJXTHQ2cdFl+Fu2HA
giLPXUtOh463N/VR0zHWI1EsbJm+9q56uHx3Ur1N/UV0AyDzAnvA0q6vWSJOOPKZ
IC3oHOVE6VunyOFd3eLf/+bQsD5zebi4f0FgXaqsMQaP97PWw2bsbJJf9RPPTW2B
bmkhYc1yDsIgO77wztA5BAp6MRnASLJPqCeaLfnGUXRx5qaDIhlAA0WbKcUxQnmn
4OtuhY/7PJdAueyzxdl+616hC+jkhKYEoG3OWYeWHkhhNZCOuq0ZT0pYJTSbies7
5Ub3N14ZVP0bXxAg56BhrjJNtT0im+g3L+ivPpZBJxQ6ylrEEeYNiwP6aeqDVpQd
NS5bYoLa0VChkooMXsUlWnGp4NzXQ3KqbL6RSfBYySkP+86loWRhczzdk27MDf5T
cEZLtxMlRT8WKd5XHy7iHojVmPWRDy739m8iEj0zxFMJUA4ZNS3nDk4U/a0E+oa/
+36XSBhW7anmesek+Cv4LZsuIMZXg1ACMUtQg6GiCIsUg5RyDJ4ia/MaoA/fjVbK
O9XP2fA/3GCKySuWf8a3pYc9V4P4tA0hfF1pebomiCfVbX4zPadiSH3JUwFGX0HC
VOXny8J+32Yor7Mkv8nNrDemuuSbJg4+MBOUKt4+yu/j8DIGsUMjD4PrrO1cdCgb
DrWzaykODPiNCuDzNwxljBm0RCGtde213I5qVkUidJVY9ROQxAG5w3/8U7j5VRb0
aUr2bFX85x1fJd5pz1sbQUqBIA4JBVeft34mtRORjs9wbLWhUlxeB4OIu/O2lfn4
tx0Dy7EF/CgoPKLVYKdwo6+BavaYqqpW2wDKV1hISLw7cxbSdsTM5B5KufBuAsax
OvB+STYg+XeYekbwL0xnFDkywX01N27yJhmEn8Idve3jwpFG0uA4/ElfQdyOQslr
kbe8ujaLY6Ms1mS1/4AnQXC/Uwsrd8nX0txkDlW+APGjv9Or8CAGEGWWU55iwPaI
jKfTmpT+qgPZjivJ82RhnOqXx4CqVmsVQPW3GY/K0+rkaNObPYe5Ve3SeC91eFgu
PM+FOLXvlhJTkj50awysNoIQITJEkDRdhhXj/073Jt0knL9SkTk9qzWOMLYZct8U
iJLy5DgOLvhIyoQTh0FxiQEX7+4Uj/l5x0ULXUhvLetoGLnh4JzdhWerAFeDeJ/D
BMGZwib8J9Qz7deh8oI60CNdxCYfWLfpse3pxU+2ePEJF8YqTW745tDaRMeGX3gU
60O2fHGlcmYjRtOMaSS9A/XqEJoKPj7VgNquNnP1xE9wIamOekbL6gqcPLXLSGgw
yr/CqqekyIjNG2Weedq8G8upjyvVGafwK5agkE17t3Ru3+Yjor3rk+i+qkV3FkrB
auWgXj3aEk6plE9cL3lEG9ZdXuZiZE9j1G7Q5budB/2jyhKmA/Ck2mQPM29nxeCs
jDN6K7hfNzcmRy535Hny8OmFbzytGo+lTzo1CL3UUbPUrahafWkCEw8SBwk6RDH7
WytwE9kO5M4AxSHUshS5XpdTGyRJpsHtLgtt5tIvIn4ZHNjWdo74y1vxTndR6w8m
3o5bubKrdt1AKEccxtOe9NV6uEObFWQ5CkSQuvDI7xk5OiGLJJfaMIn5RfhtnWIM
fWbhefT2QTfS+Hto3Bta8GL5HY/VQIxPupex2KEPAptmB9s+Yh2Abz4RJdULdvaL
pIMK4QBsmYg7dlgEXLeTNmZMEAC4P/OY3B9rdloTcg8A6jylAsYz97zjxBLaQE0a
O4J5tCPwsTz48r0Ww88gtEc1MEI1gvHVa/nuDm16aVPnFm7uBSC0OBBEe9DU+JG5
7xnB5w1hZ6BUCVo8aFlhpLuf8uq5cJEvnSI08yzc4topv/52RWu7X3ndFXIIpQ+O
gwkrvF/40uNDNjSAqDYqae58FoIFEcH4TUtum9Fsq4snOUAgQHIy6W9GAppTH6Nm
K2FVLOZ0CLhj78i95E1DyHytAsbZXF+Ovf+ZOLY0IlH1YTg3M2jsUAtXrRi5nEFp
f4/hLGHpG+GVmLCQs6i/55GiENDDQ44c8lpGYnzg9qq49UXhT+C9WHXHfRf37lou
tJOPuqSizJTcz6s0HQ9T33HLJih3Ji+LrAnUMLJZOEVarZaXbDP0xQ9BUO+lUGdT
PZSsDgEZIL8WMm0vbSce1dIaMHhtzpQqQmJ2cAR3xI9TmqqBROTnD+vZn9LibpPi
KkRiMwmydUq12qjPW/EpMtpWc9aFLd8D0ZsY08qV2sw9dhJAe7Fn8OR+fK8kSKrC
uwZ5KuwxSu2D64RK9hkg5Iko7kxyPPJO4BB3auG13qWp04b/a2XO2SL1zQr6gvxy
L5Gakqb5ytBUjHDkKTJ8ySiZZsDrip2eZIUGC0KTv9XkRt0ervODYAMnHjN7b/zv
fFJMOXIbgDxK4nqD5JBXuU7QvMkcpAQ/3qATTowQQ2AGdCx91T7eIocJ73K2sYWx
ErEyo4TlnLaIDAbCD+HQ8XXYjXM45DgKBY9F+DOrZJoaAXLAH10rRcDl3jPQlqiG
8NZ2NHALdNMD5xaLoJFV6blbUDBunC50dDkeK2Nva97U7liOEUj/TlJd+wiG2A79
b3ZtYd3r3i61u16at9bzWQput7zvxbWe+6I49Vo3SBZn5S+Eh6NCo1FuCQpQZVfd
ByzS5xBvqsCaGxpErHtGo4lZYQhEkf3T95aBprL9Acd6hyM8y1KzTcMG+VsGIcEy
T3Ro7ooMchUiXc92qTtZ+C55CO4qJz41EW8sMRHVAV2mM2NbrzGE+treQ9n7I5ZW
bgg3aUeSWY3hO0aZfJGSoJvXYbPrhjQ3JcMSnax9Js8oyUwJkwv2RKGs1eHxPp9t
hMhXKU/beIgvIYbFuXE+J64IdLGis31AaSDs3sw0pWUjxSZd9dIyut1+qILwoBZg
7uiLg9R01IaAj6pOf6ES18z2UhpZFO8u97/PlsnQ9Ug9G7hYqv2oxzU8vzvtKa5M
1Y5kcb09qONdSyuYpwDK1I4LWcLb3PPeHiXXwEUfN8u9j2v9dgDEsBsuv/1LJVGr
JILDB49IBvKehQXhHS9P98a5HMAqyyUSv9KGzcdE+VE4nUVQG3TeAJ9iIDqk0gAG
xVJoQmvmxIInh7Uw94KHoitmCCL1K7dbElMTwaGpt8SSTThFc9/H8ISml5ef7dte
b99Clt1WjWBHnLanKxypMBB11jsjB51aZ3YeiEjvETfGcni8fEnDP4CkYSSK6dtc
EzXR7VJYRH23jm2Ir5Ktn6j7bqn0R23bihyUFzqw2dXed3P2rME0Xt1y2N+j0oMP
0FTplmkM5/kgsEEWGHYWtlI+LxXUKCrZf3kW5Yaakmdj8L6SI6K1uHuhH67WCQNv
VYBbADSdSWVTuOXFUw1gp/K2ET0CaTjIkPZryATFul+f4zWpBXT+u//fQ/YAJbG2
tfegDKpAchZufIMvzOlowoixYn6wSI2pX9e0cIgHxDYYmGDOyXXNA0aavhA/ET5y
Tay1/GMmmnSyymhJ1zfDiltl7gFuZKdn/4Hz7q67eZPZBlNMtZLewKqdsbG3MPp6
WtncXdBgIdHSaYLLuKE/QUG0pmI5uStW6++axsg1M5gf5jl3Lzu2qtX267t7KHnt
FI+UZMaNoS5Q3W3zbuD9mYUZnuNqTpxhM88GO3k3/iQtcy77oQAxQOgz+SdPLbnE
hUfsty4lGU4YanXX6f0WCZ7LX9jCX/LLZV48kI7sDQlhhEUcDkbGrVqdWhpSEZ6D
LIzN7rov0Kegt81sKt8Piqt74YKmlVDyrayE3eNhw7TjBeYcaLURVM1F4d/psZ8P
FFAPR4JfmTgD0UdiRmrBxfWiPg4VEpFWO0YMOX9RJlU8hvuSkNs7Z7DL4bWgiroG
vQpPqjFuzAXrmYbNNvLWlBABuRC/wrMeu/XSuyeckp8JgwFUxCzxjL3NSSiY3tza
exK8JSRb58hsEJOm6sN/LLtJ3Moi4ohDWH2KJSc73ge0Ig41557FaAhdVplRr3HM
DK9JqPKTPLeowbeFmQj7KUMLgjE6+uCHJwti3tUH7oCMRC74KWScQ1MYuCLRBLUg
WaTBJaLEtvu08jdBnHIt6oe6qlX6HaXZ2GJTsGhnnpVfb/Q+0i+QGGoSGM5aF90L
X7Bk4SW6iXWF7NJpl87gGwzwMvTmvHdvvi4+pAtd/UXz1QO6cVtDVcEglsC+HSaS
pBfKmCXEcZS0WlKT8iidEcUnDeeXN7eKq+tZtXgX0A50jZd112CyWtOxNGvAbr1V
1mQimdkrRRZgN8oz3b/DjqayXBJRdSMf2GftpmsFgYE/Xg638edPV/BKViRAZXls
z+ujMbhIUO6ILFfiSCjKxD5+IiiioQQID4Bqz/s059O9twLzkbfRVPmnfPsoA8ZS
/MOYz2JGet5nub0Ps1ote8nxaXoBQ5gcXSJYRyDkRnYo0cLrgn6C+tkZijXHDDiY
tzfUGPOr7SyM7DjlY18lWRbGd+zWRTZFkXqa2ilvMdPWqstb8gpZMdkrDa2EG5Cw
FmOWLOinJcxDgMr1RlxvoaHLTJDWbemyikccOqUEMmcI+h5vs9Q+l/fP/xbVzGZg
SafbpWDvJ1wUB4o6vTuqZEXKOOhju+eiERJY9O5zuvfkEU87/exyieYl8WvvDETh
2/U+HCrLISLx4+QIyzd7EmWzgQfcI+cNkjLkDRjxAzBJ+gPk+dzS5amcBZIZrI7/
XRi6owXY6JuhPQpxo0Qo9pCkI8d2i0uWXxfR4cBCqwNKJ/xvvhF3RfccESsvUe4z
p0/PSWsbanYDaCWexQNT8cO/Wiscbj+bvWf/CPAjqYXglz2bhLh8VFusayfn1l5e
3neVrLDUtJlgzVIuZqluczh5amCYEUwUTOqTjXq3/HnQKh+nBJsgLZToJwPvbaM2
Mp/5X+TdWPdYwdGEScw77PUiCbrAdtzRNE5y9YU98hU6XKZBoKDL7Ob5opprwJ0H
I14HNBxoANkPr0vwtlj3mtOTuWgFjSmNcZF0rzL73jeqW/BTzqCaWuI8Wsphb+b9
xrr6dJFDQHOMyxdXLWWyE12UhsdpKgD65WG4xLnqR1HLphVPJS187GmOFs9MXNj3
jfYYkgtQ2OjdIet09YoWU/QV2vK2JYJleQHIQ15O36XLSmK46+l4vH2zfo/NSL96
n/9WHnSZwusemswznjacuQB6/HH2YKsSKGgwd6dE440fkkCVXPwu/nODLEhbNnjf
tAT1l9/BHK3Osdc69JR2m8UlCpgggIgH1yyzu6Xzw0kHyh8Gam9hgXxGvK7mHsjq
0jkX5lN4tODNI4HXxvC9iq146sDuihXvJ37bjLD5c+uYqYwGiXq2PH8W5M8y94y4
7Slz83MlvLH1oYR2njiIAW7qCxJ+ptQC2bU5Nlp4R/uu1p0dtHfXJrLFsUREArEI
MPzMIRpFoYaqpT6ZQtPWUlR3sfyNxVldTyrTvp9HW8hK8wQ9U+e4+LVNA859+nZk
pPya019DHzXCNQnRUplbokBDBxdxzXF7qH68N5zoRjPrRzWf7hRnhDMFMNON6iNd
PaVGyXQPLmbaNSGGsAxmktkUnusW+M16YS+8lmO/ClSSox1E31z9T5BnNdrOSbfY
l8FzSnF36EtTi3neoRC8n1DNoaxeTAsoU5kDQZgJhLtcEZR3UTGUzcUIUVNcG5+z
Ab8o1JLoNMnvQwy/QGiL0PFZfxfoy39be6ycLiQLeWvgbfHWHAukZtFBINTL2c8Z
XTcBZWXjN1iK2usic/TYTHxzMR88NjGGriq7qaC6Wq0013JUpA65Ub+T3xOkYTSs
7HNvUW/fJGZtmqT63LwSZuh6AEB+LkzRz1QYuNq8aprHi6WR2vbKXU+d2jPwgtY/
jep447+d8V0gbX6dBghN5zlc7eUY1sSK+EVivaw+OPnTouJCKVtKomIt4QJUZicB
cesT22hxGcoirk0/DDcw03uXBu+z3jchxcwOghfrU/xKnGJ4upL4MIg+/4zH5GEg
6357qv4jQu/xiDeauLRuVFwg5A0H1mvJ55QmubnUu3LAdISKsdFVAkaux4Ec6riI
A4ChJBJMWMNYUgc+P3GNAIWogXt3ni+DjvlibwC5L5LAqxuGwws+J9FcAyP9ddF+
nSXau+M3voXyRmZYiH2RZGx4y9YvL3KcBvMY2ey0t255/3ePj6tdF6TYa3JW1IO3
hGZR7kQPAYwMRA4whEvJnLrDPgjQa0q/6hQYOUy70WqQZPwoEzPq8M2y8Viqt2hj
cVcQQyKmvtIl3S3Z6+nrj521t3h+gB5jzlIOJFHcqyReyEdSF2qsqF0UO7J0Lzwb
6uIFngGZiaG0v7JsIKxmf5r5C9z+TxWtcYMaYg9dhtcra/p6w1gD9hIhjPL4RUua
qqnpObduRpoM6hQMyWeNzqNjrqptOg4Z9mxm3leIsM5ac/k3Hn8zx0LcRZVkZ4ZY
LlGyvEJX6CoBqpqLmqhKW1W6/11OhI4zItp5/IvDRjacM01ndBbviHLgq0kJv99V
QsTN2SfVLBJKA14cYRRHn65izRHu8yl+vBxUaL2Sz3AROTBgqrSDT2FlAZMlURSe
A+EGcKOQ7B/bXm9H8lRxU2xuyris4bNQnZdD+3QskSrV+IKaFSwXrmkh4euzH1NX
`protect END_PROTECTED
