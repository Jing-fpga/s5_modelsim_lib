`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RF8WEuiHKMhS+MvJKAE65V5/4jWvXh8WnLXScnjLOmOYCRRugoO5SMonu+1RZUEL
vbpTlGUnJomoeyEnWxj4Hv4zoQX0eDVOHGu0l2IwrzX4W5pkaW8sq885dlQITeF8
KXiIvndb7qWL5/IxJX730+pGSCES1zXq1juK5j+lsHisyJRr5bb7ErwbxZU+N34T
+T7oM72uDS5jfpLRH3n1iK4KD0gMOnOuhZu1OSum1rPs9HHGNAnsL1JqQVOm2i33
W1QFwWCWH0COy7ZX97GY+tNjoFHCvRpssfnhbcafiugprnbUJgfEoDLy1vPXfW3g
K7aYQN4itBNMtOTChyq5gdxTn81QYx+pvcq9pdp7xxYUjljMP04Z5QKgxygOR8xa
+jlUf2/SiR8AhGEf3wcDb0bR8qk/IdphX8OLZf+OCr985SjTx0S7l1GLvKZWSH5n
yj36K1k6r3qWTg3IUn554d9ZJAZeuH+9MrKl0LFvyBxT5dvrvXuSgj1X2LT7ciJt
bIJ2pensSPTCglSI0pkBAPOZ1svpWOFKS2q/vm1w8Oq7dwXyqsi7DqZuxqUlqRjQ
L+Advqx4ycChsOBotbrpdNS4hfVNHSZdoDhQYBZwmW0OH/rrZA10fDEyPHabkFte
KwOkZ+Ab4FgJ95fZOUX6CkYL8w2MbYUOw0LdKgp/wz7GjiLU7WvN9KS2iTH2k0Va
QNYo8SY8PcZEjGOqj5Ovc6hlvUuk5glZ85J3l7o+whdx3MID9Or7aqgjzn91A4p6
AKYUvp/xq1TGlrZil7Ql50FsT7JkmZ6xp2iz+JEdE26Ylm6kMzrbyrDaV7YKjoi9
9hmPFe9PNGgXBX1+VSM/00d/x/R/EXZYDgr5QUf7qzCvWgU8/3LDbU97yUvYySpC
dTWtmm88gMlmW+f5foLZlG8WVRWhcPxHIJrM8Ntjqh0uL1oPGip2IVpi33iLKCXO
WJhzjBV+aEBDfVXYvfj2ANODV7WcNlI2GfymzmVZv72OrHCOxg/iDLHFkvSd/Ahl
O4moeVvJur12dGE9dAe0/Gv0Ls6sV70bwt1XHDAFYi5alQvYAwg7TLrtr7OkdDm0
en+c1H0F48pvxyB6fk6OGHMwAbPDbDxxX7iEHGp98w7hk56V6lrxh2C3nGw51yeu
GeF9k7Iv60OzLYbY+TbWivBDyaoh13WftoJcA5C/zUfhCaTc+wTyvhE4c3CBNjNy
WhEPoaKWkeSM7wff5yzr8kvZ/5r7q/CQ3dtTzvW/9P4mogxslnB9MGG7F0HQGnLj
bSd6G2BgegOQ0a7D6sca8MvdGAMYA0GbUSPVgICk5oZLRZKX2Uanxr3/nqgqy04F
AHwP5J0RFKvOPCnJSNbciecQFYAS/q8D/RWCRT6t75UcHHPTJEKNfQ2op862AgG2
CYsXVRW9Osnq5HWU0Cau0GLdA2bDXX1VwzZ/SvjlnBiYIgvUQLIzqlRXrSGPMUcc
dtqRi/vlPdofXxC6jQ8WqWdjw9LThDTxFHUk9mYw8/uSeI5gF10NpWHXObK84Mie
LeyI1hFmDpH1cuRN4zjmb81gcBG0K/v5aL6WZga5djLHw+ssjcbEYXQMriFRKmaw
9aY8WcbVZ/Mprivys220xsK1R5ngE73BmQfvdLNg+/85+MnIhc/G8zh1CQiYUzyC
3rWKsI/Vp5Id0fy9ilC/2LKBJ3N3cVjaHgk9QLqoDbKSnTlG6K0Z8KsqnjYI084n
Hm5opIcMT6rGgDEeYezp/1DSlk4wBXGI8BnaTgENw70uclPyaKzj+bozotRF63iD
keETWwY7Hlc3x/gT99/G98om4gIk51o1evf+eoDE5CQ=
`protect END_PROTECTED
