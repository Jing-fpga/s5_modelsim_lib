`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TR4QTDE1fAmWL5S7whGgC4LHAk60W4CYWw4r7kzWps67iMeROtbzTyw2ZtBZzCOh
pDJlrRnKRHNc9IAw69ot5blvBMZa0ymI8NtaJjvBxWu6+8vRR8lw+CzhGP1boLJv
js7fCdvHft8cu5uvVz+qbfKYX5CwAUBSv1QkbG2dzCjNvoxi28a3kBXS+ItVS75b
rYsDHtZc4LWYQZ1L9ah/3/eXAPq87gIlhDVMKI5nK/ZHRnbIHo9GjpGqL4TxnzY9
9WDfoPIHOVzkNxFqKhjRwx9ZenJynPZ/tmA5q1C2QltQizCE8hHfMtLQX67OhH/E
jRNN5/SL6h1MRLUcsT6xts3MiFw/NVthjsEm+jg2JziL/i4OiUWD+vZNkQ+k8mru
yX8q2Zt1BrBH4L/GLm/atgTdaKJWwV2+8V7VcZw+D5eg2+AzSUbqhSD7wR1L10ss
2aF91/dzmk0TXsvFqki7Lty9ru7oTx/Om1DAzRshcr1VAc6YtNHhvBemzyoOpjDi
qssmEsL2ucz9GQDd1Cos9KcX/IGYJ1fXWgfBJsmrgtTbIZhayTb0SE5zN7rO1H//
quScG4j1bdRQHZ9bJenCU2lDtd2QOdB5Zvf8SVAvI9kt64kAewSRrwe8vLrX6Ndz
g6tsJOzKfX7lZPILt07Kgu+F4ecYV8vIHuFbqfay5E3FDKVEosmGY4+gO3Duz81b
DnJse25NsPLDiIINB8zX6VaHu0Ny4pIOrqHeMEjywNoy2ctL6A/LV+04xpWpQV/K
yAPelFWHFreRIr3kFblbc6VEnElju+GFD5ZWgvyPvAFzmLM/Ol5XsP4D5VPphaoO
OOOnG/dkTbVSlr0iKZFzGStHnnk/I9UiVyM47nxIhrKl3KjTkdSdB2gkdw0kSluo
5WKfE6zEhp60hOLU7se2b9yFTHhQUF5UWI+IgDq+fi87bObcJUNlPMvo0YGQnc7b
PxWjjVUyRlQf5cpa85fmR6CFMBzTx95F9/DR1xs2brtKIc5MQtYmop6j2lBYm1pb
mDf/wjefO8s9fV9DfLqohsHSK6SPg6x9HQJMz14+G6QzEL15JVh2D/fepX8cGxbz
Len0jh37aRdkGSM5f3fv/yPmSl2Fg21pTOZxQBB7gxaQrXbH18tQAI/CeH1hlwvH
qhMYUhA8clUxs/NOvZpALWH1bqxSGMowFFCD2QqVbQUzp4PRDK5KZOYSJvOK5vmR
rUDwYIj6QtgP02enFOmHoFVh2M3vN5pMnzqM+JmerTe8/47ydtib21eo/wXXHg0D
Gp0GKDc7qBUyEoXPsztSJKuen6eiCbi/Xi8RhHLNJIM=
`protect END_PROTECTED
