`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6oMXFY3g0GlM8nYkQqWIP4uWg3SCpEvDRQNt9rA98cN8ads2+D8veWEDbJIlYQ9T
q5h7BVOcHapLuoUSnWOmMU/uKWr13COAY4wEC6A6MK/hMA8dogtEq7gTP60DrJjA
gi6ApkQrS/lBAEeaMQGAvUIhYAlCR0pbHAAc4C65j0TDwDYDLHM6GlHuwJOdJXNm
1Ziu3902Lv828gnrUqVWqHZkSBINJtm9zE6qZpFimFn/QibrWOEfLuhgY7vj5npI
QBaZmfcTJ7H1fUoe5Viw3VO+OWN7TECCOoURGwEw5HZaf1pd1TccO4/rzoaDT74Z
JrZpNDwcrmoq/jBIJkMYdsd+JeG/ljZByzqhLpTWR39hCYaAaw7+6vcAjgxIJJgm
R9yPnY5tNCdUdnqCU5RbTkdagJmfY3CskiW6Wn5C7qLV2b4lDHBte1mat/pUlrW5
Bf3lYPhL9fLc3VLyTmMJbodJCvmJA0FlXniMDVhbmeA1GlQsPARDBm4lzbqzSBu6
rpLDzrtkI6i5yAzsGYkIy7P5CfTe8H3PcetwigtQJOSj9rQ25+j+zzqITecOcI1u
fI0u5uOLGoHwViVmX/IuJk9PWxFsDuiOZOmRW1vLDaDsIPc1UH8/7SSwz0ljYCZk
z8CaTmUF7rfhIYVDgppeXEA6kFxoeVobwbRgrgufzkz4QXg/EnlchlqdbDwLvJ7Z
7liUCOSduji9XnLlPxqKf5gOIOXruX+I93Coq6Fm1YPMhVkDF69xtJXM1C4GOqE5
wVnk/ZThls2LW0C/YWl+80G6Y9NS6da6WG8eYhRgPCwMqNWNbVHs3VUHYyLwQ8vU
eqLez4EwkgLG010dYn8twTR+Slpotfus7IqHAklOajYGnCwpeBBLU9RLO0QcbTdp
K9eFwwlQhSQ3rugIOmBg+LO8I8IZOiyypZvEEJGKICkZOiQMYPQB/ob4cV85cZ2H
OdWWvcwN/391OLkONduim59X3opzjohQnqbV9+EeyffcHji740dwsLlv4U22kcwL
Simo8qjHvM7gtn2Esen3Jk3ZfNB8IXlAerplaksexcVcUiriYs/pjOi+yveTzhxv
nX8Ib1l5ktzGcV7rU/dz/t+HmOmG8RsE/u3aQpoS3cOBPXb1LHs6NsT9dvf/wsQg
/NeAHkan4k3kHtFC91h4Xz1o03xZKgTGGTB7QxgCDIEPgcKcSodX6Hfaj8WNEYOq
d822LidvK7T/jghInN0ja+yIfmSMxwqzjI0Duh0c/fPV7FkqD6vAtk3d05kEMgmO
yjpLv5xF0BKqWJBX5e6VJQzOUNbfHuWP9h68GCSwmug5/2wGTqPDim3SFFVtooZZ
Rf8oAP6QXtPNFWsBZB8cOvHGG2G/nmCl5x+63OmRPBX/f1vt/H2r8O+mmSpN+eA/
UFSUO57KA334yRjSpRbG72QFuHHJ16/yimd5VRaYtmvOsvRsAzZEMD8Z7J+6xSQG
pXTD9kvIkHjL8r5EpMpdVImMbVYMPPGA62+qcQZpbeEyzD10n+NIUIZryXevLAhW
KwKzaAaymbTZnGeJUoGscXQ7Pa0W0vZxrVCSipV1eqOh7ZWGr+DOd2bNpyEcAYdK
hbixXw63iTIafgIMFbrpXMfObZqw+Biluf0/9jUITBwpAAGP6oOO/UDdhg2Qj31x
da21Mx+Kw5W2OcTLANrnn4OXddRYK409mC61lIsFNI1jlwJ6FYJ2vPtCf2aBC6VZ
/nCLm3DISTxC0aKn/Ypk+cACytHsnzOxa745KGX6+yriBi4KM2sRVBUl+N5a7Lee
MsFO/WSXgeRNvr5CRSauP4ec98LqepGtgQ+ZiWqgdQjU3C49okHdKI12cUKk9ODX
8oPAp3W21sPR7w0SJlotEyvRUbaQU9OaDQFF7ruFoPMAS1m5padAOReBPNcgvAzG
GqjKr13Kc2TGhRAdqYinZQ==
`protect END_PROTECTED
