`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VnkTVav2JtQhOFHFdyb0Q/meXM2wbtY2R7pC9AMhCiPtMpPgqLBzpy/8aKkWLeu/
jH+UKyoqyz9O1hW234UVVd39PsfjEnflvL+RnxiptfROu18EwJPjIy4pPoJADQ4H
+TkHHGLn+VU9JIfyzBqC757MBa/um8Jt3xUzaZn0vGGqrycJMmEH+FBjNtswuza1
FKMgeOwtPZ2b6BMC9ZlMhEpqs+952vXtRi4djXMkD8z0vnstAPFJMqF0/cEiLQ8R
+UMghmA4xwmBz/M8pWc0LbAWrZmb9hEakK15mwQyxY9elOKXphuQ7gyjdlx2+ReS
XI9WNnS6gTftBzuLrdGcb8eeyXXsCv1iDVWB6yCJEz9E4l4PBgsHeZXeo+x+SpKD
g1OkSJILY3b27MqRdv5gee6p7NNEnG4Z+oR0zww73jjKwrqI/i+1c1uKo0dfLVDw
tL8wJZ9/ylpT1G0i3eqqft0SjOB7ss5J11tNXW6YufO59joiVl+ZUY7DvuYiiZGs
x6loDjCSFFwKMtI0hfqLCPihggkzzv/JPXKSPOtIvCUU/1X1ypgI2L8MKskmxf5D
8iIlSNHpcASE6rDZ55P+9Ow9bBGpnevl7V2wUlArqE5AJtFsJSLPLWbZioNyOyoF
8F2Or6HuWn9+hqxeGx9/AXF36jIt1z2CL9/ODXCB9hPD5y1weRoXzjFejji7mP60
v0IGwUHvLwZVuKHVBJug+VQKoVL0IejRoZvXpH+z0M0cWx4gY/a/rXpae0uEjbCM
hp+CyNYAWnQSNOQ7666IxxRApRaqz/2IvW8wKcaGy08QB1nEOsCKmJX66C0sqREj
gxRw4uSCyK1cLwbwwR6WrZ1oFwK8FVMckjwKpYJwes5PdLzrXdaCgkIgxEvjTiG7
1sz6hWcYuQdyvxcyEvE41BMpgwBPUf8NboyJ0MbD4x0MfMHTl4xg61rKH26vJ+IX
0xgjO3IL1fU4y715MmQzFElPfrg4cTLfDVkTxvvHGYI9ZA99hFtMlWmBFiMVT5SA
yPqikc73pe30kWKIo80nC7ClVJol2VY5ytcvm5dU84e9Vl5UUyiYIzxPiIj1AlUr
IlqQES/5qYMc+/LnUePtqfi8T2sim0tyt/06De8r/iao+Zxm37Hc58VK/18Xj7IK
csylLtvLnv7hwgl6PDqJbjFffLZAJKAafzIRpUbLo0vP+vIKCJg90cqKRDnoS4e0
jxnZfV98FzKyCADgm2sszTBLF0+ih7fAGMimfC1zNvfCJsFZkW27uIr7/6yRG2kd
eG5vqOc+jeAlHCeGDNH9T6NDcXvbsZryMUvBsNB2RvVCOrj+cCQaTY67wnf25wYc
CLMprHIlj0gYGfcNkrBTElnqpydLYCoZxCnFw3V3vvEx/IW1Z8wM1dOMXCJrA5fK
qxP41085yc9hHp5e4TsChYLmOOhf7NJ7eaP+pFD32KlOfH4W1w2yFn4iygpe4snx
HJ7lHoqM5eUFpL+urtgg3e9PeCZOazbQqGSA3sKtqwDsvU/6ucDGs8lUePZT3/s9
010lPrzCLX+hlmXdTjd0dhmQvJ20RzKBUM+vRCT8bSm32dHPLx5wvyPkKVmjmhkZ
4VYafpEvbxodXuuaSCBais7ZtcQBUYoXmJ6OSW9E3Kavf7aD3pRuIkiAEjS51eGd
0t73BMC+uWlx1X4AtqBqcMiowSh2skmw8WRrK3Czniqni6wSvQJLUW9yOjW5LZRy
eF4Pz7kRaVLaROBfYFF3Pz4s09XsOtFbBfDRXA+Be62d/8sL/CiBb7D5XVde2tdm
V5HfhzKJw8foVey9gAJTI502uAr2hn/yCk6xlZVMFETPosr175P3soy25b/dbj1M
Q9bGrMtlo8Aj8H5iHF0r0wsLZLCpg1V5sTaUQn+Jc9YkplNMNxWFspezfytqp7MF
NtbbWTEZXMDx5ui7jdbPuhJCSaYpvMjne2aNYAs9fLKO6iUd3EeLqfrsavcZC5u0
B8O8nGi2LHp+IIB5RGhwbW3R7cNlk9d/Pjun5eel2CERssisLkUaF80HxuSil7RO
FXlpf13GDxP/vTewMEb3y91iiblCorP0m6DoBVi1Aqwc2sYIHRCHu1rvSpH5BmRj
fCgu+ww7m6JTZk7xoGlxawq6Dtc5dpj7Xekpkxxokgn50zPAoR4SL36ADkGqF0co
IqIdGVzLjBcfMN7vtrNZExRIAjZDLWXk/Llo34xM22KfVT7IHrpmB8lHxaqbLOsM
p0TK2eVszwB7QWeNKi+UCRqBeGMn/1LswsZgw7gv61ypFTMVa7zVJJ7Y203w8aph
dHyK4DW1krpq+BYp/IVq+P6z9s0FWH1jG1Htpj5/qc6niil/Robvn5NXYc9S9cwA
dbXEAjtTAxI4vH7mDLx12MyJ2L2MImjLFHWshf+lJWgqOJxhNSlpvijFd/Po5NQM
xXCymSCBA+NoNF1DFJY7qegFlH5r/PxzatpfB4etMcr1KHbXVpZjh5TXxk5ZO+/e
NbuiXDzO86hrfTg3bTFaW2DRyNLr9uPvRiQWTRe0nEq/EKtJDXMbPdJyxp7oclgW
czYjhs7p+hk1kqEfhk2b1Cv3vK/QUBuZGonPMhAUPfT7EJVrlSEGo5K9/SvQG3uf
3sGqW5PJB2ptvLQp6bKx3wgoFTCI82Z48WBiqErqVkUOA2sZRuyig006fkWBCe49
yf7KS7+wgwg5LK/xLcrOcllBYU+Hc4IwMr1/XxMCFpEiZAT53vcc/AkVJbTnZTUZ
f/depLXB8LbpRt6ctF8o1nbtP2nHTOqAn1G4Z8C04m1RcQna9i7d6+XE7NrU5kBB
KAD1xQm5MHRCaI0fmiuuO6R74R/8KZ5NiI2gx4zVVCD6xaRTBSaSTUKlqVQmgUOs
TGA5AF/9HyUqDSIC5wmKaQ6h0t6ijSol0jruEu8EuEfAI3Dda7HdTTNfGdVp+Eim
a4427izJcZvX9owaok/xvRaXUVLSj2KeZktlTYmboV9od2J4EKqnv0n5zlhe5lUj
m5DjEIrfTujUWrj/ZAoI2+MG2ARdp7RuwNmI/P3XnQb1WJgK9LZx8QiD3aS7vewD
nOU550fQefKtdzxO0JW/kWRe1CDy2T+bRyzSbQ819yEojAw/8utKQs943l+M7Rt7
O+O+A2uoRilQrqeQd3ToSb61ewxFMBzDlmW78dkEuTx9QupsV3VKswemgRsa0lcQ
b4w4HqjAp9QTSWegliHfPP0/7gbHu45F3BHGhKLUrIn03Ma0IaRRqsbfBq/QYbvH
eBR3CYz2kkwlWmTtRSHLeSb9zOKSLiiml00B+7HKd70=
`protect END_PROTECTED
