`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zSfx3YKlg3KIlwZ4SSfTs5SQt2xfQ/cHcMt4OTK4srq7sMUqMUIphAIRIRfTTKUS
e+ZPkh5HrQ5Giw/fXlrhGFGLC+ADnFgQHlf9G8NcKy+jAdzUrIG7X7meSHIESLFq
wLZzOTmLMsD6aXYxaEd/E6kxUeff14achccefq4SAQ6UbZbJQMce6Edf3MN9GLKb
Ni88G7W21zEQmrWCf7U8vAwO000JLtkHIvcQuzJPWcnUp3sLxBRbhEPQecrL1eqx
8ikwgzElapEZWC87z6tsPSCebQwlYAgTvceCpqm4NEd+90ZC/UwZSmeoeaAYMZBq
orvy5EOCEnI7MBjSakuLYfcs+PmFt5tnqOosCtoryX5IrHwSKS83M90McFKUwA94
ykyML4XIYB2241eKS1qXrStL+ZDxZHeczvNdHC046OXrFL6P0isZunC9Y/hdcScs
pUTL7Ak0mPV1alXL3KcMwqRo4yuIq3y8JAi1A+YeuEJi1iG0MkMLk8SgFJvGdJHD
i7pcNHoJpbHm/aGYwjhhL5ZPYEHeDRQB7KrziX+E/TOXYukwXdayP5A5eFFx9ma0
Tw9773DvWwWAIspuZhpYGRrcsBN4IXj8BqRxKRnUbabr20tT4goiVksITAwGgit/
uFhKiaeBVx8M2JoNkVx2vWTlL1XrdGJvKNPIidjsmwHs4pjkwyHg5aBHPvDLDoK9
u/4PxVOQ0u9mLFu/2ozS6V9583o5kIJHOyoXyHs3iOSG6oSnjsGAV5hq4Y9mbUTt
8m2Q+ISy/Ac1uM8rlBFgYWBeQuG+a6CPFf6hoCKeFah0fbbrbS29ybzxzeKl+mgP
cGAJxN86D+AJd3Qy6s+TYfdTUufSSMUNwSscWZ89ht6FqGJGl7c0FuZEoRLlmttr
zejTENLPTrlUoiqGzVOu3PnTSEfxxW61lV52cZ0M7AKFBIu2wkbDb/NoJF25j/88
4iL2j0nVXHOniPZtNc7x8ECUoomm4cD5DSCgOXBxzmyT3a40d4joERStO48IUM/2
3BV6rDerdyIpxvJj9ebvRbb3v1eC+X51ijyrvq3r+oCs1SGxTBQrl3NEP220y+Ln
csbyjuAnV+2p89gYJ6ZsakkLxlZ7rEH7pXcMl/c1P4KESIYVb4d87Rw3Nv1hJELe
yZ8Wt3CoBbIG6xs+EXSIBpXjR5t/yzJC3UXGULGkQ2S8VEH32dWtiAVuXg428w1H
neXc6fBgr/Jg7bAz2IQefS+VjuspbpTEhEEsZE1SpTZGmHvZZmnenE+w3x7b1e9O
osM5AdcFf/2IriZFUa3STjfRgZ8MBSnFr6uKmbSLLykb9GrtM1S5KINe4PbPj5hM
Jn/nIvOYRy20m7U70kmI7bHsaHFTyvaKndsY9DcpBj+GeR34jFEBA0Uo0p/b6f3s
OGxxFiGKKgOXkDUZxfycDrSUPQ5KhpgxuP7cpd8z4BQK7tPi9VRhY2jmH5IR71qD
LXPQDNuf+RR2GbnQr2kC/3HH6YnOm1iFTH9DX/y601WY2JMKljDbboaQMQXZeAvf
TM+yuwrbGaWbj9XkMbfqwhcx/nsmPdrobPk8jJ9yuAQDNL5mczLW33j/IuqU1oKQ
EwyltUYT51B1gzaaN1mld2xs4DnQ2Nq5F8WhSc+I/s/HmnFjAk772B1GWUADIACQ
OF07kQWpAuwZVEZ1rd+09KHQUmfMHeudxuutW9uTwykRcjoUjolFuzLoNa3iSEr0
mWVysuqLO69bzaaT5bN6kmtNYXjg8LpTV32Ym6wJcrfnsOAV9mAnkOppGEE5IZ7W
qYrphVIU6DwwVGbI6ujmx9YMbbYWSS/jG3UI5bx1FS6IbpmEy1xh7vPPFEY4AA8B
EQpdIPqfvb84aNDhHsLfhfJP0BYNmElldC6PfzXZufbrSUravPXqJYnQXeyzQ/+N
XbQv/S7U/Xx7ev54Aqad5un0bBgttE+c5DOm2VtApuBYS3vB9SgPkuKP627eGiHZ
snean17kP5q5LkJ2u1Y+b+wNpRbKqkYY9zIbdHAorzyUiISdvyunCWGxS9tGyZSD
XE0+lOOyqNnq8XKTxXyEugwJ7xX7ca5jso00YjAF822aXJnEoGyLSbOdGwqxDHpX
q0s2tygZf/YEOfnNkfRSHRpc7+WHAPI1igYJa1X5PA/DpXons3tvtxPToAOY/YSq
bSvH32WHrt5yKE5wJDc/WJMzCHohvVkFquCzHswIh+oXe+H0PgVpKilQQJwkL7OX
Mb4MAu/Iqk+eNkj4UitNl+Wm2441MlrPclc7hPrh++2J7oKKmY6Uy7pRlbrLbMaQ
fPquPDz9lcGPdbWyJHVvOHefT6D5b3hvhQ7nfLzH+YVaRADKAKYzWPMRkAVm2dFA
tSiD9WMhJqOWa/+HPLXIuLyvVDQxmxAUH8FfXxQhTLtkoSr8wJdaMC+RVraQDO5f
Q+P959RcotzVGOksWwNA4SsSLfk5rh/SjwmJ+Cf3+yMxWuwdAgxqQpVK/fKsUla9
/U2YXIep7Vx5J6h/dK6VFLY5slDpNzqOBujyz8OlWwJeQwPIAaKaW2k1psI1JeBj
yjFyWceqZi/+LeTujiEjjbcnISOlrRHDTN5Lpe2h7D4qykzhy9hjZP9+Ce4yM80M
HirmxfbVu+zHnRk5SjG9/C9tiw/xebZWNOYKG2TCNW5trW7rSMxm3kCsjUMsoDqT
CelbL1K+2MqGuJrHN4gZUNobc3wPaVKCfnsoUt5D7RuKfBmrF2UbKZpvf+pebG6x
Yn4fHvNZbFHCwSbqm7CsbYs/RyAa/Yn2MvF840joMmKefDG+r0QneY5KjAV45UDF
g8970MYMoWGX67xnUAq1ao4RG1yPRBmSl38nM7X90A6WKZhRB5Xi0ZTM85wQCv5v
doXdGkgbcws71yEA3WrfbrKsvVNTRclWhPtmaLRveDTITYnWd7ve9i6euinJukI3
lj4W6u0DiwXwWZ40RwetBnZ1SS4INqun5f8bIJe1cAgVspdbvL+WxspGwbMxLcHW
wJrAab4R7yq3kfmh+OYC30Pze3+5Oekl2q1KaoPHjhuw/2iQ5pOQ+WEq5M+AeY+X
TcX18mKB1QpVKUb3ZFuvTXtOwi4anh+myG8+QidNJ2ePb9jFRr3sFfIegd+R8Ywn
KTazQ/b7VM5P782sa3NbhaijowptfPattoSt6/8c96gi0z/DzoEQKBx/zDhMnoVi
kTIO/SSghVOcbX0D6C3qGOxXuTmnr8aws1KcKzxkKFDrhDcL1wFnHcmMf+T/hNx+
S0BXDvle90yPvufOS6LbMGqbzNdUkyZ55Ggc567SgVwVM1EhpgMVxiFtuwoEKgJ+
2NRngM9m8nfXle/XQNTSFlJfElHMfN6eDJNjdQwKuveP3MjhgWdQcIbXKMkrLIJG
peCg9cHr0M/Suc+3cKiQWbXOmPw6lkBKCWVIAP5+3Ez1rUMzI2Qn0qehIEJozrXc
0kSy1XzguAjof1lqIC+6dN/yQuq74coYYNYrOK4ttMupdWnbY52Ohfo2cTxm9wcn
L3eIr3njeOIrs2uiw2TbMoDg0hCcAi5Y2BUE17biQnvdM2xDzMTWDb35Z8dOggx1
0MnH7FireH8E/0KIfU73zoIBUCnVoqBeh18RlDnfQpvhSfJu5rY4jDc29ca6ER3t
OKe5n9Fh5oWLNuWtTc1T9dBO8mWLMfpD/sB07O1cUUJv22/ViDpQ+RPKWKofwpN4
/GROaBUXYSoUJuHR8BInoOWfH6yhpE7ZV2QvzJk/MjKquwDm22EuCQfApMFQfHK2
04U458UFLvmrBgoz1gshS4NeDARYV/w38DfCyn6VSarTEey4UuAka3U9MWX1nOXb
42iHHEnOrFEURFAdOPR08grFwcsEwI54RPhc7YcI6OkXiN0OrKU8oEPdJVVnvKJq
eYkVjyOzw7iccf42pt7F0ebng2GPyIZwFVld7zU1ISe2MXQbB3wtAIeO5jT84YTi
HPAhkSdgygIXs03hagpq/ePQLHFTNsxUgUN50nf8liEpO/EI+ALXYcw30aixUWDM
iHL5igdvbQS/sBMcwXp31D4hysHgURcwEl8rj0q1Z+v4h6AYLoIvyzLR1309F6Qa
KQe3JZoloYKp7+DgaN1XUt0Lu1AYxakpcQYGGkC4HglF8Noh1mTI1X65OFdPOZDO
JV3uIpUt/a4EP+1D4Ilz2Rp9WmSi4WvekbAbMr7mVHYGS4gpTIEXUOjR1BKtPVEU
Pdnqh9lg6ZTd//maQxa1vU00A5XWPo+0+aeJcl1GnNfI7ePvUR4k+zIfiDZG7UXB
XpvFXqANodpIzR5066m1OXmLuFXjXNb1sF4JXmpdYR4tikBZndhqSgM35/uHRV+x
ZELTXBQbnNqTImOsrlOQ5QwQZD4VATuTPCAkKnfkEhGGHVHLVSv8LCdFJ6nl4vDs
Fj/rLG8iesk+oQcxZMk5GYN/rKhGYCCbW4d7ww0H0vaDQrsaW4FvPmnlSH4ZALMa
Uxh4C8ly3jiV6I1f/coHitKoeg+VXV7Q064wF8JGXc5joJKpd/iZqSVgkglyGU1H
s/T0qU9BJs21DMNQ/KLH/rT6yL/2646togCR9zfo2jijBJcf4tSXAgHQcFOiAPKU
xLZxIor6F2dwXhVLmI61c3luAlswLie52E9HyaCTVcZqGyNA+P4YU040yqzPBgyr
U1bAO7W4jpmjdVBbFis5Et8moaKDBFcNmEs7YScP1YuJdJxCTD0ulo1LFTVcAPs9
s5IvoPOzWb0QAf3i3oP2GXZMbXq+25gMpfHFiPTbmpcOgxpam1q/ZIF3Ujb927Gr
4amqa2cTL/4D1wN4K35zDnyU2WzRBOJZnpz+KZlo8Xk/1ty86u7/w+OcKHOnOuVM
k40SZtdKHPWVu5FvMC5LXyguDJMw77JQwLnNRh+xMfedAQjVqh4/71iJG/lur6vC
fcI0sLZRvD/qMZ4HUwp4nd9dMkESF7oDy7D++/co5MX0KH3K2Zw1ZHdK4zYEe7dB
eOh5T3PL+aOYO70HgQE2Fs9ZgUu9xiUzj8ERS/RFcqivHWp5UBg+QFJeBzO1bj7z
3kWLwgrRlg4PIIKB88EOjJ7jj48mx4ryAT2zCF0qwiR0JIJWCJF+KECzfvh/CSQn
2aNDtj38voBzwqayQNotG2OIwCUIbY5tsTqAoa+Ui7NtI0TmG4+/Fgxoe7UayE/f
A/Asx+tZ0rPUqrrfuD5jZtqH8SlxRRVQ6Gg8bVUy9NnBLqCj4rQcVptbvUeQaIc6
YbUwE9E8cTbLlvhbj3y8F9Px1Cvq7HCyWnsVE5n6Ki/TYdqryPwrJkH0lYydv5R0
J2HdcEN9wVSYpCeTzJlxeuqwHlmwjRzx0LibDsSpCw+8oL2Zjlfl3y4L588SoZib
vav1pSeXFC9iorETFRRT8hZCINUzfYY6HP/5h6p7j21gwo4vK3IKMS3a9jwf7Nd9
HTmC3mLVabuBXMMX8VQJwQPE2S/1UTzY7h64p0OCgyQ9V8gaSgbs5LO64SNN6ox9
NZZkEY6jShltNg9FDTzL51xnrPzi4If7hCaTBxM7TnDi0pP8fV+JxEAxQD1ELB9l
4ecT4uX79Eu6tr08Pc/7mJB2DT6MuX/MwtRM/gDz9cjYpiyFh6ijMtlK7i/vurEr
JApPF8gUalqcaoGnKc1W6NrOr3QPM4rC7ucXNLXGE6rtJvBfbUh8umSyd+dUuEhV
A3zaWtlbwStoPBvDHDoT6kfUem17NrX6tB5FZqAP+zNzDL7K+Zs1eoeFefolbwqV
gPIeflHSHo2gweqxD4UKHOxCZM4NVphdFIGeuq9PLg7GjTmG0Yq7KTcXR+AgfFT9
aZUAk5UAus2CdNNEy7UmKnJvNNej7+mVw3FdcBiMhDKXDEI9yw+5wuNpcLbS73to
qiYggtgpdkbvdPRI9ZS85PDyl3HH06v2p024+x1x1uI4hsfMdyIqjmxrhTSCkcXX
dEeWXGISlxgvKOTCrkY/Y+nYSDJjvCbREVq+c2N9NgxUtTkYgzLAKcJIvlqaWN91
KNlun19hRhQMPej01Owv2Uf69hTVcwKWI2l3IsW1knkpFi9fTlA22mgc2zq3qH/S
QEL0XPcI0a8lTJOq5Q9lBddJgCDj8DOP7EhW6OMZoSeNpPmONTGd2Q+Azy/8FWbH
1dBENNXQVPgfYUNGG4Q5zp9X7uCglX8xPqxmE6njn/cqSFKWdhcMmgYMcNZT0bIy
VPyNRpbZcgsHIA5nfxgPhyubCad6TE956iF7vv4kfMO99zop1MNQnN1qmCaivPHf
PAHm12HPWuwzx1PYWfxCTvmaeT+JJ8YoISjvJmOYwd2W5VPSBBjvbjdgFxhjnIHb
qn4rhB/UR4M5WJJTPGYlec/elFq111v+N2QmA3UqcvjAMzrgweluZoj0ijmfO+k1
b/68ZaXLoIo1JFpxf05gzwl8DGVtWLCnGrr5QpW0hY+o0Yd6F5fdd1VLLtJerapV
QiE4ZW4zItwJWeBAFgNpVKdt9n/FTPv+jfVQoJNoyQYxoAV5YJbyQnIxAE+m0XhZ
R8ByjD3/qFOOXuOofsbm9bS1iil1vbeMkagiZRKpywRtLpOOwE4COZh8DBrjpMqt
ddH69W+9NJoZ+Hwgg+I9BUius1gqLtoE1z6b9i0cvuM60MjKBHKYZSl+6NBl3d6K
3GPtUw2Yiw6shOsZqY/pNu52wIbHkQbm4qHe8fnyhYSRl+2byVeW6pw2x3ZoBDG0
LJKGQVWwIaWKlbqu1Etgn0iEV3RfHFIJZ4zYnUK+FUGNAJ19YcoxHBLhiMsQ4beg
eUplrMOgYHKGgGkPq5ZLakFkxNiPN6NvzlYr04FcbqceVU6/vnJZeecC/1oSRASD
ZKkeqDjqYavtJ9cnK+TfYWhhbhtaES7063LFMQK+QRNDXnKPXZaTLuTPRyUeF7QQ
zHRm9SYxmt+lN3+b+zepaN7bsfO6oU8AZB09eo3E2OjvHJ54adbvNqbqmF3DrG0Z
ut6Fce0Ax6lLG7SxToQsYuVmYiYOs3nF3PPg9e//fN8ElZewLaH7NJnwCb2ZiaXk
nKbxSgGsRGM7R5oPn+gwJyW/j8hGlA8/ogmxNI4xP3o+/ZLBS/gSSKp4y+z9NNzV
Nf6OGZ7IcYK5OBhg5/YVQR/5zq21ASCaeBK8fSCpH4fyPSBdgbUCr887LrXPtH0W
z3ah46QmMtHJ/MXWt5fLCecd0QHGRT4/fiuoZY44ZPv1QHxlBXg8s2J7DFkK+0fH
RBl76FWCKfEV022VhFOvbcH4TeRhoUMenhEycOtaio1Mx3CI6ScCuuw/Egd98hHI
uBM31Vmytq6gD4/Pa25rsQrK+2FymVn8CTZndmYcbCLrLBm3XGoL/jPww+fFUZE7
ScEjEMh2Y8TN8CND4N6STZxsQr1jVqd1++D6EDoTqNHVFs0v69LE2HeJ9bofT+Kq
Ta6PsJ5pGg+sjErynbsh3YrIb8tRkaEZkojHscOrqYlODa1BwCwmP9lfNc6qMhRY
SQVxQ6YcoGt8SLD+e4yZFi53V/xNaYo0h7Pdf9N1i+yeVgWTxXNYu8Q43TiyiIFk
N7gBP8LMbY8lry4/dvVgWyHjXP7c+lnQVcx17CKO3jWEFGHNGhU0OgW+PDOLAGmL
RECzz57Pxe5rWlNoNX94mvt6vUViiikdZVB+Q0Mtlg7XPqMwE+rV2uy3wa7Uupfm
gvETG5MUAilSGaiMIsqjIMEU4D8gZVog1Tjv1k7sve+t7WNmzKtpEHpkC+AofiWZ
PeJYg4q6El3iO6knOVi9GCiPkXPxOBgkVfxx0mlZtxxf6OCUp8RfL5U9Xy1GI6Bh
WRxyOGfBv5x4l/k7f0gt02gBt5KtlFsTL+OayPULDlUaEY/H79FPRp1B3HGLBzaS
aDE8Di33GNJ1/80DWDjQozsn7BuIHtOA6+/kjQWwMmActU5O2bJ3+BCq3NbUS//8
0XDuhIZHfR9gU4uWXw6YOStCJYgta+B8Nk9/M7EJYmWKDfICyidmuquwVEPFXTKz
Xaltc6sMd2hiORLyKAt8UuACxklp2pyxUFHyppHtVrd8zYWfiHuyo/7DeIVMzXBc
jze0tmIuHQi6sjnKyaq1GP3LtqRJuSaGKZ6pxCThBp254rmbhZ6OaRoYgtSsLGj5
7P7Iucu/PiSCEuO5X4kG9dnTGUegc5Lt33bp+M2e4e7SVlz23kBPDUfWcgYuxHay
zJwEnGGtxXJUgDR8k3QN7tHuce8T5srhJVs5ZfoY6pZOwfegHpSU1W8BAjGJuh+D
J3P2B2a7Nousdd2U/bhSjvrip0qMfGQXoGd5Kwy3iBOV8Q6NuyAHH23aagAfVJxj
LlEyXP3PyUFJ2ieZyGR6L+hYKGlVDjlF/uOjbHMz9HeZBh9iyID9azQJHD7MqTZv
FqL6bc1Q2c9Iqe79qcAjwB+sEJQsPM+fJY6256A6BFiGA06tXwO7YFT/xwTFxLqm
H/rL9rKM38mRuKYqeoyBwb/Q6v0kadHmrrnmX5G3bSTHRYgQXuzIm8ebDjGOSWDh
FQvKPFedVKEtYBRCUPmuhqT06IFNHngkEoFJfCXAyLg2EUJNHfsNNxblklJWwsq6
+EsOiWgDs60DUfRf2u3Y4W8WSBrGS0johBvcuEiZMPaQBwcy9nmVOeQOxPWdDlzA
pMxxt77sVm14+YUKVt9YeLSztOWm3vnuIunWGI/BttboV5/2v3vn4juqevdLHYxO
/x6pAz/tF43peYab1LzYzuhG2pwKEi+o/hNp/3kAmQXJm2ZodvtIIrs2P5hGZ2Dd
x44FSNBGu+o5pdqTSS6ix9ePlFLhHhfM3AoByGPOGsXWNoYifjZ0xapkByLfhYIa
+4u7QYockDrVEJemR25hwBKIPrYCjx8hr6akXGLdvTjc7PnWtgiD/H7YrmNAtYL3
RO9o6JTXQvrfk1CYVWNCHBpasey+qtlnpGGav1yODMVw//x+TNPj73F9Fx/SJrs9
9LZxVEoIx4TkABNp0K0tTCvlTgNVyUmjHrcXLevvWgqkqanIRMorF8VTSlkxJCTx
cQxBEraonHnJzqMhnt1PcFewU5raXP/tq3+G93KUgPRBahcWjasWR7lJEgTzoX8N
zUxlL21WdlNZBdjafieRqiYrlXGc3F3+HZw1hdigUJ/Apiu8YMN3QVYcoPJ1yBNt
ksIZngvM3Xl5WvEb9bBuu+3BYJdh5hoqiGAkH3VDyUhJZPJNdwSmgTaRhx8OSATj
yOtucfGX4nbqTTu8pW9UKNN8jNwOpDy6oiQIaeARy6ZJHddJUhvcRsNr/8YKDKcK
hu5TCJ8QMQV2sInp5LJctL/eJtaKU24y84DNkXxWV4jiRywXwx9bNsHToskOJcgg
57fWtOv0JeIKVylAE08xyY23fSVSCej1eQjO89C850fNoFGlRrmAeY4ZZw9V5JZL
AYabXjtgk1KBKWY2bVHDbrz9KZTZ77B6bl6U38ho5M2bEg7OyXL3QXygoV5yVyMP
+x4p3p6OORi2C1X4D3Dei2+VLBlmOP6gJBn2kLGJ7cJGEof5a63+oc7T6km7nRsw
osWXEJ6x9z5UbFLqmIlFncw/GtqF3SVPT7bU6H73ukb1fiBQED0pzWaUegBfGx4h
3XYB5dkQ6FI8wJsokaQGL5NGaUpBiI3WM8btWHT+5jedVflnZ8U4GvQmpXgPqsA0
6whLD7NUmi7qO310UfAlIz+6uJBkIJtjlXvt0P8ClrM8X4cp+f62NTHnmZnW+OJg
puPqHROiVFVd+gF/2rXAOp3cY9es0v+sd6CQLGiTWQ6mW6NDC40POy74V4xcO2pN
feF7dpzBVh82od9KQzzmTIqbjczW2OOX8ZZ19tbyttN5qNTkBG9CSIrM3jxTbQSK
FwNwEH086ka8BscuPo7dNHU9LAFjmbiV5PzvyYRXZEaUy+98aP0Tz2sfYHj6YW34
GIajqa+ZdTTQeo/r0YMGnZptbyjQfngdjGZewLFi/NpjkZWaKuYPRm5igjeJ/lvF
yozdVf7Jf8yNoLV7dThor+AuNLSRcV1TXjde1/4VuXl6q6qGwRxiu8SLZBeE5rv0
Ioi4DF/+w3gOQ3Tfss59Kku6A5AKvEkFmvbdsdctusoLx5XtxElU831BClJU8FLj
+AIXUu6TBAOhis9EsXXDyu7R8sDyIj+gb9bhSWjKVZGrkhK4KOs/LLelhNp2hpqc
tst54juZVS6PGQyHFof7Qo8fPgF5dZnn1xVUlQDsf0Tvnc2qtUlHKFCjb7ywlqRQ
EnqPFVPtbs61e3iRoTnw25s7dtnH2WrgqBl7WccSZLOoa81vICUd/KGjQbWggp9J
/Rg3gGG4Ue13otG3P13If3jN+03LPnYSgz80LmJzYH62kU80bDm4CMNO4GKCa4iP
7MrWzpR2Yja8px0vD0yYK1VsLTCpKrO23H/YxT6JCgZ1vg6snAlGaQ2c73/E0fZ0
HggiRicLD14VLkF0F9cy23n4D4dIlIfiT8bbMu8YXVvz62KPN989sxlYoIm3KILP
cXP3+Ofniq5j0Kxwbi4EfjCwqf7d1gCo3KYLI37eLHMa7qsC4IePeDq3ZhY4czEC
EXOFrbb8AhLDRy8CUSRtPjSRet8ViG5l4pS/F/g2dzul60Mh5YPr1P2lRxp0YYeH
pAyyZKvXfOJcItHDdHSbDdGkSIXuyJvmJs6V6mxBhK3e3YlVviLSxkDDPPZ/4O+W
0W8eEyoFRyrd+wZuzrdR99PcK8VZ3H/osLO2d8l8qZ2brUEQjUtyyi4wYmrzFyMX
Gmnu8qHvJQmn5woxNvIr54YuiJ7gR3/x8mn+xdNYdRsqgUKr8ZE0mD164tltTNkU
SPMMQSj32WMAaRRl1Sw3hNfLwao2L319EH31Xt3lb3QBGAmCaRRiNLsG5W21wtRS
78nsW31h54Bnj3rsnGXV2BIAryEpVRu9DzQwkX5o3BEnPiOqlh6ZqMJrKdpH2SBs
LeReJCTTPbMPhMKxrvWQa0izlKBZOQq/AHl/ob7MlSRIf8Fev/mwfzhhfNZw71/K
L9wHx5lDhWxJOyeNGdNOnKyJsKZ46YRwKE8cez2CfkrAf1aXITBGXMUr0ktcZCDE
bbOYuBpbetYvv3K8BwXyDrglGzNWgsFRUi+PvuMEkn+GAWl+Z+1dBONuwTrC2Utg
Z0ygtbWJn0dktrGi+mAx/dp2N61YS/lB8+MlDgtA30yuSrQ570aKI+iqQrJmR4Hv
xSnXsfXKsAvZZDw+PCq9HGCHrSiPCvnG6gfzD23vW9T8MEvO836OQ2/TABIIWMx7
L2cJuOEhYEpTiCSJvY7EX69TvhxDnWVEbhg7Ltd4plwKEcNOid1t79Xxyd1K/qln
YuznhyjgtkDH58+gzjQbxGgvG3HllPe5O6QAo9zHivnIHZtG8g/9+WCYc2s5rvVn
iDVSjeC556BTVBJIgPkwCCEyra9eyWJ85qgFBchppSrPNHUmnfoUOD5esVE6aScq
rm+nssccCOKAiOGPA4IkvVX8vW3UYQgDlCz9gHGnzRwGZ7Tm3kuC5xHdo0deUQI3
jXTd1UPqw7wxosHN8GNqHPZJA/iWQ0D0X7ImW7lf0wlUZWEmybPfZvIfdw5JCFTw
6yY4n2oLfqcnF5Ep45XQKpS3+pvIPFectmgl5IzYhbQopw8VwXMzlxTyd3msspR7
bRy68fkuwPGnk3HAltbljbfN/oExIxvUdNqDV0a297BF84uA/XR0nxv9y6H99KvK
7iHbIgNu1H4CU+yf9iicNQ6MVcOflz3REIoGNTcnYVqa+i9hUu0ulg5QhfXUn1qL
pXM/ysuz+sj99S+Mn48qvdHNgnt2kzcqaEgqcf//CpVrIwuWo6nDHzQ2X+H0DIyT
U6anIX50O2hDPc6OqRdL7YnUFm7spSnEPwxS2NNA67TLwvm1hjlLjUpL2f18Be0t
hFQlHk+Fwdbb5OMrhPLkJrtyCHjbIld13JfADb3HINha5vsRq6w1DCKqTIuQsuCe
57dXIIFTD2w1+zqGZaeuCwpVgOlnG3kCTjgNZMWycOxnUvc08ff8b2ig7EKKqD80
MshbiZw/9mdmGoa7Vkr73+PDcUg7fw60oAtoLqR7R3JFy8bPUVG3qpwJf5cBGbMl
vIhwgXJhuIN83PU3A6+wiRX5QouDU+tFVc3/hB3iRMfhAV5Qck6i2iWCS/6gg8AL
tIq/8EZTGb8PPboalY+Ny9RS4LgZavTN5AD/iCPADb2FugNYjf8Hv27ZnQL8ul/W
VkgIm3r/9AIawNj+/QM8bBXuAdyN9K5muZXuHgBy3739JKqqPXe3ged34UjTGvGm
t5JiwXqCUwr+tx8XhFdzWqafgI1nrg839XBQuU4Zk7cbN0fi3K6RZSwxBlPQK2Af
nfdMGSLVAo1MNhJvh5Hvljv3eVUuDDs0+5jVnj1MIdkFhp7HlY084eJoNcCZeKnJ
JN3kdU1RFOlx/jZ7rUNCEb6yxk0iF19da8YYYy9qHJswj7rdSLJ3Ft2nk6cY7J3e
B9YPA697og+guYAoPwckUgimhwWElFHtasMQoqAsd3Xs55joUletGYsOSLalsZUm
ICX8S3IxzihV7ePMtUlmr12waoYR3LvUoiLqtRgKJ94rEJVMxFQCmurnsDp/FSyx
m6jaJEk1hbWU9LhK6ZULcV+WDtqMeOlbCKdFboD+Oc710sgdVBvPM8Lydjy8KfHu
elRt55rtJMTofpCIAVgoIojlcOWlaaqL0HhKxr60/addwgeumrdgGnnjvm+2BI0a
mJqx4lYLAWiwLo9HNIU3rpAHHxWP4Vnkv18ifQEPVUlGwUNwykHMzxv9UEiJxsp0
NSqeFgHNpwCp1lUx0DQIDemPoF+tdbiqaZ+bLb62l+MnzHNhbTktDy1YrJTiQmZe
Z+YLQuSdTcnSRPdnvV1Nhlxp/fCzfh1NifuGu6+791+m2H4v/F5IgylQeg8vGzdm
pFyXS5z4E02UnD+xd/UZMQOikHpNT9AkpUS0XeryzVwV1oCtzdLsPgyMEdNn+YZn
LU7G25td/rcU677YqIuyg8SSUEdkOp0ZueesxJk+lUyRnib20wTtQqE1k9FL6Qhx
b2rWkRhcAcOsnNWlGP9PuWUfetR0AEkLgLOkdMaecyi14nxwXPTZmkwizb1JayLP
shFsc+yYuhmkM/bTJxIirzyKZGZyY28sQmn3lH9y/SLQLO8UbXheXlX41Tm8qco1
ttc/lYhI1W7SRk9AS+xO1QFBI8sxUCc0oHuesiGlWImwh/X+7AbenDrj09J9rRIK
J+WksWqEsOaR/F796wGxawRKVl6YqHUibaW+dChWFYZjBqq7pwvNnntXVOF9sov9
VzKs2gUHh/pliMYTBcL+T4xrfmR7m+KyJE8vgscQWj++q8YT4pfnn6LiPJBnj8yz
2hrtxWI+9P2b3u3PdHPZlMEDTptrUd5nOg9SoSIyECZXKiufH3YQmC9mr07RIBNQ
ruGK0voCUvOIyHyN325lWgwWOz5QTz4rhm0XFHwZpUX0Z/gucCn1ysPW9PwlpzKl
VDFUUhh4f1QVTVW77L9mKAKGc6U30weYzV3A/ceMzeXVzvQxnp5IBEXlg2UDfsYd
8uSDgSc3mdCEcTvCt2BsQWc5UtHTm+9Z4+6wzOAmAm1H1hW6Sh3ptJxDl6FOt3af
0L72XVksCxkf4o8Nbmo+sk/5QmGUrAHcWUbgXq4ESfQns6rDStiaw5Pw5a4Py2Cc
NmCnW2MhlBig4UCZguVmDn6bdYvQWzKmYpKVT5AGyrsLkimG0MW/jdnyb88AD9sw
EGlyLmsb2oNXR2+BUma3ji5EX31SvNXJSzY/H8zKOFAEIAH1VbLBs3ZYcjt9QzHO
wFRsHAX5y5FVEaQthvfL9Q2zfCC6i7sWgY6miYh1gamjR5rXMgE8OESESqGqySFz
iShMUpYqiD53qemWZH8l2ctsSVj2xXZcqjjaYEBfB0quBTVpfqdx47gBhkUzC3rF
mGSGB4EVThArwKJ2lbLBlfIYPotGlKfidLyg9BvcLREtljgmgJeCDhm9vL/AzJe7
eKBJy9sXQlCicr+osOhp4uJCtG8H0oSNCbKg9jwis1T02QqVimPL/AuYYSGpkXfo
6EhzFWaTCUjST/UksNU+XRTv32zP+I8xE2TDPfJiTyyJbyVONMusu+J0k1aEvrOy
4phKV4LMweo0KBDlVIKGm2/Hj3TM2ajUSBCtprNRfvgo4aUOfW5fxJ7bhko39zA6
2mTRS0qW5ceLhbLtkt7Y4KqPRs5ccJbTUFTN3b3zlscH5aaf/md2kpzkkLOX+tlM
WzbFofWBEt9a3z9VxDRwLptbY+32OTp1XkM/CKHKZDXs7cAy8wKbMpHn+axYsf1L
rKIw97VfznIGcyLHj/dciw9KvVdHWFSlmcz1fRS7BCl+J0Vo8MA5yUhlD4TfDAGq
HVOpFgotoPVZ+GczeCQqPAZ2yqascH7aLEg6fxs/WUpREY6rA+kxuuOjxeWaM2nl
v2Qoxa2NZWobfLz2CldGdob4N05/kZ7Au0wYGeufMkFw9QX1AsbiWzCF2Z4Ix9Yb
KtEAbx8J9T0fSeP6SoJ7qx/OGu2UWNtnJZ1CJKrERRBAqrRMcWMhCLoII4tjT/Sj
vNuEWOO/66e1+ZQKcCJdYe9N+yw+QiKbqulAX5yQ5UXnmzy+orBSSYEKNYKPxMYV
LpPUb53UYN0WxOVxBGUZGPhShxG4n97aqRySqUeoLV21pSoqwUmKUNN3naIqx/Wv
NR7OI241MpXkiJ5nezD9nrpe1kyw2XuhboOGPJNmqLE1600SR/71YgxBlFn/AuMK
DJUIU2QeuOh676TQZcKXrewUIhXWIx4M7zViNKBQzX09OFSY8XWDd4JjqMXDmpGu
cd7BkGtyoMt8RQ8x8IeYqKB/qtgfQl7C27B2eh1pvR2nRm85rywcOVAr1b9QFXhv
uv01b0I9Pgpviot0nfuI4EC9xPME+hCLDlNjzIKmv3/eCsOMXRroZj0X/OpWKFGg
7BYjSbnhBN98RxP4rsGYO5pEz09kHBKyHhZG+dcYqUUgla/bHuu3hEidytyv3Yuy
KCDcN76LoEhqtF+hDZNPJHHdkU3Hj+NKvGs38rESi3QsPFDKeF1e0+eNT/eDOvY2
ZcP1GoIK5P7UjgxWTUB9IsHg66OMtSmuJXUxla/007UTgDjxq3vIHYYg/ogpvLZy
rpOpt+67wO++VpYJ5tU8e+ml+etru6Q0E2TNNEzryo+tvppGmS4TTssKF5w4b6aN
wthhdjhEZidpzLUx9gOKE2duuO+pJmxOU8Xq764I3x6h55o3vFOfy5axrNPKzmG/
RBPlspCcAXqbc6wZxhjHnIpdVHzrPDU0adzzdWJYeYYKx7QmDVfh1BtYpFoshWqo
aHRW+GlN3iisS/F+QWn3STBl7Oc0cQhm/zFqJzYGSt3ccO6NI0AlQcTsqQf6mnM1
lu8HstRxTcK75ls49ZqTexPD0C1UHa0q4NQlGyHKUXTqjQdsZUkXv9pVJHAbPgvP
6+JDdK34+0n0Ie4liiCSVGcPqMbJGeIT0ipbp7jky1lpjcPxMdv/WzIVT7EPJfjk
a3oyUJ7+Uhj1d8PU0VNfcB4SYPBojFbpzzohDMPgTT1XNnbkPWtNNsHnZMYYeKo5
PFIL2ZZf6WH40pvZA7A7bUDRy6LS13+hVXpKGUBCnc6lWR1Q5ryCvEVtwuV219lz
4IbC458Q6e2tu0RnC5Rzt2gCJDvOYB84wmF1uDUtgTMSI+OY1qIYlMvpiLO41DdH
pJdDdoetGck8efsC2E9Gox/kJ8zJpdif7iglsqH0CwtbQjeb4rsglBagvHsF2Hoj
34gcRSG56rhu5MtTr8OwSihhEWMxOnTzzQ+cGORGk+yq9E8GmPqCZc9hsqIf3AE2
OUEe2tmAD9OXNutHbvtZk03wmEmLTHAldPZrUpTXPSR6BYNP4bqEQM9usXY1qfOy
thXVdhb7UGj35YHaUdLfgodjsFVVNM3ZykC+YoxPoa8rsBhKpNgGJIJhLuWlm8h7
Wap9Ry6wfp9WR/E+GTWybAKYriaY9tl0YY774g8IPkNlE7kfqcZ/FAcjLgDiTVCn
CukqxNeDjdZOn4xwXyK9xRLgPFPGxAmQb2nnbjRLklW6/kB91rmX7v2s3+/fyFLQ
hLFbcE28UEMaTXjJHWEg1l/xeq+7eQ6RMLX1TKJ5a7nKxNDoTx8FoCO42GUQXMbs
0eipjZWwjn6Avr2s9hGYGL1tcG/KHwZwntG8JbgV6Q4PvsR0YLHT5xNFWPbhJMMj
fjjeq2iC1SdxUKcaypQFERM50251L2c23p8Llyj5GXUpvyFR+OaOi3LOkS4iiYDy
D8Ry3Z8HfmP8Y1XylSL6obFxl23D+vioD/yYL9rO61YOtWZRUNgEnvPdjWFWaSzD
xowLeywWNFd7OX71d3ocQvtVDjdB2DrNWTtlyDTNM7fej7y0yFpqysoDDjp4Qt4E
PCtRh5ZraECMF44XLiyqR8RCyqR0W86M0rqxvFSWbpJsYqnkKXidTOjczZAbzjeh
cRx/I35QLVp/0W1k1XItuC7xvH1lDJQZrTNmiNoz8mnPyk0pe64NhYpicBlCsXu8
SkvKgf6MTSjjbwR5B6HJJsuy3UHlTMXE/qBaa9z85rbnklTYH7VrpO459de1ydse
ejUDTVV8n9Q8QtxiK8z/qTINpPLo02YXF/NUj4lFrgZCaqYtxJvr912Y5uZA90X3
OBtYXw40WqLZEyvzDdBl6gAzRXAEFM/A3Dh26C669Ly+xJQxmHcDQPn4XTn2DcM6
0PPjQrB9dFfVTWF5RJ3PH0jvXX2w3l1EnN+Zrc7kxMtF0Hdh82rx09l8kWhrgoNK
jYtLZp+mlPgUea4dyoRBZpPyEcDYZAWyW4fP6sBF4a+IKEZ8v1PvDhDN5g3JXUOP
hcnJQn5r4q0HVCsoTCdaWFKupxBdMQej5THI78vNyI/gz0xjXrLZUNmy+5ompBwh
ZzbB9Z8/v7xeDf/eqDSU1eYn/Q97Y0JCYgUsElaYqu/GtUl8JG/6BHeRNSiTDVxo
ofo6MaxwlLNozvov0zZLyoMlissLrIyAYx/UIyMIfdSClRiY5ooC8x5ehWTL8lIL
KMfn/7ijfMsfTncRd9NKwg==
`protect END_PROTECTED
