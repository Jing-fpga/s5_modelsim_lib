`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HWggEkcYTBt6+gOzhlxDhmG5eT7gkeiW+rMVVQDQN9NdBpRoa59thgWAnAe10pwA
ap87eUeBTP3uerWPV/Uw+x45GrHyzKYwaq1KAk2z3p04bEDMwTLbku/WV4dGC/u/
8SmOywZjIaccf7Zhtkd3IptdpMTvGt169wJ8Q+2rv8BkWG+auJcqzm8zPRjq/nVk
BvefYR6TJfY8W8mw0+zZ6OWgYwqfoDp0Nlhz9upQpswmfkPceJpLoiuLsKqhoskG
q1Ms0Lva+4ISp90zojdSY4oyUpIvCs1p1QG80NWv6gSMOTGBMgm/LfiutZ20pSw3
6+0dViP/uFsABsKsh0OpMFxiCqrHfTJHonxv39tKxxItvBzsodqHIv7DQMAi/AIi
xERZlzUF1kQqq4fxLRa88RupQCe9v63k6KS7+dn6bwHu8LktnBIl/DDYcdvcE9sI
XQsUDcxV6a+LSu00zMKjSeRH9XOkIGC+Zp4fquYzR6sJALN4IwoscMaY+x3daXJ2
Z13cZTHuCRTqvcriq27odFdRN2fKTU2jaBP+sHUjOaY2do5GZRJkDBKhJhBCpE8g
vYJHZOmA30Xfe3EyO0Y53TSidJIBIso53mum/CkdhwRcnTX4AzUP0X8ijFYubrTx
GOGShiihrsn/R+CxFAE9rnVjYrITOJ3MyBopMRo5K9QUZG+jndPFuXOsIbca1QFF
c8jQ6bUMW8nHtcNiDtwmE9Q0yPWu/gLCGOnonEv/6WtIQ+zfR4wZ/2vJeZ43BvB2
dOoP0MDWDl0qg5/B3V+lyQ0WmKXn6/3WCgZydNBqEyb8xBHRNbmpOq80Dy43TOFc
2aQ2Xm5uQEG5wfX7zQM+RdGgg7g71xLZYucEZ2X3H0kvfR8i1Hs4g22RVUIz3kSE
nT83zVDbfm+MBWlKRWo7FLsNQeWBoO3coQ//hYYH9tA5gxpaNilL0K/YJyDZf+Tn
fxG4BIHA+HeTbI7Nietpt+U47PKiKtqnEGpxyc6M1EzpqjHx2lS1vpTmj2FsFF0I
xYq5rrlCgNvmC8PsVjLEnYf1AfnuK8WAUdfRcAEjwP+ZGMGxO0DgcshlmBHnzLdn
naBvt+Wz9t751KFV7rc6TBRvYc2C9a0gnueqQA8zDOO+7Wo2TgbkM84ai5/PQpLA
sK+zSAJ07JDg51VGp9GGocFTiGPd0xGszNZlivHP2QI5OeGNagtP6i9AYlx6hHqd
7SP9zd7GfDjq7pNAbQY5QX7lwsExybcYlV2KZjnT2+GgHc1RN2gAavcS3yhTiiVO
GWJSb+UWCStP4PyhQIZkozEHe19XrW5jRFvcduKfz9JPtswKWJzNP1/LDG0Uaozb
qWFc1s4UmRLnxNZalzzq33H/L0q+FHK6Kxg4QztSsaU4iXeHvhahIktuKf6wTxff
uSGXH6iSViIpiR5lM5tqNNwyhrAv1Gtrj44iwXA3+WMZHn5OftjcOBOuvHadDWnv
J0hiC1R8nblVsDAXkuzJZ1wXBhG315fPClTYZDo7UANGcAtiq3HRKGm/2dgbdJ3z
eG4V4DqE0pedkM2xMFT9YaQQdAepASPupJijZqYZ56/2Y8Rm+tz4VRy2F/ppILt/
I1seuzonI2PblePMgK7qno0MgycCUXB4o2zTgXihxGJ6rVQOmXCF97mRHGF3EMcL
cZzdLEJZqfDzB/2YrBFHz0Jk2ivHOJDh43XShaOFwdm9LUAp7DXNvesiqAkUIhEG
nd+Ycio4cpZ4Ye8AAad8kOWIqUk/WoNOyLPMCJo8sU0OmS9Jo8NYTW8nlSdIR3Aw
J/ZamFWq/2YfUa8l3XUixdxwMJhSMKB/CQz4PtlJluStPXKBqR6vosofN0NYxsgO
jyirJLybWkLtV0Sqqd6TYFJBr/R0npPxe3TCPgam1xx9XcFwPyT3B7G7e465qwF5
q8VPdXMXLIRUfNsCwM0z2kkMV8qGKgqhfPHVsGehTzJXh8A6kNoUiUkFTrzCwugU
G0bPA6NmylfTB0SVnSCQcImi1jn4mXQAf6HgIFdTwKUmYIh7SCFGwLdv8vTe6m40
61iUv3gGYrWaXpEhpz6ZxjG5Fxmuw8Wr6ckcva2QzUti7b+ZapCs2PYG6Mx0oUzy
w4lS1UC+NPnLy2O1l9bYJvYIuCW+j9f70yx500tDPt0oSB/x5feJ5PGtE0m7GYBz
zOOmfUMXlhgqyKy7A2ceG1bR8IktquTOuLQEz/VspIthldVkr8Oa+VqYLwnfnrZe
dudWv1gMQzWOb2wPK1fU79zF1lHzGlQHU9LmT3NVMBLsQtUnpNJBP3gtAEYA6tEX
leGR9BotG0FW9k+9rGyo6SGTC8Zoe4/ORbRX2JbWst6pjPVhtI4f4EnL7k95kqF1
axkEV8n1TWYzFh0zQV1ZxiIm2UgaHT5MRuMzMNf79iBC5/HC1BPy3SXayVrmieo0
sM412+NtAjmg9uVvV6r5lvaO7HgNaa6cSg953z70jxDyGRCnP9mQJuodwjDtmWg+
rrYCZh9n3FFDK1gKbjmCFh2vCXz7WpusSMCSbGOqIXvz/b/CLWGR93ekIsrT9uKB
1ju++0AU4qlqp/VKuxXU9/hg3cmq/7fS0AEf1ywyzDtLujgRQFuVX1Rz5jApUuGW
Y7i2uFK01WvSuFj69pPlzwD85gGQqOYna/mSJtLiH7EYfrHA6SRl866FJ36XfCzO
5bfIkVgIjmToccHF8j4nSG7mh//F5Sq9hkD/8gLPFtx/G4GBT5WOYGZs6XewtyVj
AiIs8wkjGKnAz3MDY9nKcn7U9ycDmUK4CW1QrxgUdZ6h0SOAo+nRKv9vI3/X+9mY
scaHjgkzpzP0V0Otxy69M0DHcLw97qxhVWkDRuB9nVZQ1V5d9llCd0OY4KQJA4m1
PY8ArK6mnxent78GZwWf3hbn17B1s4kjSWX2Ja2SJo9F1KXhu/7ecgWf/MRs3hGx
gj431IWnFl2244Z8oRlsWS26CfCHah7MfwZbtq7LJTf34MAyo3C4w5jh1eqIM1ai
hsXH9qVYCNIGlSGoOFlU59hxEKGbDu2haGfYqmdF7bX/m7zFzElcRzTyL0xHQoLp
ujHZgA6oHGFd9UhMT+TEre84KfNEJVF29lInGcPGozwckyCXUmbyEMuSWvX3Ryzv
OpYoFwluGM/iKAtM8ir973wggmz0TJx/geCJfGiekFVre7t6nRueVt1UPe7bOMoL
VfHfJ7SHMtEUH0G/do+FrmlE568yvc5Xb2i4fikfS96Nz7/V8AynmNKd/rQfL+Iq
/GXxzfpWvnDlzSYYA2RXpsxKMOtNerzjUPXwn88w+2QfMIj0gZ2uvHNS+bl1JL+E
eDJo/zI08fFEGvMloS0V9lUfNrozwFovc2aZi901QhAN+9FGD1havdMHG2JPMTyW
e6wV1nc4iE+sZx2PJ4ei7RG1h5rUI5Az6psX+pTdpUwQH0z80ahbUA84/1ojWF/0
KA1t2vbC/1BR9xPnDQhP0cQBdrTqnGqi7HTocQTLV8DjNsZag6y/EoFMM+yOGzg/
b+91btt19TUdCvY8u3l5aM7/gctWx3L4+XYqb6WsirSnYQQlUk0mVM5peP3nLU3Z
LtAWxI2DrVb+Pq0rrA/cDCyG7RIzuBW7xOh75Ut8MOysLDRT7Cc4JFFE7d7SAkgV
GqmY7YJmJAOnAE2GS8J2eW+UuxvzxJUkhV6S0vtw2dKPfh3VTZxqWNvaulJzIJ7N
Bv0nANV2qomfWOt9EYPqWz4tkUpDEiqnOi9HWJbXT8vqiH9WkmPNR1QcNjyPbKH8
bihJWaQGLYL+s3qyQRjB7jHRepJHXuhmWROR0tAekeCqoHfa4B5Eeui8SoLN5Q+c
xYMskh4/etJ30Ags6r2O74PnBt1g+b56ptljEdsK3x/K7V67bqOFstWrdch3TYnw
ikssV/tHAGSm8zn8ilV6dnLw3DU4kiLWTzcLzPphq1LrXhFvAKhvx8WDsmoWDiWJ
Z1b/APjUDq+YZ2NFR5Q2G5gnY7+dZayR3iRdJlMOxCs/yJFtrRDRQn/hS4cBPIfP
jXO4G9dDdKJ46LhTACc+wnWzI+Nk3L96MPvq+uUhu7NP8ZOSZTJ0zWjmuJXHnIXs
0QlzvdXx75/pco0vt/bzncvXwfn76x8hEarvCS8Ou4MdxX7pc4jVsaEFdA+x+vA6
UhUrjgpO2gJWB9W3HP3QJTqCM8+NO5JpbuwtoaMwGQ6xjhAeMepaj7j33luEdKg2
49QI2G4gU3PuMZyRVVCI8VT/obgNQvladYE9EjzG67352aywpJcdRYqy3n3V/Gk5
y9q+8LH2dAWq+rQRbQxLeGAFN/gNwwfrtFgVKzp3AIwZSSXA1YSmN9t8wenLjKeI
sh9iVi8GrwTLyqH56veYu3UXKhexhNct2/ZEGQdVq0VXjgprFkkem0jPwRiqWA8Q
IHYF04ECQfMqzUlO5GLWyvKB1fmbIbJQf5728aYOfxhUEZox5NJwbR/ihCbi+Xal
2wUMoVXdaJbh03YdAi405ybHZizHpYpTDccaKO/7Bz14DTQUh78FQ2b/NNubCsc0
25zHEmdziqoMWb8PkqEP+9tXig1LLTLydKh9lxvEswlxzUTq013F4mkW29iq48dq
4S81FDIL7Fp+GyJPN9U+Zrs426MUjVy0fLt4bgLKNAf7saYztTabDjIAuVo2OyUe
rNXNENvmm3lB7FBP5QTZ2aJ/88mFXvKY7JNe0kSvYzAxTbK7GTmAwCuwTX+5KM1v
NeyhrWKIt8xWm9VeTQBgPmIQiUwx3mZWj+rZJJ99e+kz41O9W865B4aiM6dMFjLm
FPM+AQ3BvjJhETQjtr+VlVxiqCbCUdWrJn4V4PAOVi0VYbUEGHMTWOTdKkll+K+p
AqP4G1cJ4Fxy0EmVy3wTaEOCTTeNiFjkZJzmUXWDiPgj7hAKkvSMZ1BHDGRiZbYm
DhluRZuxBf4hvuKkI4tQ1oZi5WvrqTH7FftXch2eI4kge/aPZ5G65Wi4CxSwDE/h
Vd4tFNzEtaFb4VjI2XbYSZMcXEHYBGLw/A50b1xMEljmxIk25wGGPy82/Frxh4m3
EVmdMJkjgANzL7EQCbxxMEoVmhpSSCuANHYlTPPH3r86akTyFekqhKM4lNXjEmw0
YKX8CaDwrUjW0bgwV05c6+qoitRfy0gFouKLpATzdADAZ0bV1NKUXciostpChkRH
kk2aM2I9u5PeIvtX92+eQjmQQYtyhGeytiDyeakZdKzXRW5+u/Ch9NwXy1kstQwj
SbtXgYbNNYgeClTcUZZevF7NBFGd47GUuKqfShV/PRDWJdHOSv/iWvV/xRdsu71I
hUZopd1LuHAa0+F8RMp5mAaqBzbD2cjpagmnHtDf5YsG9f/w//mFbn3KwOTdkKGE
roBokzCGi4nhJVUvBZDOHxsyr2vmwo9HVqIMyXaD5cQCrIJxDa8+GF1v3D/vbjlh
FGu8L4JvS4WchrTzAxiV7GN+fN+/Gf94J5iXZ+p3/MCS35L+zSFbx4ipOH0u9bT/
oQY1ap3fj/JjBNqOutRU/8uFWUk7CC2EtQdUESuHvjHYqpJwA4ZtorjShj+w4t88
b52++RrSz7AX+Bz/rdrr4qNHdnD08hlzD9Iq/70kO1hfAGeU9KuGUiO6arU5UrSD
CyFczjQQ4w2SIPD6S3+NFZVFwfIRzHFnH8HNbVamf6r7cD07Eq+aYtc6bSrloL/h
y2L2DERpyEE4c0s9ebzgTBtu6JF+rO8ySSrLTa+uJBg2v6UUTKSYA4zT/X7Ddqbs
4RH/LOiS5u511qd5kwmY4ZBNvC0Zvggjqj3JFtglsFetf8Fgr1hNL5RigQzIrR2h
Bv3vd+VS7CsfuH+uvsgSofjVc6RAHBZ0kVk6NBH2Wyvto2/Ijh6OlLZGsk6qqu74
E7GYw5IDu0zuk9+dTpQYdU7IeafKNj1jsIHolluFkeq1lAb+u8mg5q1To2RbegcH
6aZEtmcOg8BIXrxcB/oqFFb56RIBbzHeHmZs+31wZXX2tgT5gyXHyzMFcuYxAkJi
Rq7uc7STH9VcTgKIfOWFsvIeqaTxAGE1ktTM+PjYtSFJPtvZZQOJbRu134dt6ehm
PcaFJA0cH+iuZLpUizo9UuyC+dfbeF/rkPmTvQA/rOOSXzBjNE4jKT0/BONIf4R5
jaND6Bae6iSWs0fqCLlkDjk4w0p8LDOkGv1Xb8Ynsk9/KLCt6W3w1jyEMySBXApJ
Q42A6YtQm0Rr58X9FohMNWbN3gl0MaFu5KinYCvnSuU63+8CbHSLk31Gkb+JnepW
orPSTKlChrb3oJG1eYyqR9cygsLBS4bZRchI3D7MP8R8xoRNDevSnf4NZqvkJGoS
1fDDZcXgEHbOS7kUHzNtvaT90LgaML9rhEKFqZolpPXW5s41f6symrBILYz9StNH
Tl6j8BG0A07DkcsnFCs+srr0Gk/jS9Udta3ig4EN1OIQRQql3pOLzjJ0qLd9l36O
JyJkPj3l7gAGvCYaz18HP76GEqE6INKlYoLQK2rpqPXhxNDnO7GDvdwqcLBCi7G7
b6R1X5s4EDOwgNJtBUuAykumiPOLysEDej99ZauV86PeOvjQtSJXxMZSDoMCZVHK
T8SMEbL1Pdy9FPM9pogX8wft2zKm4cTvrI3NZn8BixQYW0+V8S5jDe1B96y9Avia
98g0I8jZiVLMqr4w1xwFHh0dvNSZtwJwNfX7WQ3e9NXaxriv82CdOYIs3Jupatd6
OTuYAeDiUGDxeXpxEOITyJea1OEZX3DzWWjkfQNe/JRRUlGcU6vHBM3qkq1N9r/c
3CUZtvecUvq4DJLCL9tlRrliTnCqqATR7g9I1V+P0yNQ564oQgEOz8g3J5GehO+3
Y4zX8zWFBPE5zJCBS4CPNiTMsQs7HGFzx5xSDAjddYtD5DEnJ8q2PF534il75dGV
FpzMQ+nBU64HUhFr4qz2g90yvTsallLsQ9okCA9+QKNCv3jP1N71vMQ05uvpZ1c/
svneLCC41S36+oqcqlt+RjQCDpPQQmJBXjmJK3F3ztIlwNKD69xHtw7SGOJflOqV
lJtuBZX4a0HYmfkfScaeAJbz24y2LHGobMz6OxhA4n9mfTIYzAPeilxeaagwg4Yd
94H2BSlOnjLU36VwTAB3YFzgjGhrW1Pe6ADf6f9xPxu2UfLBypUUPXccw1vpoJqr
v32dTy2MeQjBjRWazkgS7pmlsQwJraXXwgByAtsWB543t5GWhNGejMfaDCecIxVB
WGCjNDjJIYFfy1smUTydI3S+TM4AyGZmeB0VVwBJ6q0wn3OLOngN0t6KhtUGpEp2
gQbl9YCngFZvLF1VH3pyGWyYiR5xHbVZTEOF7wlfOhfzOb33H5aIaVNd8UMiuTBD
HxrzCEkyXzNQBGZ4O4lf/umRen4DT3hDKAkldblJUR9sPvadSK6KRjA/Ev/t5sQr
tnazPQTHAhZAXTm5WgR/jPy9ZvmcGB4srAtNdZ2B45R3t84MafWM1bJ7duU5KogX
U5LDRUzsqcojzW3p9kcE5M6UY5o9UQ9Klo4HlQYSXmAhKy/oK/Jky/GhEHYbDQqu
QpCDqhd+J7pZwOiHT7iLz5oPEd9mQ5t4jBrjkMfR+J6XqmHyoMMtVxHAQ71Kg1Bw
OdshJzuTW5BFvhMWNBu+NhT26KycfGzVH2UcSuCXlvyA5pI2fjQU3Vm9q0e6YBt3
F0OOQhtLxHuo1WuMO5gl7EiHWpYMGv84Ohrm0c+Hx4gINA5dxZA4zs2wWBYP4ozq
DAOALFjtTbX4FoTi8ofDIFVW/qDLckGWidyBff7oKdg+//MA+ZZc7zprM8N3U2JA
aQuwQ8v9i/htClZJ5KrDgpkKJcYAsUFvMCF8H5B++DtP3HOg9wKxffpyLFgP1gbN
WDrwzmoiJM0+H5SE/rn6yP2iEK+UhA5NyWbMfjHGcXsTDIk8FCaekULkQYVr8IO5
KIAyVVeoDyGl6nx1JAQwbZNyB0LZWNVPZqybKk6NEN0ziyeZa5jmXTAUBiVQhax0
BpJDTxUQoXFN0qMqptgoyXSnYsDZW1OdERrE0GR4GVrBYXF8IG9tm9r4zzWRgS54
Ug0jfM74CMC+u41n277kJBEjrWjqhxNXK/psQMb/SpbZX/AVUoCv79pJrWBKsp6h
A7hVDQXtHgmPg/LiDDZEJDkZi9fTz5M/UZwfBBkR0duv2zcQHNFiL+d9UCgZY+x9
m8WaTxnpoTOl5x9CmgdeZdatmPW/FPU2qNrP0go3ze2tFGoUs3+jZWwUgH/1JZt4
rC6rrNuvDA7e1HxIgsREq1v3oHKXUnjlfpJA+B7ItVlmpTqGpL66VX5AGp1R+ZLL
U3u9RPFH/PSo/A3gqssWQR/WKyYO8L8Yu0KGaXQtI7Z0fyo2PsukM2+pIlua58C+
4wkbZ5dDMV9Br+hPN9wke3ffcSvSzEQFaondTLZ2tmYHKLp/BxbAXN58Nvkxk6AF
2HFdpN/A7ZKOrOxoAX9oH3zvQYA34nrPEKHqSCvWZ9m7SHQm3EgtnIidHxKfDlPT
HqTU2feJEWmghrA2lOgOcFKIRZOqxb8l4DOYoLhn4t0h8UTK6apuB27mJ5SlEFNO
tXNU4JUgXjJG4YyYvAPQuMhjnBG1EinOMKlNna2XEXhi2pEmUKnnDrwCYbOY/cZD
PJbqM8hRS2n3aqnbd3SSZbBfS4S0b508xEXeLQGNKsK+h+Ax7zD/aN0qpUjnpfdZ
Ql5zBCCKpb1u3nUM2vfGWB32JfWJ/7+tzExCPtZWzoB73o7/GWhTKUSvVuJmM1aE
sDBMrHoRfw08bcRnuN5rDOuLu6kRTIvhtu9Dpy88pBtns18wL581o1XrsKyHvs3m
i0j19OjDcPV4ri1OFdrKTMSgBpO/fZDRj/K6DqmSYVlKz5MGy1okpHi+bjy+MLaY
obz63Bg3RY4Oty0hZJf350RpDV0dJAmo5gjqHyRA1jKga39E/fYqm14nOt2DlJaW
b+IORuv/XDkUSd41qBqik0R78GpIHRLp3BPbmtQhOcXSwEZvpAW9J0w1QVvdJgz/
C6ncJ8xinBfvhuQAesoDJ8Mtak/5/AI1pQNq47THHUSjQWa6nJvVD5iDzNPr5ZIM
QVJSpZ7uyW8R8TvzqRXbzzLF1eWgNGK8ZUvG6MSo85+G0JX8rF/xyyQWjaEVAydK
im9mK4ey5QZjsqH78BnTagSjmB7K/rjiuyAks85HjD19D5M3tA+FfIx3rgeutC18
Dpm9KPs6cr7OvyQzHYtV0khMC3zpV4fSafCIpVfP9diaIZnWEKPNqwNySFGreWX9
yNxOGqJV9FTedYGC/wBwu2mc4Ih7md6kWg29F8139CvGPhg+abFxIIwfXj+esV4c
R31Mtpud492iA5zDnfdHp1NpsXY8Zc1LfRRW5B+294SIdrif15GCJUZS+kNDfO6S
fQLpIyvhjJHH/QxQd6D7tdvlRUyPm6sUtlNeQvOqsQYpMd2zueky+1DvWlCV82Yx
VVsiBMLgupHf5CBwuhUTT97M/VMCq8Xjs8mvy0NAhZKY2ClCIIsBfgVIM12XhiXn
S1TAy78rtXWz6gajFgR2hXjGn89NRA9fIsOpwLFHzjMDbmip0TQdEVEvpjiKr8YG
wXe5ZtoFKeEsGNbyjWZ4b+FHimoSvgDbNJqcONTpBIcA6ffsPWSlYPOie0dIia7r
prRou4OWS3v92c/XEy5uhiozlbahdAl4wKSb8n/U62RP5m9Fpk40j7xWU5sH3qUy
2kOmip3fMu3+2oC08fwKTAJuFkaPEeAMS4vh2cKzPgJKYQ/5JlKwttKEAHdOfP+9
+S1FFLVmusZuQ45BwHL2x0tptnfiNs2kV5E5Jq68tKPFMv6fVrhNnkDltIIEWfpk
Wr9cbA2IWWR3RLBGlEv+c884xSx8FYSnT/Rn3hOSYL6jWHn0Cy5qJhrnex2+QhKe
dCGYO7zZ1fiXkdi0ohKi7rxI0c9/9J5aOe43APsDMdHbsKtYjA74s6aOI35gsUKz
7MzKOBIJMb9Gx+Vovmx4dTkmhS2mL+l+MwEmNTsSi4I8HxsQRGeEtARAM6wLf8up
JIa6LpR4A/cMEYCie7yqVFkJzsTsnAiQlLlbU44XLtLWpfpI7KwCmmj8ZFiIWcjh
EI7JU5wiV5Rl1SrRzhhrwfF6pWftKtl2pPBxyV4Ny9CMvTlw9nP2kFaOlcvxUWbb
4zRcxKjGBMO/us5Pw7tnzW2JjyJIckKNw22XxSqp5MWAnM//S/uFHJ77JmbQeZIY
RPcfBk4eTJESla6JbaKM7OhELKkwJmF13wBuqjqpPTzmB1QBuV5whNyWeEUnOvir
GvbTfvl9olIfGiSfZ1c54+PLS/CLIs7CubJei0dXjYNAwA5Vzw6/kkwwIaPDNzvx
LhG3vf/lhTRcQRlM9l9QSuu8D+IlzyP40eGIODJuf5tfWjEJaVqnuTqGjE1SMPz3
76JCx2k86nolMP8srcfAGOBaUgvmFUIPdnE+ZvLPk8X9X+wtri/ecTxQt4Tcg73b
B0o9Bj7jRFf6+C4PCy2OE4Q7iBGkQB6D7W5FoyQeW+MiuxzdLOFtcAJylkKH74Ip
IwDDt/CJevIFHunuISgraUnPTJUuiPKw0uvdpEz+eH2YK5LJsBpdO9XANXuig5Lr
AxuhkbxP4eUg+uTe/vrYLFtarxB8z3u1BAkrHdhsj9oOfas5I3l7tDE21N18s+/g
zqGMSvgd3r++pdNJ8Rc0JVZbKJPDawSvuG7OEh58IfpTnSj4eLeni9SNmVEFfa/9
NIbYY2CYLGJTbfmOiSU4lpymhsoG9zXmV/ceBGmX7r4Ik5lWz216pJnaONFlf33w
iJUtVE0YEXhLW0Y91jniZcHC9U2ostiFxYS9sLdcDdhXeE4VCJrEtqNCNUIHwy+H
SZVZOIJGG5Yj7f+yWCUB7BFOIlC2MyWLRbSyh9X49HnhaOjwrxDlTCIui4T3Em77
GLuqobm5Y8wvSxZTsPIFZwONAbKdfwG5YidWuCJ1ZigKVl8TOPSirFlf9+fC5Qp2
UYQ8PsgEpweOQNCqvfVBUj26aKN8rl4OEUB/hyNF5EThJPk1iQW7orGxIFD9puYx
Sf3aR6Qr1LouaAby6VWJ89AEeNLhXKdtx9mXegPJWYbzQpIH0ow0uOy/9kL+q3Te
jwV3TMMx2YopB4U3hQhIW+OAKyXpHnNGG1HFUziuEKyzzt39CqZjVtkIuPWjG0m6
K6z0eW3qwdHU5oemBVI1e48D3kwOconM6F66MyodVzizppLkbvqpZsyhx0pWxin7
baJE6M558S8CE7sBd10jCgXet0BxjkkKAN9YFqaR1q6c4u+EINb4F9FdTAcWYMD1
cByTmg0Xzp12wniFa8c0q9KWEeUE8ep0k4wMzcSfjMNabj7RNSr0O5k5SPyQ/TKt
47JEH06Pu0tGcj1Se2pynDFea9X/bV28drsMZblhbgItuIAc3Zh/bpLL6/PjJhxZ
okCtfFHsk7YVgbaYtJCMk42m8dT9OzpLaPkZ2D2Dyzyw0dkxs2xDxj3cA2J8O+tx
NfGB43knz3KoINQgVRPyzVznayTns8sErFkUSykLWerKgps6ibdDM/7JVa1xBbVQ
B/U4YKf7q6Y6uu5vpValPbqCKunGYRHBF1QS30zK+L6saspQ8mJiVSRjNUK63c+K
YNscZ/DD6fjISqe7pKr0X/Fc4RaWzYH80eaB8h8wqhX1dYc/OcJqzYjtqbFI7VmT
2+Ue/3tJCdbiKXvyWzOBiZ5nsbblbsr6REFzs6wywWX8QQwY5LOgxRVDD7LVdLV6
J76zk4qwF+FddVgUchnmaAQM2EfAM0tpTjhrc2wBX2rwl7yCHodibvGTFAGafXTV
SiSZmE9yjFdR1CjkmHPut8C3cdxs3FIabxZ9AtS6mB0+8/JFfQggBfGcMgTug5KT
/PUjdz3G2llSU0pyLwVH19Ag+tjxGxD/klK12vxhaDoXn7GADQIHx9kHkhrgNS2v
chhMTIDsZp/GtLnVPvVJnR0qi7LpgL9L66mbpJL7Tp4tQUdYCLtt8hUMlxVe7uzg
qfz+upNKsxLFmTIov1XNnH2Nq4uyBf8Z9mZK1b3yZIprYH8kzQ5RgsorQC0OytJk
hukQzuyupf4ufft3PQlDxteImBzQugArzLL2o9aA53F6wM1fPajoqPc72iQfKU2A
ceviyuxdsp7zanZFMUmdoon0Bq8ML+mhxrVsGDd3jY6x6TL7SBkvzjrrmIZYh5P6
BI8LQPnPaI8SJC1nB4rty8+zZI226scb/ooly/QYLbzX2ITHenkCX5UC1Ww6ALhB
B0Y3Ek2LSW56jREfxAh3y5a3RRHydfyrQi8tCGXs/8h/qPLDUm+dtECrShY1u+Cw
oXNTmY2BC0VDhZL8GT44WE6AoGBI6jjZtZKMPlV8LQtWgSxPjG9RwyjszvIEl4L/
ybK3k0hA2pEUNq060C6IMqUEp5HFVjXLj+ywS6OCaUokVjoJaebokeHwgrD5+hwl
nlBH/2XFzl+PA8mkkBLG+4Jt1mEqLKpUHw+kf3q3iIn6ZvM9ybU56F5zRfo4QKV6
63E28wYOw9S5OZukrSqpqaDPAFXaRqywx29Dh5EKK6JWGJjko4Skyc4+TWglmvg0
ImCJ7CpVbHLOb5z9U3S3GrEwtoikv/s2n7wi0d395nzUlaTFX8ti9CCYTsYvHmBY
9PRBSM1538reMMAWY82jKGacyP7wcOM3aCI/xGU15cp61IyKESFqv+gfx6JBG7OS
w8bn/a+iChfgjNnjZOqrtG5oNTcVxOUKp1QeT6bMS2ZkkcFl3/Ji/YtzeC7Kk3mB
pJqQPMnTpX0U3o9aRMY1lyoG9VeH88pHDIYC3BNBY5yOVaCkwLBTdRjsfS72CTZa
Qc95GLtCdfumCz3t/EJhl8GgCB0qMbHIlkp1suxL4N/qGmQOe7tLE3D8JaxiuZv/
jkS4e+StqZPMGzTv0BKbmdqwCBmKG9uwTPfErCSP2YRAvHi0tSQgEGxQfq/LNTSN
/ef3oOiv0z1mppuI28HV3mj8Zz4RZiLHY8pdGsC3HJF1r8weVRZAru04p7LjCFKF
WySqIPfoMFAYACny+GZn5rmmRSI9Mz0IE62qwv9iafoa9w6qbCZwEL+rB2XF4AUJ
blwpkcpvzfcRSbvSH5tIQw+EobAmjJPitoi553ZkdBgKoAbCDlf3tGpwtWPbvejZ
7eUjojA2MRGrzHeL0UHtVmWxWh7Knduye2yt0u6QqgPqGvYeRwlu0SoZ5err43e/
x4xjfKA5I3dX7kYf52Ep664JPbsw+Q4JXXlyGbxCvgbWErk3AsjcuGOok6oGuUhM
jKGgzQeBCJQvTijFdT+Cvigw5JWNtx6yjjf+LnPsKSFp7VaFp5x2zqEbxgzAFMhc
mcvCGcHVFGhqWnXXUZglS1JthSLMKrQpIMcpdb+EvtvY5I7QZ5OuPma0beZV/SIf
G436IjaXMWl/oATzt8fG+ZrOhW+bTFSVTO5I0px+tJKOZsK28B1hDdoz+qE7rHOK
XZPIrtdFw5Ph8ccAmP7eUjsfmFVQ4Ae1cRApxGLqYnQiw6vwygXz7bTJ1JWGFT7k
IOsVs2z9oUJUOFOcu45uVjHGfnTO2+qTD3vAM+mWvGYTfkapGqdFV4wDt6v/gPhV
u8luh5CBKVyroRbynxoW6CYuCGTpBVDhbPoWNj0bfVBlLpJl9bA+tTFHR+v0FnSi
QppoGT1Mcrj4PWBEjOLYXI+PRHNqi5Tbm6bb0601KLXF6m/3tLhC1fHAR8ypE9Cz
RJOKrJcx6P79YTI01yWeaqzYSE69VCKfrvHR2PS+UIX9pp0ek9LnRomRE9YwqA4D
n3HaL5WA07TmJNGZ3ruodaSPqzm6jrhUXTyrP6NZEkDERv+xLIeWNXOta9eBequw
jLa1iMR4VCQasiF8MhwcVdXdsCJ4w8DRN1ho1JsSC0xrm2SN5GjD4Llhb90RVpiA
wmVMLHhvAgF2shjz/b85KHpfYh/gDLoE7sCN3WV9MeNP8ao21X6J1r+ZrHe/+FLz
R8oCme3QYozU0vdoc6zIysK2KQoclqpugf6YCzMuAiOnSmYZVMFS6TIHdmT8Qd7s
aH1JpLStez3yCV4PEVo2HdkjEO5P1B464g3x5V7nQztpTA9GlcJXN5aFu0Jaoyn4
QuTkAlvYenYHxZz+m2eke6Bgr+QN9d6SQD9lZtTURbprSdIWm1UNwsO57sAe/qCh
yHy6X6GeXQRFrWcWpjl0ya2Fh6e92UgEqPdjE2DKQeuTgCDZwrv5gWOIaPzI/Zgk
DcBB3bwTUgT+fpCa2uQd9lMYfWeB7/+YnnLVOLEOpj4Voa5wXqGU0pu2jjNAdmM8
iFB7yJ3zU0LagAlhEB9/gxtJEsfgq00RN3AlT1U2BTkOy5C8k64VojptJhctgQON
kMuNEzZDwOwpuSR65NgOqZMEI3QpoW3N4c217PLVoTnuQRAbvU6kKwHURfkpIOaR
IBaWNpE9fucq4bv9PaJHTRTrkPXiRdzj0/bEUNVTnRctpSIEtuKeodSkzbUdsY+1
UhmdgMNDuwoHRqEF3YAnxi6Ffhz4FlVtHXDCM6rY1XaYGAhvcnu/rU31KTfSX8dz
tVuO+FUd6c5t0IYkca8hIh89m+YOWHKMvCOSRp6dFQ6DdPttGbkyNb3z5GlWupiB
q/95AJPNAG3wYsWOoww7b7ByzT4uic5mqto9xsoT92EZYmbdZAAId2eOvFISOutE
LiIhhltT2p8/N/7IownGGSmNkmDzlNvqClap1aAXVmixQ8+7mDv2PFB8VSDvNGD+
dm5BgUDLWVtzRNcIA7azvaMshBkwPg58UD49a0F3P829Wq4SYFQWDfE41NHse1Mp
8u9yZ7mQBIoQyO1np8VDIGV5ksg7DAaVgMSiRhJFfwfR7ZNc+X4jJ+TYYiuYLqgD
0RPs+nT3ZT6QzbNy4a5y0rcM19VH3FFrR2hqw89ACybL1BsKPXv0mi/aqLA7Dyew
rR8Dey+0pZZ2MIIkCTl5P21nbmLbB4vHMpnHLov/QmycC8718nBj9WZcm1Jl7At9
72rNNxEDgEiCfu/krU37Pmcg7mGk76MIo4Rf4Ql69N1CQDnSn7qHWU2pQcXvqmOT
CxzZP3nSmSKEEGSn62tvX3Yc+KjWPH/hEIk2nPuAA+8KI54oCblVr63jzrXe9R1h
xNnBPJ2sqHrIKXEnVm9hghPSHeyhHiv7Q16JK7lytq8oZ/RYmIUX8I3l4uO3ByD+
FzYOFgranD/+5CifJxmx7Uda6/cyWb4L9X5MA3ngiGCVOuqel92bQ2RKrcsMoRdG
vTnFzg6eanMJ7C3mpmturydnb8macOb47vQelF5CMSqHvVld5pXDbrq6tJY2yard
juT4ceRwy1/BTvkaA7qiMtxCr9PO0LM6iyZhbRvR1nuUeXC42K93IKA1aE6/nUIx
SrK0zkD6sxHsViPn2pib7KKjABltmSE/trAT3iBeDyfRwhvKWVtsItBOnNE8GuIl
5GnusisB5mdJxZ80VwRgITQuykrm0fc1xpgOgMN7aYMvcIuhguQMIZRLB+hxb6J5
4M7/yVrzPhFO9cUvQx7m1vHQij0tggH4jjc514sP6TY1aBnfMCNb67UqO69g/MC0
ulb8jp/blUvJZatDLJZKg3QrZE653TvrRCMxuV2u8xjRdl7G0VNploWTTinRKQCc
+Sn81BksHoPZIu0d02Re2tCGjwc7Z6IISwn6md0HHGo=
`protect END_PROTECTED
