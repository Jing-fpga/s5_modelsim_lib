`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GeW+3dNk2W5x0D6f8Aejb+UMf9aE+CbC4f/n212Z4r0eCqJxQhY7y150nDqHx7SC
Sa6q44LWwULNjwNqxEEGS6SlZD8prnKkdBeIMuUQAFcIo7uOCS4Hd0rI2aBwsgsl
OirwS0SFAStFZGBuQO/qmK/U8HpVcXvEQpRuhsM8orRq/MaNh4AkMvq29bYUeFmY
01nlkyXsQP2OdpgbBzmu8CiGeIPUcyOCYEe67Dmg5Ash5xhIEGo0d7U9d0+8Ybns
P5krluiuUPZGpycolMHpiZaoJzOB9KnztPVF9f6OFqgUCHhLtHRISPOwg9s+EjJB
1iGGJOeeHDWtK7jUGpBh12q4VDaOkqPHZPG7P+W6lxuPH7psr5iO22YjghFg0DMM
jzWBQYdEMZ5lF5JyJgUprAJDmu2A7FVFvBQ9Jj1DBTydy7XciW2tLzjgIizHQGus
lIbqhVZ5EBBmTHx/40jYeI8RwkUEkopJP+eqaiCRPRwVBzk41sRiUdbWToEJGqDj
7bz69T2jxIeWVfKXBlZ02o5WlennARkO/B+kwiEDh3cDbiwzOsJlzdx7fRMLMB34
Qte8DDCBXT9xmdWwc7to7wN3sy15yU1yo/kquUS7fejD2HPdvBWEwhgWaEqvysht
jpY//JwmGNvAqfO0Zrent+VOLTWDVnFWDl/o+IRc/Ai3XhxzmAyPAh6nalKY1kHD
9gYTaeB1TTgzOHWMKJ0u8JOQc2500Tr6Y/2FWi6ecyOBG+6eq8cQxpVZU9/WDvfP
G9n0++KIS3O3iLk7IQnzPLYgTZCqWgSmHWbwbAJ3rWRxcCQHcX/FRtZYyt7rhyRh
6R996CL4g1MSsKX6BfH7kgFZHV3iq5DyxVZQ3pk/pSx5yqhkkk1jvdwPNn3BesWj
pwJIGE/okZvxqRLqWnctQ4FaB38OF/b7i07LSZUbJiN201YDgk6Ww9OnyPIV4AGu
UpR50xr2bTPnSqdZtYVP4+WSRnSDBr5Kno2gQq5axweh+rRufsPxr8z//j5+iuas
8xP3O37jDGiA5bIdbWis0dSaJhAYd2Db3+uB8ak2aEp0ohKLum8buPKMHa8l4Gys
OFgkkJUN0nJ+Ab+F+tpOeQwv2Z/e0SZzrDn0bvkc7dU3sli160/B9aRrprYGWxUv
nLTk20NFb/g4kWxPs+Tgcgui5EO5es7jmRhOqsLCyuNX8NAFDCJuugjiRhbxOA9/
GyAwSmFhRksepJwIS4Gf5CzbOKh4JTBv48qaa5fJJ0HokEaweAbZGhoWQfa8jvXd
iked2jKPi1G6+NPRTUCNi4qnfhPUXKX1JZEb2ABjJM6JJlnr/Tl05b4k/AWL4d4k
dn9U15iokNJ97cr9lzAqSZA0UbX94eYoLcCvrOCBsHRDDk+FOt2rKnF7w+biD7GO
epHQbOaZlGLsNXAtUe/6pdRSE0lUTVyTUftZZ3C+lbaWza92i6rzpXUyKaw9+S80
nBYDcgRJ5ilfhhZH32o6DSEOJy6GVa4oAsueYlI2QUQ=
`protect END_PROTECTED
