`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JSFzhQ5tFdhXqCoIl45bu1iMdq3mVfhHu0xFqDtDYQAt5Z9rTOphmpKUi/yY1rNS
vVnT01VaL9XIKc6BnPoyT7zO8XaKfWFO+s85umEYd1Z8MpJ5FbkH9aBzqIVRHZiZ
wP95XmTuKK3+TWNO5Nz+io4J4BSEafVCLFEGz9/DzD6OySzwAIYIxaTeN6h6aHWe
1Gc3wcpd+D0UHlOLjpPxZYx06tD5yse+JajePU1gK9/j9xkN1FDZNikKMXJLt/PF
fur5aktLFMe6oQE6bLr10Jl50GdkCy8b/X5inny4SW8Hj4sBGIEyNEbdUQWnPTGk
BIZUicX+KG+w6g2ywMGALu9R/EbsDpjDlLhTuV0JxvfUXB29nsPr7mWjIOiZuteQ
H3F7qrYubfRWHxtZdJEg0j1WzrjJWHKivz3qwhW866rEEQycGY99EKQKLitPFMUq
2YM1N9jSZuHL1uk5IEM53ClygZYTLMH2swCXDveSDeRqwsyYgwxPOlC6as8026z9
uC92B7URHU+lDlZPa4PD2zozfwDd5ma/sqG/nFcFQYpP/Cq8ak6cOaagd8+wWwZk
/Ik8I/1gBojyrLcecDvncZ+I4UESGw8Kc8yE24H+dZNmO3FSKR7R5C5gnee/fxUI
anDgKcVkLCkdcNUjok7dCmMFizWQJX+lrZGDIgQ7gAlWTL9nTuZWbxhoIw6omebo
kzbQg8xZiJ9uZ9laDD66oke2SbiZsStiq+9VdmN1PwXPhCUFDHW948uS1G4zACyg
ejY637YBLXKSwjsqX14SwDwcBwc37zLfL6LYq1v4BarPmBrQiWASFIQ1f56jTdpo
8gORHmGq+jNovAh4zg32yi13bNzFLa1JXJH3JxOl+QRmdGB7uBFHfZRS4KVCRD+9
kNzHQq5z1IQNgDwB7lynv8pCe++PJSsMlUCy46L9olAa0IcDksslJQz5wkgV3Nfb
waZ0VmV8u/LWTEZOhAtJgOsL90Ql9TIp3+iYbdP2lfvxH1ppRqkcZnPejh/K34kj
WQW7lO/S05SWEocSiYr2w5DN2SyJn+iSN+11dGn8RZJkmkBcXfZdJY6oJnJ5znId
AKcr9Aw8xrenI/bR2v2m4BOocfj3L5VTlQng0TxygArlB73yEzgVXi8ysguqGW/B
qP/TRA/Nj6GrGtq2V5T8n6eMooIJ0HPPN0Az6LYt9YdstSYUQJS6Fe1pcxMULt3L
08wcz7Xbd5CrKAsKN+IS7LL6OoAJ9uESwJtfpY2Z6PQ3dRbw8EqIvoHyf0p68dui
dgLQSdhgOnEkkjkfGc98PLmcp0hMAERbd1W9LCo3jPA4ebUe2/HV5+6vN6HIzruE
iq4XkoA2gxBCbXyR65tsEsmPHpypqAsoudjY7sQaB5g/niKakbqFpxfKiLsgEB9B
E0nLIragkrLWeEzBmG8q/9AM6kIjGxtutoAD1LXM131wF71Iiq95aGomYzkX35Rl
236yuI1a6IlBlb+2+T8v9A==
`protect END_PROTECTED
