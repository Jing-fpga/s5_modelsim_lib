`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VDm0KccfPs7tk9gSuBIYW6+Zu63F5W1GrBMmJ/TU6oaS4NDvduq8W2FUj9l6E6Df
WE2bigjGizQMBnt/bsxMflR5GhPo+bWFI21n50j6DdHYL/f6Ybcw4yFgpRq2FICE
tYoqFBfg97dNjKpHq+B4aVTnnTUKx8ExE8r5AXQybFTiI+lj4/EJQ2F2Zp1wnYpb
XUk4kIpGf8sTwaBmkPfwHwTqr7YZ20J3qprhzGMnYXVeBNX1mw834yvG0p2x18ZX
q4Iy5nON1kM4oUlH0ulWV12p/kyLx7FZjU8XB5LJ/PQoypArOiZEXOt7WQtNhaSL
+2LhBVEkVxk+JSnWFmZ6oyUDRLxU/RNd1G1mmSp3o7STGOsn6/8Ru5pfXTJ1FFCs
PfGRWN9XlQG/UWYhLUi+KUBNuJzzvRy+2/iDj/ozSJv9bECFh9hIap9sFJ46afYy
8qhHxB7spOzJRy3CBK2v7w7zCDp6D6LLo3cuu0TtmyL+25Y6UOLZbdgcJEBGy0nH
TPVZnnKkPaTYrdtHIfOFDteXtr5m/DZLOuM6phMNfUF+4Z53Wlpt5stUxhUa6TOy
pgU0z47seNf0oGe3r/dCZ55WAEzqDJSI55tm+Mj7Dcu1CdwcmMLY7mESAlc7e5aH
WUej8jgvOzLt2WhJJdo5Wv5dhy99MWVdB+SrS3Lh40CRefDEKo0tdvvC9Lqu9SmK
B8EbtW4ZS7tqo+Vx1Yn0/TjmEJvEdYVp2vSOOCpj/WBrtimEeryGTDITfdVlElDx
n+lI1L2JdVUqW/osog3PJAs6r5w2mN8oqL8uxZ46zm8hZIaE5mxXP/p7oJlOLl0/
MYj4ZSkTAzGe002hjbsXSSofqtLXDVIl7iJNBdG2sSn/rVvzcU3JC8VXKVR3T7Ha
OW2hKzuzRrcvWj+fo8SWjSjMQ3SJqZDvP//3GMfUgCtKkp+sONmxe51RlhAEVAV2
5f0/oB1ThR4YiywOL1/yfh9BwABtrPppMd7VkoL86GBTiao6QA7/MNWh7SqSZtBF
7JfrHzxPcM8DWbs9Cys7k9tp0HhRZNFL2AOmhThdLIbjxd2fUx2+seYd2odxZ91D
nlgUm961+Y12d3xVfRMJrYCRR87QT1r1E3zViAIXeryiMqOhC8FpcE1CRQA6ACDw
LkZUB5cTYY2PZ40zEV7Pk8ShZjgVM8yQfTIrYRAlJiOG0SxJAoYuiZVfEG1lUCZa
sK4VeumIjD8aCvYUmlMwfQGUs9lv0cdhLBBIqoCmQvemfMuLHhwuUWn4jiGvqZry
9XeB6EOBkAiWfq9owoLt+1QTkiPbdZUOoaw9YuAlIkUBfVYl9VS+VnDshE73wuFW
PeSHOvEedf+O6wojkGpDnjVvpDd411p1yKdqVV9LRX+OI1VSuwE9iIqslBfeVoNo
eok2t1G9Z4rHVg6hQ5J8YrodfYoyVhF1b502vrBFvtlBGOVVLpUN3gDOIyqLAwUV
Vwf+R8ioKsqnc8ShTgjjOapY1+4Dvr3AefELZtAAWzJaxKbC/8SCXz8p5R8Mqa7V
cuOmdo12bVADGvpCmWJMK+AuMSPlhi7YdKL8R8CinFwC+nHMjzuYIDGwAUYwT+d4
dPHEttKJF32V0WQMI3JrZ0NbwIHzDMbt9e2h3vgwm8m/svfvlTUzFbBEKYbVDEIm
jY/FTsI04tAgWDLR21dYPH7/0EOfTMc/7f7sx9xflF/mMP4IIGTIA1gK6IaXDcoP
TTCVKJrO+GUgATf6oCp40wPv6UaK/nHNaaGGed5v2BRUMXQ7Z9yNK2RPWxAfm0Xd
67TbCbmO6ur5A+uubylpUKLP+x+yN2YPlnkWhzGwy/KTe9tdi918LwGVWQG/2s8s
HPfTE31hbR7elEnACQ8juxQkFiY8KePh6LoOsRhqR3FoXvlh0TcV2MMDHPgjDVq4
V02KQGP/ANAOz51rMeGDqcVeHjm1W0PXJ0qO6RJ4A5ENZ8Er7HBXUkIYVz2cK457
vCEC+wfw3+veLRDjIW5S1hEfOy4s5jMYM9M9nuTrf3hBlk7P9zIBb8C2LDCt+uJ5
Otxoz1Tm4Qb4PiNkqEA+Up4YCXUoJSGaBUZ63BacIvWYh8UpCxAxg2NBcy2D+tQ1
3IqBXQ8K7IfeqsQet96nB6DrOIy0UGHdhkwSfTGosSrajNn02jd1L1vkLXDwvVnQ
GYQ+v5UTz8LOWamI2sRsQE5yaw/qXaV40dEkO1SgGKM=
`protect END_PROTECTED
