`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0pEXEc6Cy0lPxv+vhBk9zEaPnF8ZCqfHzQvyf76YRlcFkzL5UHcSTVXEIwyVvwUv
JqdYswIU0u4Sz5MV6q/tN2Mj9mpNRM4l+lNdQZCIOhi8Bl3+MlPIBfRl0KqEljU8
l/344x7+vWv4d2v8V7IW9ohHcnJ1GtpKliDl+0yWZIHY3C1EKtIiBWiVLdr2iTp3
yI6MgCY+lywrWmzK7g+V7DnYyhN320XNPvPCPkgbvIpPWkdtw0hHtMopW1CgHP/9
wd7JhN+ZRf3P+i7vEtMz+44vq7wCjSNaCuUzXC4YTRKpG9qICiaS/idZ6bSd2CKy
lQ8fn2fG3kUGIYCJSL2/4xsyaLSK62SlZMsKAJwU+HgmB5ALfj9p4So/jF6bAsOS
NEoNSAp2hzhJ4/BIAVEN8wP0vj+qkHfmVhDM5Ev+NgVOdRNw5HEzSCRQWs1FSoy+
IQaYdECVFq9Wj4mFuaaMRhVhFHlOYXUjExj+y8DYM+yDaPICtjkzDFxLTWLp4lll
U9m5vEz2dyy3GjltWysmDnrPfA8TY2WrIVgr1VuQFj22xcq2n+3BbQpohxrpmGoi
qg+2t6/C/HL2LNXw+9HxHsdyZC96pWB7idd/oyoHYjLby6LDCIaC1MxGRa0boPT3
mtl74RlZaJoa9sp3OOQwX4s1simZLY7/9cF/W1gtnf4qN1njs3pedp5XS7QhF2PN
5DuTo8GkV6UDxaPcqpE/b/qRMiOic1QfPMAL2Gf+O0Ozqi6TO8AEBB0gt1OFOLPK
HWpzuytL0fY+n+wDJZADjAF48o4ecS30aqri1ZJW3rUKv344oW+yUWovBsgUDqTe
6nF7qtmJFL40U1bDs8+4340eIhWjxGDN/UONboX1OTkB8mAKyDhmkqgiavRvR2eR
JH2aUHFseLUcWYjJlygDGtUERYC4WkVRB2wKOVaDHuzuPef/Q/Bp9s4igBLoJZkR
FUx5G0+p7QV1VI89gBM/QzMRa9hG6dCL/btr8zIPk5lG8L9aoRQbjEYTzlqFtHTk
cGYPJo5X3WJP0fn/S9iTHQDZiXg61KLN+YgHSiYlqVlI9LgD/3r3TXmgXOI/XQPk
yLBsip8WdlbMZN5fXb1ZdTJIOtjrlb2RO8QaK73SQPCUiPeFGWzZCloUuLxWl8cf
`protect END_PROTECTED
