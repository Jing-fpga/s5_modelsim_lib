`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8cYQJyj8KxKsqxFHJWpXYpnFzguV5ddelH905FayNR3qlEMlU8bakPXYJoduKLu8
fVpafpyfXjzVAi+NjUrvEmoX/Yo5NNoc/CHBZrvjf3RDEpcoq8h9wHgWRcWiJ6M5
FvsVjiWZ7dGYr8B6e08YiWfkLcgohpLZoePyLHAlItCyrVSstNeU/2AK2E1YiT9o
fvtfJ4nQKAaSjei+hGVhwA7dqwjjEWyeOtJzz3/eoEWtuBy9a+vzfeeHDIOaeSEy
dDrPx9zLGSDaISPtORYMuuXgjfhpnANigAW67lKvk+TvgwQi7QUzCP0AR3RKXM/Z
4AxjtJsg+sjNEVWdCOj44RL456THGVprAQezX6HGIqBkBcLfyCDT+zYPHAyk7o+X
Fd5D8ov2EmTZ8TT9ylOa/JaQwUf9u8NBbKdNamDR2Nz28NIL46Zhqks93PP6ehc6
I1i08AaZ4axsxhbsSwto5Ck/vmYZzMVmuhnBtFVVrMjK5k2B9PFdx0bHYfPCQdZp
In5CU7gOQbiCy5lo4fXRBSLf1ZeQPePoiuLlPyx+dQOoiiKvpnTPAHYrFp0BijK0
xYg8jXxeataj1fT3mmGlDTHNbwFh3Lr9u8GPK8orRsrTMt5qPP30ZNgBgjHt3ET+
6SrgmmIM/l8yuuTH5/QXdkksIhB0JkM5gKE72dcU28jZBvLH9voZrdSe8A/KjTyB
m+JuBxoPXYUBYJDQXSWXKcfpqnohE26HFDpdiWq4E2XkaPaz0JIYJRETTXBrwnRg
XAs/lKE5hYGcQMVxwXGgjsqTXaBgqvuAYKYJdoulWALjZnsmPKWimlD9GVuTDGTy
KfALqGYmTjsfKh6XBXGPjXsepF/hCMHJwC4bHsh/MvNZ0ssQaU8K9xsQCinNKa9y
25CYgbwH2XQvgG3Zu3Wx8/+89PB973jmjvXau8VxqnAf22OxYIqcvgFgoHxYxEo1
Jb6ZnR1w9VkoN9FhFG9XpZiT+1k0Kzt2dXvqXZA35s09/kq+sXwU6xEy1VWTW4Eh
hMFQxgwHvxqZKJWrlQnASoEsKryhpNv2hbH67azLzssF+aQyzz/UbrO2tsnoyNM0
5f8TFTdkD0jgidKzhjxmtdWdC2Vc2fq9qD6pwHvnEjaWcDm8aWgExLMc8i++pAK4
/OTHeOLzhv4AtA3Lve/HN5Sn/53GMPSAcDhfR1ya2Y7a6X8T3RjJ1P/QrrKVBYEz
W/tTvlmwz+r5/rA+9pVmdFaxWQh9+78s1avVPu1oWSL1J1F7X3ELRqdZzCg3MZ11
NC7zaU+sX2UjLS3l2h8mp2GurQmH31LVgYdDS/BL7dp7huhZD1OkS0V2KtjK1L9a
uA5DaW/JdmiTRIt4sDiadQ7VNIzbe/qmr83ifBIaqnkJ0kqyV/YmJmbb6VcBlI3P
ppXgXdLqJbeWvkbs4pzz++8tc010GvHR9M5iKXsHXhRGDLeh48ZSwZ+XFbdIPapw
PRQ3XDXHXQTkSYNf4X4rEb5HpUEfEAs+xmG4uTny9yDJyCHPU0GqNfS3sYAALJu3
lBm9liXq92hbBe4aInShdWCtjMh1kOqSquSbiPCUgOrOfRGibtn+GFeTrHhI4FUF
8VPcOMKnBQSaIj0p5c2tmhfG6NAR8tevRC12+25y8eqmA+TqUxgN8iKqDsq1gstF
lWo+5jjG7/oMjHsa2Lub3+TwJZtl0QLFaG68AEJyjkDs4egGqXbPjgjxnnwX9GeN
OKOhj8pZc9BYjAfNWxXTVmpmKigTFuO/s57dc5OgSYDpW2d9whFolKCrjTewXZCu
Wn6Ty9DsFmunKTS+aoD6G4Xl3d/A4vX8kTum68oQsjIeb7p94oGFHTcb/vfDJ7lq
j/dIXORPDe5hJXzkoQWlp6JPqJv9CRFanCpv4vSnvjLhM8oLxRbeVBRzmdr9spc1
s06Hn64HPGNlNaTAExlsvF12iUTXG81uRP788buM9FkJNuPfxyjoLGQ/KxA/MKjX
JR3OMcDX8nUau8maAvflz0Rn6w7zX6b5UmOWcAkoE10ohzsaBIlZgjg3qJ2oLaeQ
BzUnicmUwUz2T0OaO9ivGC3C24ehvVx4oByiKrLdLX2rzE2ytu3sWMIsmXqar+Xs
vinh/tgG5JeO7IoSMwD1b5bTVotkiKTiOtsX6kN/XOwcnsqed7DHUyKR9B3gUyvp
tXvk4T/l0DQ7zTxR+DOC4hzUvGdfl3X9ch5jlh+xTItrtozATzXOs/ZTg5Cy0D9S
UcrUGQlJx/93KTmjRIit5jA76d+u+4iNw2gOkCGss1EPuWMsmX4jRuiJ/6uBv/Ef
DUF67BuMAcHk3zdF9hGh1BAkVdzVQvwT6bJ/2NfpsOGO9Kpw61P3rEoqTvUVCSPG
a+R5uiDGCLKKZ//E8DTS8drs0OBp/tM6RFr5SjSz48B5mLgJbc8oB60EEuFeb68P
mSpR8MHrsWnok7IEfGehReQRS5yw9y4W0uJ1QWotOEBFh/t51l9Vpn3OL0PbRKUD
j0vnfLNsm8WhDFWc8c5ar7O1KrGeS4++2KCPAXe/QIZPRaC+ljWUhjMJ97dbqeOz
xqL/RrpQIj32VrNx99o3j37cSJEwwIWbXNqhXrRdhfe+AjmK05QuEcYeDeL8Co4e
y2pxnzAiKqOYrOJuuBPc5FNJ7mDQqq/WfZLgqWbGUnZ1GwZ3G2SITKpwxBlb0k+i
NTg+f3cej/j4RCWwXWBbJUtyIlLZp0ys/cJomH4tUYU6fCTw92T7x3bGQ1SD3FEl
`protect END_PROTECTED
