`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VGbT9o4fgjjIub3HEQ6r5DFhlJ0kDw8jm8MsJl1p+iAS+fAJJBCTeTPF8sWUMxWK
r26s8IliCRfRmk+20RhORP9AgB6g0hFo7du9UmYT3F9KVfEkUATTTkH/5E4nO9+8
JOa5SjWzz3BAxdmCzpWinjqS86hTjlbSponV0iwq4aOGv1InN1AOfVW5PPh33NoS
ZlrhDAJETK1MuD51Y2ZparIt7UrQsDbdTxr2e9IRGUcJDYtyX2kwOsmK+a7gRl3y
mLK0ENvPE6KsnUK3zd7CEvzbzDgqujwNkipAlyvf5Ax7ElFpVjIDOmk0kBYUeqFu
uu0AmELZcvtGNLP9/3LnOXpWeT8Btvb7gzXT8hjwmZ9fBS5PyzPvANXEUsZUw86X
5Xgi8oyeW0JEN5uUH2bTO5zou4kTOKVWeFOMsTJn6vF0WpUA8xLXlPjcYvlLxDFX
PMhbQRvwkl5dnyzB072uhY30vYl+PkPF2OgrViFpf5NZIQgPPNvnPn20uGM8h5SC
F8437df9diQSle6dLvqRi0Mswa2/ekeIEPMk0SZ1Sj3t4yCTCyQuMq5Uyj6YATQt
SDg6d1ixISnTSlaZzRDqfH/VKdCMitT7xNmb1VuBv+G00QF1fqV0kpfL/CYUw7aB
JqSZIhXBWlZrbKJ2IyCZvIXNssGV909xJEm9wMLegi6wjhrho59pst+xkm4IMEo2
R9/YcEtJK8xTdudka/0Mh+xi6WUE3O2rBS27+gwAOsuzKO5uVx963QSxIXeSkXTJ
6syzzFMT7u+D6ujna123lsb3FijMSgcm/T5PVBZhfczKC8fCi1nx05TmAR9dNjSH
nFMyVYVGxfDeXWh40+CUHt2wGukXArg0lkxNmF8KuYkCy74SufDMj4W4RY/RGSIL
7CkWufmBtRZx6MdoiEzsxOEOa/W8927xrDKqMrb9ifCDqW3WhERR+etGglNMk9JL
K/jN7Nqc+2EAwsK/bCO1OO0oCEWI9608rjXKigPB1vl3QanMb4f3mxzZo9oP83NT
Yr4VvypKXl2mYWxOJfaSNZY2pp+O1FD5s/6YplS104xqlf4G792xhpFMxOp5GDEb
nzPlrxzfYcNIpcJaxBhti4YnEp599NvFoEIZEamP+VCfzFvA8O3yN9LWeS4iAJ3L
qrhLBSGhcQwb8r7u4JAfQFiHhosABILZJPMivrVqeNrjh5oXEnQFCU5jlT21H4dd
FejDgxP5uHpYf8f0ifSIxlZjxYCqxJIu3l4mzXIxoP7bf998WgeXUd9kdkPcCr6+
FeTMFAobWH8LnngV3siDZnT9ZWIctk9x4+4dLubv675MQ1+q7egR298zKNM4eZQ2
ZjWWIgX52xDAlfbBQXRo+Vf3y5C7shQQeUX5iTP12H/1c99sjBJrw3hpXGjEF7b6
WT+m8OvxpdfiZvi53D0E2TTSyahbLgmRndGwNiLm+XeHxLerx4cy2kvEoHtT26Wb
8BNemlmunravLuOcfOQ27J/xHEpxMKkTRIptKv0S0y48YGNJ4vge1pM4GXmP5o8/
hp9oQwXvNRt3Fml1oy9fuHOpNAXUYjPVC/bgm8RxZau+UG4J60c304DihuAZ88Jk
fa6jP3VYuTzgUMaWN9hNnlgd11DL1Rr9xor/Iv0m90IRN2w3k8XINAa+AFNZbkTF
xjUg9CjQuNwIHcEU0GYgB3BmcFNM9p7fRvWhPNQ5e5XNccEPlSD0cIF4aGI2HIsZ
oltSI7Y7cAhoDdoeIZPhdyTlsfNN4Eip6+/UYNxserGO8tvOQCehSBd20Lm1jyXb
7kGzp8n+8DBsNRYnEwbLQ1IkN4ueNPp6F+IHq9NCFVF43iMIo8PWWwdar8OVUw9M
g/hOlGgvfswc2lIGRAKSs1rc8doGYWVNGV6mBAmkiH56SIr3raK4LsCT/J61h3ZG
GnCI/HZL0Jy4a5jWO5OCTFdPpow/guuTGD9cW9oYBOL0JrGbXQrmwxNKgyr1bz0K
t5XvmT33rOTUa9P2pU21kS2cb7UUGJsl/sDqD0w9cN1zaXB98sWbGcy8/uoBlfMt
zjof2U6VGgOTZp7D9NdDb0mvaIzAdOteo/gTLqkiz8DvJ0R/fcvsyGWlq+TqH8mq
RlU84Dg1bgZmnxw/oJJT+o5maudDCz06b70ucoMouGmVWZyjyD3svcUmUbtnprZj
eLQ20Bnl5CI1p0bBjt9NKY3ZRDgz2KlDrN2licvHh8UgvYsZshmzZ9W6p/xLAioh
Bf4kRh90pX4VsFI+rSYWnxfvBpiSTmR9PqA7Djx8u0vv3jZvN7opjh/H5CbWTRHz
/40OvVDKv+og1uOsygzDLMKrJjH8kI6Ckyu84psnmkk60iQp5Y5856awC5vGJshQ
H5E23+iemycGuT3ewh7Qjrp4Kfm+Yp4akvmKaDxfVTuU5mL0+wveE9bBBj8uO1i2
290eMygoBhCjLEnndHjkKQ==
`protect END_PROTECTED
