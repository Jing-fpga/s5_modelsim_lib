`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CLE9ioImgjSZvbfynIgCTRjqMS1ul3r2ePR1Rnx3GX31uXuoMKUYCD3PojBrmztk
OaGr1v4/6oetsiO/JS3Bq0yEnMLru1Tvumm+U6LSAMVIV2Ak2YWPZfqRja90NjvG
XiCTpB7Og6Ng3M3UaBBXKuXSngPpXDan1QuzhQEFUphf1hUHk55zA10U8MViCIqE
GU22+aqOEe5QsZ+qhAQ6cf1L0QRxsTcwlI5A1JjRvo3ACHQhUuKAfk1lMObEsZap
aEZ4iZb7PY9rzMcv9G6donOh7GDI0BqjcQ8MQfGSUXr2u/uySSxha9Fi0dwCE5t4
bnBOyKBvr6Qo7120Z6QdSKnRM1MOE8qNsAygMJDXXslm8jg7xQwK6YlecdKjaPvy
lF/ILPs4jqqZJDodcUdksh7KnZ0FZdOy/hSGhgsXRtr0Y2AlwYDcdZFo9yoW/eTg
DrY0/jPAttNSbjLLyzO8br/XoSuFOA9NeT6Qnxt0EF942adGI+pyO5BVHQWsH58q
1JLYVe7Nfd7npnhb8wJVJisGD+oDW05LaxFeMSjF8dRI9georWbr2YVxbtfY9VWq
olDiqPgO1JrkCzgxoFKTn0bOkL20gHq8hRrbjFmzoP3Ho/J9simtb9s2b94XxbQc
/sw0yzdYs9NWZhIJZR2QMFfiOPSSHJcehSwliTwHBNRA2fX4AeuPK4A+VWpQiHNg
+497xZmeVVvTC3BVgIaqaVAKGSTlI4omJQ/s7V1ObpCUQuHz5D0cChR5ekBuxswx
j92CQJY4e1FpViH/QYEU2OAjMmIkUvSvpmhGfFgCrSOm1JSB64zSQhPAQEJok8jI
1bRy6X7KBwvaevBhSHNQgbxdVSD+zh1mncL24erye7NmhgTZD6D8LrTWp7zpB4kU
wHvl/TlKK/86iaIggjk2vF/kYobLFUyCZwu2n+eJi5dQTt0vEDIN/M+AisIYpgJq
Y+nGp3BshHAioeVU+N9ZqjA7XHvXxarqdlKi3OHjmuKXBD/jGCQob/0xph6iRWO4
pwx9UhMI8fI2UZ8zzkU8Hbc92HakDtMK6zbJLhkuRmW4F0tkXjqH/mSoC7c7leVx
yob+5FSCtoLQCzsgUJZUYsaqpMq4nb1oRlEavVaDHNL3HKHyZQVZFXUvBBmMNdL9
UnEYs4zatjjDyp8O/UzlgaEoNqxfG0GOzr8672xTZbfq3S/kaxReT27CoYSOvrHK
Q/vpChzuerUAkCvNU4PnZ8MN0jp3ePGbN4a+YBfNlFiOmNBwcG132vJjyeeFQghp
21JRsosR+Rc+FVRqQT+Vw31Kf9IhDTC3MnXaZV0397RcrGb4C1tVKqDf60uqbr7+
xMsthDXQg3BGC4l2dejHpWBDVPTHj1Tu20TTT7UW4Yu8/MHoyaHlN437OR9HeTkF
lK1vsTKvl2RnXv06XfoZHO/nyCnPH27rx892RkSq6W2Zjt2Cm0sToyWF8uIctgsa
zgA5Mf3buKMW9CAETReQgLIT3q4n+auRV3oMnZIsEaTI+KrZHrMhg/vQ6wSSmjLr
GQsAAykOT5dklpOwbsyAe8QHTz40WXySyZ1+8xicyAW8LJGx33OXXS2vZFmD+kD0
u035ejU5UkD3fPubUKVY4RtlEpGpBgbSD37wXjaT5+tk8JZjjSXTbfnp1ESbwXqA
Pf7gk4jbiML9jIsmH4GAN/urylbpb6dE7Fawmx9lQ/RVuWRKvDXJhl5jUQg4inqO
5YJ68tecK82BMaCdquN0iY6manW9paoekHbJPWCBYAwMvUKlmebopJQXdvHQKyd3
GlO4X3YiCReuNjrUXFYFZIIB0+wdntxTclbnt2x5FEbvlrHqXQSZW2ggEMsgWIl/
x0ESwdfQkSLHlOKGlTPqYXQCInZoczQeoYDg7uhYzSdGXEBX0yFyTXY3SAX4xir7
UqEPwDFaK1IVcTCfi/6wsgW+dHeO3aX9K21ieeuziLCPMlS336EmVzVCV9fr41oi
+gF8X4BUrjwU8CYtN6xrDIiR/PFpvG4SXVddlDwsqZ29J68rZzFI9eSrERMy42CW
+Rn5wVyMwerXm1lR4tEzWvigU82Jlniaw6so2rgM49yH+ylVhjDpcUw2RWXEbVVT
kwxbClae5yTl1AxY4ISuWIr9SPdqNqIR+revP8s0LdiN4I1wxsGYL0Ai0zcVQHcB
L9UYsKJRYomHF6I5yFdddXFqTBcQa9tWZDgOYRKGgx47Ze3XGLrtqv2JMBo2gptp
y2hJ6bBKWO5bF93b+7FVY6fnX+1I23WcXQ/Dkd+oGvbSFTVc/HfXXUrh+zxgAGlK
RKooDO7Zh/455t/95nh2GtokIOr0dgknjwwiyNTTgo06YfYZxfnY7z3E+R4MIXVh
xCxipJQ/rzYE6+8FWN2fvW2/d6Zh3I8pEbu45+4qWpdURBdoRdGlLsqAy/ZnV9IR
HtNSSHYMFpSlKf8jwjfv4c8g3HYAiwawCrIoyedYDfZ+otNQuECork4/7svK4NOc
DV+/W7zVS7JgIDVdhA0qXArRgtTlWa11RjRZPfDz23RASRzRDKkAClWSW7RzzqUL
EP+mJVgSQuIFCe0bd1+DLLC0Z9G8lgJAor5lewnUlBtv8Gi4hsNqXyO/3UEFNctX
ahF8nNSfVE82pYKbRe5oFQhrHkcVG8TUanDzMaxqOk/spnrsDyGyqKG8kMJTIWEv
GIkQUQ+GZcj9rMR1pOf484gTCEuu7T6gq4dN2If8fSXZ9nLdhi0O4S7kM57U9nDZ
9VhTO6KC57y4ErJkYQ0MCSAuEdSmqVHyLLR1dQAXPAUXk8FoKgQlQ4BMUiQE3u8J
mloRO/sNT4ttiV77aw33VXsgSDSh2O3UPFtwP5Zdo09ziK6E+hP/IHEQRRaOkr2V
7gjhr5LaoECf8IwP4SL+t+CtT3uy09jiDYl2jy5E2b2saqfmSF+t3jaxTx3+GuY5
CAfv/PEjNLk+nsQ1gMKov4eSvhDpOe9AoIuuadKWoiCAKyLzhRfMZBmxsYBzYqn0
N50Qf91YCnDwuSMjKAQUkgjfqIC2jJ8a/h/T0EJHXHJDVUWM0kfTUSKS+VU9FkPt
nEoVuY3YETVic0k3R71PEfUxirGY5E6MGcgMb7BIqwYiaAW57EP/GtkOBjoMh03d
6syr2xqH9t6lXK5QkbLu9mWgHdYRzK/4c5ZI7hBkBkrKEG986E/EwAk+bw/nt5XN
7TqgWrg248dn8F4RQ2YLrb9yT26PyO2GegSRtQzgjH1Rih/0JdbyeygHkOneuo89
0dwBRFQ5AAeZAwehIiaI/ilpNW0cAXBvlZR5AQ1rIZr+yi0125enSfBvSa9n60f/
zv+/+aru1w0Zox8hUO2hm+e06WyzXzTKazZ+T8WEZ4RYfIzpZAB6lLdk+qTejbmD
Ts0Ks1Vh5cm3259AV/jhf1BZyAAltnTj4qFwLqhKCCMVJHPR9LTB2tW3phCRHnaz
wm4ygQSjnbamk5vqsJ/BKfm6DwX6q+5ibXz6Cf1+w6LvhOBicU3Ppg+Lyziw1eW/
ucwWf21u8HdLT57xQIEcPA==
`protect END_PROTECTED
