`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+4Ze+D3KP3CeYZ6lFUdZP0HjRCyL6TQ8iY4oKJDQl6xB/snIVdK+EpvljE3Al90h
6oa+PB+A2IXEVZZNDM6ZxWnXFBA1Bgc+5SveeK4CwVt9FNrsyqPlTGnGvFQMmGyJ
Hi9HsGeIdZ+oIBzbaDXg+x3KwblkjJXYZT2cSZOrviNNDJ5CN2p6+/smRwgRUst2
4Z2II3/xt37cuBH4IJmo7sxCDUkImAJr0uwXg3V7C0uLbYjw0LFD2l74ch3FRGB/
y/KsRFWFbcQRQQ+DmVro4HmAsfFQCCsHcTnAZ4lVm56Ar97FfelOCQYE3hk9bL2i
K+S6ciIvZOfM43GrU5LF+6rMJF3W/NvIaCF0KQeDuVJYzPGYu6SfCy6zwq2v1vnJ
DnudWd6yvwMxM8X0WnLhTi0LAjGTa0DrZOfHPMBmIISBPjq4F6F/mUYO8MV95pvd
etzvkd6gSjLnSjuZo9qmgornSn1DUmzsxPOMjvKcE1E=
`protect END_PROTECTED
