`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MM8aw9sur+a/4oBdzHXTQqSr8o3qevI5leOnTTm7H3hIOb2lCawALjj+QaWSt2f2
4QgUlwp8fkShHpFmG7xWpIQw+SX4SlIjmNt9kUJBADOGoLo5tjN3UjAns0Q4zMFQ
anipj6ZAUyXvM5W2j25GWzfkK0rMneIat+AdFvEhWfdvR/qo5X4L4MZjx8WxRtoY
Mq5OtILpbXS4ANOsDZq0uvhkBrJlWhJKR08S1OzupQyaTVpDTlNuh8M2U6aq90EA
+aIJBCxJna2SuilnlnNIG0tYYu33yhqnE3MDIYfOStCHi/0R0NlDAR2DG770dMW7
p9mHh5SjWQJOeXqT8Jjpdjw4Nqb5jDfVRute9WdQLChbnmsr725Da1fjMsF1zhJz
Bm0iWq3s2SsKF95XNPEcpbQ/DdGRCUbYm/eoCYaI8O79V+pnHrC1hFUALp5/I6sn
s2O2c0FxreVWU4jtRmycoXqaQKCRywEUKbZY3WZWH3N5AlPEGdvUjgufh6fHygAE
ffSbflGj9wIqBTkU8mSK51vRVHf86OPBBnMual2rHQKxpAT1QAt8LOY7djpUqk96
8regK/mhxJYbvQJOBONSzboOPeLpT8iei93Dk12V8RoBSrT558TT9jCcTR+6m/cZ
waC1pzIa3hr01CUvKtVO8lgb/6s04/IiOye02iufCPa506Rqdrm3vdnWZeHNFFFQ
jiROZJz55LX5cl9sFTd5tw5WJKTKD+XV4UQH2KG6vqiSllnVjHvRYsHryI+/4Uye
Jwg/RHA4p17AVDgVrjZpuz8/wP6icMWejrvIc1fYtc9P5fH2+L82MHq3WGcCeTS/
OohXNT/Dm0mVkOLe7PagFO4kVXaZbwOwVqvXv/SyJqliBQ5o2cgd+4GKQznwM7+l
bBlilJCJYEQQd16oByJOsgjC6lgZG/sQhg8hhwX44AZ5GiFm1CYBYaEB3psEWsHI
/pQ4b6qX8H4o8xALmNlDj+VnXnVshjr/M7nWG1N9U9Jh9Iee8XDEHn2Jiswu5uEQ
g81UD+woYCgjXiR9FofmmXzhqDQfeJCZ1uH4F5p36K33RESGYPTEWerPeLMoAyuq
2rh0iO2/sDTbyfDK40UNolxPsClB7fVfPKRzpZin27HPc/R8IvwNQ9Yu4f9WJNAa
xX+RSw17Ucc/UEJE+LFn7JZCD6CXyoh/eiEPRuEF3n5ipZxZf3BzS8uYarp4vio7
dx+S88xjxidHiy4UDIfOrZGA+k7iBgyOwASe9Zuh+amKKVrjVI76OAqrTOC+axBS
kIOa+k6gEDaef8i7m/sy2YaFGDntLHRyNno2nsG1q/sjQqC8blEwGcBPGBojB7KU
FoMizU/YFzXB1jfRg9H80U1fBLqhCluGcK7SXWLDmKDuhL/Y5WdA4EiK2AVPRUlA
oLXO3kx7QFBNQB4br5aEEI0W7L0CTs+i4CRLvyuWQVju9JWyZPfjmKELurHj+riI
9m2gOb8/jDTxslWVBe1EScI2nSf+7eGK3e1k39u6YlThiinItdorRZLtkG5u9E2m
XpC7zMvSrcR6yMkCWDQyDlXJ175lUdgimTvpEZy3ucvkAel7w3zX7CeYiAxiWxC6
AuJFcl3vsqa7PyoJDDfTv45T2l3Fq2tluDkwbc0D56uXb5OMr9kwSzdNnqw7TeZu
cGUybo0DkLCU9YIOpRy6z21250Cxtxwh7gU+0+KaWbDgHRs1V/lDyXCE4m+MNW+h
ES9FTL2FxJN5lc/FmcK6/KSXLkwrKxcapkNLdzHfswFxgV1NhzEFO670TA35493l
e18M9Cg+w7BhX1edUd1fAuIbvNcci/xVVdwmp+e4A6Lyj0ZqBkwLujzSn4jD9Amj
X+x2fUmg+1FHO4LiRlr61D3Ydp/u4Vev1mj0KO+CQuxdHDwft+3OjdAaIFVeJ449
oAZyeIZtcS+SDU2vvmePc5Sd2s6qSn0GKeZcWc6nx5lgpyoRqbJp7BLBeW9fK/GN
RH2+0gNQe2t33l2SgydAy/2F5msH5JpZfrQj1C0JsDEEJyT7MpqtvM4OUngjwflN
pwdnaFOK6LafiZ9SA0rkDzzp7L2E81UFcdYXBZ/gVx6Tnyl43pPrdItucVd29fa/
fd4Ev1RcowBFXdtUkcLyBSKmpAjfuUyeKyzPQdq7sEeUC/2ybBZJH9sZ+WJ4eaSW
r+Mdc0JxhnsDKD4uUFdkDQ==
`protect END_PROTECTED
