`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
apbzPpFzDa07mpihATKJNQ5yaK27pdu6pTkZ9JZMzRoi7/WFYTusykFT+xkNBYvE
xwoQBm+HTe62KBAAfbPRZK0+arhKalrtcRIapdn49nsdoU9+KEgeNDvzysKP5EA7
WNyMqpS+oPYjb+ABmngy/6+jqvCPIcEqjWj1gMnyY59ss2sxn9V0ZiS7R73V6dU8
H++n8HQa/0Ej6C4nmu/41ymtRVYGaJYH2lfM3S5KGvuwBTdM2iJyfRN0IHVYpIi5
ZbyaAzVvG53EXZz8gVLszzw3EB5wFPFCUDEynP91H9hrv/U/N8Naun2ogIJeP+aN
YtyB1c4zeqze+UMNQRdVZirM/49+O/9B9kW/jYlVvxwpQz1N8bxSesvDUCcDTKHu
e9jQJg1UWmrT8oUvli0sOk0HGHQV4S+Zchhzg/NoRXCeezbFs43MYJfji9np9HpV
2nK7nb+bg+ReOAyB3L2tgHViJIS/IBbh1C3OyIPtbKDTj9WAtYKfXHbCIB8BWqWe
y3qCEReVq9WwD8hNg7cdaeEPJ8bgtRgVf+Yw3MqLaZ5y0VyLQaNx0qLOGgKZ0zWL
G+3W1PVP4vrTIYoFNIl82CIXYSL3Wo4SvxxIwpx5HdAPgrH1XCEigFX3SGd065IZ
35016zymGLMezXLGjZ4bOXpvqDxeQidzneV5L1N0kVy2LRQYgvg1Kfn1jtbF0svl
2BKN5kWlNhjdW3Yq/5trmQYkHRcA4AViKoVurTfmRBo3ShL0qOlJIaC4Yd/oAnJt
t6+dOywEWJ2S8GMBWEMTTsAzkgCyg9OfX6cQZi4qUq22uQtVK7EJtGtD+YSWtwI7
33kCUbL75e3cfnAlT0zNsgyb1Pm6WAj1SzrhOA0ltWrDSa/CB1VsEcnsoibVG+Em
MhuXjgzHIxUcpyreOBbJYnFarB7blUhfxxAotaxC4HJl3HEY7H42eY035fwppx8b
Npu0Dr+93/yM1PwXHBRik9FbhDTZJvWm+6nYpasvFhD3wusKWhlz8EaEO+So+kQd
qmUfOQkQwmUOaySAOOLL1bAiF650A4Qv92xTyfkn3luEzXN0+rwSQnVHnQhtLDbS
+MSj24hPLipczO4pBYiLji3TziNMIwmZ+e7U63lqtuMGLJutUqXjmxfZAKv8YkcQ
+fvpvcF8GzuHATdjgm8ntjRfM0OWT0XnysvWsR5pIkfMfmGD+PNDIImC7IZK05qR
EwgkZTb8QgnJFIzXwx+dus9V7EKDmrdxVrMlofO3qU8Ml68DOb5OS7akKZWZ4W1N
OCh2TvHFypqrc0AGslDQfqeWZHN/0ZOcuK4zCyTSawmsSgaKPKaVvuHSdoZ4LfFI
r9mr0T+R/7rNX9SyX4CPqpSkl/RKJU9Csth02LdoNKiznbYeronc8HrA0cISOoBU
Vg1fhKk5lqcOeGV++jjvfi+bPhcoB23gJFMI79xvvHuS/0tnVoRv6bzSh6zknkBj
b8O1Ih6/QRCc9XZCXYc+Wfe0h2Zy9wmGLYrnRmrMH96GciL8/AOgMrIj91F5XeKb
BJ/nOVRzgitl3tulC01vdCTa1fWheCvABuDf4xXXS+a+INkfAbQYoOeeSRhVWOVu
MnqIfldFFdfX3xKch1EjRi+06pihTMDkwxh3zjXDJ84Bu+QbPgvfo4ms+eN3dm2Y
26rWC6bBFqOc+Htv+s8ObccWnVr04NbgsdyUGQn93QzhslHy8Db7IhZ2YRz59Xd7
4ifr5nLuzSjkQY65y5xni1XJgQHKo/rmZ/8j/EnwZmg=
`protect END_PROTECTED
