`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SVjEq7nX8Q6PfqztvA4losia0RmUNAKH1ps2sPQ5JkLdPDeoyjPPNqkee/ussa9z
omh5qDmrw1bHbr3CCHlERp9h/OoC2YcplYdqQptFceLFC1StnOfYKLOcjDNQY/7u
xElrj7v1J52SJ9V5rpDxD6BnYITfMtzhYihtWsSarXaaSKIfsH1bxV1EzRlNgyQs
I4HVjT1zEf2TOLI52cSIUHho30ix8YnXjA1cDHqFP0Cu7JUZNRnUOYz1FQb/8HCj
U3gGuPXZgy+RBaf5DyPLMhOT5YQ1OLa0QbIzL9OMQqEMACmFQvzVLZzZzlUx50MY
kGzpSLxa784zYtPwexg5Dk2NoM1fLwhc1nh2F6zkii3leq9/ccRIFGmHT1GItf4Q
3X0+/TEvPsAEhANwLrUEyI37iA+qZtsEEWy3o0fCoP7d6cgt3nRyx9VqjfZryQp0
OGmi3S9tdp1JYKOpawNRl6wI87rD09p4eW8l0IAbheHR5WbfOMSt9MUe16fdXzJ+
XKugeC3C2nyrjVabddn24MMu3zJ8PkZIRx3F5J1uGNFwae54TmWS28GxgkXWic77
YLXwgOveabirbSrdeJyjOtQ5WLCAIzTYMra+k748phmbhjOBByV50B06GCva3SUB
gg4QPc4LcCtLeTcRQjec6qRU/UHv1opDeizvUK9KV6M83ntTccZodVdfm3cdtZWi
PsKIfOvMxOd+LLL4KjDb6p/zHKa3892CIHDiG6htH4Imvqj1HbOPHfH0lAD/uKhq
5dNFg5htsFJSFZG3xDldHVCgAhzyKSox93piU88J90iMyxc8ALG5/W7aYmCWUjYi
ik30826xwYbvejU+KpT6LiBfDIuCh91Fa2mY174qYvJ3c5HvQHWlBXarXwpw9Uhz
yIHuyX9Zxtq9HPn5VUTHPVEc+xbzlcfOYcPlRWTztCg3hYpyPINV+0y2iIHvI44G
xDCSui+QbGW9P8CF6cztgmCmyqwU0+rlE13tkFS139sXH1KI0OqZ/F8XmFmX6mHe
y/M3QTaaOPouSSJtm+vvrEcnjAbl/hCYZBAHtZbdlP7eWl+4x2Z4HiBgkLHJRGZ9
u5jD7hoJzWcxF9q3cOlhGYDEYPEkOr147JVKo2Y/6JPpEPAmFXtBkfJuarr6C8RA
mV2eUO+eWHUZ394mF4nbPcYy47yhuZLyq26tQIFb/arUdSzSzV/4Exmohaj7LS6/
1DKNWNW85mREqeqYhkqdHy7pMfLi35G9YICvH3ioyp26lYtd+NNLE3hyDQHYIOPI
F6AKftuxftqiUYB+foh/Qdup7AWbs3QVMjAikZj2q7AlJacER9aheBrL797TfXgy
+WWdX5kwel1kwVrKwNgChCewjUv6T7PxXrrL1T8JCOk=
`protect END_PROTECTED
