`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fd16VjKKc+GwTtOE0l3ZcNKdEU00rjF5T8xF9TMKKImchJpTNDdtXyy4Med06K9/
Qom4zlLS+ULDt2wM9TDsHVV+EU3ClUnMZL/GLuD9kUblNM+3TCJ3CIt0PmTxeVm8
G0kViA3FZStHXoO1451cp0qXs6EjjKy2ZDQJM66xuGPRRIyUEanCjtKW9G2VUBTJ
M85SWdcV0ywvtVl20U0e7NsHPBfwwISjLnJzUp3jzY80/VGDjFWOAa5rhnAum/R9
UBu82DrdNNErIb6uNbUUpWznbonTS7Jc0PUc21W+MJAqaQ7zDUxIE5PfLuTh++el
eyROD3wIfOMgBCS0nZhT/hBxD8qWyWCzCfjMh0hR6jOT6tTkB0PsxNNm5v9tCnk5
AOP2X2V0Guj//aqsDMdFkIiGacQpJquOMYZAwLVU4qdMgQH98qzbQDc2SlG79zcZ
HNc/TWHejv12FgSQTcPhDpCFc/CXpb9vCRtL5GAebLNtEneu29lz306MMLXbSWTC
jYTUqr3Ck3UIH94hjQggOwRn6zQUjh8ZZkNvyPVUSxN3IlRtHFxUgaqyThV8TPxf
wHCoYaK7czVj0P92WrliHQQPCyLlATHVsETP2ruX+efk5zb4BrJ1hMWe9f5N1jh3
VOzBNy5+fcVzciuYYDiYlGDIlGUMQ6tKDVd6lJlLzRX6K9DTNM5aD+DSnyFZmurz
O76qHycNeKCL+5LlUUoE0ArawNy3ZZN5JRaBZIqgwlJ5psw3wKAPTrE5ZFVZcE9D
TlalpxDTfrxuB+i02VX3Ex4niq2CP0Dg3LttQruP3IXXz5sgxL2tcmTA09qAhlII
sOkcQVbnQSkhswH9RUSCbDl6+VQvhT9r2Ro/lRnkl8UfNMfcqzqCWcoX55wRSpEM
LhJht47tP6x+H/16DP2O0Nn4XE6yqUrVkxnBR0JGOWetuWZbGWpSWxxeJQPsq2iW
7KxLTNSAFOnndVvm+uwAL/dYO8tueaEgmQFrhLamu6NMqTco0XKX0dLzsrZ/ZIKS
hf28xrKn5nHFCxyBgTkNt3HHYpQjFBybVZswRqhMcmWfmMkdiCt7bWWG1j1wf9Te
BKjhjAlnS2dTjwS8F0MwQ6Osn5a+Hc3a97abn3NsYB3glG+KgRwBqwYQObyFxKNz
sFz3B4xig1ZftfesLw/KkO3uMXIEdqdrId+9VA1md2CiejYbjbxyFsC4e3F2Nm/v
DyIr3Pxe1cXpzcuHG8U/A+TWS+atIt/L1ZNp41cY2YcEIULIzpMCS6IRFv6tFSNM
lxEr0O2tKEtppiZ+ktm9zBAiFQrSCzW+KPFxApUhsupQnJEr5DcVilQKM5n9WqTD
DwRlMEI6IP3KasOo8A/mS2rhgA3mqfcg0gQRK4bMe0OPYQh7nzE9wS+LTipLCqEV
1VwwEJdcfjJretbM8GGxoFjPD3wcGo9fvcowyljhsnFHVExSWBNHFoNvSJ54KHyT
wkeM1m4HqTwwJsf0thb48qh7EeiMlQuQvqWAQ1ovk0QcYMHKO4p5dVbAn0oMPGCq
gri50n5Rt/V88zmfsFfaCfI5vYsuZlvt98J1j7qAD/0xpCsRdJe5yAODUMyVRrrA
f+AUVNWk2bzsnrZrzhAc+BeQ3O67Eww6HaVpnQ75PHV+ePDtFpdYTWmrcx2OSSFR
eVdNkItoWI6BaMnE7d8FH3XXbWFuZpI5vmmngeqaaSlIW5t7ZSB+ewWJueZ5SNEx
hhPU4eQDK+d5stBNFu7g5Vchgb6bUDQ3prrwPBKbvHC4lnOu3ivFXD0uLU+Oatns
IBBkXlncWNhg7bLJTPYb3LBeiBEqUppmkXJPWZnCtNkXE+QR/p9xLCmdPIp9kkm9
jxB/Ophu/mf6u8v5fMRrXHmJxeQhfQs/cp67J+opQyn7H5sFvlGuY1R1SojeqRzX
30TN9BlHLdhFl8t2mXZB0j5bAJutUul37XiHyWpNAYdV7fJRSZKzO1YpS4AlS3dt
Os8OhrGQkGhXxTXc3w/JlFQHSrpboRhw/x9fAdWiDtvPnVRxQ7gTMckFJND3oREg
FJOqzq6RXy3R8XZc5gYLiyYighVKbaK0cvqB5thaQ7xXG0ClzdAq6sZs+sUd5MA0
NWmLP5XWEGp3S/L4GQQltPzzasoQaGQlPCvcOo0dfTxL9dNXE9UuMRxIQhP4ZOoj
xIt9hZ/G2GgrSIWXFgKAke2MxgttT2myuEqGiiB1i5xGLE3tlwTCmQSeigX2/4QP
E9QjQ+YsiIi+8c6XLSQot3L0CLoM3PmYzXnzeTzNHpHdoqCzpYN7Ph0FwvPn/fSK
rCLcVzH4Di42X8dPNT+qwzrPSGun+f3Q2Yy3B8Th7YFQJKbZFgcIsgFefITYOy3Q
LaQjH1bdEUs5IRWPaJwU4PBSL9uLNsKfeQEd/hoUNm6C5xiyJFM6x7v2HSFQjvCa
tHfGm0YaaFYY4YH9FhH7CW5Lvx96Rwu7L9P1E5KlsN2D4ZbFBuUI1DkwUr/odKWJ
2NoY7x/oNj+dXXAppGENb72IkkmLp5eJ4cc//pY/8sBYuOeUcf0UzoWrh4voDZVU
`protect END_PROTECTED
