`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7hRFtbO2LkccMTZLzIHZWudKpaZaYDJW3diKRKDx1lI/5b5ZlAvQVDewQZzQzmvg
21CyQftLs4py5Jq+oHvwd/g9FcKAiXfe6sX6gD7aFt8HFeCxRsZSgPKjVWBMMThK
SP8aiIwku2ufHkFnR4QK02iltLNBbIspgdgp78OMsJ+gpdptHdUHZXJkEMCI5RYW
BNXtLhaCPhvhSE5ZrB2lLKxtMLf/IVn/elRYREJCm1vQRm8T9arm4wwLAXHJjJKK
bXPU49A5TySSmZEKq3JyEvx+8fHZi+9/e9uCgwPzcvxhtbgLEf8NDeIpfkB2iqb7
/bsh7JhLZG9xANXq57G4BHn8WM+/qAStCcjTCOn54XvQenc8bsfNTBB1mAUgUPX6
zvQl+kzRNixCnU/Nkl4652u0j8q9CwihvRB2t1yIaoar/rJYO9u0PBbsCKbj9bNN
Ps/Wsyz0z07SQeWh4BXHdLr7q/pYlvtndq78g0JdUKXUjxKSAEF1VbNILlyS83ez
5GImJ36TDxe896McAdRmPotd3MCASsenAnGZu0csMFmSG1P8lUy3lNWq5hT5pGER
LPFLEYU0hM15LSMaJypDKQJS7N6c0/rysBn4QPBAbyxBGdKCbhKo2ikSS/R+LO9e
IRK09Qb1iU77wcglN2atgvH6j06inhXnRoJdcsSJS+n9szKxCwt+w+9+cwFFYzRH
tmsIeVQD0AY8VVL1/KEon7mnZqYb6gHTcvF3WA4ih3UNUugjDmDZzLnNnVGYyE0Q
WXCCTnN3QK6xOHye+Bouqd34oBU9kZLYqXc1r/slsRtRb20GQPhFbvCc61VbTo4l
sLOqgIg73RhTCLecQGlNBfx0hSEjvNBbsds+iLyArcLKu966h/EMn3KbGkXUwdrQ
MWW55AjL4LDjzx+A43VdE1bD53ndda7DO84QuhV0YlmAPfOJ5upEipC1wzy2/qv5
OGfBSClKZqlt8/zTVHDxUMHz+MRe/R18YwghN6syv/iGsdUoE7gJmoAYBT8av+Ab
1MrFkveMrUBozhMyBxza/AhWDQizRVA62HnaUwiYu1UjNXNkDWuLV7keUJZYCtrq
1Ogc4iBnJJPUExKSRu1diq/JPIqf+XKVXsKX5CpB58MYtMXkLybUt6WQsczFKuBj
Xj06uxVLEPQFrhxcIFF75DsTr7V8GdiWRkWwSy5z/Rgt9Z+oXPM2kLKhqt7ujBdw
QPX31YRxEHjiSVvG5KmF1LfgWBcn976JCYNG1VhP+zYD6nFIVHLnoapVP8silOtF
sG0+/Aqw87mDrjm9Q9IYtUSOzEkqdyy2TBJ0TC936Ss6tyVQ936HP34C7q8VhY+l
KSRNW8zEcII9DAx+dJNQEK+xNsayms2GN/mSTRTh736bgMKlICGNPX0vWMoZuHJD
mC7s0n9DvrInNglae4l/+6s3PcfAgXkocICxROJvEyk5nwyWeb1QVdUY2I4/F+lS
ryijgGdI4q9w4K8aiR8bGVuGhPoJQ6Gix81QGZFxVHV6Rw1Garzb7DKPIa7yPdDe
IDuyZf5Dg4mYDdgcjd0coC3waAhJnS4qtRCfgype471fVXoPHfbaVj66cA95dkz6
Jdk+QnINqSj3SVLX587KXTOF75ncARHIR/+JOfU16RpBEqFWCu0we7au6CyjmAMI
RaA7OrJV4rLMgQ3pAm03mzPDYHBy7a3/8zV3Y5VAVMtatDKg2dZltEtbtFyplsR3
sBZwphexTMRUHvIov5tIfjDu2Ehd7zaGul0OzNNVqZpZcItSY66Tl3AC21LperH9
FwtWQNQwSzEqmo3KaJ8oOvKJP5PLbedrRV/xndPy0wScAiWI5FHGtHU3/R+KVHaK
J5OcbzVeFn5EIGo3wvdJToULps+RhblbUQ7u/sm6v5rFDXNL+zZXJRQJRhyddS21
Y0gzra/BO4NckT7P1urrXSd/04r3tgbg/6DKRSlwJL4pFWPGufYvlKMLWCFOaS7E
4pcr0HVVCgJUrM68j6Cez8TSqzRZ6p1s2wqonWy4FhCUkwNJWokyKpiST13DPEDQ
+9Vyp+1j9iOdratSFfBx3MdSBdjrQOCYDpcAeoNQAZSULGYrgvqZ6sXOBmyE4Idk
PzhjTbTJ2twBRdlqnHU+Gvj/ScDSrIDg9wAS5AQfnAzvb1TD/roN1AM9LtHURh79
b1mCc25OyVb5vf1lRh5SX4ahHU9DliIqqSTXa/bM8UnOonIC8afEjGwlf5piMnmK
F7VqKEqGYgUN5uYi3lfAWDafSvnIJswlAPoTuydTxC6BWc7gQRoHONaEl4ie+3eD
OMS0wOE+PQ4r9RX9MrfIW7eIVtCuvwVcpt+Yn6msHkbpl3n3zzi90YITnJMOoFs2
ry6JJjzY3ivTAfc3j3DBpCvpsiYptRECbdaPoSNh3SBQPNtNjK3mAZfcnl5AyqP9
NhPqq+FmmoAOAZOnrWGRNcdYPcM03xC0ffIQ+OhB4LfJoJYWVhach070G9BQtQ+r
0X93lJhLTaxL1b5EbpAD47L2Rq/hZ+qggE4VbdChR9coQH+3nEvOT6z//PbjcP8m
0+OEahWSdUi0EefJSDaE4Fis/na0Yfd/25Yore4Is3LuFL67itlDK8iXj51WjC4K
xu5NwHpkEleMmlrvxPNP3+G3gmRV2R0w/tc6CXwNPnMYVpzD3Zfdq0+GHxSN7i5F
IN9JIEbRuxTBuIIw5DWbpUScvvNiBQnMajFETRMHFk0rZINShcVVo6j78vWt7Wig
6387Sk0ZaxunTvw8y/pDtAOaOMsaH0wubiadybOvB5nq/4DrvAiMzsutSylUmsrw
yvI1gV5GGjW0SxG8cQhPM5Y5VBddwee8TOJ4pe5xbCz63QHl/SIHJOKRwEV/lUT/
PEdidKsArNNfu97rf14KRaR3IL97tNe7rcV0eMpNrjWJeGjr1X6WZl15k8okqDPx
WVsKTGyq8ypimddQq0eNnDNJsiNUnIxZkgrX0jAFwEWdxTZlP+W5NgQmRsqKV+rs
CRuBPFJdLqxsfSgPK3DI6VFuLB9sqVvojUHmtGTUtx5txrMIcxJgKp46xwm5FHkj
FSgHCYFrkGqJ+XeVpv+8XLR+fUsvgotS+WzmBzvFahuMMWLIX7pCnMNPkCN4KSBC
VVQNGB8b1f8Q7+NaCg2Fq6I+LXavcmZDTwUzIoFDMJGuj0g3IQ8tXPxGVE5SrLuC
b6vqwhlx70RelPR1K/CS6b1EzDjAV33cTCv4jufUPcojW+i3yd9hba7o4glTBHU8
UyIVPrH8GBSOof0gjioxRPE7ID2kn6tiRuvgXlUBuV5y5BUUlkapyJWqYfHgWXWx
I5yia2Ks9EmAKoE7E3zMt//dl77e4ulXPnKEv0EvexH8pn1MggwZAA3h5+zvpOpy
TdAHIxGjq115yZ4xzg+Hkwi8u/LEZX1uTZFJqgtqKkGP75ZaP5eb8JCVbNAueZgQ
7mIWipNXBYVGFX4WWOj3Rf9CATXqowgXz+mJqVf5DLnf2E/x5zJjUG7qb/uRsjAW
G2OxPoW5syTDIAmaMhbGQ7N/Aq6dIFBnQgvHM43iw/lhJvGHgdnBl5SD17kp6g0D
h0KNAYlSHMTuXEisJabCkCWAy9+62YCwsXyr/5obzh8RNZqImHBZwfKCnNRIqKjz
N+fY22yPx5+jgSsZ0x4+UaEe8sPsOSNksm3Id2cJ0lS2ack9qlyjR3kFgxqqG208
ftVg325ZQdxBD4d1b2/FxBZwJYacMorf2GhsQ2gQu76lJzykWJa2ksWexf9liZcZ
ZenFN5pUuekv9GzPI8saaiVN63oYVBiJrjqmDl6lfkUwGiIC9MgafQ+3wSH3YCfI
Jz93qcG71lsVTuGyBtKfQSwDXsoBwh4+9LLACJ1EC9bmEN5vVclDGkrEN2bFdXSg
D6d6bWTIo65njJcQSYuViU0899bSZXQbWz8EuVxHZnkHRr3dmT1uSFsHlNuq69G0
THY3z5hY153YORJA+cB9iOP+9GDTqXyaw2YvEeoXuVsnpJItDCaNPyLyfdo402pW
U3rB5HhwkYJZqaMAetjlv5pC619oMd8YnUT2VFOXAawb8fcCRtPd9KcMlMTrSHsh
c9OwpBZrFSoLd1/HrmYyis0D/yycDobKGkHxJ3M/EMQ2ha9RFop9b0Mfn+Ut4iVO
qjc/r0xTbMwqXEQdBAkvbMdU4wtMQpmAdirqGa2eTaT6ayIbL+Rr8JzKGig7LmqN
1C8+O15ZlaSXO+8ihRmrJmzoYT2+3VGgfeIKEl79fUj45/APVUkB1fCE1R318Cly
1Pi0/Xk2d4FBAu10dM12r1wchQhOJfAsvYXE2FfAQ2avQo8ZFhX3+RJYxf69pF4K
TE0Cs4tq+6YOfXICGiXSciDBAHREHvJEWMzFVsFIAQuGzx/PL6w9wjIn7kLzyrBJ
i/2O41mYucePZ4hfMN7Bz0tbcRaJHSBc7RUYdjj1UBc2vt+gMVqNgxUgMg2k9Iz3
ZTO64irhQ4tkLBFBsQRU/6LymrSxxGIxIIYALtUqar5kmsgqjVEnK0f+wuZ2XYPw
t5fjMYbT4PEcUgIbG262z0hF30YuIh8cQ3lZDSUZ6xqOT53bmtplWCyJ95hiomWT
N6SWH40RxUTxyf1C3HYodYp/gzL5Rdk8+0EBLFcZWvY=
`protect END_PROTECTED
