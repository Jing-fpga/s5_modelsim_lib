`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lIki6D+O/y7MyUsr9yvLQ+AOujJuCJ/j4z7Qwptj6S8mejEwY2B3J+hUJDySexuR
JXI6PwA+/a4J16XH5G3y10hZOqKKJlB6cQpzoG6pHuMtm4Ks3XsIbjPqfuJiD/lO
MyCTh458Qz+wa9lb9SydiSfL6suYQejM0Sce6C9V0D5E2YETNTSAZykpHHhjoN9z
3twsGrkSBtejR3kIxIWGsFCgq3Ko6VP9oEvRjRbeDsFEmZXb9lrugYcR4nX3bAo5
E3uB+SJfQRbi7oBjDFH8QLZlnmO3fJt5EnfNK4H3X9S83OfzZUGXOCl2wE5eFTyk
jSJFF2X4QNdVLlSIEWSEzfx9vQVBIQ1u+2wmnwLqAmyCwXMsLMyZvZatgQbRHf5f
z7NuWhw6LL+o8o73LFNzzQZuDAR/uvAh0BSWEr4x/wxSzSuq063Vly/amZ3mQreB
Tlf6Kk5aYYzoz6WVxScvs1PuITIFNOIVuHhKCOxBQttQtYuvP+nq+mvNXwg9UgHE
556xJ5rAWIhbEblT0gfvwpIa3szCeMwk99oBBVc6uIViRL9I9ruKMjr7HCZr0LOi
dExWNay61W84KA5wphmpcoDe04BCYsFya7joUc4ptEPw2e7wHfQadb9tyOXt2OPC
7l4bdh1Gr4xuJFnadTc+6cY/rDfw/XDkGxJWAAdzgWtAiaNmwsj/rnkBM3uZQqa/
hDsuR/ybtPBthzkwUYw70Ke6ljBS0HZRfdBRxAZ8SNcub+7l4oeBQQ5FTtuNY5Pd
H+Z5Ycb9o98GVR74KBzshwXvcdV4DT2I4JssFytZVMGKKtDHA1G/8wTVqsQ+LMtE
X7npTgGPZ4MLduXXS7c7tqNCq+pa9+KFMmeHJfzf6v2s88yVjvakbR9gOj2bPEq0
sHUyTCNUoUn15voLEb+6AGLtqIEhgBqfTGjbVYzb242Fx/gK3UrGdaI1ss53b+nx
VhReofGHo5pTzjcHGqrloeSWAzUvJNZAiCsCxNUD4jzj1itYnLZI37uaxGmqPSso
xeVraRLEgBq+JnSiIqeqko3YYJLB0h9U5svH1hdQARPrnlh71d9gJcVQsiIzg2qT
GfPTdUTfoGoBf/wro/a1e3kbxQOQplz6TfxKOoD1OrrfwuxUuVJE8hXDyzTXJFpi
sm5yXg4z5Ls9fBk4jpYdQz84opAHZWxgFUdtkSIS8IgwTXVIUVcXBoSRwhsIVfmU
2A12UCNqc75m8T/iTAdMM3OMT9OmOnGIj9EFzii0usz6/X0Y66lBxxr3lD5cb7bu
wM4IQdolqavUCb+GGrsAygeWAu9Ghf/Ba+d/u5Dr+xhyk8DE8EVe8uaWXNtxa0JS
vmMBtc8PHW5ijlSYQosvheej9rLCbwxaoR1Lcekz8KXgQduCvYJVujWPez19FRX0
hr2ExT1N4ZsyART6huvmhEAUaBSt+Dv9zqydK4L5TaEV7ujk86/m77FqPpstQbNd
pDti5FzdAnfDC4ZP19WtNKOohpYb9xB1dlljoKb6kPa5jd4Ex2J2yZgNEytgFzNX
nxrkjE79MlaSZ9U3/L2ED4GiJQReFxhqO/xu0sWd15LjVRkgYDNw36lBEydPV13W
9AcxhSlda9tfY1F+jprhQavr11AiGU/yjR2z7uwqipfKa/xc3GkfrFUV6kc6BLs+
0VaWNcufiTliz4lyRNv0bpcOoSuFBEZLhGU/ZH9VVUyZh1VDG7GUHfbkE+8vM1T1
SwAOem+tqDuhhaPCWmU2gKOrMl7/lUK4+i6r6qJ3acZ9jk7j/TW9uGX+gaS6RGak
bx3RoHKZt+UlSkvDoWT8wqgZskqAi2bhf4gRgZbJZBz9aq4Fsmu1k3VrmtM9YJG5
/o1/QzObzxObXwHIiZ/w6kdggjyZCXyvg5K18p9AvSdz/ca5kEtlaVT+5+qV6yIa
QTbGJ6fv4mjIl99aCN6dXAwq03T526szbYnO89LhalqIag6w0W7YPxjmt4oewIgM
wdGL3RRY4v26nHVyMBv8yL9/r3xH+bvBxNPh+hIcrUmpGcbw1+SqKGg/4kM7Nujm
0bggsJC1DffusgqftWexVOAt/Ehq0WZZzqBfAVfix+/ejrrOWoWNiBmOIefUWO+H
WtHYwckaT2qL4z4BoyvNb8aaIOqz2d8cHdxBbA7doI2hkxGer4KMrVMXu0B97gcP
dZ3d/AiLxcL3TwgYVHLsu+koHAzrZ3GvZwM7sk3w4yjFNN7xjlJPUHAkLlAW8/0k
OrNqs9Rxf1j2YLBj960FLt9kHAAiYB4rM56WoUnawcngnw0lkwVtNWDZYI5w7gJ2
SSYcaL230bB1J6z0Q9B1+Ojmz46pkd3bynGwu1WsyQHElTEuSuFVVAqW4PzoAoMo
vCi6yPmhMQ/wcOpR0qt/nOYUfP0yjayoFqLxpD8VdE3n6iv3K3vYZ/V8rDtIaC8B
6QoTmXsmoP9gGZlW8HqSe0ENhq2IAG2Cyf6W+6qWHW7V4jsMAM/aLQ8lQzxk4e8t
FiMgYnG9rvzy6JxDUXoV92CvpyJVWxDBr8R8epm5lSjlPN7N5WdYmLVRObFIYXsn
8UcYt30o6zIoM8T4I/CIypIyyOI5340vySkru7JFk8L1udX5ZwDTlPJNXh3ID5gL
yfY40MlZgYkHccxCKju9VFKH0eZL8OFDAlt6NhQq+eWpWDFNF8qtbk/MALuFO6x0
i7GDf31c0QjDsJSSrVBHUJeBgvPVWSV37lW3mOrEyamnDFwriUrDybTrLLV3+J3Z
45aveOFfHMKpoJJljbVUb61DEGfWg4CpMRsg+Gu07w35h4k/ouuObogDVvTrUyoQ
DSCCZfeEypWKuzWGc28di7+RNg//xri8huelmc6StF3jni1EtA7biye5PbykXFUA
b1zY1q1eGxIA6xcV/FFF8DmzuGSgHBN4Ecjm2s38QjwaHei7syvfFIJuwWajMfBg
UQlGqmdVyZfFB7tUYAut61vR6L5maLCe5NdDCjSuWRKx2vb+P5lqvCf9GtPuZWpC
pYbG1LZc/df9EYOrKvvaRFKWlHLfXgr9EXG/cHpB1FnwDIXFO5hWXgAni3F0jyDD
pmcdD1PegjOt8aD/JYEKl/J5Co8UnAM2KRU1+HXhB40EjELq3+C8GjGrk7msYqFw
Pbq9+MEbV6RB3TvHoEYIWDKVY9VVJ3S5Wy3eSareE3iJfKvE8ZjrV9g3dZo0RTh+
2RGykWF0cYm55bcfKyvIkyu005FYmMW3cFqeMU01WVHURooW4iwNbhcovHfg8WLb
+mBHOgvyI4rwDB5a+lE9KyfUnV6DziKaPvgfZ+XoV5+S6Eb3C4urW7ISpUVlprig
PDLQlmTlZzYXzUsLxJUkY4sZWC3s1toh7hsdB9CLsvEfQn2i+QsJs52kBZbffq/0
y6bIO7tbbnEfeOE69ffpeYT7y39XC0jvcYYwrCZz1/VCO5fzkrkqD/dUsP6MwvyO
C57TEbQDT9l5HFcUFrk1govarXoj9F6vAbhoBmSElqmL/wUoct0AHF3lNF6ISiN/
BZJlCwctKdkWAURCXnroDKZr2nHqdOwYOfeqT1JvQngdEWd55F5lTpUO9oY0R3rx
J38NniTGIZlumhauzik+n6qXoiM4hVtOESpAOJGjPy7lbgjLsSDsDPBQMnpul2u9
9Dk6tKzwBB1qnEzXhLSqnorF8nAAYW0dNTwNWUxx6r5RQQlu75ztuOqDppsNn/RL
/qLSnz6vpbb1LaDIgRxMExOn/GUCcGlCjEYU8Sgia9rNt3McZCOYQDR6wJworGng
c7CjEZajo92sYmqnFLC/1xFbVf0pwWPu6jAFKCIVT2LUREbL2qu9h/FiHsjx2iJP
jk+oS5Su+KGu9MRjza9DLs4I9VU1m7y0fna+V/psMTguR3QLpwoLLyBblmDJK2Yi
rst/6awsAPnmAo7wgEVpUjbq4dcAphs4PSzZwxlIOAY6AY8OslJ8PG4IN0gMuecc
Ssc+K4DhuNECI/lItFC3CLxT2FaW6ZedU3VcjdDFtZWrwiA2oTOkR9ufCVR6t14B
fD0Yafb5gHgNSx9OHPK0zLmFPYvUTYrWHOKMUGx0gTW0Eof5ss82mun2t/f7k06C
snzRXs+iMp1W1ZXGosvpKV8vRQJ5FsSuklc4WXGf8K6gOlrbAwf7AwCbN39cB/5l
biHbcgIQ2MvXxAI5jGRuCntyE9+kLTpqs5y3WMuf4cilrpwMBmW16slc3TKqXlL+
UAI29BaYll3Hh6eoD2cO6TBI29gb06n+tsO6gsXI+c4/wxAeCq2r+Qf6m6o/o3c4
I8Bcjv3iXPJh2uvJxaiE3lFjQlB4ZfF+Xmt9FQ0EneBINLUc+Y8ruLbcG4oX/S6h
Dtac7MYohoDL8KkLsFRpcZJNYIRMek2O1mrWkVh+0EHGxFndMh/eLSliy5ROH9zg
42Z2szzWnyYBgJIoGL9+8XJ4wIRta7Qty8SqKyenFGINlPQFycc9t4l4TgQGoaBF
ZI0ijuuZOKX1sBZAOsFP/GtbzbQIHP9EaB0CwbrJmaOlSSoeaZkCd75mvhNnxQdy
K2zFVXXTH1Fm1B+yvWiVZMr4aPU1TAb0grt6vo08tdz4WlF8ITkH8WwUyCdLFvrM
PQuW1TbMovIR62Ef8r88PNJiym0Lme2LDDHedALdAE5wp8xyT6jpqCUHAGafoDd7
jgNuHcZFD7IQ+hTd9vDxvq5e4v/C5pDs2EJ9/3NXBd1XZRulhjvizDsK+rEXt2HM
l2NJ1Sp3JH5W+aKSQAX3unXAgU5sfZQFdTmER4oaWvRPfTeUjRaaPREqn1iEDpmc
uihN8m2a3ncTNAE2EnAdZfjONJVlZH6tK448qPA+8YNTLInXmlWe2GJvuGj/WDqu
ko7MzNJTvItrIOAFyzoxgBMj2xnlbdmfE1YZHgIqUo5KCd2S541WJuB3Lkxh6ugA
wgsVuUEBAKDZcXGQ1iOmLw0MFYSrXjWcY1QjW7t2QY1Ca54wXqvQdLmKhbVyGHwv
qLVJWyt6cLup/yRwG6IgGoMwqvM0AeQ0I++DcPZ5rFSUXIXd49Pnl4Om4OKntTco
BuKFmviDeXl29p3SAJzrvwz89FKJgyThVbB2YlZKN6qE9aD2xFR9yY1FSMwW/k8f
pB9xf9xzf4+YlwBks/BKV6BLDtdzBileFrXYrbgESRroxHSBJLhYFwzwkPpWPTGO
0HgXehg446/iasDUZx2Wwso7UXHNRSBL6yToQEi1t/QDT2h6aihgU5fYn1RPqXoH
s6zEwE28o0iktERVZoBL6C04ww7iOG1mFA3xKQ8ywm8+3UAYmNv++sFieSrbYNEl
7zxKi7DRif4CLEvvpfcXm/bVIHcCKT6+tbk5sAyhurMqOq3xJ23dUS5QKm7Suzd5
V/HhTRzU0+5HAtLsRLNOJVTtP0cPz3u1hJMNXGGJqC2W5WxzMeBqkSGdgAC7Pd/J
po3Gi6nhPeK3kap4y/Yss6V8Xx22aYXOGRb+wwAL2VgTaMnRIj2JxUFbiIFuDVVW
1GT2QhD4Q6o5RVTmi3a6m7s37XlplIOCR/XjUjpB4ST4FOgj56iQ4UkwVDjfIQuB
jhAxRtj6hka+L2VQVoLUkIt5lgkG5aI0tHRP6wAFGjoSDKzXhzeFOKPTaIZ0G7mU
eqj84vKnyFzuFiyLGVst6aTvgPEFjTOYb+4RmOFpQIlCXtianamu2uU/HKx9aB9m
me7kTknNVm+mWrFkQ2eCWd1kswDd7REHlaPMXL1U9zcLaoaKr3ZhodIN8ySENyeR
KRtVnoVjQMd5HZGOS85lpbyReVe5R6KmYf4o+RVtGTbyopRit1klNDAQHODtoGib
f0wW7MMAZSVhLvk+1hJIEawZr6zjhSois5GyBzyOZn4FKYAriT6eLbKQ4rAklBZ3
/elTJOEr8HtH6GQgUhqfM8G8eizC8H+ojyhRg6R46sww8hSUJGIYmQVy9DlM5DuV
7IqkhdTSwb4VRthkrM78wSX0pCFkKqEVzeTMET2FE5TCbsEeAFFcH39TCarcuv5W
cUKZfj/XWVEjrjbZnw4mRh2+H1GmlGf6Z+vL2whlH8Oe2PD9y3qGVELZWJa+UFD7
Clz62zrNsaVhqOEoBEucjcMyax2yQbVi/GuD/1PCmtVxDSLYvl1gr7RpAm4E1PJk
lzf31DS45I7qGtVHFSHLF8N5gNyatU8O22Ut+inu6qascUKsw2qCtoom9q7rkl9B
pckNe8wge8YjFK9/VParwf5n+ApL+TIhOQGEnYMSkaXKNGDJ8UN8+DR/OP70cAe/
bJ3QPWNJO+am1FlX8NtlsSUIq1twRe6yrd15IbBcLAOvIZ9IxWxl33U4Jxqa2UAW
fs6nhbAVvHYqBai+JuC4hfW2ENWWjrhfKFhnuQkQLZTOmMTLu3pdoKQAwLMc48ea
wA1oIjTAqqyMkO65t/W/G33ldGNpfmbZA+ugz5nDu8F1tmVP/3x8hH6gmj/uKUzl
TsCTPbACAoulqTYWvuxpkWDOXu/C1TYqWp8FPncFyHwmvJE1f9fn0OQ+9g8/Z/Jb
0gfw91j1z/uvFdAsAaL1qTIHMj0Ny5YDeNhuqe2CpoIMCvweCEJ61lDyrsuOhx2X
HqXTOuhtDm5u2/YLYEGnDmvoyCf2HjKwSXW9ZUOEX8Z9dwwXURDe7y7DaGWBTj+c
QfiiveNhYnRQc8HCd8k5b5OMpdcVfFuqZsTKHrdIxmPS+5S9EzbW8rVpAHbsoYc1
Bot/itQA4WmTa/Pixc9dh6RpPEPbG2sNRqnYjbhvCP7T354zJR8Fc80uiXa8Twjc
byCcwSp8rD0KcHtBWSfpQ/AVoPRda9RWhdhD8KXJdp1swd+KX6jBhRTNiidbor/i
vpJY7+9vOOAS/2ivTV9gPn42qsUJjKVn20nHiyRSxA6ltedurzYIQXnZqFYFjopL
P0LhNpkrCalfDSH+YR52ShMj0QSQaKOUaxakAs4z/Hy1JYeMhb2RC1Mxby55EN/L
Wr3EmH5e1BVu+7aGWDw126eT5Xfdj79h4TXD3S/ZW1YczWSWl/P2f70nyCX2geF/
7OP0s+xsvL0cMvlOm0VKz4RHVynkPx7bCCr3aQ5ZnegVVLXde2gZbLdy1sWrXQlJ
2JOrWZzMJU9miMdqS6+f5BzcrHu9Utl/cA51nKHRJS15a1eqnf/a8w6PuLlveW4P
MILRFsJICB93VZOeiokQPlOotmlKyf+mUtOAeD3D81lhhGMXr50Okz0hhWqO96yi
NuP2k9DU94bRsO5abTzF6nmyOHWnU9ZHz0QQYha7pp9OS5Lnf5aHEUKpdtDDh9tt
JlPwUY2swmwg6bleXwYwgIF2CPRfh7AVrXxPu+rxM2RpvpbNUnDlEZPDQs7blvOu
l6O9vDmCu2EMJFAu9f91Rfju/ZkFceRkEB5Z1wYlP+yYFMkCe3Pp1BawWe9XDQHR
Ymdkql2244QCEmcVRNK4hUQdpEAWiesuFeGnCUGE82RTAIwJGC+3x+vAG2hbKYmV
06gRDWcCzmyvFJ4lF962aP4pMOZfXmbIFcVL3/63WfqoUaQgCyM6S/iX1pC2KdgC
iY/wlzJLA0baVMqw1G03vtahILy4NJ6q41FrGaHdKm8k7Q3pT5WrHgTUvqikuQ+7
GviDsVde+4pgQy0gjLOnD7m05q1A5Q1DTggh5ukCKWcf17lpptW2ERLGl200GNBU
iKZNAfS7bKYHvymfMQ01xitO21HclIpuQ4T+GZByua8zlGXUZyM6y4eFM2vyAPoj
84BSHph+Pj4HY9+LuEw8WZ1buwMKHsXwxbJQ1U8uWifGqV94xcdhj0xh1bBRxl4l
IQTRuhSMi9E2vkSkYw9Sc6X1SD5lLwB1UR3xBwGYxbfQ7XkUEHlpwWjo1WBFZPx2
pmVIyvSxBmgU/JCHP28XCGg2nldDdnNF3XIEzqBDjRlpsJZHCLvnw1+A2TQetcAI
o7HbOaz0OvIP1J0ntSlC0B5mTpR188aoxRmu/KTEf5g0j4+g9mlBYAP8JJkJ/bJg
+Rx8FPwCZnx8FrPm+S7UgHcxWtVDhRFGTfhj3MHb9NG4SO0cId84CbwQifSa9dji
QjF0XlfVmPGXhlS7zQrAuFx/uTQAJlYQYU5BLoozMy2Kle2ZnOf8PMQ4noUiqFyR
t+WxezFYXXO4FEIKZlNbfb9lMoYuO629HnPXUSL9GOHzUO7srOtcT9mD/bDri0Gf
Jd26bK6e96aEXB1PEbWR+FU2MNIW7roYdCdyZG/5EQJvkMsXOSKKC0OlbtZtTWpc
7GbQUTqCHojjbZY15lJfsvJKktcXMipLENDtlCac/NfzT8bt5WSG5vPAH0rWPqdj
ch3nPemO/Z07V22rrVeAfBEZ3U0q13cs8eRSRDIjPssKGzveZUXZwfHZwomXFf2N
BP2P4snAbEVXzBlA09Ar6eRaT4xnsRnZdHCZLrr0QdXVYLHS6KnNXeYjlI/lxoo9
aKDYVpn1oY6exmHdyaIV2IvmsAqCnqCE5jCvc+Z7GlmVrGA3JMAq+rVCI1dlpNT5
NDXVVmqGFvjuJgt4aj15rZpE3uC5EAbvBCZVt5g8czF6HXvQLq19NwIdLA7uJiw9
ULb8gEFasDzpQyjYB9wSn2Juce4F+XU5KEIBvFaHR3NcEpWolorqWi6lfwGsfQpr
uwnLg5XLNP3rL0gnLNzVPoM07+Dw01TTd8rRpU+EqrtB6rcFYd+H+e6ed4bWwWYQ
mEw9Rr6RLJsU0ner7ZPPO6/u4XxnvcQo7MqIBDoco3t8EBoZFshZ40peB7dc4X9U
9gnOr+Mg1qAPKMduCNYnGBXTinhY/p6+C0QQi+ErlABgzO7JNQ5b1xBeO/6CpJuP
jlaRK4QA8yTFl1Mx3gY3MSIi9cz2yMRbrhmbZEakPLtzX82Hc23/oI5TswkRM4px
G71ixLCdb1N/1sosHH6yKVH5aUZL2ihfZX1ATFB5Q8d4Z8VCegNE+KW8mNjQvWpj
cX8obayPTgqfWzytpDGh0CQmp6pqd++lZyf05ixSfAAN4cQzZI8QZfwchKz7Yn2w
j6FHds5mCQ1qCKihCSakqxCvZWWOSNUk3P/rE7Ov/p4ZVr1H2tSzWu8I5iywbsTP
qWD8nQaCDZl6uPTp+O9yPoVRHyJMirSuhVr6X88TiQElItDVoFEw3a3ML68eGypE
mE/BQC2IQqg+6BudDOvp8tKvBYHKqMUhhcNBuB1tO794NSgUtCrwNe1B0tENsO3L
x649UQEXJReVTrvgNBHcW3nCDyf8TgnsfOvNY36syKBpUio4KAosE+v7y+7KUOmO
MW71ElhOvg6bxLkseqWnuacRffgXy5mwsdeIa7UUIjrLot9sywt0Kp/Iyf8sYxG2
LVOwHBVb+NOiQcBI60u+r9171nOC1g/NQ3kVtOEz7A+/5sPkRCnNAuD09eZ6z5p8
GbtB47lQDZkaJOJfP0D/wo2I9ebnDLWq5ytpRj0bM7mmAeAv64CG0wVILBejLmba
DUh92wwCqkZSfglbfbpnmH50lNe/J9VnABu5A13uUhEejW4CTS/sjM7t4CKbaG+w
HBfkvDESdsGRfZe7cgp3bhTR8T4/F5nBR2yedmrTPq5CB4ju/pup4WJeSTMJvUNg
cynu1wM4YO2wF21Gg39nQ7fo+uEc/KX9etnIyEzE8WExl00+DPghkOpCjmj95DSW
UScysrET2MM1CpCvmBp5uGnHy38tRthJqOxtNPsOMIJVweLEkuYLPe7NXK4THvAA
YA/VR2d8k9NLqXCaeI8ZS4MpVjrsVEyj4awTvc28ttJ/Zh84v3YzBK5Zwk21I8fx
gj7QpUGIQBYWX8qmIWyPz078p7JIrQvH1TGYNYJ3p+vcjsEeYu7p1G80L277XctE
1ww4TS7k+LvreI984fkiYj6ejLSil0Y8bgo+D1PP2nYjI3lMc0D2wJA5NWUSTZgu
y1OQT4AEeb7/rH2mClqoBsVxC1O0AR8IgryWnbxuEshdgoLkRlBGF+B3YnSeyDAC
rifZAnj6RRDiTZsnCuKO+AjXSGrPkl9VUYYA0gF48I8AmZra8W4r9nMB/Bo+bwGY
nDUebfmFYGlvFLLFoqkiqdqItOzwyV3j1IUaik0Rn+3NTqI3Byv/jAOjlEQdR15q
x+jY3KmKsXBZ+R0mfitAEb4V18CvkKPE27j74fc7mhZk8ZYe+kVe+3VtkaQ5O4Fe
9kO0ZBp1MmZ4mg2Ph3Kf5dl4icPHML+q3pSAsCcPFwvldyiDngiAILMPvQQTfRpI
1eMeQOrXd3uzGQyL4TQDBrrrTFE6MCQtMmP5IfHYoEaCO+rgrLxfPh7aQZNKbSrz
YNGAgj/76Ol2oWfqYx8hik2RBcOn0xQOKJHymur4uXZqv5zS/DZt8UfpqdV47LGK
7MIPI5c0f7Po7pb+bvonJkW+MQjI7e2piXK8BXzNmqTQieRVKPF1whm16JvnQsAH
/2cjs2zerYDcCb05IscWVcIlt52XggAadjVznQiFsXF0+Zo3tfArgDlJvsMatPBS
TB6zy8m+4CavZsljRicgZFqDOvixn//k76wVSMBWfEgwKliQHzYCcm8lrJh+B4ob
K0sRQ93dZOQBdwOrwzGjaWV2dpDruNicf8zvLC5jGooAMnUF5P9+FFlPnHqOjVIn
IHR8qZzRWyumH7z+FX8Yx1dGL/y1Gxf0gwWkJh4o5N4F+buuOIw2D2lR3g5D7bBR
pGkX9mUl+W8JESLEP48yU2VKa2TQu62HFU5HJu2/qoDD4D2OZojBxGEGHurLBIl+
xNw53qxphHE5SpXV/3eWt9xDIlHEPveKAgHt5FnTw6wpHbM7cY5GRK5yJNtoCca+
UFiR6OrQD/sonJIE3YoRZzvb+AkA0w8aci0TdZysB9R/8YEarJUxHLsDXsXuHmlC
CTZj1xMwOi1xQqt66wdef36IuqqFhDXh25DMdcs9lZsB1l/loGuf4AwhxjWe5we7
zxEZjENjc888WA2QdqD/+hrDmFJJCdOroFvsNF7Ix0BtO1VCcuv3zNK2O3t89l7L
z0egKCOCC/d7eQj/kHkrxbhuURFzMBGZ7fgFtvHA4AwuvNWQ+jU4+rT9bnc8ieGB
T9BaNJZ2aD/lVPsZ5RIQUxAZFPWf2DUhf3lwAGOj+Cygl/diqD8Db8SzftlyB3t0
WAkAt5AwiefA34IcahOXhqK9N0KMoaBmVE22lgO5Fj3SQ3Ssy60qTd8zN2iBfxUG
9sj7yaWcuRwgYOkaVRx986xYv90zfseRoIvvgjqav6RdKojFYVhOFlIT2d/vcUav
LwBzGgpiRzk9DP/utWQt7jul59nd/OiWT1wIv7E7ViFp85o53gvTZ9hFio2/9V6C
nmTeDrspzP5m6jNLUGZmE24PnrLcF7vhFdvsBRwQZ1APIlBt+mmXjKwlbj5kx3S6
xyP3hwTYMc70yDomdM8ygWwQpsj+B+y7vuolLxdY15Cke0hHBMojByN02WovADg/
HUbPNM+TNQP0PzPnPgBzlFThHCkF8B5ihkfEbnGkTB6LVFYEmRwMCOjF2AuDHsrn
kL8WGla4SWZFhN4pvZ4kcEBMUiM9w2TERVecJ9fM72CGS3kcRftjIJVczoDh+XBJ
BWdFldGPRBxsrJM5o6wN0Y2HEdkNXrBlK86YMXekjtaybap38LFXr/Ra0fc/hUhL
mE/m+Fm0Po/akQbybXxP/EuEw42wOGrV7YHozYSB9mr/RgsyraSDpiONEY6NevKf
HsW+4Rao/YjrYbu+3+Jjh7ajIGGRNTs2R6Qxo2O2GbOYIRFpiU05X9lNs13LFDMW
DxwQB7+NoZUV5L2jeRXonLUrI38Efg64pAAAsU0R3fWeAh2WB3Gb+ic0LhaQYRly
kIudczOkWNjiTetokZXODZjqSijkp8UTjX6zzZOWKhhR8ZcddNui8Gt81WqPZqHs
J4FK95PklAsn8YPmQHpPLZ5L4W7GEv6fwlPxaGw8dgA5esSHWK0SOFtPP70zpRtU
Ir/NXQdXGNBsuGn9eQ+6povNCviB2yKfaTRBp/xmy0wcJ3168WVUWp+0ebhZOH9z
tPxG9QYuQ7ncmyVr+TvMox2szUQqigMe57EVfCg2efwa+tips+v1zMdNDOhvX5gw
Q1Rb+w+AvRTq9CZpGPQse14GlWLiBieXSEKOlxVp9xyxwLpToalGD58oIyZkwFx/
wYcKzDwUdc9fzEq+JhXUcj2BgwnIxWM2ds+Ym23u7uyyjejqn5C2sFUX1W9Jlr80
BewIvbHmm7PPh3Ggm87kH7TPGGT7dkynWVVFp76XKLYFnWozXCXAJUR1fVFe8Nty
TgPYemlaJY7BzY+xQ6MYI99VE4YVjVAaZdjkRCm+fiF7PGGAb0flXUT5kKvJat2s
6gATaPkHmLu9NHOiE2jLZhVysTMaZvDjtxp2T8VYgdt+cHfKUT/vNRIOnAwxguif
isjab3CuIGbYjSmthaRTpqhM1KCqwrelDXz1zZzd2wG3ukZLxWG5e+JPKq6obf/d
ymFSmi+ppYa9V+ihI7hvroBm+1h3pOIWiT/SXv1NUIxCmXgEkMj4bem7o2K0+i21
doouhUmDKfGXvYZ0p6STAa9TxBIsWZQ5om6QRsw4un1g2rU5hd3uWp4khca4fbra
8T0JcVEcp//U2XJ/fn1FalJzysEUvUYuGK8XD390Q6fsklo1+IJGIVmj7vmNQJ2a
wVEPQ31bIQKd4g53V/Bae0Rqy6yRt4o9PEiVUVDwEj3DeIFBLlbI0/Tddq78FdUe
h47xQRapPfxG8MhVK3RKc2yJVN4aoH+M1BIMXSH2csqSC35dJnA+Bc0PyW7QxiRx
tol8Ydd4Uj2+e9Luk0KHVk9LAbI9KSjJGLy9SpefweJu7RTcmlS/BhFEppK8zstm
cem4mf02FlcYPsGCQ69Jig0A9kOMr1xbHB+0QaNMO4xfDaEOoBeP7sTTzIUEeiUi
Y10jl5FrcDSizDH4Vb2RWe2AXtg3ahqXNx2NRyu9wV7IYLy8aYRfroS0nnmDzXUB
OJDZSg0EkNA37CgpA/Ilrx+uNnoHEs0i3srcM26+WiWFT6FpojzRldeJqhBETuNA
hVPAo7CTfvMVMzjFO9QylvwSODG92tVU8GU3hp+oJeIA6jhJmXgancjwrVzI53Wj
ZB/1Vg7DHhxJ2MPd/G0bYTHE+BM9eJHaJl4vBdDBsggogmur7TWOraBAXEaiwjjs
3yai2sdGhGu8lOKiPD2sPAat381/tI9bg3oDy2tcjY5PIbEr8Dc2UFXisO41lxF5
1GTLsPKsTZkElCnIRPiSfdRhBn6fDLsUuxSN0mpIkmfNmRX7eYVu03x11ZZlDvLs
ukqnlx+egAVRhJCSuIfr0mJ05E4/dwAYrFstEnpNG3NzPkPv9rpYsjBJPJx2eztn
71BxnD/gLyxcgoLluuUvrcHbUkc9gLK9EedA/rmW53Ww3QqDurBI1d5kYWk13cMW
SqNr4hPkZ5D0+QbA8w7gTDgQkHiDHbvvbfndOlt6LXP+TBRmgxiB62s37yvnMgAw
4BtUmBWlc2GZmUXsYWQU7CD8gC3/u50yythywGFisn8ES6QdRZ9lpYZVhCylwsKm
y2wHkaLwLV5H1JVaLgeOsaB+EF1mdzVyNecRPjB1zFG4GpFUmC9IJhJYjkwiteEa
9gf6DdKzXfJDXTdcT8DkJN81BwlDxnID91afHFiVTNc9RoOcjqGSb/VFgfeotV6N
WQ9UBV1eYZogvvWnmh/Jbw+8bqXo+X58HcyKwXSAQZqrg9PP7L1EAcXx5Tc4//gD
Q+9fM4wtme+sMnCe7EDSTBVSxr3oB9TZLymn1ITQf+MqZK8PNY71QjOp6lAZzr6K
rDZQ2cpQWaWZ/9iQDvdzoG6GPeIXDV2cRKEIl6KLRdXH2SKulrtmEzWPnKG0H0Uy
LBKHnGBgyRGddnLETY1ZN3ZvcCPfY5PyopmMmKR/JEjMo1KkXaFKjEJs/DnIL4dD
K+a5dKjDQI2A+kh39byac/UlwiB7OVBskXsvZ22B8XI1Tl05X6l9O7C1F3pvfp6f
7x6+f0J+jfIb3Uindxt8KI6KNYCw0WQYiqbcROJZFrUeo98wh8wDotAVsztDXMYz
6n7nhhD3rW8OBOeSkBCT7xZJpeJt+f2vaUE4FWHaHqVRIjRZCk/A/F96HpLUAukL
Hn7ymMJQERLSFxLISYJfGbXzx67xeW9xn3OqJuzyoZzTrWxViNJGCcUP1VQkQtpy
rPNZMK62duv6Y5UegI68B5SWh8e2BKt/FVA5UOWaNjtS8DmwBD04PglMbvXizVId
C5GDUgZgHyjgGQ0tJOA8SkhqSDgasVkGBrcaE72am5e/XaJZ07oYwhcfAjM9WjEo
YXg+4wmdD15cutMWyt7vJiXEbkyh1y0o3+K4iJd3VvhpQ9TBcfBUMfVUoEEly+Xi
A1kJt2YWigThWFsPgp2i6cBR4DGsOp2q6Qjj1iLy3ckYd0NwB7Rs3Rl4pHlVEeTN
6jseoAV+C5XPYllI2z4UbUlqD2xhJLJVi8ro/AfCNWaUp3CW+M5E7pjX+d8SeT29
sYPeZRtw28PV5XGaO6iSgFeHSN73eHjiTzb5GBU8FdPvjAJM1KztK4e8uY89fm9G
AykVXwPiIj0yL5Dws7tDleQxAk9oqA57FYUdRY9r9ADqi7ulhdz2H0B6yz1t8zdI
ns0qDSTpikYNVlhM+nhaLmGryGrO7BQVTOItfAvW1FM0gztYygA/G48f+VKeyjWY
+d9/8RBtlwiRJykC6TYmkj2UI5BSHQNQd7DrI8aaj8W2Fgif30IT7I5t6pKmKXe6
eilkVyzRSiHvMzdkgcSoCot67uaUILFDN2H/TdjFqzWCGS1RtxrHl4B5l3ZVAO/B
4UJ7MX6EcID+0GrBN6quSk9ldK64rcnX3QvI7Y8ua5LuaEIs8Bv33hd2tRKHF7LN
dMhafJk9RoIDjAmfKonxyECGaoYb5ylDo+U3GLboXSThtYPWYHnAK82le77JKvdG
5nLhH/+q1I5TrN5Y3YvCuPCLBw+vAtuuhJly6+Myqmspbr2ofRaJYCeVpQggURKl
7wx60tCh4M1fU5yYSQqrIKG5NsnLp9MP/yLq7I6A/xFgkszrW5jTR1q/+K/TtTMQ
E2ujJ9DctLK+Tus/aT5ieFcp8DPGsll+izIqi+rPvyFUtPJja2DqG67esb85yytO
cnry3TB03ncMNN58BlZJCjQQJ/FBF9h6F1cm4eHwAbeCeTdlUpp7bAGepKSX9Rgp
QVALHfto/9rbsGe8NWwBKmCav+GiEvgaRY8p0ToMc9dYWnx9V500CScsDvnMljAc
oPkJPc9J1C0kTU++DQP1pMQl3nVBzQGvpAkAnK6Xgr2u6FlQ3eczlfudGZ8xVxER
X0wgO+UOGE78I7leeFqm+p10uiLDf3yWG25Vo3OMtR+qV19hWplCLKQWzbmuh5Fc
i8NnBjztw4nupSVME7lEsOuUWxaXyG+bsI7ENKHSrqxz/lftPG9o2GNGHsxAwZAn
KeTh4S3EO1x3j7uwfsjcvPfEpocXc9ashDSWUhdb2sDwAR+li1Nc/TgqF3mo2j7E
jJUEo13jHKS/ZHwRoSKuqkEgGyK398BKCxHVo0GeIAxDLshY2rRd+3+OV8cVDK0H
zfnd+DVXyyVV9Y3Qk+pfhFlN6A7ZMb4sgUex20WqtPz1VVm1TeDoAhGuglXcdSNn
XRtqUPN7y0HNlykNsMv52RFTzELsLL9rmjJYckh151tq7DPSYKyUgSKrvhSwjDr6
i6WSS9O7UjDsEXRf7qT29Uxq/PtfiNVIFssSfPZ/odsMWofZM8r41nPCktz6jkMP
cwbdxLm1veWLIYRPUUuLp5o0hHyK5nWkWCQkt1hq35+62s0xCqXCY8mf2NlUoy/g
qONamsw+So9n0HHm16XCR2RbXcQCvckTn9xE6hGzPy+z1b3ik/8+JG2/Pnpgqov/
wIgZVgskpyrR+emqtkqBTi5uci9A94pxBLj31arAs7mpsXmUzNx3yxONy9Ah5hDd
7ZBCd3vXmdgwW0eViel4sdpruEqz/cttiQAVcv4nmHEGf3YYuFWc9ePwUsQMUsGc
shXEYmsIbevqLlQWujQX+osVjXFXxjGINsu5i087q23K/8urOExCqW+Z4vZaP+ND
vZ62ueMreKC+sDslvZaVcr7eazRx81VkgjIml0+JbQ4GfvpQBrUCKFYYiUzWStDt
fk5isr9TXrMgkNCM6vU9WxNEsz5X05AKQthVZmlvLBtoQIStOgKTC3fRjshOWEmn
n9/CZunnkg+GK9pJxolHhAK+7Fw/osJIxt2cKh+ZI+3AS/6MiooL6+xHHGryQnFX
7ttl/UWH1U5JV06g/obPyWtt7kP1+opdwyQLYwJnTvWQV++AUVTCSEWWpXrcW7p2
6i/HC4N6nqDYiVh8MXtZNAovFPfR2ZHPHZWYPHO4eleRKJad8PypXnKjcV+inHPi
CaZg4OcTSesdzSAt8jXzCsmrfF4aoA54jjbc16KDVl3iWDiDrble007/Q3svac01
lC5+9NaaAET9ejajvhArdZBufskLSFRg68WcTF8uVerlzVvu2QubF4QV6P073Tg7
HBoImrQcP/gNttjE/RKJBzQv0iSGekcnoXp5zgdNFqQSSMy07FtQQrBldFGBwFC6
DZu0pfP2VsC4Y1CQsprAt4a1Kjmik/Kzsf1wiTbWMsxp7rfJDon2QJCoRvuwYbUK
ujTL3SsSo7RjcJJzqsOfcNE7QOHBYzYX9t8+OsLmwe3WUd7h/wolN+54wH6xnwz2
qRARtyL9wA+RY7bJoOBPdHiUhQxawjT+P1M4BSpOIPVs7/JEYaUFcZavD5BCuKls
bez37lWlbcsXhGRKfEG8Xi+KaSIMMdJagcrZnJYOfUE7/iJNnCF5BcLNYfNKcTvy
Ec85qRl9ZofqBajvy1cJ09pI+OGoVKsZ/rly6H9rtVk1W08+PST5kjvyBxs8O2vU
xMhQ17/yiGtDb5B6DSoZ5nGiaNZ+XIXSI4rTXaLXzfqf0CWh5TDKlanaZCa5gc8E
zYY6UPhx9LuTbywYKUS4EeFCZLQiBfF+jilCruNrNd4hvtQFdN3/YtImILsDS1Wi
Jj5kHBjGBjIF/p6rGtHR2oDw67yX8De9uR3TG7G9AMMk3R02i3f/aC+7bFoMR/B3
PIqO5HR1pcyQXwwED1KnpJE+63SnmjVL0Mc1d7W7KvEgm49XBEZGDr8fL8CejQAr
aL5EzAD0UKMSyiYty/pFf6OZ/dgk0PGXXCVffkKTkp3yoUuBvKyOe2MCJfw1CycR
EtEIRXmj68BcaF2IZwkR2MauN5NZYAlgpeK7Rl1t6sikGO26ZE/b4T1H1DUqz8P4
wK6Hstsgdf9CdyKNH1j3OPqT+g85PIcwcL/xEc3WDCrqS2oFIjqQmPgm/YytxilW
+2ZKNatMMso1D/eGaFXfAqkGba25a9XKVhL0W98kazlL++Zd+ARtCedT9EuXbUXp
dOYqERgcbPX1EwEbAObjPiiaslluDbRnVMP/eYjrtDMkHNvQ00C1mE3kVFIaggPC
vUz0CPnpuZRJZYq4eTuqPwSPN4XEcuWzeymOFdjlu/TdezWZdgt0rdFxmioXGN1D
eZ79oHw6k2KME3iFWNSmU+jE1RHg+PaOOrFVVi6P9E2MtUGrKFQydQi/ISCD1YQq
hTtlYOIGWvIZQINIZ3Q8PaFJzFbhEmOYGPz1l3FYCd5uz3ieZhNuigHCDzkk/Wkg
vhPu4+D70AHkGKOFEfoCEq4FyVUFuU9grFdwjvejqAWxrU+G0pHeriC05hhgVAMB
7TSF8/KgOkceIIcGHqDv+/KJrifPw49TfY9T2wbPcDYu+J8J2LyyDt/tL3T35Qj9
gR06YHWWMLAf854rhstZkef8ghPp2xfnvBAm/fGxJAC1Je7/okfbfWZ+cLfpyJqH
H/Ydia9QKwX7SeN3aI9YOtPNT9qWkz6GpcdCY3Wc/Zb1NMA2m2q1rNzb/cnPzV4F
Lb9nrHLTTjUsdxVy6JIqz7hCA3YSeKDQRjtAOX4SCgRIRNaZJwcun1crP5/BKLd8
beXwt0gYR8RChbysFwDFysoQ3zCLY0gguAqhx5cr/4tzhuuI9qX2X+k8jkZETEVN
B/GHA08sL3F2s0nNKlWJ3yjLIVdKx5+hWMYHfyoUdnZf6Jc+nOSGrzqe3AA94HU7
GFIhRLSAOmAIE7FbH2eiygeaik59lbAse/XN3pkqxdnq0d7vDJCpgNaJQlzVVrxS
RfBg+Hc6XDEdVsbyJCuSAr0GEysZXeuAF7d9qpag7UFws0IzUiSktRptU8eTQHaM
5Js2X4Pmgy1rhzU3ojwF2SkfxHPmoPGDtxuZB05k1IWdmjvMRkh3+XMpBvtnAEm2
V8rCTdL+Nrj6ijlEKdTLgPxXnxggx4L5AQv8ssM1ihsRMbuPZncLCr9TTEbcJRDQ
nVRlAKqyqHfJJYPx0B6PGUqQwgTyBEnPa7zm93n0Upa1HedKvPqlqhGEtLI/Kfpa
Dk+sdIYxR3VyvPoPRqOb9hkvTSKH+FC/r+jVoSBJPs0ya8D7WpJ33xQCmHpD7emv
a6u+f+86qG1hGlrDWCichJTJ/MZE9eBpOR+tirT4CsHF0Cc/4bGlhmpt9gA0xe10
/xwVwh3u9/p/HltmkJm1YVRfPo4yUoljVgppLVmJYysJRcdYKwG31jGVeVt4+s1P
WjOm+fNH5TaufNWFUwswxWjNBrpXjEmixSSHD0U3SaoQ6lIpUzY8qJ0Np0o+hWTk
+PJl4eFxdQQz2dxXOiPc4v4kNAUexrXTnFUyulti3UzZqqraFQHaOj5Cc7Rc+8mL
Em/q1sD2ugyL+MvxAXlLweHCJE3zZNIF7RqarATe243ec8r90Syii6JXLyMTnN6x
wSIvkmQ8gTFzWoiVPQZkYZQMjUL3NuqimFXKdvOx6jxpz4KOu3KGbNriSoobRYEA
f1wF4agSEtJqQJwmX6jo15u36v1GvYvdCk4/G5+lGl1cuPl5gbfWTyOtoR1zdIye
YIW/WnClXsmTuEg6+HZa47w8xNkQCCgF074cSwBauagXHbfVA+1cL6GhUvKLG2cz
2Fy92zLK7KCXtry2wg5YFMf3lPKEFO6Bn5e5kGk7TOOY3Sg7ch0EpjAZxIxjGitD
gHWSkJIZJw2SpQxiB6MM2bJ4aolqJUABWIF0IwucGlySEB2c5JlUAHPB8yPzUJLQ
jg4AJNd5GQMgLrOHkS1zpStAEZb5BmwDWw9orcWWkyxX2y03dCRoX3M0vGpDlpDZ
Arm2SLN+sPl/O2VB068vc4I8ze0S8VIKn3Mz4x2hQIlPwfqWlAhaQZllRS9EnlmC
3lVeQCyq3/n5uFlFMCAIZ20MeoQaE9lz+SQwMAogBSK3lDupZVRsxpNbOigZ4Cjv
Kj3zpNKKesoxxcdTxtDZliqwyr58DIP4cJ+CnM/u3iy2GtAiYgLi2if8SUgewKAv
5oLArUjh5zdt6OSLOWgxwhFiViaQbbDXOzcDPH+PJKIH/8BqycVWDuslh8pmSVZq
RH2f35nEEepbW22EYpb0W+4kMuoHGhqswwxqzX0aeMoKkZWIWtMhhjUCa4xEVDkU
7DldSoMyyZejxqLSrpgXqGSwkvfOUlHMP2OxI9wgg5BIRKM363qY0WwGBFS4Nath
Oq8pYUlO1wmnrZakYp34qbVHRuoUn9FJsQehO3wuzzplE8buf6/1RWUUm5fhGFks
Co2X4jaJWROjl35af03+3BvML3c05Ml1vgwY6WOM+GuBXRy0kmJTzvCj3TuISdUg
PpP7v6pmHU/RRc676s0VynTiMtleNY0c4UfxWgAItTc0Xw6bEUK6YbfwDl2syjjK
j1TcDqdphkj5siBWUnRV9ZkGHf+4ItXHM7Ki5zskThLZtqDajXguIadiXnIn5OHh
0ctjQZUF/aWzxrY/hL815WQ6aXkEBfLJtHFNhbB9DgLfsbEl7xWOqeGkjMz8pMsP
rFPXKEA/tVOm95V3ioszy4FQL5Lc7grUtMz24tAPKnHg6NExEz+BRmJr7cp2iYR3
GdTry5jCQ5T3byCo70LzhPyqmkvF3HoYDClDM9oSYEqrZmd42iSORMof9th4DsTr
2VqD6e6JEr/fGEkFuk5UnXWJUxgrjAve/FzZnfBJE0GIhzxN24/VziOmk+aWrplu
vN1U8O5RmmUenlSKYtCILnomK/IXUnu7vtAN3ize2X+fEK461UI3M+I0Cgt0neP1
IsFtOb74U/ulv8U9F7iaKUv0r3NYt06v0uTy03jv/3vyV7Wd/yjyZWbVUGFmDb8k
99965g/X9PFdQofB+Y1Dp2DRgzToaqXitm3AVRRtJLc2+4VmVISeLICSGqs9PmXk
K3Xri1Nyap73dHuzY5Ud48gsq6GLR4EuVwBmzc1sxpmEtnqJ6OgW5Fk3GcnxJGqU
sbZ1gBCe/OP1oK9pRy5pwvHW+jE0tWIOVeLSrJ/SbVjGq6kaDDYG3iAyJ/O56V+u
x/AQR6sBwegF1/B//l7++FYE+zCxNI/5piK4fnNgKip/lZy00CrBKGAWOPiHlcCa
lDGnS/57CG+ye9WTXtlJtWm7KI93B1liDAwTw+675SkdVQPg30PXGmEi5ST+QjnA
02qkKpHEanfzd7eAZz1XrzMTu1RfnpvBw4g1Ki9JoPa0azlyXSMMpWfWf8EwN4Nb
k67E3w0a+7tS1TUG76YmxXXbfpTR691PN3YYLuomrgpQjTStI1vOp9pVp9u441Hu
Vr013miZ8lqtS/s04fkaRhIUQcgJCdN8fNj8WEv8lDcxUEsI5gMJLSNUL9ZcmbVH
6mbhHo6lMLIJfsR5wsSycXadgr+KDWbLqtJLLvKJROi8NS1SDPOSQ/JGh37auw9E
FNVjQ+SjthCsjJDDiheRIaRZDUgz1OfQYVY/T2VDwV8NhkcFV/ZIhhKEB3YpJ4y7
+J9O8btLML8sFsCm0PQlfCtdfzpKaFtkxyqQy0htcRpJlLaBCKUCQBIAoqRasThU
oXj4MGW4PxuYJp3/6vYQMiPqaXzNYdg5cGj6jFlhjcfB9o+lS3F17sv5bA7uBmVj
luU/anGiAhl+nZndRap9eGMHOcyugvnpqu957kpUwMw74/Wb16/fwbs1035j4QMw
elVSlzLnPZDo/vUOiFhp8+tTtz4A7qOAZLVPAnHCKBKt8gFeph2kA8AWFQf8XuLQ
I3zN6Pf+8+NWz/tyY9HvvNZ30rlycxNy56ayUqf6y8873COZKDE0tCBUCUtltS9y
5jPV34s1g8hWiT+seFgXhG0DiWqY1pt9dFsTFSVUihN988BTHqXVQZtb+v8v0O5u
lGa7N6AADh/8BNju4kOOBo+JCTVSGvEDKdgJ/w7Kfs9n0QH6CmrEu2AJ1wDji40P
L43QmbJP5jot521BPJgJof8gCbGDuzxrMDe8CNCEwEZlmbMvKL0RSpM02Nbs9ZHf
QNGSqotPe2JWi6ns020ra9d2nVNGrtbkVOtNqG/Tbi6bLGzU2oNo0UBGp9BBoxgz
zkuVRseHfyWvsdxHGcaXKXMHE2nZgfNz4i6SZfUDGH/uq9uwZtvx3sTWZEIRnbMT
SWH5jwObEtdoay4JswjIOu5P1ZieonvRNjyqRRYE0yp+Pwmc54h05LSUGMDs592V
oroyFxZ8fxhtKo3JJ3oTxJeKq6EqkOHGm2paSzWDsZwkL/kE06kzIBWAm3Ut2jmM
B9yjjAEbaRRVIiZkFiFSSe+thML/OsGa7jdl7vjEXW7JG82rLuyiAtjuZISreazf
Uv2dyefBpOkqx016YRO1qtjPRrMntWOsLjiNrP3p+x3jCde6i/xHyjIpCnxn1Sf7
heFcgu2ILuqhNY5ndUyBJ0vEwhvm2s6CRC4gdChnYfUwnrwzudTFINR/16BFlBW+
oj2R7nj58NkP5125HUqlaZBuYTbIHHdRWxPMsiMAjJMuMPpsqFfQRu1WGYXiNTNr
DqqgL4oSRz+yhasqO+F/wrz3T77SFP/lsgtG3rbI8ZEVRppCETYjMKMAx0qc4JLl
uyYBpEpoZvmXP1RWGoJULKktPY/A2wV6yC14cLwEJ4T7aSl7/CbS9u6OJNv+0ZRK
Hp9/bpBEi55ZbgWo+JjrEC7kVROx8Nvb7OM19NmdvNGRKZnxU1a9TpMYm6IGtOyh
I517vm0f4zZ9SIlkTvStHIDC1d4z7fWW8CgCFyrPWzZzpvG2ErVlyfvTw0DHMwiL
s9klQi2Rypj1Ba7wm9pjrDjCtwoXyNne4ZxG2Pr9Xn0nTC7ZGEOje2AJNSh3b5fj
TE82RmO1UBrf0gtxgYyUN1nfFhBPxo/WN86n2kRbwqxZCj234RBI599Dw+KE3h3D
oerB58RaSnIM1HuoiEVQj5t5dUz6OZrfFNx+C+N5k7Gvy7FCk9KQ1NJ3AXKsPtKs
Ln2SzrKfyqEFdVIdBTajVDvOTepYfxC/IIB2KCiKdmpBh0J9N+Z2b4+mI98pDAkg
q5lSoLzhOapJzBQHDgBVtp995nxpQF34sfrp346zBrBIa8i++ci68R5XWXHP4x2x
SUtneOfU6qX6Q8Cmql8R6uKP5TpV5Lg9FKifCObBaOBuuOyM/NIFCYdrpDo/IeaK
Rv7mYSAlAZKmT5HpxNBRJsmlYtK0iFuDykHxV3lwdW9xNGQUQ8Y0BUZ/BL+tFtpI
EFTBTSwUVDAbMUyElqiJeECiyZPniU1avkaQHkdkuXJtlrNX7mxB9Hr6KWWWzQHz
fXdm818x+It23Jazxv7is8cE/C1G4Le7YdFUltLasipp8/qvBDBhNKgqGKdQtjnn
QtNyapLLviORdEVz6nPa1fHEBlcugiRCQ7ZiXJdEW092P16dQYqN2apwF2I4Mmjg
vuqM2kAhl4QliW6sXkv4kImkKgoprMc+URlV5EMVym4Ibw6Opzj85yN+X0jYPS3O
c0fkdUvTP29eedz6cm9GgZ0j/tZwQBrimKQUuItW8OUahkLsVax85Hd9++bHpA10
G2OMDB0FUZ+P2XqALYpzs8050d3pjc/p3bfftGTqiUEhD7WX3/bH+nG9n6onG3Tr
i6DJtE44L4/gu+DpFvS65kNzER4L7UpbcSorUkFLHgO5aY7LqQ0pCcP0tkPfhPoJ
2StnXHCW0gMiSJkBuai051x8SYC9OBuAhvOysdMj3TjK5o6NbIqt39iSy4SbQKtk
zxbEOsdFlDQ3f9dJRdjGVWI2IeTFC1PkMLkc9CkFXPTt1itf9ZN9wH/QO+Xmo4R7
fWNyjnA4YSZomVe31cRv7KI07wkqMV10sT5SQ47mabYy5UDk+79rU1lt63RkNOiM
don4bkh1t0+zTRxsgX4QqbNzXP12ImMqEsv6xFsYbDQ3JK0aEuJEaDbXGN1LtdGW
+Ik5QHm+4hjZeKOSUm/iLKwUxP5i9qVs+iZEOpVpFxsqVbLRah5NVAQ6qHOnSUrI
Xh63VNymh05r4bLfJZ9jFMGdsjky/W9/OBH6HV4cI8ac9OIiHtWvQbwmzotgNjT2
K+4+Mk+1wBI1i4LZoo9KBxGsQdZTZkMnbT2v3ekxvw+866NY0uxEIbGbXezWidtt
TiRmUh/CCcb2qff6EYsFayPJPF+3Lr7wpgvOzLrzpLeMdCAayVtHERIeb1fLQeAn
hjzueuKpynzXf4T0nf5Lsp0joGAZWWARX+3UbGroChGYoepMGStV+W/L5afhayHp
jqMSuV0gpqURls1TK75mZVrMrLJR3KoehNrXjr6AWDfoTva0vzCUN3KaFGK8Wi3b
sv3nEzF3WcfAr5n6x1IitZBBs6D3YDo5vHpOGiN/ChmD/dZv7igFz/zTFZE5f5Gg
qKhOJbNbMkefDpJE8aDt2J3JwVU9ZQ2+i/B9d8yHilPNZoUBb6cxhckSCVtzl/eR
AYjnrZMu9iin6LTepAGS/rHTazPb36qhN8xcmEUuosBtXDhcNj4LuRHLggSmRgsS
p9xyfOp0w6mXaPFCHNUo6k1BOOxUwLh9gsWJKsz7wKlHcnPqXwLw1fmNki1/sZpw
Kqd9kZQt5tEBKkJAW9NxUZgXjJg4+BprDEoAVsQzrH8n6Pdv+S+gZcWMHRDDlSah
xxWvInlF8Mlgb4V4z9zHKnCK9RiiKx+t6Unvc7mG4+A0g6VpFRXzuRgCWAbXrnYu
/R7UFnyYIPZfhSsM7E4E1O4X/3ioc0sr6uinAJmYu1/Loj7kaJWljDbLMVmlbXzz
M7ZaWkosH7+cvgV8Krcvtxj/sdaPFMTWW5F8hLltfA/TnU9J0B+P5/RSvRJvvOF+
USxuEwN1SXYq0elxYNirrlCFkS6g8wzfcfaYhbKra/szM5dqveIAduUyW9uXyR+P
RScWK6jWlT/4GkObNpdllNx6Hhr30Ss0etkftT5S4ctUTv/CbdvlPiLxNXu6dfcz
rGMJqB6sKtbgQLElo4f7Zy8qz2TsPJPVEZNei7FfmTFYCPw+GV+j+G/7OqqFtgCV
xx5xhmj/pxImWu9FOvO3aiT1lTBq+jcIKDXRH/6x+VWAUk4oNvbE+UPb+c+19lzj
raFDWROf17jNxdVmscyWTYvgKtVakEHLWx/Hw/OpxAkp1VNTq3WF79fa707sHVBE
Z1OjajYjdepmRcoCLsdMRWcEivWgwSMRsbYQw+07sZ3rDJCgU/jfFUOY7gCm3qY4
/6leBw9Jk2EkXCiQe4aX8vwEG1eUAan2dwGjcyMsluR/jJuuY9P+EGhURjvt/DjQ
z3r/VYkMToioCADttMlsJRZ+2GQTdv7K4xijYiilffcd26qZ78kJOgIGPRYUGuPx
vpVxl8mbnk+Uxs0+ijuh6QG0wOzGXHlu3dT5MXdC2hdYpTbcixxFzJfqWF+l9YAT
V+4lg4vUe8bvVXSwiXKodXM6unAsp/mw8B9I3SVQ9mhFoRUHhX/45zE7LgYs8YNW
4UD2X/S0QZii2Wpspaa7VSXcprattgG2Ku4ftpaZsL9UO6/yMp7BZBEldS4naB3K
wINIvAoTH13xOFxe4MEA0+nOQwyx/KhKHnkDtGWQa8/n7CYkdruFxdFXNHItM7Ws
vV5kRn2SWB6nAqQZFx/4V2BJydtphRJTh1sdo6vCYSHrGWz3jO5/npCQWCuB3Iap
D9DRGFwE5yJw9M2wolVd3ihwWsn/z0FsvhtWm7aa/jciZ8jfACUhNlDgdFoO8ujz
v7ju3z/xVCgExVA1ujpWcd4KLgbQGoaWH+lcbxRGf8fV0gaII4K3aIsSTY1jPuNT
cgSDv0m7zsdjIxTcOuN4Rk/yr63H1MA8rIhUEdfNQyTsGmWxOTV3850Z6f4lnvU6
mz4u5ZAVBo0oXVUH0hX6tKe+OHzr+PRvS6CMBQ5ONyf4bpWS7hvvC0q5C7zUtQaF
P570vZbSoFpadPKaRH+bPQnMv9oAikHNUkGCX1ZOBbUDUe1b++LLH8Mi9+Pcg49A
Cs1+ZFLvqzl4DZqa6RA70YBbbIXIDfki81FNhMZyfL+D8az6sh09Py5Y//XHE36H
vTUCQaHuNeDbF6wvijF71lsouUK584C+J2445ECMQ7eoEirXqhxlpQdUMJKBGmno
x/0BCT8uQ8Eg/coZ0s61IBxVBUU+hioQGqqxuJCM5IuLlWQidnqhgpIMl2nx5f+H
Ugqx1ZAHyunoSOuO/cPY4RixyIbD5MNpqIPk/fgkD8cMo9guWbpaaHvVrOOws5ld
nBJN44IdveMg8So+ClWRfoonynpFw6u5KFU8Y0TY04uwWrFWoqZafPESaYJP16rM
LJrZwcoWeeY2RtHOETwAbrb3CxIK2zmU7+Nxczsyil9B50yCk1+MEaWg6DCcPJyP
b3JOtmaIV5FhZk7iN2taEV7UjjRWVnoiwAfy373cCItyFxhP35dmqquuBMhU6GGJ
8LsUOtfGDjww87tbVWnGoD/lEhvplmqW6QYjXQv3B38vEAMyrLzCv4+gIbt5AJQP
QxYpe7y+VhVDzbce0JFKVUoYOD8/SNsiqCD8dwQ517Ekuoc6hLtL4kXy06hc69q6
CghOUATTKxDvFaFxUjQyZx9rcb7vu/pKxINBaTg4YCJ+oNjrRMigiywvIDgSDG4Y
2X0zCHR2Z50QteSm+A1qIIBqoe+TndBYPD5GYaYKZBFMPHksJKBb/LjcCsSitLc/
fuwLQpHSG2NBbO63M07IRz86TJ1cQH7wwAHpaMsVMGVeTbu70s5VbQolsc592P3f
X2cnop1sKCc7g2+8odItnL2Zd4uGBVxZ0inIDD+vexFuHHj/1mP7Fxr/faRtwwoY
GGdpmCE+IzHBtjztKzmC4xSdkW7LvkG0TTs3K8BpQckbejKnofQzZ5Np8VvpffV0
Bf2paZw1/0/Q9mH8Fh4wSrpgHwkHh8pRKxBZpPSkK4phtgh/YJ8TuV/NB+nbrz6K
Rn2qRvLItFhM93zgZpn64ABZMioD/1fij9oLLV6ZuG9+F52dMiudat0yDjxJ72wl
RyJSiXRQL+A1V8Oiu0LQAZQjQvRSElaG0B65xB4YvIqY3SPIQOkgwPOY6ryEtGwM
NJLOoO6pksXQ+gcpKrfJGxRon99cdvEx6/TmBNXDWo0rwX+ubKxmO8VjAvjAMtoX
ezXE33j+Pw2U9afUC8cnhWygL2+AlzFhwofde7rUp0KfEtvmMvq6pB8KG4RjgtdF
bUm8/2tbNn1egRwoxrEekSHgZalPGbpcSuIQSAKuLL6AM7MVAh2dGcSZY5MwwWrt
z6dRKJDDx6geuYojX64qTNNuNBjC7SXqlzF3t57zhRXDoJeiNhWPl7cWkt9hnrF+
VnUK4WrcqF2SnPjvR/+65x4bzt32+KCUZNbp2uf5XRyJFFjMW4gXJgKqwv3Hl6p5
X+DKVQqT+988wAcykBbgp6VXXsdlVp/e9x1hFtkkBt6l0hn2MDSerbGDHZ/bJGZJ
i8un3qiXSi72YZ/o2fPsvj8TE6D45CDZrnsvNEqFmwjL6jqrdn8ZmvRZ/S70P2oE
89nB5beF86HJAJtP1aj572ReemU5UmXYTviaUnT5sy241uJKVu1NFXFgKdwDdk7S
eAwRn2gvuJFV+bdcjUNCsGGKy414cjeDk7gWfJdkX3vyhniPPRePhJLoX1r11jV3
E8Q9fl2DnzWKUzlZZQNkWKCI9cXnhgLydsV47Q6f3ADOXJgRuGdoepQTDyAm5d5I
toN3vH5Z5SNCK6dFbiZtb4DG3/1NcSoH/zOcmqy0y4OevmHr521gjKm1d3Zu3Nks
WTQTNwC4UNeaxCj0bx6H+cSD559rpBh/0Xn+7UuIBvWX5R/tfERASCz1NJqTAf/9
NqGCoo3kQdLKX+zL+bnx/0ssTV1fRnEp2SToYbw3NtFqjY5wj7rGyiMS9S0gOjbk
ylmQzVUrTyfZdrzc//R2vN+igLjWzUbLx+IQNUc8op+rygvOIrdtMKImSnLQkloN
Kz+T7k3T9ZwI17sStOrLbFKIGbERUfL5WRE23mCq/Z8C8OfmUh+w1mS00iY8pTrp
cnpqS/WCQLABWDCHDFHWuYuNStueo4a53A0iTjszfzH9B4NTEJCSGFcHtH7Xacg6
UDsOyfFc3EXAs3/MrpgxOk3CEo/NMvXe0aiXgOraojqS0ui0fML+dzF6JA+hRTac
zItYQLaSrvaSKjYv/NGjcyK5MBmuKW7ofHcw31SM5d8ONhhxvNzFeUjJKMKanzlW
gWvyi58zGOYjtOsBJ8xWsDdan5JHxLfGXzRdFBLHaCQ+lJiTCe8WX9lI6DreIf9+
hAfYBQNQCCGc6ePD5XH16nsLFLd0ela37nTM7oWYQykIFZ7C69ap5kc5GoQaE/hv
q2VbCiiHHClygyS7TLMu1IgkP0Eg1/81qkjC8t/4qhkAHpLZR63aB7DjCRpmVHYa
NAaPMDwOiGnZMFuMoqaFzm8/ddlMLYKhoynYBKMb3sWgGsLaqXWZQY0rP68IQwaL
rulI/LClLc9PB27ejUF52AbvMvrTPBQmcoSxI1BolC+bKyvU5fhZ92VY3VzTLKq4
eqLtVVVMjdnSBsRwhVpfcXmaYn+/LSUQ5f/nfKUwDuyDjQ7j1l8yBG/PbjG3Di2o
aw5XWGEwM+mwPLtm9f3yatOIJEbgBPz8FlY9X6Wk5jBTWZWpCP8bnTkZ5UCB0CNV
FsSWhT5ioMAI/gsAyJlJQEEuTjxAV0c+DGh3PuVmm2xVvRMCu8LzzoniPZy4+xXu
+6JrW27W1YCBHm+r2uV4HuMpcF34uTz2t3rOHetUBT0JHduJA33/ucCjthLE0UFg
PNr/gbgZGbn972rF03nEIduWLn7nE8RKWo0vg4h2sToSXmzCpQwzmQuCl+YogjIc
F3itRxGDzLV1mmxka3eS3f2I9OCADnq8UqlwOGbdv1VrkqQh/4L/cJ4TA6l/Kqgk
8rh2UWJbBVreggu3tetQoSPk24k8oqMNDFxKIQKNyhfDLLCye4xYs5G0qxE0IRL6
6+x8VtB5V1DWhY5J24rve20zR/ImSoLgwEcMAwnxc3eXuH03bJviemTvdbovnM0/
/MvFulQ3q7gQJsbqPqVqqEm0PJJTBZlyUkjmsvIAfMCY6u5nn7/7/e9ZqkdmOuK4
qBfv7+s9DenuJPcbQaZoDLlBVCsOE/xEIrpfjIjiYPMs1LyFDYGjbPD1j99ttlH1
mQDXSOBaonVogBCzadQCHZnAwfZW3nQs6Nx7J5JbXy9XOGbEng5aoXvWl0YQ0nTZ
FCvErz/pZR7Cod5OrwhWSNt66WbeZhcLEMXvG+Wyc6jJeWF/0VrLaLiG4JymVOgX
YtnOfd0dK6MX7DVWo3IMIP/JPYlJQDmv1cF4qMMIkTc8UXFoKzUfv8077bjSPKPy
j0AVGALUJd5qJJNHetCHE4buKBmI2ruMWVZ0Ml/J39zar68i8cmbQ5LlRit6cbwX
MIO1o6Jln6WOkYaYWdwxV8r1f7k26QW22RPTYIonHIUGgRQD3cFj41ofT0kglzJ6
fTozv9Afr/wr+zqSapmDtEeZ/z0DQ0UPIYbtFApc0aWYz00H55u17j1znnpTVDpk
ukbYuF2sVHsyAUozRj7mSsgN8S9WCU0V6J04QyonV/bzrUbBMNm9Zel7nmdoNjBX
fys5PmwmIPLyKwD3Eao55BgwBIpiF4a3C3j5EOApwhmuevc1fyQGjJH+FUNXsdJJ
G8fCD4D0CMHq23Nboj8Q15aK0FZSAlpdfFyEW3LWQn6jyrwq+GJdIolQ/df0jlq9
WZ+rdRtW7mjuvqIYDxUJ4XKzP7oA47H2eYCQShVhODtF8x30lRev7nz2ZH1QhH8i
vBOriRnsAMvpJaHbQ8QbPJ4s9Bri+p+rXwtwZKK17fqKUVo42bzpOiWlpUDAdKzR
zZIGifblZjcPCfL5ePUciEFOEjopwQQ0qe5D5h76ObTNB6MTkTpS1iv9as1tdRq1
tm3Qm5o2409arBgYMDc8PgImNosKDbutBcGO2BY+WRHai5XjRvujtzV2tgssa9IX
Ld36fppRaQA7OpyMdJ6VhWv5NWsmh+5C1Z66jR1Xx19lwdCXUx/ORVlbUyu6JYVs
TQpdRuG5EWM1qQMl8rMkeGSKm24dxK7rJLkHGNXgBFD4ZZepcIy909mbVnkG3++/
8BEPM0VNRqmtINjsYlmsOkImyUYaDLQPm7tk4JisrsRDLF1Ot7WHPPEGCuVGrSpN
S/vg7GmTOEQTEdxVMA20f6RQ7tGJRgtB7K8dEzC39oaOp6ClHOkm31J0Mx26ijwb
+eykiQ/w303QKG1XaYlwzRf/QFczwq9vU2LXf660sZhGUeu1XQRgo6YDbUYY3qoB
ewqGYDW3pkupfZK1O9WS2auiWrHdUiiU6UhEk/WEAeDGCDRKV+O5May45GGU3bkk
aOJyV8cuay7JzFssM9G4ujddiPM84my/GwZTRjAEVNJ28iMXsPkpQIl9oGfibrKq
6Ptt6yarKLrBC5KHrlQGzM15I/MNqJgZ2/4kEPEHQDv73Iz38/sP8G7kF5/wpfr7
BsicO81TjBkg0Ai2XTLDrZG6Tp1Rd2dD6DgZ9/CoZjDHkgQjcw+ByB/AxBdSnX7O
6hE6fQdNxE9KCgor4HPVSuDNCpJkVAzbsuqy9Lx1btST2H1mMRIb8QQwBlU0KOr1
EwVWFdYkH/tZDzoLoij0wUKM3y9Hoa+qkqniHyflM5ImI6Z45US0m2SRz837OevY
kV9LV7w/9I8fZTX4SEvhC3ApOM/8m/oo6UOlCKqqTdKZoV+ICr1aE0KY+Y+PCZ4q
lLsIxQsTazDULN/+of7l5FzhQ7DJJNzGe8kOTCR+EOTIVZFmKbBFpwrf8x0hvAzC
6+R6wX8YW2LqqJXqPwMgL56KCwKUH1G9xOZDpzno5GrCY3B4fLzXHoIHHdJwrW4y
AlO08CkiHNngepX7iRb8+aqDix/d8QEz/Brtm3qBjSc7sj6pZ5+afWKkSkMTGhcv
KvSbfJwvxudaxCxfA6QEjZfAgiou2lWCqqPVnWLAou0KK62MXlq6uQqY4MrChOVb
GNdsZ1MMW/bo/Ko+55mDwzApRvT5qg7d0twXpvJSGFURw43cq5CUnpRmr7F1mpfK
UBhIQmqXvzCZUxp3qQJjlYnaHsjmtKZ25OVWkpOeeLPxt6BMxsncG2C+kLZZd6bA
NO70m8MjpIAY0FFMlqQ2xEFO7Eq39QUezI06dTkkVoCDmUsFAkr7XkvQjrpUuxhK
rs+1rhs2wTAIF0KlVfXvvs4w8ikwkUfcQ9neSs/tC1+BGtaRsIkl7woPbz8GymsO
rFBqJ3hXPaEGzFqCr668WL3Q0N2Sst5e/IGMAkUkKt6/xhkax3xwsSl25yPEgYqg
qNi7xrwMcgi8RgmrbG42qWeDHGJiNBkjFy+1so1b2110vVzIoObiLDT9CPb2svKD
suyLPnxNV2MdxB9wKf9dHlCDNAXInKPntZJGv5DAVdfZIDnTrU97sDJZ/XutIql7
LvuWt36irGvM5c8JKQRUvSzzFV36Cuyw1Ts7R6Y0OvvkGy7pFfnstPdjKdEdYV0l
IG53gb+IjL3xecxkHvPXDGCKvBdj9URIR6XNs2hejH2uc5gBxYlkKLZ6vW9dV8Ue
wX99Ey4Vty/dQW2cf7kVEM/SX3zv3KgrQLHU/TWohgjWz6QSSxdrH+i8vEMAn7Z9
eDVmExH/IoBp9exHBCDhejMGEOGVTzIH0SuCx350kugdN27m8+YqUniRbC9SGubG
ZyOhCDFOMDAnbsLgWqixH0T2JNRpeNCrdUEt4AEreXjoVZH4jEUEcCDTSj77mhFd
d1kuq0adbtlK9NkSdudVF3giRuLgWd8pcHhQPiQdDAqpncUlRgrbD2mYbpyEI9jq
IieFXNe30hso5L9/D6sx6SOIWKKIE5SmlBy/O/hWj5yTCZiOwgmonEqwR5VTdfp8
TbB3VWjAxEl4ZngjAhvClLam0FpZwCKMoH1bFVD7WPVedPpL8KZO1kLoUUvr8A+V
GxrwuSwqI0CRceAMPONeJvTedFNlPS0ZfVhnWhFCCOBJmITrcx+6vr9kv6SVnPW2
/AkEXr2YhpZUc5UeSUmWJAqxitHY7MnVyikPT5zjamWWCAcZraaDTQ5C2F6ru/51
NmZIg0H1N0IrClvy12EWlAdLu9C9cL3aiLSfRYSaePY4CpPnZX8kUjH0jI3Gx07D
1AnlhdkC1PMDE5MWAuUBOXL5edfiWrjHJ5wE9x4/BXfPQfxJ9VF4y5nMWrEr288h
UGHPbD3bpAPHTD6fRHjcBa52/wcLD/1bRg5Xx6ta66ZMsku5J/r5Vsm82C9/rOUb
1LqKjl9CQr3O2GlFhjlLbh+CRQlXFQGoPNOdKqOyOIDC23FUQef0L1fiHGQwz9Id
fcXr89PtYXpu9zv56o99H8T0TVOaautSpIX5M85PokTY7j4RrEdoiHSrC99HXnbK
xw9vCQu7oznQcBnkKsvRw7BjJd1uao2Mli2gW0esDNc0BQM+HQUERsiF39ouxh70
ipNxJidDmzOxTUcUkgD6nB72jOqQIxWMsQjnEtJxT4sr5iPvw2rjE1vD7oUUPX4x
m3A6Kqhqvz/tNhZZmzPFk430xkmck4+Xg3ik8F4niR/J2h7dzS8N4eC0gp7CvIka
KyckhtW+YinDiencKs+CGe4ycDKDFQVwbcpI2rzbgcamcevFOb88P1PAs4QXvuqQ
GfcAbLr2s+miI6x88SCaNFffgWpUWEQcoB13qmcre2wZZCKcNwhF+DoMvuCmO/0R
GsmWLVWuEnZwD6HMSEpTMfUoZet7C4BryIPE9p6ScnqddKHbLRRgt6q2UHpnmXUK
MnYnX/nXt4CcMOdJ+VdnuyM+YP9P9AZzU/apUC7DXBg5gGJ6BuytjSwLB3Bwukyu
d+g8kmFQdNoXPMqk3X4iOrY3O07BOjeLJ+cltDFLMR1EhqALZxPPAW3oCx8KtiTq
DefXpdvvaFfB0CyfM37k0sVWu5cXQ7XncuCsKwpYQiXM355XItIDLVoYqWq6zUaK
9aISkU1/7l0K390Rkbvp2nyilZnbCanM7Cp31TrH6fPYGSq4HdaooJjWHIhlIsNd
vDNiDG0ReaYeYKVodPHNaEo8A9/Z3+AkNcVhbIsiPsFztZrXwyvonMTAwYYHoG04
61YGT5xsKk+XeCB9lzwTllsO2uGNRrN9V4NZjPIIBIPZ4xXtgq/PFKMVtJ7gplYl
eYu4BofLpxc9JCVpZ6h189KFUbWU3fc9K4NZxIKVbOOV+CBx+mj0745/iUUwLdMZ
cFJ/DgATzumM+LtgfHu8Mn/7LZE1X1aclkzFimMvs3JxKgcXd/UerQ3pmCRpadTh
Ts0TzhW4UbLX7+/sSORyzK7mcz+lN+xUHd470zYlE3PyAhD7HkJE3xF+YGESh112
SQfYWQ9CgUZr3T5MAQId6LsgemoavlfAEIHr9TfuIgvqAMA62SGH4aq1UpYrPnt5
kchg9whOuLPMBhrLk8e2vPHGzUuyRcf6niHqHJVSIFuBHHvAIGaz6yZeZKJrtXms
gjyZYaOZiitHDWD8EFm8vtuNoj7isyftxCAEAvYMkFLAHmfkiWER+fA2QTGbdKHf
obXBf1kkuLhFvawB8ZuXEetLhCx0tSke++cqNxR6keX23uxCVUkbTKUx1LhizOR2
Z7REXidrcoVo8Z5PNhDzkT0H3NwewiNAVMRXsSSuNs6idyz8fBlEiekp0j8vS2jS
DNeH1Z4eSnkT/x1riIrCCaVXOKZZnAjef/c2zIpOHT/Lk/kyHxxbCLxtdyNyQU5V
uWKweNbnl676JQpZcIj7koqrkm7O+YmMhyQ2rpDK4RUTxz4suyxvN00VElM/W+I5
5fCS7T2kZPO3PN+JV3vFXVE51yAPTK86HPzQN7Vb7NaN5KfQ9Uq7V0263lO+hV7u
Uz+Zev7ds6IFVGFZoaJf1MtQb0S4aKQgxEmzvmy9feD3kLE5vVyxUvqEkYxLLU4t
VE1smoelrezr+4lQhjmH48yfcJ/WbJzHJXGgYUj8PH3gHJ5QaGT5tpKez1L3PmpZ
85Bsn/ZT6ztoTk49MveTCui9g1sHVXjIpftVmZoeY5FOvV51fHjOmbch/1ih9NoB
OYfCANBXBe6cEhrURfm+GJQ6nOyPE8G0WtZ2znJXDXqozAODCcwKr+EllXOExaM1
yVcJ2kKui8gF3Ybll1+R0wC6X3roXPuRO3kJ+hBMtifUN58Yr5lkk4D9NX/2/DYr
qqPoz3RIwI/SJ25za/MmQ9X4525qdrJZbBV1l/tWMWTDm5sLiWCAot5cDEE2K8z7
eR5AeVffrfdcOHqpnKDFbsIQ8rzWLPPgNoXbCeNvPQF8YPIZnEtlxh0bxx/wLnWx
U3OgMf+Hm2vFJ+trE8r+obQTP1+si3sYWN98hJ5T5JaQD0qhJK5THMoXlUlLdAeI
hUqSnuLMRLGJySVvrIzQaKJGqONpMp+SRnkpRjeUfam97QltuWI0CsPIgw4wbDHL
QoRrxvRqILPZ61ZhBNI7eHg/0hpqMN/OP+vmMi4vx1l7Z4AqJ0wN8Cdx5kvm43Zx
kcRJyudTdAl2P+H4dQ7LKPalSgxP7aFhoWt9KmqhjoZPQeoz44u3D87h1EXeh5tX
1ZT/gyi+puCg/TjRX2qcPogP2zqQFCPCbugow0QC0PGPrrHpFpENkagEbvqoaBGV
/GrzMINDjjL+t/+qriiHsI9INqmCbxWC7IAWM6vngOychbqHttdmdlUlrcJKkTIZ
T0YPD0W2eJHm+v+CU9E4yAT78z8LLN6jrSkn0uzhc1VbhQe0D6Hff+0aFkWZFM4f
YBBlo7IncRjASPSbpiJ3Lzb5W1A1Rgg1E3aMf050KvPR8X8vFMLj7TplqmJzN72x
tfiLHUqd/THm/cJhpIYC7dJZUSeALljPMsDMnJIE3QoNb9wGlRw5pNSry1jHdxRY
D3HHdKIJ6sjT8bsmSpp6jI7o+hAN1Fas1/7y9rXDtbrFp5UxyV26e5yJ6iMDUTdq
FuDjmIsGLJmUI0Gtmpu77EbipLLJJlka5z3medgZLFw9e/eOnwOC7JSEw8rEhTI7
t5hxrTCJYPIhyjl1gEK8FXbLw4atDCi0T1Gk0Oy+0VXm3SL05DMnOkk+qnktEdvm
Ulo5uK4yrMpbMSZnKkWq56eaIs/40lRGOrtT2qL4WZIGSTWKUUEPqyiJkgbfqIdS
DJOvDznnYKTWMaY5tcq8vZB1fVfuo9+KxA3wjOQ862zOWA0XBTGJ2yH9BOKGT1du
joZ8rL9jUOMfHUeHQcJ9v+rDrem5GF3otLhqjUeg4J1Dl7T9abqQn5I65Kwo36rS
TN3hAYTPFOHoBPOJrwfqO2DSh+Xlr4V785GuDevTyCbpQUcQs5akqEeA123Q5MFz
Z43nghqh2Yrq6x5VMMYsX8A9Qn6D6D0kgLR2QMg4PqqdTuhA69sLTe3BrAl6g3OB
91K3iWHO+hqHs81nZU5cXjoGFMYEQH7plgKvoHtRJcUVlw/v5bTw/sLnhOotRRIn
2cpbxUd0u37Pt45AoW2GSElaCNYhsqjqBCXxSLJmYDpvNeTHQWGbk5Fku4GH9k13
CkcMRFdfiZQvM0WvqBeDgQrGNdJ/kmSL42h7JWle8t/wyLzTLUiDoN4qKgeJBngq
4+KmcWsgyJdt2boCtqyA8gLFzxlzaRwvPxu699K0YHxlTD8t85t+tzcred2IEAFz
nVnC/6Eisn361oOacQgtoQWcqb2qchHUppH005w23iqIws0O+wMpAu1eV2I5J/JO
ab2yHDh1mxI2DhT5wLLUiqQOArrzvYhykPQTFUpwjRBpmjzxxv0bX3BDfZIJm4F+
nzaZ6fKBlnUbZaJ7P2tXLPAuqMJggPEUsQlTFbCE/xnVhMkqbeie3ZNcP3sue8UA
bmaKya3+LWai8kakuK5ac6SQq1GClDN0O0xHk0IYV3/yUmEBP9F+jUFcwk9ZUgUM
dDovk2ewyXEALS/htkD+7zpxd2UQqLmNlStMpAjVyDObpw0O5OPTzJ+cnekvsT6p
srT4jzbA1vqCEYOAPfA6zJYzrP15uaAPt7yDY6QRHS5DAamINfCzW9na26VM9t3b
TZBOjp3ei+KmCMo628ssbj2iFvC1i7gIPkrT5CI0pUGfSOMYl/IV/xcuZyleLX98
Y7J8JYIrfSpVo89v/9NLUwK04G75HfXDOZFcRDASNASHqGL/SMLcEo2fvVQeGAxq
wPVXnp4qmzVfik/jpbcSgQiiYhe1SLz0r+NNgVSItJXp7zBVOG/psWQxUFkF4anX
k4hA17mEBoG63pbW8cfvKqfyMQAD5D3wJ8IX3QL1Ju+t1WroVxWbB6h/1PhXw0Ap
apbPZMJj1EJK8PTflZLgWgKnWZWymo/i5OS82+JWEkEIwtxAaIn/nkIGC7mFlsdj
i/0kxVFeUc36vN4kvHCYcU1nKJsx8ZoJuaNG0qFGgoKCAvwykHYvJUoWrOlvc9w2
5x50/f4bWHl62cJtCNEXsjnEw/KzH7nBFWO2//c72vVHiVLLwCdBOV2ljFyAwJBM
ElizYB51KLOnnd5BZgba/zlsXRKAYWg8RfuEobBgI/8S3Qa5PtShA/uVALYo/Cai
1BXBHoiOluuJ/u0r4FN9ecmHNJZDXsakSOlrd02M9Yuk3bHGvZ51p8BlQfwzaBYJ
5Ue+R1ZFxMIER4QcHUVDkB44xTgshmn4FQjK2fMkJUisLO2ZGYp+IKj6PkIh5VxM
DCqRthAcBhIqKsigsQZMrbWfAjOTTafZpcteNLd5PW43H/QRwERsoz9x5xHoUFQ3
qgHuLgC0QOfWTNkdITR+eaQR+WBQUWJBtY7mK4uy5fH6nGpP9Me8oDHXqlsdI5Kq
yPK6MCWokEwhVI3/SvFvgssUoQWwM2aLpPqvD3BfcaeADo1GyI7c0/pMKpZjmz1i
pHW2vmEh/tcSEThe7JwS7aLkueMe1LG1SQ616W5XsKHA11J004cURZNUn8Y6MJte
NIWTC2dtGtcqSV9F/eqEZFtniDll1gsv00A+nI4QprSQJ4FRG1W377SXod8Hhljs
sjYHiN4kJFOUOCCQu2pdfumzl2vKFtuQnk9i/4o3eXCeKF+9+Pt0io098GKn9FAi
RumAKiUBrXKynfcEXu3Xm7HPbm4UwfGesto5JLL0qCBaaGfTLTytW1Lj0+x5tcXe
cSa9zktppI1eK4dKABnxFIdec33v5v5gthU6t9NkABcY2cMsnDUNKNGlsPRR9xvQ
bVkCyIxrL+Gw42+xhnZ0dRVs3pku9b+BN7MlbfMItdahA1Db96HFKGkfEiJVZzYI
J5Ip6QLRvAG99eiqz5HCp5UGAif8QUyV48U2WQwO8KI7kBCRK+jfFRRqvqfuPjsA
Hxp8Vod0ADDwC6pd6ft0tMd1Vf2dfIFktjPH9ZfJB0wJ79HX+TMP6Jx6/dD8wAxB
9k+8vRjpWPonnEh193UBYgtwRmUChbWoe5UPKYXo5nohcdbmuFsqvsfje2VdcjuE
ruX11ysoVed60nrrUdxlSxykKg/3kd+tJrcssbSPtO/YMmA9xSxWKktRJ4gP69TO
WVKE2ZtuiOMdtQXQF4t8FOsJpQozCAXOuGuHXuK85FhrK763UN0ezgLRQPS8qnxq
HKC7vvp454mGeOuH+Pzl64fV86NBsuNiO2NXUBc/CfhfC/1YKnhPxBLVcKKz1BFN
62jAPEV/ACLFkA5wx9O2m7w//YcwJSz5bwCHZOZB1y2baInMFq3fbDHDhbKez1gb
AqZX6MpfQ4F6Ut6pJxszZjEpmzuER2l43/F6UMukWa8pR3Ri1sHiQCaFfNh9PZnC
/MpeXh9XyJ2chitQImyI9l+xiq1MbwObjlnpbaTooWoaErQVHnqDYzmnqx/Zg2g9
bpvbuoVsdMJRHJ1Z4TAPIBufP4vDzI60Ffu2SlWEhRYNHOJVeqD9HLUoH3zamt0w
5+k8yc8d/pXu6M93wnMQtj8a0kg1AfSbwfUerBJmDsT/L9B/3CY3zYGWthqSwgyU
ux+fVFC20ea39P3LaSyWvb5bZt752C9FQZZbfAN2rLQm1u6zBQfxygkBlHXtuFPr
cEdySCYvj40MTNKa5mwXhohwCOkxnoOlMnzACtt8k0H0qtHceK2OiW/4vKKNvNcU
U5EcZAg6Q5gXMvqzilSriioAISRXlemZE7YcjDrhqugoLt/pQh7Kd285K2ejar/0
fu6L/MGKrcdW02zOPumzCuZ2sbx+1xFVGiWpb0blnU3qgB6ilpQYapO1WAs2N5JM
oPKWKmILSeID8DCAcfaz98kecpEoIvKtz0bNKLOLeGD/SF+BifLuLGVx4HAIw/ki
+HYjZTZAwXqwNEigEX/cZRqgClxQ0ABH+tIXhcRa+EGIPRGwT5/QDe6S8TiLnoyZ
Sv9OJq4qlo1qDxYWWPPj7LAd2O9aYtYOn2K4YOAGWyzjTPUQUSNxnD+EvBN3SOpz
4EmFg2D7YupGngpcoQLI0pA+EFQGxzeAVr2Ww3mq1eWdo6H9Q9/ChUp6z6F97UbN
XnFfEEIIpLcpLJIMOO7HAMFNiu8Ln7WpSbrKlMYh6XFu6Lixim7adVK8NvBsau6F
g/ybHvYzMmtnxRZ0wK9Yap9jLeq1ncyWpT6mns+NOh/YR7fP7wYOuquuKm+Pt3yr
tEvIEK8xLssxQmJ/J0p3Xe58i/hCe5SlR3MFt8GatXnZxeNhjzfGq6ccd/3Z+XJQ
ky2w4249W3YAHujannnaKoSEj9qLA8+yauOdk26zxKkQuccBHfZV3LDILJzBommv
PhPH9lheXdQtdvau+5lpn1HQHMAIiFGdgpn6wGR2VE35GK0wEKC7UTZCffirpGJU
5pLmlTiVwr3mksmTF3d4oC9JITV+vFF/LtJIXMP9tapDa1sDZ9ah/FKTdVMg10mO
YlSoG7gLutce90ffp/tIQdq+C4eK5Y7ImGiadJWNLa2gSSq3Pb429g+t5vwp6rTH
yIfG56Rwl2sko1Hmq0VyYw8paApGp6KRDA8YeDDBV12Ox18n1CnpBZEjhEGP+GYO
awI3ogdu4EXivO9Fp+LX3N4RYHsycfLk7RsgplS8BhRMCx+qCBGGW2otHUWRRtuf
9njMz7gBZktvcevdKgiw5cbclDfzUUBFLtv0UxJcbGrv17LfQAsBqN8OHEd5Fo72
HdbqZnZwJE5AiYW5vdpAHEfQuSoHOB+iYyy80BvNqVLCnFHdUD/BpizKXqi94bkg
6PvB+TA+/OY01YPhrH2yEoqSqSPKI4WCAhFvZfgAWXcSxRQy5BCaPPzQDdPRn1ce
UkMClgtd/agP/J1GVvAsqO0FO5HhERF/ze5dMIQK4rEq8k+Dxkq1yaJe/MWr3M0i
csB7D4VEL+ENb5kZO7DYK5P1mJ5DA826bucrbdWGgRZRaEG086kxq7sIJlZORKwg
rZUxwasFDgP5TmFltmYSE+L+vfIOFH78MsQsV9bQZS2jfJdU3a9ZTX/YRevWaf0I
TaLPbMMOFwh2Rsh9x0Q0pSSfRBUh6/L0TZuzurGzs7fie84WZWrIvqLLk1mAzOsU
RMtDJEYIzwUwev55lGJ24YkCVgPOfKdtOl8oUYEe0uJftNxaRrkUcW9xjHkqv9nn
aicosNQtHxmUMt4F+3mEJHJ/oLtshliUDI5TuGfOtztXlALXrpxzbjQj4k5QHqEp
+4yf03jlpbsf45+TASgrnjnPonSykgRl1bBZLPqH/lbFYlJ2CtdizP+VSFBDWUl3
dJoK84Ym6204Ay1sdo52LtEt9YpYWbXbwTdWAHtiVajfQqSydX+rtKFsdfcY6gqz
bTVEWb6Hw+o9LTLe8WkIXH/llfi9Ybn9S4Dl0K0R7nBT1kS3bc2XZWRtooTioSEw
vLPF7BpS+U214+pPucNpjJ3/E50fxC0qhFDBpaO5oxkZHtPpMRRKYIzznTBmQ4Qu
JX3tVr2OhVcRw4ccG5eTHm61UJ+ndNF5EBTEMQ2beDp+dbGdpP9vj+jS+lgcIz+y
T2dgikDHKF+s92+n6iHD1F71tsyOGHLQyqWNtXH4Ewp9HvquIVV/tAzpi3s/MyEm
jf1jv848XbLCvErDHM2nluMXw/HY8LBPEcflzfitf42tKGZvQDMmUbrTIowIlJGu
T7DOeVQHxVnN2nii0UMCbJZXcL/CcBbEddg8NajrYIq5ZLUHOWGhuIu5NvXMs6nl
jrHUiISVUZG2jpJ91Q+7IYatErd0sr7oBBTnQ8OmZMPXDlw7EBYrw7QkOq2Or8lP
Lgu+xle48veFQfPR2/j4ck8nd7MnTbXU2144VGkBKmEbdmamA7ZAqCQmZMYj0h7z
bMEvprvsKigV0c+8pSxiGGa5wb+E6mtyIvIQQmFTKEpTilURe9jGOeDwtfpSq9ej
Dt/LqQ17/M3ItULQG7CTxk7GHtZWQ1AytHCU6xvFHKr042Q6namExv3FVSfgWN76
D+5SlY4aOi3FuAbj25gmRiEXkamq7eUD/CzlLHhd3HNoI1Hu1XdNC0VB1s1E41rz
20KuYLqgOKQlRPWpQSLcSRp/fn3G4g4DjN8aUZjNshXJ17j1ZyOT+5Z9IfUfkiX+
2f5/x9zb6MjDkDL8ct3Lc6lpZhmlyckoctxi8ltPZWyZFX9LQ8X5WTSz9pJqqxDB
`protect END_PROTECTED
