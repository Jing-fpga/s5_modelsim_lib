`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dzZSDZQbAMsfUmQDOS8X0oC962I2QzwRk8LdITKEuGzUa2JXzQnJ7ORwF7pdSUaR
LfStxNtGFqW6owIaEzXo/6scROGCljWxReXiCt5w+DNnMHcXbTQ2cHM7dmBMOYJF
e/0jveF9+5Dj1h/heX+DQ+B41r5iemSmQ5UFsT/zctkhSFhGkDtTu7CSaK3s8mhd
zpdZ9dg3GAuLWdBTf17Tx1T1q1oYiMeXUjWVShnpPs2GrxCC4bdRIMe1wVgVyyy5
Byb2usc1gSrobXfyJuy9wQWe50szXNCmaldi11PU96qJD9JL8/z+LQVvjuRuhziR
pQGaCq3KTVGNJwrmNQF6K6Mmd96kbeGDj7VCNOUPDNvF7SRuktQnA4VvS/k+uzs0
MoUZ+iEuLjd6j9OcFcuJjgRgXvIAkiqjBumeNwyHVMQdi7+L7oo8B46IRnWdd0jv
R4vYvJf/Dp8K3a3IgahftfHUPV5dE8WFEZ0hekSFhtE3d9KDsHWfD3yUQFX1KSX8
hw3BibwixXIm+QRXIg4wsCoYP8sUDCOEoxE8lTTZ5OR7vJl7Tags2kDC+wkJx+I+
6UDrlbiRF5whnG+I2QcLb0XMJDpEx6RALiRImIjEGyuXkEYX5nYBc7WZlO5iXwRO
dgUQBhMAF9wY7moZnftnSuyucSUGMvDddemSlBxzu/CtI5OJr1dPqEJG1f1jZ8OX
hky2PIyPAKCA7GiLyp61YM25CrqXAQxh1neWCTDwS5hoZmlC74xcTDUP0l6DUaAp
gPga1IA/MkjC6RFp4loE+FZev+cD6wyRFioBY1cuIBVaCqiolKZgEAw4xCoykV2h
ZPqEw0ZdDj7Vu40yvyTKBqrAsIKrjsHMeyb+b4///v0tfaXQCYbweY8XBVguzIDV
GDACOyPINNTGZ6Y8IEPbnWJ38g7QJDcg9aBQoGKzjjKnOwmqfbZfwgIeiDRGcAxp
D2J44Z7v1NoFH3ILR/nnfqF7M8RO4n04ERAdv8hhL+U0+orBAjFK4Wxs4GKucsd6
kibgw+vW/D+INriSEMZWhxZlkhSPDrs/NLFPu/FyN3IhnlxfZxSe4hlzPaWZCIgQ
Y8M59JF+uFttc5zgxErZg/VLabGxArnfxGbm8+smTELOEQYGT8XM79YAqv7xqrRQ
Xpi7LBofzv/UuLisJ2gebsS9ZglvX5ACY3h+nX8BoWdHy04Z1KFHVxxLqbEiMMCS
/tsKcnev6s6+1HfVQoAL5Gy1bB7hhgwgweS4qS/pQ4C2mWwh0jER5zI5Vu/G8kl5
+kONFfryM6jkYyvAx0bw8KHNXfbak2gc+TiQc0SyN3H+vkhA5H9X8WWWK2aPjS5V
qMUiWJeV/Usu33tPuxkrk5WRPW+Do3Ri6ZXv+UN1JQCwxIrMqA1p2tSSQHkypmTF
MFKc3QLpQHyfrXyfExAZKwsatq96yuwyEbUNCykUXb8SmyagRv6Wzb1hue7d8Fsd
yNm331NI+n2wMtReKFWLjHlITn/0xLD9FhxnGiA5VmsWzEhNqYQUXaJiqLYlehfE
fj6d8EtEpivFC53SMZhfIzgNVYQYbTfT5u2wEstY051qeJCLTWZQhTSObrYH5PtX
FD8cH2nurO4GrPHppu18MwAWVnll8i0WMHL3fl1sgjyFdXAj6q+pPi2GUWURCODP
0RsQQ2P9ThzvD7f+fJtoHEBn+qBPFE09agjjhLCbM7VHHYSOrghH7mr0MEPFjwas
UBMQwnbDd4Kdz9U4FwlRtwxEtgfZcMx7N8reaWMJFG0lIq+bqVwxtvHwzaGSkKaH
imtZyzx9IaHG7l/X+TbpWGNIMMA31+BR44pa684szIZCnJHeNUaJQoi8Wiu6ZwCI
FNrf3fYOkUSfJ+krwh7dE3s22kwbro8a4YjYVhQy/AB8tBSP5PaMEWchTgI3mItv
0fB6DKKz+Pby8IlZ27fsmkHYRwYgjzUTLYWBK1FybKjRSLvZo91kM34IiVuCNQAE
zj+1fP65ubT852ttvZGJI0dGKjlrgdRAmaftPoZ9gJXToZflFgwP4Ckf7L9op4ii
+qkCe5vgQOY/uORa+o63OEWe+0LxHCTj2ga+jCvIp313rric1xh1rURKfGh8Y/AM
0oHPiDgtp4ZwbgWytUqjcehJiSmRVZT39xA5G2BofWc26yK+7Vd+RbnuXkzn7vcT
i/Yz+eqO6UpfRNZh3xzVueJoYGsfPDRt3nmrLsIoO+wo4jeCLNyk78p8mDi+QjIC
21yzfTNHONoTW62wzwCTM4770Rw+imujSDhaXkxpuQq/A07MXs32XaUjnx0IgoVV
mSo3hr85Z4oOmdeHmIjLxmTnsHbWdRRXH72KBH/WaqdiGFkD7uTa8Qn45NspFXOL
T/myndoMwUQYi10t4439VmQyqH7BAzzSOH0WWTecq8gBizauov9DxDbG0OF6Zfa2
wH75rxvLTWo30aMRRv+IINJrpLpsqxjjrCVVdUKsg2bHhI7NhdO4CdJmtwoNLj/K
H4wukDOcMLUy3fmbidKAkeEMUKkJztyB8s8/vcBRpEp1Sh6Ng10lyAn3CqNoYRlQ
hGZI82mbHkSRodlfMidHPuATXe10DRIUkNEGK87a/vEez3g761p5vqqN41VyY7sa
D+Fw0lylwVIjvahMo33w9gtzLQYX3ulEqyfNV1mFxJ+XGWaut+OYJv3uU9c4FESm
K2WNKRfJS/y6EWQ3eEqpxnCTo3RR5RZnMYWU2KdcBBDxYht6BcpC5k8+mYM/JulI
kp6r7w0Nol9/X0n1lggJm+L8oOdV1ai8DjGG9EoyC3nZtWR9dVhhthGapxXjkps9
gogmRDgJOPxwmIWw49lUphyYLwvsc5e5yi2NDG8AjvqTUGz/Na/t94lOA/7M8V3N
/8t1DcNJTEev8eMD6yjUGETcl3/aMz5QXnbwhTL7wCj+LemjoLCDK3iYasYQUum3
ifgUWp9D5OMbydB55aaRdFtkgy76r3XThsRNZ3E9GWbcz9PBD2PUoORTVmwWXzHe
MWgxBj4D25pinnHiKm+Kxw8uEey/Te2J9uMmURaLf1eHkzJPMRDrrDtfcZeJHO2a
oaSjXgOZ/XyA/YHMuYw3aD6d9zxYxwxQZ8belFdu0YoSvgT+3+6pEPBp5Piy6D1l
mnmOAVk6WMC1JiWhjaMeXs+WqlZ2VY77dslnoXJnATGNlbMWJp3cs5wfiIMKKdyv
/sSgZOIDXph41WcjSkk2rkbcGAZltLDh08HvvmNRHX5K//NxsXfKwSzY9Pzecm/o
wvmKRCIgcAbypHhoEQHLuq7DBQZPyWZ9SO3R14SaVHMKOIMrZkF+vq5mXODbkR22
fgXgjeqgsitjAYEZqzzrm4d07+KWWAtVsUyFVdoxElKZp2DUiAo/ATD3A2NFoQvs
sV0EpAkYxA9keP1kGQ4j/p3nPPpKSqHTXBHCOYMgM0OJyqdZ5w6XgSBCcC7YPV1A
E7rjRgxa0gq5l3rbpBEM/QPCJLQfD1jUwE85mjpSH1DFQVrqcCRBw5VQX290Fkqf
VSj1VzfL+tSWISEb5OQ00qdXlbMvSn2ECPwenaXuTovPPo5Wg2qw/9bAa7CFP4oL
VZJQWrnUPJtJ8zwupP/TAhmF4w/wEOxQz1RLFYKy7cLN31W2FjGWGQBp0k55msnW
DEVVIIO8qBEwYKQYhz9MdqE4iYr5N/V/F5cOCtLOf3RnVokMttLZDAKfqWlWUaZ9
IDsQXNJUd5YPgcPksvapE6OLw1qALGOm0It+9aFeUmxXocw4TICjAzohFF0rt07n
uKkHVHUgAkQ7NuLj11Nd7cRX8XOCwy48wA84+LwI5pMaXh1cZCER5LTINNUUNW4r
6JTdlGq82sHmz4BBiBumQ0AGCJNcA3IvMLqXfZlEMi2y2knlVNNZLcFVjXMe/8WX
V612RwjtqLJhcJuwyzUI2AVP7qsGanEIAIy5BiqYCIkfPM7kyK2P2urJSqyNj8fJ
crELcTHVpTOjurS7rFv0SQ7t+hwrhrQ/ZJg49MTv2UkVTIq8g9TtFGUBwjISr2GQ
SCFpZhwNmhNwwyEVstmhduXAIiqAikSlyE+RStKMBJIRgPlhfEO/1tIm+o3yhRjo
uBg4C4GDWlQ8OqcDJeuRdw8cI8vjUF8XJU0VU6GpK9C1vDP4I/6TYqFhkbZc7lB2
Yik8S/VHFPkzug8zEbjD/rpzLUITHHh1KMadiTCaKSCKKo+5sdRJ1Fkdmb9JhnyT
/p++XyfUagPzJcbSoK3f935MluQZ45Jw1Aoqah5Jf4fj9Vev/Cam2pna6YyOkArz
rbjPXxxGsHnMiuOTbngtVn6IkHRPtgvpWB5cQ/o66dPDRZ0QynWb6kNI7jfqNCNl
9Tz2ZnBVbEuhXCD+ijqTBr26VFOHaAfd+EnrjxW4fGjhIE8SZH4LmIqC8Ow/mOyU
C5MHFN/H/jUpWvPQbqQxjp2/rCx3Fs1+pG5dlEm77oNEW3DRIO4JiBnrfHmOvmlO
50oh4n18LcbMf0pIabSgf55Ec1l6Ql5wuWTFDqLaKXBSsVoSNe4O7MIeA+JyyMaa
eMz719lmzTQ86Tqhr0FxAxh006oK4A/dGtpq5IbN1pOXqMB/aDOoherFtLN6QS/p
eY+Phz68zWOHiHfnbgN/GAEGcwJsrC1eT4WzHw6XGd3P+wUUTcHEDdrfjsqzMXsq
A5e43sOSl5QUYpoIrz4DFOjb08AFRSun8zw8JdD5f6oZn7WgsFY+/mSCt0YBo6no
3qZd40S2iJHWuAtwA6rIq9lRu5W1IAwVU7otTL9xsZNFEri/21slzjYG3BQPMV3Q
pC+RhsAHUXnR9w5JJ0q5SGTuRFxiDtxvgy0HzjrmgQDwrCs8UoLNy8f18+BzxxQg
oMZHD40s8d3NPwmlSfeH2w0GVLtrA5w1ddpEdhb1jeevzjNG5hGSR2dKV/S7/0Jj
1eXr+i5MT+ecfvQegbAmHHgjjZ756ZAlrNz680GeWe751AAPhi79c09Bt27PyWOJ
+v+YNPxfw4mKVWe3bwsSdIHwRnGTqhDpsF4hS5De4M1FGrkkWsHWXH1xgGWt28PB
ysbrWOaWpF2FZPuhguj197zl+QdPzNVPcwz4T9FrgqnmRCun8oOAkmyxCqKgXCMx
8kLICBBPhrxZxPX5Rv/nyrtRAM83wFqlypYNCi84I5yU4vZh73EzqldKhIq1e+AI
fUFkk7Jvl/sMal0u8rSrl1G9FfHcdPSzBWw+wFkOJFTW52BZ/obvwh8+twpyA2JL
qk42w3cqK2ei9iWeL2uoPn7FXtF7P1i2vzlGj23EjN4o2AzurlTv8Eb0AMQFRLJY
OrJrSxy0nCjDISDSqVrFD+lDiBd8ut0GBwLlKk+j9Yt2yAPj7p06gEGagJtJPu6V
xYtdfNR40AkjETX5/JZB9n7psMZWHrz8wPLN0rX2D2hcmGgT6FnjnCsaWj6d0QbL
4kB9dP9xMmtJ6ctTiEd4r82reRtBx4ft+zgo+0Zyd4+k0i6P4gONlK5TcU1ELGgK
hFrN1yBl1DAEiO7NNhFd37VOa1Sc0eyW1LxWbnIaKsvERCqEz9aF7DAyRGBd5Vp3
0nigXZJ0DdEAAVGJ4gCXamuQQQz4s+mB0xrzbWq887swT+4vvR6DlzFm0oBo43y7
N6exbWw2Oayw/wCHhksXBNQA7R5pFZQQnqMJ3xHut8+Yx6TXC73Xl2bM6j3DcUVI
mAhnFPN6R4ARsLPVMjeDlR+THxR+leT5/paoFpqa7/VVaTowRgUSwMx6UEC8VE1F
3lw/2SjnA8t0W4or94D14CTyA0myc174le4tU7PeMXyYBoMKhNd8MMLAGY/jcuWA
k+yl5Gsc+Iw7Z1/YW9RBoaqBdyk+bZbhDQ0kTuClqDxCyqwotIOKyFVlbE+fO3L5
RJmwsJdm5qNoLsdPBi3BFqvUbSvZAklbe2/1VwPMeUtUR8RZ8aH/BahANStmz2DZ
jjibf0mVS8pQg6sNwQ98Yn5JqQjdUxjjGu0vqNXkaeTgTrjbfoKgxp4qxyyTbCox
81pVczSHespywcLyXS5AovFJjir5Z4xNxBOi/LCgjqNNb4JQgsojZ4+1WzWw5lbm
S0sEzyorKATIqoRTUQZU/z+Gi99SeGXfUUbgqC8UkgTLQpULQl03OgMW2MuKVoHR
ax0vgYmty2Kitv2ogEjTMO1bwZw3zmq4OBpk/nsB/QCMfOh/AVMi7RFdEFoSVl78
rMI3XZLCoDENXCcYGKVTPBl7uOg4k5E9/DkUia1Nasuik2zjpZ2Syoq231jOwoEO
yhFBZFIK9CtpkZyvNkTsCBMBpEY9dsw8/+ApWgAdu+urGv/mx78MFyUVDG3eENBb
GMmWLxM0DsXCACl9MQ6wQYQueoafE48DAHDnmM/JsEnTNvk9W4qcBrHiuLKPhqX9
tovIazIpWY8dOKRtF2VN8mVUxfmbcE9uMgJeo2Z4T5Xq3ZpjLuAm84HIDJQQ1JLa
5bQCLBVhC3BbNCuUreemO3nlm0ryHNlw8DYAUhivvqSBRqg/GZFiglWdz/8IEmoA
N7QOR9HeeAVeDzKijIae1xUe4Gmz9bkVZB+RC/uwgZcq3w7/x7WE5VEy+hvYTjkD
1prwQzWF7RGhYJZ7Jp1TIJbtfIyibdFinpDjseLOCJvGt4VE1NEQcAC/ts3H91/v
`protect END_PROTECTED
