`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H3CGcbCAOTffEuBc9dU7vxr4tgJqGoKa62CQTTm+9YHYLC6EAWWnLGmLYa2JXZbM
ohBeky1zBLMinJCPLZV6oUGSYFwns10X8Evg5tEXKt3rsAZ/Q/HQVKCpktl/TSJZ
ZPGI+59y+Z0Sa77gb8b4MzhC9RCBsiDiinereTFQbpTtz7UErab0s+K3BsQ2nUgr
HJ4kXleonGR5EwA9Hhur1MsBFUWByxxjxiwh2NsTvvjk+ebfDh08PJ343A4Cpv2h
QYkFP4PEvveA1NQ+rPoJR2NS1Jj3z9OvnYfTPn1Jy6wYXghkIQR1jYskxkpaPpUJ
mp0pGbTDnnOGG/5WVwwgDLBSgY/oEqt8LnjyJc+Fdr86gfR4ST+fPeI03EOOyiFY
qBi3FEx6OUSOHJ6YaNLB2Urx88v0OwAQmJ1WQSDejXGNS5OdN8Hu6z3Qo3r7uISp
wrBfzLm5FwxwTv5lUn1Q7uH3rIS0E4yDciKlFc87Osz4O85tJd7YVgUmI9WZak4g
B/whX+YAqXxZLGL0S6UkOanbinDLc1I3wsO7mfNjQjJTq1FEOs+vldct0JeqApNd
LUSp6/Jx/gk4FRqwWvByXt4jCSpiYZ9/liMO3TPaOOcRFyibjaHmNXgeSE4UkOh6
Cj3QBvFgeP+Fz1U4tauC6dKk/dAnW/8mO0GbKmqS5Bc6skIapTmzgpHL1GTmlcS7
REEh4fxf6Pu6HD1zOYGqq3grD4R/blgJc7ay3u0cdt+tMgBVz3J01XcILIj9T6PG
Nk4j13a+rnAmF/LzXVw29Afpye1mvFxpLSHmoyxemZVmm15gC9EqE4r+PAJCHQUQ
Ijk0NDMqZa45jxF07AJfdpd47Us5YqhxzyxQEDNgY8LwEkMSbl6tAEilVrvgV/vL
CSzdjJleNnGJT3OyBzHGlJtJBD1NjTcOcZZNCikLugNYbZ3fZygtO3CKoTMsUUzE
/E0QH0O/W3Hx8d6w+2oqlb/ZDPHVQyAH42H7D4LrhxTBLC3cbQmlLCsKsjtgbWRJ
rTpz6MfEtmatlkLKVKWvEw6NPMvps+7KocBPGOSVDBbeMwou90HldYovUWnUibgv
nqcKsmYyLg0aSypsjJJjX05eXmbYJ5+kq4R/9UCsqZpqgpOoXaS/nCjKyKRkYoJg
KJC8dLofXPliOP9WY7/zxK6afkFP7qaBdLYEwy0JcW4T/KDjwnOmd9IPSII+YWep
YzA/t+ff9g/xamX8dQ2wG9xVrK/jnMQWCEyLmvcG/r2kPnZFgH7dhan+bAkqn1da
X6jxp2yaExMwNugx1dr0DEz9dl+kN+ELrixU/NNgOOu0I+Y4TpimV3prJCIKXQrk
eYor6Z4wncNxSvZ+tWiLGqj7ob50VlzUE+kmwqVinQH9cmgKuVf7Be4XwIEI7kNZ
90JRyfeJp+ZnWu5UVvlLoAqluymhMWtbGzydsKwIEnrYSXMVj86hdSlVfdkSuiyf
INgr2yyW999F3Du3wePTsYxank8uH03DOcwlg/EaXMPtYhnARZe+hwyQWcSt0t+m
cCLa5Ew6ZnCgCou3BCVVi3oxMuyYrObec3LgczKr26UiJz1WQpMn7PdDdeHbzJtw
csb2t/5Zy3fkdz3J1GIxAqn+KDkgje71g5br0X4joCW5ghXUtwe+7eGXe7zh48Ni
dPj1IpTcSAgWmzakWU3PR6FoM3jWZdQV/Q33KtUGWw1bajlYP6Acv1accZOfZbyJ
oDV85zJ/01lt4ftkVDa0zBj2vxfoV/jZz8/0HQZgy1v2WWSKcQ/cFsr6eS0wlo70
GGHxvBnd0SpAyrzCEUU+YOcISNpVbrupgXoAzhkQ0V8BHeZCXc1lw5wNUqEq6JB8
f0rjXDBqOU/MTVgW+OjqRPx/gG8ty4CUpRTybd8rWv1rc3QoQ2ttUYnehIDz3yYP
tGdTiiMBRfYzIR3/u/vLpjtgtIOICJWeRLhbJueCuQmLlb0XIYxrc0mc6sjRd1PG
jCg/hXG4J2Q+7vdf1Vp4k/orFbjJIPmEf1SX8RvHpBGEY8E1m8FXnaNUwonY0/1a
rp3FeZRNdZFeAtw5a8ywuv0Pc3QuyHF175UGN8iToacLw1jEE9D3/joGl3h5eZ0a
YJlvkvPu9cS7+gUXh+rg/dfcmdIrqj7nxEoQvHuMXjP6/0BNJ0b1LeCK9uPLqIe9
lH7QIePVkqPNhPxzmfWlXAE6fWJmbctkzN7UqGxhldCE/Ck6tpA0hZTloyIcJAA2
ZcNpCrP5UR+2lys1BxK5aN7cdA9dXLMRTN2GI6Ddf80a+kvYCYn8fj3bPLR3fXeX
66/IA7oX9zZtatyET3QErfPq5hLvuIcnDP2nUjYbcRccqd65lrptWxaz5DUMWDEB
Ea3v9mXpSSRPIVf3VV+AlzctSWosNAgcalEJAbkLycuA/xoYA1q3dV5YifP5RUEP
avF6LK5Qq1jFJ5n3OhL6TvMidPKi4DNoIT5UMEGyL709sJdmvaSg3R5Ce827qgnP
jBi+GSbAdltfJX3aYGz0pkSwhUrQZzwWLbpqr443Z4sZ0IASEmwORzXgS6RTgaZZ
CtFPVwNeGRmGxCQvFuNT7zw+r4QCWvhCF8+ITXJzOKph9b9KkZJoiPt5mBGO6iV+
JHi09dfAkkdtB8JH/+spODNntcvzkJiZ3JXaM+73YXLXaturjAFpgFThU/1Fr87d
jyJ1JqbNqQYv8ps4KHTkTHUxvFhlr/oVYPVt+z7L1MakObXhZJ+8YHu6PUKXjWKZ
pKC36EX4Gm39Q0E07FUKG/aX55JX37cvIhTDCcUrh5OkqdCJHDo1WqJlQTmv4gKr
KVGDbLuABEg/21pcZxDb2LHq132MN7SAmVDqHj3QM3FKHFMq10aVY2+CxRhBpL13
SXsH0uyu91rLAMIUc1+pUuD14CmJYoavrRjhIM1F2jZWo6e6HwrZCvHnCNvw/os+
Gak6k3nVMpLfP+8cPR3PCUrnqsMSCXfIzl8VBsiQt1nt6RNpc/0Da7CM2lTmJMre
CoZ5NcA0TU++LhjTPEbNj9zhjnd33nw9zr1ZRVaUIfM0G0S9ng9re3uf5Swy4SP1
zLsZklhyNWuIQSdroKs/v45pokgOZpfUDKPGx7Ym40f4C76o0SfjnOd1MjaJ5iBz
CHEXyaTpXmd7BI7TV5P84sm+OARAOfqukdHTZKSQf4ZWm1HdKnXFvndLYie3H0L4
vZYxNBDRvK1EdGJd4fv0DfyFj+0k9BS8G5wGXl4gEeHebLnJoYSkiz04sh4tk4pr
68xAqSFEjmXfFsKHVr7KI2D6qAxJf39QMfbxskN2GPe/MhbSCm11nuL7XRFxYwPk
dJfQI3QJTXLAuoYBv8PuEB9NQ5tJPw3FpuItQWmOf00d0+BGbFG9YBkZ8lqWUbdr
6DNJSsQYMyJcwrGL6SLcfzmiR4V9asU/VupRzNMx+Jq3Kbe3U0HpykIzzH7K43pd
NTBsimepp1aKoRaflzL6hPKlK8enGTYnIfx5SyCl1zJ4+/VRW4jmi1TMlzSoNGKQ
n+F/oQIRiOuwWwoNsciDGBQpYz5nzcdLw0+Im8ZGV47pmjKpiPNGSt59F7lUSqEK
QC6LcVLocBfFwk+gg7IdSj1AZBzTZHgtF0jdmXr1t+i9ijE1osHpIT40NHcWshv/
QChmScBk+skMX0tL/0XiLrihLshEzECwcRsGC4i2TsJg5p6Bd2R55JMDSp9ik+6I
WK9nB5JYwIC3aT0iD1TVMMF649pwK+iBPctONeXfwZqZ7UHcEGD5689gGYmmOq7x
xSryA1hLomIOv5c8IUL7DpRvhiynhkL07s2I4guOAcUM/BkTSwofuxTczkdQjOpA
vwXmW6u+rc8IG6/2lfVxp0nE/IdfRp7/5JYbKpQ+yGy6Wu51IWR9zBGwVpv10aQ7
qQaYRbwAPVuxg77LH2DQfq5mzfUQARtO6KJ9SAXog5ek9HwvonGZ62a0s6xiqXJ7
hNx8ntIpMDDjqE5fqIGw1iLDBndVGBd7zPu18hpZg83Kn/MDlc5YtnAVr/PaZQUb
Ql8gqR4PShT9O0LAWjsYvEhHWcrJUsScwyk+raNVJseT4xbijax0YWXJoXGAVKYk
E8hcDdyVRPyvO8XJYBiHmHejWG+eve5GF2aDpdXTJBqWnJOxCxOQBwl5K4WlFZIm
N2b0W+aSTohdvHc6oOk8uQ==
`protect END_PROTECTED
