`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w9MkGSjpvgnQ2kEfz/j6y50NjDgOOwXHcRvPbomXGDGiGbS5UJ2vkqnl6bJ5srwF
EOg3hunHoz1mk2k6RRajcG62YnwZW4+qT9f+A4yrmNeSP3XOt1M/pYJQCJOyzqMO
7UeNVnXPOYUyffzdhcWNXmte5xESGbtMdayujO+pfEVWTcurFDBV+ZyqbhTtxAyj
2gkSqGlcOr9+44+hs6kCbaYTqandH384WhrF9DPbatHVbPyDL0ONBvwI5gRyoek6
g7JpjCi2FgJVG3bBfIFaKD+IxkEXmm9N+jhxGVvPXhyl1T0ciD/VeACeQjcCCa18
FrFUkeatPB20v1yduL7RSdSrHz3aj0VaiOXRXXokt2XyXLpHSGreX0L1AnRKBfdk
KHOBxZCKnMN/KWebdEOrB/T6Ega3YahxuTmD5Wb7FIQ1I+1meSPuAlnPDXohO2GA
HDcENEOnKSP/GZoF1tAiaMtRROdUFCnD3czxfFD8fsDNNTUS85HXjl2cCreDvn9h
aZiKTM9PAOkF+qzyiAHOyWIRDhbtt7YQg+8R+w0MLiHpGaBEyGtcMGdag3efBoxY
wLNiZYCet0y+TpzZPNU0swlDPmaXENVQ+4Ukb40D5+DdUHkjcwcvTGseQDNaBHAT
RprOduCOk/2ufnZayZX2kM3vTzE31GOGEqLxg54t3wrfKoHZuw8/ad+XL8IqkrIP
Qtd6SJpOjWEhh8BBUAdzt26D1NVhSRY+WcCbe+gs1+k1nd9nJ0+6cvLvvDKTxEE8
gw16T8T2Z7sgqvSB3qOCb8VAys8RvWJe9mnpk14N2vcwavxN6Ci7wNgp6+MIHbUV
TbZWs29FaBX4/vuj5VZJcNXLCRtaM6KMbR4bla/snFgJHUyY57jx01X079TmLzaB
/xs1lNRsNchhCQgfmJxr5IpG7dePQPF+yh6NOCac39zh6onbp84Bb9HTLnkGxBfy
6u4n35mrmGY7EETiwOolzcF0RN9YZO8bCIQaZTu5HTXq0EtWW0uhH81PKi8eyV2B
ZXExQ10xA5XM/VlqKG1tTs/ZFWl7z/dUwu4hFRP6RtcXzZBrem+nzNfLw8yYd36M
DHMtRM2/91EugpJjIj4shNHv+s9dTnqFi7fM2z+5QD3cepRV7PADOChKvP1zQw1W
DXZkp6mVu1X8lvUIZiWqgFg6lj2KeSlT29r9zJNhyk2pJ7SQcT5lt7t3Zkb7JDDV
BIl2cLLYclt0ggha1vdLS7zCTntGrofUQt8Wfv5+XG/bcnC6K2M/BVLivsCwkGSS
b/CuyWm1ghY8p90lbLTZXdQlSpxdarv4WMmkbt2sFqNXMNDR+A/P1ovcrIb3i5z6
MXIO7ILyO32nrjKznOpV4XOs/fQnbD58c2t8l+FlCYrCAe/xpgaR2jZh7TZU3NwZ
0lJN+5lnoPpknGTg/KIlWw==
`protect END_PROTECTED
