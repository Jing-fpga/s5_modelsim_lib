`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4bBBRT1edDwYG8UW4Qx8e6PXGevI7NZKvuHxRoF0vUaoj2QrJELQ+H4D0fVI2En9
o0IAt/bb5wAsDh0RSIpGU7Qh9Vul0xDbQJSv51xCE0aR+okhLgS1hPGgkHDnFWg4
ndsVDjf3bD2mfYMxkGrLADtr01t5aPqcV2e+fhiiTz5VDLzvE432JvMEPj6i1IG1
6LDwHX8Cv5B4BhwGv/e1FcWsYQB/2nwXM4GwShAt1t1I03Q05YjPzHelyTD4wGpI
0H9eD2k9vfm9zzMMo3JSzVYvBVyeb8p8BZu5qfP2JlrGqDHB7ZfJUu84JIVAgVSz
+aJ+L2O6rGJhl5JV5IMe4jtaVjjaWGwhj2C6uyqh6s5Qe86dVj5OZ350VLQ+ZTFV
jMWMPn6M9sK01cGFDMVU7Y0nRurGSUh0xP1ntWnfB1IfhD8glenZx0b+2PD30Gz+
U+H3LlaO3zrbkYN0me2up4i6scY6hBYkuX0WsvPvZU7G085vEYlvhC0KopFBpvXa
/61vOcZTzh4ZFRL5Q2YI/M7CjbC/HBB5cF6S++dXPFrbGrdN8F/UCmc3uD0c2LxX
wEYC2x8e24OkJfXvC6cv9r2gS0gtmQVD3H4vAkhJjmssxjdlXQO07QiBYoodbK4H
0bSrXx30enyMllZ43BX/iCkXsYj2EC2plP10qK1Z9lk9V3QmS+BqaCjg80LKOvYK
J6q/2mS6OGMoMegZi2Jn9JZwkQ/BMqD9D7YTPmKgNGt8j0Da/oEeM9MULjEomGP7
h68nmoy4u4vvAdBRxwG5Ha0m6Lj4ySu3sLjcP4jycqy8A8NtjgI3zqgZSkJMfEyM
VQZwpUtvQ0Z3J0jLiSGYPXgqeRftmrLSJQrZ2miEQj/M1bv2T5SXukpc/rBDSUpi
2HB1h4cexfGLpVWAUO/L/BpppUxd9hju+ehZ+DGxN0YrS2aTiRPo+ZeBJ59mu2Y9
Gd8jPsm66Rwnr8I0DK04qbdeJ0ssh91hwb8Y+L1R+tqhHNw7KPZyUY49O+Tjalr8
LBnoejtGmeLMy4w/lYQaryzE/BSTn8R01Bwfq1tIp+afmZz10AWghLx6NR8XlEct
havlHe/4gQwbPBw9TXFAemGG0xdB6vm+C9lLmhBboDOqTC3QVffLN4AJyO93gAGI
4jJae25JMNzkPMn//Lsx3UH02/4iMZrAyhGzsggrfoVl5455fOfbqGUjcuQ8NL6D
0SiB6G3hnkxdrTsU7R3LVxEu6FbTQWIfL/meUwFuOUEzj2mOAFdEpBHHjfOLYVxk
1fFIpbOaTct3ozMrxdNVo/091GBl48ulECpsDtkfdrWAsFyDKddOS19wY8AX//rr
U9LIY1yLPNyeYLD/JoUVDSpJrzdiV+196nSVOG6GGmNfEOn3JHnKxgLNlXxdj6D6
S6e3mJ+fai1lFEir7B/4uvHV2rJ5O5zXqkraScLOa56E53VzecSchap6UVEagZkO
p5ELNGTWe01ewOck2+N8YJ5tNWvhVoMFEEp2ryj768Z82BFSglGKW5kKdtOot2ML
icGhntwK/B8c2HiYQtkOfgUx1N9C7KcNjAhckndRV0Y+5a1gGPa7qGcx/ugbM6z2
gfg4ycRUC9gN7DkkuXY1TyVwpgs19VMCPgs5kSQS0q4nmuyg0lBGE+1i7MTfyQRy
9fR436LElCkb1OiLshH5+N99FQN9GpQw2B4svVePzIaSpI1cp9a1TCj4MEBY2HcJ
E7+ZTmwpQxBWssg9HTsMbM08totSTsJgoLsORH0UM03FtdNMQtoMBIJe1uDh2f2X
6zX864PZIjnBlhVjJyolSLGhoCHGapzagQ5n+u00tPsj5JIv8+IBJC2lfpfS0VKK
3eQHXRX4RZ6nXIk6Qd3keciarP40R3k06s2PA/lOv4BQNh0npyU+upyWuwr6hjEd
phW2fN84oSMf9lBxFKGiupPml4s6P70FNo6hn0sEr9O9U17Ntt6Y4nubXQpvT0lh
zOXnVu4JworUKWG5LMELqPb/le+nnnv+x3VVI8sCmJg8h4pVglia3VWOzMT9MnIT
+wjDkdP+KiuCqygE4DfvVkwVIbHCC5AShzSq2KAl7joWbvgrJyCdlfoW0h3wFlQg
Y9EWXbndBe397stU203z/CiNU0IYRMlWhK/jO68j9SIj2cBZMpfnbH8QMZNtqHpO
t1faFdQtl1EpfG1PQWQKN+xYEazR8KWIabwT1fpD+cb7aca2ASruaFSR8aEco1ca
9LxWn9EOMimDqgBq3t7wnjZ58+YBn/i/zcKwAPB+xaUj/+mLnJ8yp8nOlHqBok4U
5J15zpe+rbRphXb7Xpe0fOHWDfOjsCuhWNs+tNZJ70am4eiZ/eq93+R/kUVt0viX
qQFfpZKrrkxZDyrNgsFrUPYb3xQZmvA/RWihhyqbeMzpOVHWJ/CoaMBqEz+MORsl
5M3VbQVque5aw0N2av+TBFZRpSqW1jB9WeKa8aMSHCKQh75Opy8ArY6PcKz3y0CI
SuH3jXvHgUqSeOTR2aeBIL7kxGi8v/oRKSlL7uVm8Lkc+iUD+dEoWhAzYB6KbxtE
cCcZ0dIPSpWg9FGRqWLEFx3SoPUzBOXPQehdLEINk4pXS7FTBfrUBAN/2cnw/qJl
fwpi9C9puDvF3V0qQE3uLdOPjmnTjI2fnPeJcNPz0YaIoxwh5loMpbyavgXqXVbM
6jcSh132bZHLbkSimoe9kOfdZG1oHFGcQHchPQZHmhpBnhfvHv4nbhuJhh9vp6hS
U0IdStmaHWIHP48HWnQVUa3mUwSih4p0/SFLHnywDhErhpHMfGXub1T3NAeeKoky
ahy18FjoHSeZmbiExTfzKKvtyXrFTQBD03PGKZ9Aw8g6XlYTCYhQ75sVT1xeTgI6
Zs8KxNvshcC/8uzhVdfx4+ZhF821gn42914SIAVCZ0/aeuTbH3iAs0Ah6hnylVts
qL7tjeQVoER9YIBesiioAjJFRQh/soowUesSkNSfPbm8vxGS84+ZBd+Dmj913RZ2
54kbnns497T2eDafRTIaBh8V00za6WllhaL0cE+Wmh3XHIF1d8ld5t4IURJQT9UP
6H9SIwZ/we8+FrOu/gsjWPWkMXA7yJayh9lx44O5TxcHRAgU/diFi2dcQRDzzR6P
K5dRBmaQ+ysHFfyk3lT0cRf1ohXpOmZ+/jW7gODf6HN6yCZ2c5vxw/RQYHEDxZXM
b+xgb5t80jxQ5+DQUG51fl2CAYsqmniKAK1ASs1c8M+PPx0wwexCyJN9FkJzSW0o
BR9ta85a85Q9SNoMds4tfsQhix+8GFTddZEKNVWsZsFlF78/f744cCnBLa2LuO8B
LUhnQbIalY8U2PuLCXl8OmXUz6mdyldN/j4u2xyIzof36tKFrYbpaRL8JHMJxrPu
lSocKd+f24oHfYimNOGiigPgUup/E6/F9zDc60w5WbV/CzB0W/iQ7wMUXgNuCCz0
sz3/cDMJl2tHrvDoD0xZR+qOolPRWuTAGg8/HurLidPPmIs/7/Hc5x24HjZhKX12
/jhInPWAe5T6jF5DeURfHYbU5KgP3VZtiaxt8lGKcwovQiBAwPZ9TBVXEhPOJ8/J
iHm5Ps40hqBu6LQ+S3TRpHKeYDS0rdYTSdeNbcRKFMWOA0jYao+j5IzBT6BcnrAp
Tm+eJby8utUZfrIqni7lHo3uHvYXZFqygMhSz4u1GYsJezFDNSwfPa5u5wIwTsr1
zYys77o42oAt5VG6+qZPoLNXz7yljZwgR63vADrrKjLOCq4OoTshVo0L+hAsuNoK
I4AlxAzLscAdxXXQeNAJJ/usoW48NciBPvUarhjQAMcbSYKaTfehoxaeUmzepYkR
awU0/7eX6tQJh8mD+vbAaeyFXCILfw/sqn8Ehpgrizzl8I/BfgTORhVkhfvJPPjK
9hGgIqHHCYlRjgRYUYX9BJ2jYwuEcTskMdIeyei8Sg5TCP6liEwB7ftjI/LCeCDh
o8CPKr+VosqPsQZaXsWmzkhm6deGBWduxXgkvnpVxWw6dRHqvDKTCKtjk8clJRBg
DTbD7urNfM9qwTnYaMk5pWDz6QTX33SxiE2wfvZZ9K5HDHLuktUlTJZHlff44BcI
vZ9Zwxdlbff0Zj/2VnRcDWSeJtMe9WBfchFxJgSkDJU2zfFvhUCUUzE0izatCAkD
02P+Zf+NlWVgKyd11uWFMmBVAJaQh36z1sDOJvkaznj3q/aE2pmWxDnBVPpP54D/
7dfV0nv7LHCK5VrpIDaN+dt+F4g/Dl++RFGgAsoqK/8iH3LAJB/Ww/8aq0+BDJxd
YvLa0yTI5jnUR9RRxxhVj3ihsD+k9wcCsGiUwgApbUvCveHbf/bxJAWEQbfAD4El
pX1J1GaNIcBmpTpAsgAb47wKhjQcx8uKtiP1FY5ug3+7LIjZV7AEWGhVLy2DzIrl
n4JSo5qfeRiDyvD/L+8747K2xZZ9NvbiDiSOFuhyzXP8K2bP+v7y/nhp1Mb6Gk4M
1PrSM5Y51h8jTSZ1VtcMPQXhIYVUSiSEdMt7OyR6FtGOM+oYt8L0bD1O0MKA+v9S
WQyM4KZ1231uNaWH3VAlL2psW/AsmgKA50xwcD2cYt7ekxusYuSCIsVCtmLgZ5FN
sTOD5fgPo8iL0uBN/+9ZzZf45OD2iFBXSLngHrQCXkHoZh1t2CnvMpaw9xDoFSKb
M6NCGe9gR9WL4+pf4b1V/uJbGB7lP81vJxxDLJvARXzfsYW3r6GQ93xWnRHdxvbt
BnkUtrjQ+z4BJFHkf2BED4RVJunV117ePXBnnLLMlrud42zCkrrGFq/J/qpXWzkP
ZXzp28P1Q+xKzQAdiRu1zhFpMisJ2dab9fUfmqQ0Fs3jut+uO5a/uaMqH50Jdkwm
+2HaigMT2X1JQdfd4dj3H1zN0aJ81vqgoRq6uR37TgKAG+LjGVcf+iCSqkvZCNPQ
SxpbDnD8uss5UCSAMU8E2I3HbNrmTnIWxKzJDn6BI04/AOQVDRTCUn1ooQtuq6uW
MMw6efiyGRbIJXI/guq8snTKVvX/T9lueT1zFm1HHnu1Mm1tTdlKai8bu6/Otbtl
Mm5tDvRNpaK2Mx9vLF+GWN+40g8V1mi+NQxkzflNqplceouvlSESkJWsb5UMdCCq
DEhtCLnv0MXemvbmpzseYE9wDhsKdJ2yUHd5y6Q4cukaeYQW7pBeW9kSXVWpwsbC
m8rMTCoOWlL4H02e11GdmTo1smQiugpJuxIaMXkAzRsf+OL87QsvSjIukgkJeT9X
hTHbKoMHneitRS8cl8ycXBiiOevW7OjFxsDlLTlJRRXkpV5FDdSN+o2use0lxMwa
hALoU99RDKEmnv/PnwgCgJUlE2ZRciZ8KZgdRFLiqA8X9288yEaF0cEMMe3eDkJp
EXSRtebf/zYh9Y7SkQaXl2fxX0/WVbeYqXRxKO2jW0ZqtN8MrWz5kM3WT0IRr4ss
fMD6x9sbDf5aI5l26J2WauezwWt77sgtRkxF/NWyADIEdjDofdWWOvtsvTVchwUE
fHopLHzmAnKFV0cdKxMAzgQTBsiDgdRpoxEXACgoH/8IuhtsVGjkS/hd3fGfuKKY
kQxpc/IqDt+p5qJZ7QWSou8evpcwheEByUy6d9qyZXikfhJ9csx65rQT3kxh0FNm
vpb+h2Hfoxe96N0I/KXstuEkCB5RFjvgRFS+aNe4pmX+o/X34q+kTLX0bKGVjavy
9IueBljn4qEEwSM42Qht+vLUXxGlOLxI7rVNQEynwY0VO9RVCYAhQLGHgJCVFxNy
Z3b9NSGAC/j+EXPqnzEHPeRR30MrDvzuPu6HHXkIVkQK31u28kqmpNxCDVJrNdXk
zflrtKH2wmASNbi8DVUQElsu8B7q5xa6B5DVIa5nIdIesKS1abSqq2fzSA7WDtCm
Qw+OXNaogZpi0hrp0/JgOu1jRO0qeoBYm4pvKet52EFdq8PHYDGZ8yyoxt/xA/a6
1FlM36yqePlRtQKrl8ipjTBC4vM1ntc5XUwlHaYQwc1saMBUCcd8V+190oNy051d
jkrMZh+pUXbPtOjsb0AnoMAZrW0WbJVvN7AyKzq2CaHsEn5pBNgVute/kBMxF5N1
q0h58oq+W+kFrQ4bAk2BPwlEUZVhkksImapQaLGy0ggWyXAdsAbGlPU1AaMMsQ13
hQY9f5A7VX2gqL7S8mWTR7SFttsU87axmAw/hm9bf1vgtSnzaO8vywdCeS2YW9pW
a+7B5pHpZAkzAcQFWh6fQcCoTorIk+QmSkeGbHymw8oidqAm/EVIdODH/rU9hu+F
Ss2alaa0H2/l1FmCthbtPy86FQTNof8oTN9tGK22JvbuAT4VTndlkfpqRH2VwujJ
3wIBGpDzPYRbqqwqAUireXEsXdM7VJGN2EcbBGRa/2PEwzvkueai9Mu6qs4JJKae
t+K2+5PXRD/YsEpGljFZyMFn+HbwADgJGgw5Ez7ziN20z1Br8+sS5lAswIwe1M0C
MtyA6KaLZqdag7s+cJGQdt+83xDruQaJ7oLbMYQ26VMgnpYFU5dFrHSbIQ+Yk5na
F5XiK9IkPPGMkIIXZvmvGv1gA8KmUibUTbpkB90va14ENSg1ZXskzGKdUcocTskj
5SDqpsTLX84WsAC374T37ZlMMEEfHIi1tPEZJDIX8z2Q3b2ngxbtumCAIUQ/vyZS
7SsZOx8imbrNne93zwhQJe8lhVHScyIaRHfomdCvr6sTxdHOIbl/JJp9gMlI6AvM
V76tYNKZVWEGmqbQg3F3IT0OQ8m8u0ms9O8ydr1gw/Axgy5bRCpJd9Zpqb1vzP2s
CFXRo5xrekYcEKxQKEAt+tZL/gp7cyT691LVXkiolbDlZuwFKnMzPIT41dJGXU9y
AYqPpaSSXWGKOsFJzRcmvWZ3Ze3srFs72BVJxogfoxU50ZFZieIQYiMQtHqQfm8B
1jWznYOP7ItUgp1fKVjIeBNG6M8ZZ8A5Mirv7P/saVwSSR+mAWMbiDhOD+9noLpC
3J5Wv6zFah1xjWfnkXhcCafOpCaQukQPg8DUjIDv5FyErF/PIRY1C+9kS7hC3p/C
zGBaMBrSV8Ohnm57EtFHohR9/PdgGQ7Fjcnus0AeSHtAWAFzjh3yMiBhjF2NuWq5
Z450XOFzWNFUEFuSG++uAlBfUkqtC0SfDUJaixQ655KQyAI/1iVvafbbTI+p4rRb
KP8hDMwTz3YQbFvqTtjkm/AvnV0R+RxJAyVLNc+iZe07Ndqi+hIc880cPyMFSZIY
D3kSMQMA93Kw5shc0b4Ne9IwtQdtTsTnMo+4W7MUb0WKzI8jukgrIKpU86DyQ4JV
eVw2xOlyx/uswCIEYXDhd4BPyh8gRdXHKq4w+F4NbGuMuWfvomu+TgtmtMnxECR5
Js4BuGBwDiwtGzwbU3Tr8peYqPAIyPfUEA9PBV8hy/5n4hRCr+MWHHC9vgmGTMyy
y0J4YehGoqPvqvaSNCP6slRfFY2CNfYzBBmph/mG7Btthwg//YWgvmLLMCMFRSzA
wwSxzzmvGcsN6BSBsYi3Z22X7lfW4wSJ2JEFJgd08Cd+A5PpDwRtgu++ZkalRYfC
Iz6CGH7Fs+ImZWOXqXPx2ObTJUkAB82tlUqgcOWfwXGCkEZF00iDGaP6yj/0FV/V
gb7EztHehSnZI3ofVrgU1ULok0WCuff0m9PEwttbB6TEkwv/eRjtRnY+Ng+7NMBs
YXIlNX2XtsWME4kRuim64ZPs4/OJzeGktNuHZZq2GqXIXlapWxrDOoHBNaOiaTBd
JTj6rrzaDDgMpjok+HxNOsvDhczuKlqHxlznWjl9wEIm6r6FZ93hQi9UeJ+GnQYI
o05liQUaV0pz1t7F59pAOHgJRpTv+RotI+NvN0emGQoV8g+6fnkiF7ZJoZsOuofI
FDJierN9CKhAgeJB7vqgtTDtHLDgcqyIjec16cC9I2aUl66R/ST7DJxCpCRz7hi+
/a71s3t2z/msWEA6LTHU8TTIH1/ciRVBRwNqvfwm8kyDMBCVkofNe07JirZOedTa
IWPl71fGxH6XkAMk0KslPeUmTr+bNnuyVxTHDG+bzwrrliQkM9SsOmbfJ+H6Liw4
2OjewLcW5OlXU+Ih5CAmSTKQbERZN0stx5KVa6wKCAF8PwWo4AFPIDwtwDJRZtXr
8h1ALiA8Rdxjjt1nSbKz2+TrqSZLuO6z0jsrwHtN02oQfLlYgiTpYSShvyIsywJ3
I1ftNWZ6PpzarEWsZy8VbbktOw/J2iieAJ7C7uLYMQaiT0K5Y5BUsWx7mK3KXEj4
NmIyP6vts9EE0cBrb/YXSFW+kQfAbcAuIpyzS+iWTP+NV9T9B8fl9RalaWI2b+vd
EcrghXe24L7tND/e9FUjugSDoR0iOfrVppgHmbYEJMZKp3NSS+Sh+8IZqZ7OFu7D
uqrEmaOFlZiCMqe2x1hlqisgxPtoWswkxnP5DBQCW3+oCRHeKn8rbkCItRSb12er
n6ujHBY715Ai5SuqkXZtUJ6jSc/ZX97+fegPcWYoTcUA6Jgjk8WOaxpCntsULZWs
UzvZM2LnphitkcM7AUq1GPQR2nCnGQnaiFuHNdkejNsxXZvNIXIaf2q/TPdDPZV8
30ewyFSdTRKg1Ij74LVkxU6AMajYxg1vKnwi8TH0CNAqEZKf5xzevlrL0OfyQW3i
JO8ObYQVfC/3De3JwtIDk/JmYkw9IB9Ep9cdG0NKNv61jmYhwtRtrkfRkUWMwbef
cJ9axPF4CKusIO7HE8PNAdFZd8Ukhlb61Dbb4N5qFRgVooYozQAfI5MgnHwp4743
4FxzD3AsozEMVSMIahWJ+nKBLBlELo6SAGNBFY8ZkSXHZHYt1FePDGUZJyf1uRhp
BhBfU/Gxen4+nmOcMQ5VBLaqvm3e2vycZ/JNvElvxRSaVKHLQ9Edl2z8/obJ+x0o
P9TbE8jVeAIAjh8D35m4ijb7oeSdt650KI/G9FnnZ2NTmLCtyPDwX0DTnB1hpl4e
PAYTDr48BvAtkauhO6fHLzeYgsonhOr0bQxRTc6OeOEDyMP1FUTQ+QOYFcguhPRT
SAfMnv/YAdd7aKOnCn9KRaRIcyqMMTKUxg06y2LVArwaMEY6oIvJ4TtUSMjXKdzX
hE3eXYV2OcH5RGkLCjN3bEbpmARJ6mRZwf8beD61Dn9B1Q4n60R1xT4JVa86TKcM
++kr8he2eMOe8XDGn3PirigHLAIet/yqVJItYrgzZNngCu68CF7Q88FJKxyL01vJ
rTMsZIBDQ/VeLLp9K1RTtPr8ermciF574tz1Yt/xnKSvW7+f48KIPXzuUecCLwoq
kZ/mWGIdZ46rx/6POHl7O1ND2Lh4b7kLSxa6+sGdTJefdDC4fgHH87WpfnpFDfqV
gglK94+nAwr/pm3nVkA18k6W+h6yEHAEOy/dI6juHUewcGn8Vmlk2T9g0aUg0P2p
tSn3lecdZHSqq5bB9tcu9Uy/7WukNxBlt/4bFryYNu+FX2t5r0sZT+tFPSnOpdTt
+WM8pCjz8bRYI5/6kW2xyKMFseAxbYZRMifi2ags8niSGHWXAZTw634yiMvqO1qc
gig+s2RdNXNHETigJXTElAIBATEriToAhMNvFxrTuEdt+LlKkueMGkDzZcw6DqPd
s1zgA9dlD3eOqAbpmPo94HKv1yyN8DPG/gQ0qleUk0bBgoDnLoNhe76PawGK+cpE
1Ay5Y6TNxdYt8hJ3FPMEqx1z7CbkH39F4YDAhLzhndM6cOd5q5IC6FF6zclrr4YO
4wVf9E3w+IvLFwzfYmIw8EHlDpL+U7yHphqrQGnK4BpRYpWC3wrQi2R7uS36BfED
/l0zRPwQuT/ay569LmB78MGG7wmjtwUQHfb1depOmCdKv0rOE2WIhx8FBNufzj0S
I8LJgLqzwRgVVnZsZ4zW0Uk59Y5NmIzFVuj226jPmfNIUJnd+N/TNPPTOTi14UJr
p/ap0VyDjipGjxKTknvselv9tK4mQK+0sIcGUzKXBqD82Wzr/bjKhixsk8Nx4tyI
Fqu2VRiUy5PAV9Ug6epbt8ARZMjrJO8aTTHdbbnCvTqIZGtiIbKNTpQuUW8x6fUf
CHbkjYPUSTTWukblPcRNBghPfUGy9enu/4asRjM80xM81+OiNeFmV5vOcU0XpMX3
Yw9CrTCvjRFYULzm3UwjDjyqwiqTjLmFAu57tPwUMxOS5QBf1B8R8ZAMiuI2PveU
1H5+USwfVtIPXkBHvuTrh/sPzSfj3EPmnIU2dUP9/V78rPyGCcpSSA71xN95PuOT
rfuuGJX3vG8MBNlIJ7VYNuMt/Bdc93YfIsY5xfkbhgvi8h/y9qdfsuT/9oTFgUvx
wDZSalf/asoDLO010KqOyMBQqB/HamNOkyFBGyKFFweWtlsEHGqJpmvWYXrfMewt
uKbxtd+j0H2eXiXYjTqwv8QiEN1/TRW4PjZWZogvSr2S4XSoxA+GHeBvvDt6TtT+
4598ZSdRcM6cMgWgijMIGNxzLw9E19J/hp45KHUnN5csL48W6Rva/DS+BRaGv3HX
7gJzg407wToSUJh6sf3oJW12y1nlPi7/xwHUzllLTerpbaMmrxFk1eMjsx8Vu+bp
jM7uYPqHUikmgQWb6vKVUQjQRSgUN95mbA323U7M2UU8Cr1xFmmIBcxdQcgmmH5u
IccA+YMYHvuA74O8FI6nT09b0F70uMNvP5SERCB1bRAW0laGx3SQLkyOcjuAFR/L
uZe+Uj0mMdj6MKjoyiB7o/cjlsvtxZWruRlNQCV6OoQfq2EzDpU8eMnV9WmnKDLT
iOfM6Y4sYRczj1uk3277xy1Y44MPW1mUhMA4zsUAY8yob2H4xz0xXxAbIziyWyej
gHJW7TuimmB7MvfTdKRLi8a6XSPTMi5kC3ffs9ZUeSPLNkS27XFgwG/j02yPXGTD
E7XmgHj/KOQvISvcQje2HL/2JE9xAG7uywMCFIREVjpRS58h0jM7to0fqrxKN+bJ
DIUKlLmHk48DWHIJBaQ2haMRv0QW5ScrL+X/jaMV4AXPFfMjQX9kQSqHu3jgHW6R
eo3cFzRuAQPSvnwzlBjTCK4IQKz1KdC3/9XEXsfqVV+xI/2c5eOAOcADto4kOEEo
ZleoA70c1OInLOCe7tw44aWJwLGOuI4GShSFyyYfB1/VxSX5vYiWkk/rnhhMAWJ5
eDTvuc37cf76dfAcN5SHIqEpIXicKtAz5ygemULdPg39FevvXM11jEqzyYjpWXEM
ZZwWnx9shf0cdB5lK0yr/MTXj3GLbtU7bX1EebnKN2sQmvv0T9Za+Doc302pDezb
5yKM4TSeosz1NO9ZrAZuGTrPtonzq7F+GTNBxpGgtig9fo2qJx8L83e8vQoxEXf0
jxn/kaakHF5b/seLA3ZwbtD+RLl2mm3cSnAvQLLiCWshBbUMCetmPP28wbOPQbkx
AvstLlMZicxFC9a0lf+QJYjP8iMx6ickKFwuuHJ9mUhP05H4yhpthFqn9C8gE3lI
G4zPqmjrC4soK0GV01pMWfpp5KhTDdFuoON1Qkx2Y8LuBKgfAaCmvAmbYakdLhuU
wwj+dc1tl1f4TVHfp3KDVuEKU3ihd6+jQyL6G1TqtXCQASgkKLkXp+WX8nzA+yOG
/y4fJ8S/g/tYb4Mk+7OovRaj6FWNsifdbahhBn68mfPR5jre0P+LXwDQJyaqmf6x
NtDAzu+lNIwRb/9KySItM/hycKWfV5ED3gke72x/EBq0g7jWtl2hE4q6fLU9pfjj
kyqZsEd2ywTO/3Bp4jd3N+vdvZfW8folYkXUgQQTjKrMakq+aHHwYVFLY9EmCLGP
RIKKIwOpMGaJys/9KCSjIV7Rt3jV+Fl7PalcPgkF+c+5R/DyQdQ4YNc0lDIQRqn2
VW0hp3PE5gwapIQoUo02EYsuu98yzayO55GWChzQcSVOs1ekgYyCLTRm0y4J1288
8YIYQnN8kPXuNiB1q04F4uDZ1lBEZAW90G9ME4D7WhCSBfG/QwGOAcV0lpuKKIS2
AIKeae2LiSzLIv7nS13IQHLQ6HX0nlRceKjZl7lJYquhQf963lCtX/LtzWzxKPGj
iCaYQ+31IqHD38tzVC/t3Qz0qBBbiAIDAHDEd1sBG4+GSEiZM8UPSt6yzCfKKXP6
P6GPFfdYlT/IxueOo7X59+XecDF70cY6Pw40v0hlzczzqpInBkEB8UMhQ/Q9Pkg/
GayEbf8bSBc2tDoHKwO6MrRQNWhFLmqZOma1VFvCcjViZNy1EgqS+y5969/yTePM
Omoc88JCW6573joGf/Vzl5Dr//4UMpNgPF5k1KU/9syYza+X5GC6Hg1IKfBsp/Bx
MEhLcM0bHxQ0cjnO2p+EhHtC8IMasvAmxsQdYAIrVsCsnlSuRimh3EC5FwYjwNy2
pGP/wz+OQoSHQKr8suWJXRE7UYronjl+Euihiz1oMhpcZCYOeVNOA26jsJYR8fDx
AwSkECAUa2AgKj7YFmJUvMM6ybhItc23xS/PJ2NRaLL9CQaD4p45QpG8HjtAz290
kB1gC7gLoKbKqABlqhNE9xoyyPtxDq65QQVlGoJUpOeVR9uTkkw1xx0kGYLIywvA
u+PbGrdIaTWQGTx7ZfSDAJYc27JP18zPb5T4ItGmj3G3i0+NJJKpbnB0YYiNVijg
M1f30lYqy83PY91SO6t78IYBg5JRFl5ZLu9LRDWo1Eb5IUKkkytzNtnl+693mxXS
PZ+kW4h8xKNjku/3jXyEm/zF+vbw5dW9o/iw4G7a/odBk0RHNv2acAC3Q3eAO3uV
3Bw9xRm8Emzn8f3mx/4zSBCzil+C2aZwg12ACMTFA0f4grImvT+9S39Go20jFAVu
j3B037RkMxaOYQmORNxpBQ==
`protect END_PROTECTED
