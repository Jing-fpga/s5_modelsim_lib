`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xq+0B1L2LglfWtn67T8QnSqBoYUDWjIcBu9AzpPxlqpoTt7AqdLnPRTZi84qsf0M
w1fd/iiBs0iRVeTFJ2l9RaTXaFnvVxbrmCHzoT8cqzpwUkTKk7C8vhEows7Aryw/
gmjpHRQUTqprf0v8UOFghAO254k4IHepE+5Owar57E+w2UMVVq1513IdOH08EBLX
yzwuvb+IlXdKCwZ2QFrQjrKJtWfwE+1Wbnde2g7DxWJi+UF6n2bNfZ2/vdB4moyN
MZsv5k4U0X/0PyzpuXs99qyRTxSQ+ynT0tleZ5kgpVNyWqVMHJAWr41Zdvfe4GJf
q+2i4l51sDN9cr2zWpQEvzM5xvMYFoe15XX8degMwA8w4y3S5H2Baf8/eiRZmbtE
JAnPtAK820R4dtKqx4eC42PrBP+Zb/R56hiZI9soXJxXARVrE37I5LQ6uPBpfRdx
3lT7Y80q/bZXtfhOLpL8h+h9nH7aI/hHCLNb7o7y0WomTSPl4DYxARUWmiNP1C9V
y037fgmE3jObUiogyAOn22G/E2uyMp9W0j5i5WETwDh8qIRM2q6gNYHZfCEDBJGy
Khc1AxklxfbKJdwdAo0QehOoFyvfciWA/o5W9WDm4MAve8obHN+jRJJA7cpxWoc2
17BeE74c2uq1wjbn5Q/oQ2WDYRzOa/wxpFb+3JvjAhIzSGPXG43moH55ZAWsqhFr
mlfsVEJ9TyMlZIMl1Zm/nZY9r5GH+I/01QBSRgp0QwJYqOZtCd0IKsc+Cn4w2vsn
Q2mNDbE1lMOQ/7UQu89oWlI6rNewrGY4Fc9+csjbU33Z7Q7WUHo2pH1mCMyI/DiL
lHO716A6gv8e0gn3mY8bAgQGKSgmY+vqi4Zu2XUpkyTBz1u5TFnNX2yWfF5rXKa5
`protect END_PROTECTED
