`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C5Vc39dsKtYCCki2uLk/7POAm6BxAIaGTj9QmVpTHV2PAZZiy2VpZpPLopYa7WUJ
s65eLufJb9u0XTsd0m2wcVA9hCPlYeJ64qeIHY4gRu2QgpnIrcMjjv0DAUw5EfxD
FWYRqv86dbl2/OS+0eK278Jx+PXIkmA+k1YEvmJuFCJw0ju8+luSO/gdEtvcDR5D
PceEl9qkAqlmSjqqkHDeCWOLhWbXy2ONquVhIVCyNKZjp06bZPvenub4LzapXDye
30zoKWrDTh8GZFbsGuXwU4EmIjOfMKAcHfJesWri4cD0xK8tQK64jwBuy6Vuxfod
o9GsReGBWjU8kLh33jvwgxPOqcxuR6uQcqMCayVE26vtSpGJowEH8X0gQaZkrNg/
7PmouIKhMhvn0686rznkLYIbr+453TDe7pPSYmfHoyGvHEqYtOkkWU3ucSsRmejF
p/h7rxfx0MXsNV1WhLFcqtJJMdnb61GrVuMlTaZfI+1n52st5sc6ZS5sIfvRJNCp
lMfxZkjqHLOt7blH7xJF+J3+wwhaGwnsnjVW1JHmFpigtQ9w/vcslsQQbSY9TktV
zmvVtYU1sBNPOoEfILzCI2Sp7SEy44C6/mYIlFWgrl6J6EhfuzfnJDtFmUcNuU3z
PLYidZnVpliVBQbCQvbCOu13G7GOk9y+R2I0XXWCWZdsnduhKiCWrjv+pvm0IZ4y
av4tfyzTiDWqtUWpkuBRPlSA2etrLdf7oIbXt5rWlpJ0QhYQdvt8o6xxqrNRHn4x
UxBwBizFZQaRS98VmUwIhp0vcg6cuzsjZTy03qmFxtDgBZeHeULxyo6NSk/AcQ0c
f74IU5IhlV3utqSrBQrG0xsUT2+12OAaklD6h7SzgyuHitxJU3p9Dt16jgDfg+mB
4aNckFt5WH33PN5XlsJWKMdBOcqfCC+OV/6k61JeDbel+4wkToMsW45/w1CCkxs9
ob9HshBaimuB24zfjAR63sk22sMDe//aJHP6YVS5b/wklBR4qquWIJy+henVsjR4
Gz1AIeiX4OsOgv9rlsFDE/ttDvU+EJA39n4WxY37Lc0kyMIslYV12Wb5VtJT42GC
GZxaG4TvgSxqkI6ZPTILsFCP9jbbj3CKOw8NcoTIG4CpJRm/k8lumQVSm7Mrcj2D
lK91p25B4wMyM+E7LKNPO0c5WtwS+fXU9Zzh4GZsidToY7qvn+QFY0asMgikAgVD
3ACu/7dO2yV/46Wy6kcqvDCRN65aUMkqD0rYdC6XZE+vHMzX+aUMXslSTtR0OAbC
Fpg9IfZwkStyWi5Ue5WLVn0eVA5aRiTFTV6y3pmmcz8D4tiY3/Y0dr5IWp3utb64
AWMkYOZx08RwSNICzUm2sx98abeAEnSy4Nz8YEWdCx388jGau+b8HrdzDgjzX4vt
N76gNT6TlmHEyMG+RJ6SHNkL9gaBEJBC56h76TtwjScT7yZH7jLEmqjyEkDwCDzQ
81QQwXy4MJk688DDoZylq71xnPS284kpo9Rg5DuYx5EdK9ylBhslsjfqr9G8D/O7
RpHTVvktQTJMIrzOinUWhaT48mrVDP9D0Lt8GWp/BBmVf2I7lp99LfVgDxlV9Y+p
QA6HPdfd2uP0dhAbGAgXndj6IjDsOQFInbFt75CRLotrk9yq2ivZ89NLtlb/Tc6i
y+frSuQzm3JpPAgvdJpqDlRs6t0AabgUlln0jr7laHqAev+6/YDxI2+NCw6R9ufT
dX1ArHkPY2yDJlYiq4O07QRuH627Gl3F6WHMPRPvaC+rX0RBZliFQDaf8dN6SpOY
Bk97edlUr+qFnnHI8B6DaxBQOhLJ87DdgFJG61WTnm7I2hFoLxRFCsQilvBz8xH+
ob8K8DCjn9AjpclVhPVgWZy6qw7sC+gTnzPLqRIu0u7Q8/Q9qXa95E+s5K6x5Sv6
irqJvf0r7HG57lJAY7SbeQ==
`protect END_PROTECTED
