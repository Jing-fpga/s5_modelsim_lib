`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0xvQrSX57T+0b0Yp6jfJrGgSwH8A0ciLBshNpd5tM19gHLzWCNYtApCxTLSqa2oD
jRjl76zgH1aFvYw5FYYk0D1V/re++KzX84q/7dFAFNgBzJ4r+MCdyoKcXgm3quTm
M1bSeMrpziwB3PKx9aO+GaWZJdn94gqevYkbTDHykux8F6zJd9HWQWsrBoznTMQg
PyfdqfzVJazsIjNfFZHVxaPgTHJVyfsV5GX7A6bSoE1pQL6CH+2YUBKDm9yUyAVc
4QuG/jP/wqQAJvhim3SXFNRk2Xh0Hy2ER5566FspXbQgieUfWrtsMPRRFH8n4pRZ
z7mQYbGo7mLEmbPBp+4kEkvcgh2YxpCs7UAqiXhJJmDv08LkJ8skae34grnpNJkf
L+KlTaP2sW3G7atzotwwmM+hwfyIlbX/+sJGokRkzc3XoO7XaFcL/LzgwzkWzJMH
2UYdzlbb1y8jIfA0nypLDPeb/PlDHYEOE8ZUQqTQKu2/sVERlvzE+DWrOlIBXkXC
6iqRkS/6/BBPUDfeJKAqDgVGn3QY6+Kz7A3AmgW8yZFCTl0DrKboOXxshE6Re81I
cAR7Qa/QO9DqNzkIUuhV0wvRWozh2AjaCS9trKZoHENWiYO7/cJNgPfIuZEEsmCz
ETYY/AXdVagRekCkjcSZ+0F65hmDgnce6PAylaF6TDKpOlD2ta3uvgkAP087Qdy9
V1CpbjUDsDznnKrYFTHCjwwFvvQK3M6inaqw2C+FxNUbcWSPMIqtsvwiABDKrYlT
IDLZkCmB/HETA0AUgnJGrUhsGLIiTqu9+0EAffoj6ngU00E4IJYKf/3ZkXi49mOe
H3k1Ezz2YZscPR04w0aeZR3DAmnLssPU0EfFw2MDosJnME9vIp1KLNJNq6ouk1kG
dcJ+cV/FJ8kpha5FYPqcscv/JGaU2IS3Bc1dpUGjVaPhpMZZ8nOD7HfftvOKY8ne
2sjF5IkO1Tf7XnMDGXph19z32Cocz9XxAPMlIKf3FRJmDNbwNqmTigyp6YutM26s
W6itY8jtOEAJOgxAltgd9di1g0U6vO7P4wFkRzOBd5ZjhqU9R3eSwVCS1VKCTRj+
ZjBwUz5PHZcItkN2FsO+ctE3iwbpbl85PVtyeF9MhIh7pnhYZhpXcNoWjaGESh4J
4Qu2M6HdfhJskQWzIugMH5bp/hr1wYSuGjDHPWCPK3XpdhRrqLIJcL9F/jZYfVmK
0wsyYLr6FjZUywA2CwhvaJNmpALqjk/JMqYGl90kd0nidf+Z6KNHg7uTNiALS0QQ
kDl3Hv+RQZu7i0xMhP9ozHjkB/K87dMS/vKtqVrx6PEieIT1mmBvgVKBSichVpkI
zYl+VYrCH3bqIKL6NN5s+NQ97YNjpI9lZRG9HVV27t5rCTHbhQSLQhpzoP7uLgCa
1HhiXTOdtWt+tirgzq+kdRRj+LyTeeRW9e68o3RWuelLhZ3svy0OACQLsDDeDEPI
MO85WhS+ECQA1GOIFe5B0VRVOomspA+L1ouwUVjbDXoe/fH2MuAbMV3Hfb8oQ+Oe
+tl5RqJ4Syrns7hB3rmsgE55Uuf2s2TH2QF6sYZwGngrzDLbhAgqDgnvX9fTUpCd
CNlnVHgNJO8jP968DsHzCdzDCw1wICU7w09FMNjksZIMjf9o+aW7os592QvsKJOo
Z+olOaw2vQBHJyWPC2DfQWZJYq988F6lKxWh6NDw/6MIkuG6IRgDuRnxPVyvE1Jh
nrWtWhYHSMPMMYfS4k4yDHQB7M5LYyZHuX5P6DJIlhL/0PbO5NnK1AysuGcVonvB
iyZ444Xeqx772sDT+U0yXJ+GyyVtVX5uAoKU4TlqH0bwoBxzXgt8bpuHWGDx8Sb6
ho4b0lYnWM8JY/YDhmGHRx0/8PKfstB4v1qKfszqRbVYgub7qMimWlvFCa/5vIyh
kZe9zJu9C+OPg3bVqaij/c8Caj+WF9XqeRInyd2A4U7q0h/m7jSUcsNNsR2YJ2Jb
CXHl7GLZ3nECCofs5sDWmPm7si5FOIYCxkpoN4QkwYjnadJx3rBY6hLB1SV4pyQK
LG17Z+l5N4w9pzvY/GfGEy2AxI0N8t6BmC6BuBZ0jRlMLsKzMathSe7g4lJ/pkVr
a+f9Og9ijv6JNac4ReO8T0iIditCNMDK7lR7y2bGHgiKFy8he8OtSSg/j5l2iEiK
2ln4cyM9d/QAMjsUbrynLpUVhqVAawNzidfS6CEykLAFrYjP8f/LSHJBXBUUcZLD
14PDkRPML4MQx0TJh9STcZCqDOfP7TfQtO4k9TvtgNS5W2gbdGSsNNtyOyMl7AAc
`protect END_PROTECTED
