`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
60sL57o7Jmp4oOpfggt4jHI9Rhb51MZbnrkN2nitBtfwtIaTowTlJ+XlZmQfz2pK
yUaPQTy9uIiqcQS6PdMwuTbbQN9wkJ4CATlgF6ySy+d3R4X1G3F2JJGU46D2/P0U
cMmx1QDTJuJ5T+hwIW5NSvwdviB8bUbn7coJnE3wwIqq4iOceBjxYdkfcYMPFFlZ
Trhn8NeMrEJFRupB+L7rtjGOQWNQiI+H77MwaX1WdN6pxI3+8Kj2+UhhFoyHRJ4s
QX9S9cjLZmp5HpCZHfkOUr6737Y36lnUmAWrlttnBZ0GWiDo/Ce8Mihlg5Itz4F4
zlG4DR/BrmzNvmXZM/bR3iToLi0GuAaAjPl+9c0eR+e3x6lxMQil8mP2DdKyPZa/
R6mTzAKMVPRNL5Bd0OxY/4cdMbx5u8g8B0XU+JDVzkL/fMbWng4n9mM05Yc+glsr
mD+2rNOTmEitCN1ApEs0Yd/ncsB32C2Ouk44JeHxf6bMvdF4Cm5OkOKAWkeIJOCr
FN+e3YWxwm0u1IajZcKBLh86ecviZoWXcRDa8GPxApy/YTXrVKl+ktRx+Tcpofmi
GjXRVoJ+Mn7KHmwBmjoMTpUF/ugbNZwgFkbJU9zP3/44tWiBEkheu+IdoWRSlkPm
Cw1zzpGES3ris4FjtRFG26htgmSfMgzryNA03POg7GRT3E0Nblmq6XQ12ZZpOdAU
Sq+AFpVGG9ytvVSHpwjLCa4/Cz7lpkdT7z5ly3uVvcWisbtczcTL9Z2sjFtRH4ZP
hRg246BIcrPNyUjbJRoOOjcZRpfepjeGhMRc8PnR0Qf+ZfxTP1GEYAUZp3mGIRVU
a5CLHjh7vF3R9qQ89B3cammxvFc2zMUPqDp/vlLFzvTKnSj+f2pDnpmneCGoVSyR
xp0rwPNHYcvo7WqNys4ttK9dXZ8Ncc3wl4xu7IlOOHSXiVtBKw27YiXB9gdeQQ8t
/62SZLC5h7OxamMRjNn99oVPvLAfIdvI2h+X7Lo8T/DeYWqK+aRBZnTxFwC2x/6e
ux7ETuZbI5MYwA765mntsV27N54CGSR2u2pknA5CVDjgEXXiRC8eIY73jicnYT7e
2zybdu5R05WronDSNBJ7Os24pgQV4esNW8oAivutTZ8MszBj06DbHsVucU46mDv1
I9YpNmLjfUsBvt5syELtuPpIswqiTtNwPqQY567jae0VoqbWtUXjZELbsBF2+/UN
tNOY+5E+A/+7sb8Bw+CD4Qz6T4NWaDrNyxjN5+KUcgvcJOurNKdjJmrZicZ1l/Lg
uo4CZxVbA7PIfZ6rvmE7Kzry2Haj8WqfWo0SjxaJqJTGdP3n5XYCW59v4/uwglZO
YEIZrpn0AoNSF44vSE56arQ7wSe9qlBDuMF6puIKcZUP/O1tOd813Vcw7xLVZ1on
dBUMyqWzIf2m7yEfeSKX/itZe7V8jL2UmdAHHdqtP7EAyZ1hIexQpKuHOGCX2lzM
W2MYObtsxFSssTn5KeDbl7EYiA4rACxrwiI/OxEfy3yYeh0cXkpoBMuN0n8ULKWu
irpEqYQFToTJdLRfG7qSDg==
`protect END_PROTECTED
