`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MwTWjylKNAaPv/rSyx8eJvrMPHLkkX8RhdKpHPxjk0IhkIc2EpQNtAVpFhuvzYXT
IDcCSD8kWCRi76/OmeQxBB2ib3RKoV4X4ZGlugBkfrgi8qXXLKHTss2IzZWkNm9J
oUJi8hv3K14I9ppfksZyZaFQ4xiQz/7KY9PHq3OYG1iFf2DaHT1u7JXB3Gx+zOF2
SF/6KLY5FbmEY+YWe0ewlZ6jHZyF2uM1OcJHx4X3TjOdmSoYeBs3GhUUqxQP7Z++
+Y3lSt9jerdUD796dllWpzGcmcMHlKxubPkrUhjcDpFdnfkSOiQUBpkQDdqScjkR
V2Sl6QLnmTjmAUOi1yyDvgQRT89cKI8x5E8GehFqeF1zbK+Dvq8hTG3fF1rIZDGc
nyi18ud8pifrYHpKXsuAtKRvAF3xS+2iGsgZcSdUnfCwjxjbjq5wlLqk7L9bO5+U
H8f57TR9818fa9pDc+ScL+rpCQElXBb/vLbw/wUEjbGEUPCS/wQ0MdfJyWrK7erO
M9uLtWiVsuaY3Z5y/JzcPFX4yXbfMUAQ5evtknEC0V+eN11dSPzioLRzOTDTrP8q
+wEDLQw3KEd68/LR3vkJqoVrT6GUR6hOXtlfTtkv2tjtRbYBD7pXFtXJCYxzYU4a
HaAPNbwFYTook01NWrz/sbTCzGd2UEs3etJcUXyoXUxILOx6elPXQtUjq0tUiPY3
3A3RYOokaDGqYENaVbAOc3G9OBzow+7EMqHryUAw1GsTrOPAdDj5KT7f9r1pmH25
tRyr1drVPJ4jYfcWr8GYbYyzWwkvx7xMwbw+Eb2IpdnaXxGh2u7qJtHZYqDKrGYj
QAnIXbrwWU/KTYKK+KQbcY0rJRyBNjt4ydpfErL7tqKMrkNYqocpsmAr8OXYcA09
5/81AkNBFt3sifqMNnSv2y/Ns+txQi8n8h/v/DbKoGGMWCQUpOOBVUyrYRlN9wbI
CK2hVBjQJxTSsI36nA2EEkNndJjuQPDrmQ+GRon/6pX/svyuG2iWngRsvM4i+CRn
eNZToZIdWnqQoeYgObJL3u8x58srzOSBjhPs10V5kcmks1WvQlJGLkKihQFtIqCY
KGdKEB7H3ueN2qybMmljbmFOuncFvFlwpt2q7qtorqw6/vFg241dHa+tg72ePIqp
Gxzp4OHCC6cIG3ZlKi/VvYKcwxRD4KRw+NxgjVe30JmVPlCPdKnVCvtVQkkCtyfl
PI9Vx3n8N9s7b6dylWoB7QxeTcjM9vluRSPJsavPQWXpjtGXJFkbcoklQC6lwHm/
udUKpqjv20y7UzmQvPaZpURbXkvJBgibhuvGEM19yftVwuWJ1UtULPqtoPqLf8Y/
kycoQ8MdIaFxa/Ci2H9v26nhbtobSIojqYVs1fQOWUXFo5kek5yNhl0bWplsigUf
64kHkyAlRYaJbHg/+IYVraO81OqDt4Uc4slSvkZ84OGfEVsOL+/65ysyewOByBl3
28um3jvrSQLZfz3YNEzw2MpaEzfaYr4oOERT4xWy9NgMRY13ZUgUjfktQ6oyByg8
YfrlHdt7wtbqzz0v/rdVs6ucay/n7IxfdlenXk7bu/LOWnD6K/r8ziHQdvN9UJj/
9h01vEbwmDz1Y0LrTQhIbnsuDLyahhmtrirW1FLSphOFM/Q4wK5w0YZ1cIqUn8PQ
gFERozU7/z0nVkUtAKejUznTlLnGtPC3NFTBChu5YPfI4F3vB+kerjUAM1D3wCsn
hOnByAsClwN4ZTd4x0AXLths+DUgXAh8O0vSWHuihuaGp6Mq8QgvgnY5ktm99+xr
7FD6BjY2wntyNOF7AfRiZc7Oxx6W3eU6g9uQEBYJxe3Jc+eeeYR6pPfCoAS0d3TV
pOfWJIQaFKQ5TdE1BhnEC9HIrcGezm5PeV/eAv3pAl+x2fAh4dHGe4oF0CrhykHF
fNLxwUvHhttrP8bWzCMoiEoQoQmXEWjiIaX9Vd6ifoyCco2b6YgJQKOqMuTLZxzP
FGyicb/NgsroyHDeVt901NicOPN9Eh/rRmmgpzQRDyS9S75+VGoRldvUvyTr9nlI
Tl2i2qJY3UzUF3fz4/NIrol+NRdg5roopXFW1ZiRRKFTxlGrNFgEKU9H5yMIZrCR
OqiXSjWI2FF7QWZJwDuTNnz74UmVvJItd2lv8GiJBA1VzPeRqjSEEH8W7AWKTCL6
g+MjaQURe0rMIjybpu0gIeN0dLQppM6ldg4nyVA3OQ/BgKIM3x7pGHjCKpRCKhZ1
sfF6dCze7Arh0QnaVOjJUX3jVqzKNXCeWiUQn1ytAziuncpAa3a9Fvs70/sjJVH7
mF7yNDM08wRJqeGTc3V1khnB6RX4572LdNlyYdq9DTsP3DYy+zpk7FfBu3ElxPiW
U4nCwle8YtQgIcO3V+dS3lHtNtsV0iGufysdWuXd78o07QTrzJqYcbAwLUboTbjp
97GWT0V3v/M2FenMMspknBer6T5tILWReBKvkLoIm60LihFH00/ggWZSJDNMpPOL
v5vKM21doP1yAXaYVekcyipXyy/BSaC29XBSFCpBg50zAvcb1M3m/YFTqhtfJ0X8
2gvi86SR953I7ZG5ruQrKidXheU8wxfFxSo6tOnk4u9Rkef6M9MQWJA4uinESSDi
M3D7+eRPUuTEQesUvDMsDtpD1tCk6vlXTerxRqtMJ+eLLGuwDdvyNq2Raj+Q3Ly9
oS8McxBoj2uWVt/GUen6GlMjAjkHKe235dgymtJ2zHdCTzCBr3LMvddkRb0tHdEK
LJDIRMWczEv0LlchoH8UJiruFYrzFCH8WJ297OgfXmf7M4mX4uCViqO5s85nby+U
TSyCckJhYEs6lXQ1pFqNArKV6DZg1CUAqbsXBqkEd3JeBLk5pzvXBIPefxdBBbku
FjgkSTF+EOtasnagolqiRAhasAq9XW+aTEdk3XyeZQ1JcK2/tldlHuluvVmPsreA
fL62ZLRCCTUe+jkCaVWmX+H0eQoDnXuORQl8EXgj/6cbnLI9KltPgQ7HswFo/mLM
kJdgrzTDOE8uEByxkevV4eqX+g3HbmZuSzXQYbC0ZY9FnQXor/DJHJluFQznGKtz
vCajeFnGAiIwSn9eedYr9m/4bwIhA4oQ1cjZ1LA4u0hvdDOLU34wzBQjre3qjK7Q
AGM1Awxz+44zUXlNJ/qHzhvkSilUOqXsudrYY9U9C+eQt2sYQTAKuvpPC3WXpn39
btwajcIfAS1j7zWJXX3yHeSZZfGvZbojt7CG3qp4SLtVe+rsRImTRZKAF43r0fkm
yRxrQ6DARTca4nsNZ9i1e6J24m364tBIZdMOC91yFUFIWLuFFh5ROfj02QpnBMPI
s23HtJFH3UCA5l45JF7k7cViOnuvk4rjOwjUz05yxf8fqnSKLZQr/dInMr9+RUXN
dJlS8TwJtjY37g1LMRG4ArnAxwMONuNzQMMrFPR1+/O8qQfcePajlZgHW1sk1fDb
9Jjdlr9zxu66knJGPAfmFrrpXgHctjkoqOHLbMnDfVD/JZB7YqxaVzxXoTI+QFFC
wscaWTDSKtOZs9u3OXbPV38WrdO8ryiSs7pO+qWQvcbd1JtttbFeiMQMgmc660iB
irqwlAsD7xmr9LaejZBSIIWcaZPmhSiR3AOsbddFgZ18/Sa7Up/V3L1W0f7WE2sp
3BWyB2frl45JMQVJMcJVOZKXI+InZ+bWiBO7GBzNBAl5Ddi5yC6J85fcY3YIkO1w
DCPF1dkMbIplVpfHS3nRCo6CjdZn3duX3Xi2oaPl66fabg1vQwqMRu95Mh6Sru5X
Eg6JeIh0EaBAKJLSLh4icjWIOTyBOpdZ+1c1Kx6dpGO1QAe3PliX1dpqqLbzX0La
SfN8wcD0EzG0Ei03kg2bEC4KXWdO7IXcBi/YgHLwEyR9XnDvCizU5idcbM34ABOq
TnLaH/+2iGxmhwD7WmZ4ioYhqxjv8HAgqngDmuKplzdpUeThRyUkxOq+/SP+SaVF
9Nw7N0FogyJ0uIpH6169GTCDIPwYsBDn7ktc2oUJaAQ71+aOO5auyxX+pdoCLuC1
ZvkVyjlp6xHI4opoNIc+wF7xXgYlBBJwywhSvU34iE7emeqoJKGjNyGA+WNB2fYf
KrfaZwWisEtCvzYLmZF0moG0eLCmMin/yxr8hqO//9XXPw2J3KpWOKvV0sFG31lX
ew2ya5YTayG5GhPC7cqOh5CF3IaLRm5+ZZHs9tUV9ZDJ2nUWGj2qSj8vz0icI2OM
U05WPEviN8McvFxPJkUgYb5amUCnA3tTJAekHTU7Sgc2A0wn1PRwUhwCqTIVlg7C
BY60TZ/3jJ8L9FljRIkFv68IfSJOAQTHlOMYG3sTwREuKrYlz1M49p2vaT2uOX8m
sjdKsoeVcKwAgVxHqfOsGK6BVCukQK+YZjqEZauHg0k3TpjOujjyz6oCMawhgK3u
5NXzuNy1k5jjnUvdQTQ7NYObtVnHyDUvvW/TVh3FCg3OmPjf/9DWSxwSEBg8h3JL
oFOgY/asMg8yzVwJATzqSVakXzOOLF7KfD9LkkLV0Y/5smkHPFunsYlWwmOhexb1
pYlnaOT8/7+HggZvLX/pS9Pn6+rI7gD6gyToRDuNSAsmz2SEsGRgZfT94uUtKH6y
7yIOLR7DUukfpqNEn+/p2R/GrMG4Fbt7o7noZcesxyIjdkyJ/88a1gHd9ekGaLAa
pTN8efTPugjL71fU9X60DfylV3FP4UTn2HwQ3+Vq+tVaI+S9vd9L/OynrY2SLtny
z3McIzT1Hb+YRFpsno5FA6Ls/rLmx/dGwTRx5YkJFR5ybZWEFj+A4BJiKbx9F6jo
KkGJN5ZzvObbOfZrpiiAO5lJml3ga4bZeU5Jnqf+/uPM8/JaVkYBvFs5twwNhK9f
o1SHxa4484WWCIK+izEdJozrC78kUXYJQ7d17jC6yd5pnS1YV04cBPzDnXH8mRR6
W7mFfPlba5H06Xzq/9BU4caV5+AufPs0FXGFDj5gkA0MQK11kLvcyIP0Y7ZlqD4G
9AQYFWBF0mIMJtDk24CpADQLjrUQDlq175HZEpT/nkAxUAXxVyp5JIQMJYECJ4qc
+fuJKxnN9LsyN7ci1YOM2GWMVWjAiOVDotYBEiaFpfEI1ybJ++GAVh4bhOFcOfO1
HAe3eau4YUPCVPx4yS51h6TvFaVcwC0MsapJyVJp87vgj1nRUWLmKyGe8ABTOnIi
0fm4MA8Qwa1rH8pPNdcFdF2NW1dI9LmPvwSssxJqv6Swmz4afVz9YJ6r9QAfEPFD
sp/mznlXLOTDTW8S6NLFf6ND4+04Bc8Cw8AbdVG53NQctWJHw5afdQVYOhxA7xQc
lHp0VdIakqbwp6ilbWVO4h55U/qFV55GX9Zps/qaoXhnUfsf8GnMlFMZasxFOGUP
kmN0RA/KqazJCl8R8pPIkdYuc11MJ7Jyf6RK7RJGpUHWKJayHjIL4Ck5y/4h6/C5
86HpkLVdlzW8LNzcz1zeVSpHnDZOS6GGcoP2F0dSW4xYxnrxu0KzNW+R2sIgwM2I
HO0mxFsWanv556KUgbpvjjlVq6gh340612Nm58DIk140Ve7rkxDp6mr30rsHOUWE
X9bUfjtZqRpkGVdDKpu6WjJzI1Hg1IsNeOtD9PtLbTHeP2aFdzAV8tQdw0bXRz71
C7IpIrIJHczLsXxObFaVH2CDetrYF7SKEKIxCbAZPn0IFfvn9QhE51ma2Av/bVPt
L3XWjo3mTiF+qqgf0gq61kyyJ8q1Oq7MmpbwEyWD9eF89Jn8vC5IC5s4YlfkLWDU
EMvz5OP7apphtut7DR3a4OrRIEcg/F9jlfEtwBfRtjJLSTEAz2CBovh8POIfSfBD
eyC6xmiB4LkICgy1SbkkkT1QnFRPyylVQYfpAt/jTZzzY16ePFH4QgyhVi7CLwP6
cheqxOdQnoU2oeCJp2Llx9PEjpYWOBYmF7/0h+RIU9/NFPjYurdujiRsp+8OwYeE
6Zj8Uvnr6GjorbNpbHGA6oY+YwkAtr8cfy3IjGqPwAave9dxMlVW+obILCL4y9dr
RBiC5zt/ciikWf3FWWYFbHrKfMdqp3miAC6IRElOTfLhd/J80QWUBljeAqCPGAmT
/75H27ejw24qKBqLflh6MTE6qPqJeogdXwBvbQbloOqOvQuVUIGMrpOcmhJiC4Rq
e1rGtjNcSeOfpgZ+dzufmPEetswRgX1yGtfZhAvWkCyJTULzcs8Ek2bsv+mYStE9
eXLXPQtnaOQvekUSudvs600WVeQNZ3MYYvs8w05OxEQfQuHvy19fbo9Pa0L8ETRQ
X/V7p77EnpTtGyYc/XZ8XA9+Od81T8vUr/SiXJi3UMbzv207TFMz7fnf/ia87Qz8
UFAfkaa6Y8cztwftClmCKrkXQjFR+0dWUuwLQUQbMLHDB5YJbHjnmnOFUYcbQaOO
Eu7XPw+51qVdXriPXQ1I3xu6wYn5f0/bI7aC7GYhXY43aMpP+tG+r2MSoHQcwBHW
2XV+KDxsV/URu1umf4ApmwmfN37jxEiFTw9imSZO/KJk0zPG249D7n2PdCx6ikQk
OV2+PWboyv6B9xmg8EZ1Bh7llBGYX5w6w4bhnXA/twFy6h78Y9AnaAJXNpoaP6l7
lbbpwt8KHo9Fa2mdGRaIYipj8pcaGnYHzdCzA7l9/RlDcf1NKM9n+kkuu3DaUMtY
DyBIFSqmR928xT7YIlO8WTGybx0FN0aoO+9fQxZS0ee9CHsJ/gMCKMlxK9tV6cHd
WzpiSCg/B2sq3rNjQalrT+vB0sEjGQfnvpcZOl8GX/RNM31+2m5FpRit1raKJSCI
N1YHpLTaIt+dr864txl89qgDk5DevafwVyuknMVerFYGliZAoL/YzHZ+sPcmGD55
1A3hMNSiN+kMY3lwwU6+fa8v1H4oNpeA8/kumVVVyOM5P/dk0bTnRfzeW62ykdCn
CdQCBCviU5jSRtdPMifriAicEa78+xC3g3XNdziDR2TycWJWnlpi2nM6N1B3vrOI
945enQavx+5JFGVSBTOM0KK/Jj4oRoolIaPW0b2tt+e0LTtll2ISOKDglcjg3p2a
MPuNER9419oUqg7vEH3tzBFAUjFWPhRP0/KExOj02Q0igzcIMGF4B3tnrPLYwzDO
3b7lZZR8VOOMebICRF+4DVZwcWzvEHw646tuAa0VHuaY9O3V+F0slOlwatspW5cr
n3sm6Df92eZvx5KRRK6+k7Kzauvv9zLJ67/5oBcwajCxnU/p9tcABt53bbhc69L2
y6xZwmq7tKFewpGAG1xAy7kZezTQPHpIMZm3gwq854SiG3OCbYwtMv8HM1kJpS/8
NVjYsjjy+5tYRYn5LebBTwn7rurFB+ZP6TXNLR8Vv+Sv75k4FOCSAQqlsy4Ssw/2
cRa28BbyNHA1fh+9UdRyYDmifhutSBgwB3XeAh0Mt4WDUFgtYMdy//RSK6xTSzcC
tgdzmozD/958xlnPV4QJf7ZLRJYsRdrkJ/Bavuk5/nHsgBE0Y8AwR5O6bQojXCBq
oTp1I0ozosks7NaXHcIfFsAi4/RHvnn8iPiRW8XbACQw+d8nhmCqNaJEVruWADFW
hKpYo57dwJH8Mx0IqCIpz7hhOTWLF7Wdl+8xWFzkXYhXXFD6z6VKUuyAtO+IRUWC
aCQLA4fwX4kfXN23XWJXiIq/osJf3E3FydrxGGYFbhuDXnve8g0fzT5fF0dvkhaU
Q+d+/OGNIMgkOvzVhCHYlqxa67rG0EVr3JG0kiEwo2O5TZCnX450+JZb5Ydl7EuL
UkKsQJHiu94ohWPNzpjCOvcKfJETpZuFlPeBQWZDHvAS4S0YC2AginMWgFOj+RSo
QDWC1ytRx3g3oDaGXN2B+iDJzmq/8dWy8tIM9DGlQmb3nQyttAK13n288f9xue96
d/Oz8AHe1vhHBYPtknOlZLKs/ihcuZtXe3xgla2ISgP8b5Ocu8U9XGnD7DvnPZSk
VCNJtq3EKN3iLqOccaZzMV6VU9z567vn7BuR5m0powBwgUjUJWeE29JK2upWPrr2
qvkpTdCoZFAqQoonyXq9ZIHMvOgNdldFgV7DVWTFXjXgDYNJOzuaFvevlHufc6qs
DOv/5aj9i4PPSS/GEfw/Uz20rLEhQTDN/c4JQzPtYimHO5IMKrOXE79gPOxns7gG
o8HQXg21612S3vHFGQLVlMJkddzCL5jA0lWkrGAdsSnqX6gM9dFvS7dNT/9lImf4
FDoQ2cCnDjPqudFIrp6l0IyuVRsRhtvZBTnUdum4xADcAp1GiOBIHOKMzmMtQ/rx
wXCcf+5MhB6dLMvj+L1WmgbAhl6InxhGGvNYve9Sqp/yN0z4i4GKOAg9cxefxkrp
eMPWuFgLenH+Zkf0N7afe0iL6aqB7MnzQdHCDkaf6/4XLILyb1jU41AuZeaQIttn
q5Doa36TPcvGYhjASiU64v0UOCPniJgkH64NBOMTJMT0XeYlOlt7DOMY9ZsJQ+cl
gbrzUm02BfXNqXFMWo3RHInKhZ4zqniksmp/X23AjrypVuONB0YHfcsiZOekLiDL
DwD7AoRoAyOQmSKQC4gdP77nXpP0HevbRh0cyL50ObZUV8luxqtHzKdlj0uD49Uq
LxOXgPWeAQekRnLTg3/2gtcLmXI5Fhsb28kIrvSrwvfjoi5eaT8SdIIiIrrgcmZf
GvZJ1BcoSgl/l/8Zm8Jic3gK43niyUSzXZBuMV6SQ+vttae4/8gdZpHYR/yJ74vB
36ba45RdtBHrbcDSxfsrwLT5efGfYsOVaoqwrMnPFH6YJ9cjcTx2CFFjUg+T4ijN
G7fdj586Qk0DDOWKgpLVbctiVYX++onMk4rHr5RErnOsI81BqfUvLyv2iYBK0PdD
SC73FSH4+U+zauOfaRDOoob8hfcs24E4tiey3UV5hssNiOd92WKmJTDRJX71OY9a
4THofeQCsRHpaSU2o3aMvpm4c93Hpmv236y6LIs0b9k9ubkqARnIZv+OKS+5gGqO
yMfwvpDJFvjox/jKh/hpxTVG7Wh7UdU8nKAktLSJTZjTqm2fyxLprSs72FF1R2gJ
nV8my7dMQIqL9Bbko5cvAub/0fgI1OB9PBoDLuyNakkizPpGIzbe2bSTWZEvCsLe
kkiPSxxWmgY44oDIibeW6DY7ywPsFevosHSm5lcwetp+HV9Em/PLHD0IIYj7KY8V
BHwoEB63iRuWoXjDo+n+tLLZgjlH0oiQJrpFlCNJe0DO0RQwtwcHMTCIya/3IDtD
YQECGaOJ5qPyRiY+sZDpniB6Yr8XRGBMW3eIKxkng0dKtMPdREYKh6npftXv1EWO
LJw2hQb31Fxft+b2VgKlmEQjyBV9ciYY1Vm+EjjlDlQJEYkraSbtLPQpxrJBAgt4
IhK1LmbG2PsRWFCCtnQ4qH+n/+ZkpkLSIeyG2FksoaeAMfgcI9/F9o+P6NqQaDzF
zpmVSUZKExZgCxCBg/AgtNMrsYsfuePP6cIvqZFM8KzFqe00rGNut5AfjB+J3i7q
WaYICLxGgcykVGvT2uda4/YmtYpHv1xo7HaQUss0c1vH/3vX6Il5wu2xoiQYkA12
KvMVEDwkiHYZGvlphtyygMnt4gycsawySlaiokptMgcHqgnYE60fPy2cwjbeUnXe
e2LXw5aGZwVYTSJrDrdU6g+Q5KSrUZSuMr6ryzoTFuzoY9tlkcGmi5KAQJjo2VqY
UovY9oVyyqAoxVascfW2kjAWzUsEqd28uWOKz6GixcI=
`protect END_PROTECTED
