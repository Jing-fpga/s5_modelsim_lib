`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T5dIOQhH5TQEFooGtuNQvUxtXSnYk6WKbtWNdDTHn0Gajtf5uqyeo6MqIdj8YSPp
oBvohK7gFN7w/rbs1cqszpPKjMjqTtmgXmasKr3YDayy3C6oGAy7i4WD0MOh8itO
E6tLE6e437TJ/YsjMfawwATWXkFGNjCO8fGN6cpp6hSZpvKNsrgGtGmFG/+bTyhm
4H/oi2nASogSb2CMQ5pZybh5PB+zP3vHMGxeoBPFtocDtjxcHaAG9e+XuAEyWrqA
7GdlaCDXRH6fIexxn00QlDUsZB+AdervIYRpZurIv/IkIqsKXYH9BVK8Cy3lIEDn
RHRsDh5VCQTZ3FP5bSzuym3cY8vi+hGjocreIeiCRmUhvQL7qwWwTihvGIgoCTXE
MkNvsPTPk22ky8SC8DXWY9XGtkv9CSJNgMEuIUwGYgT49j/YVRQdqYzHVrCJRUnv
8HD4WMcKTuMJL95QLVJlHLGgDsnAZiMcsE3D1uh/YLu6KI9tUGjugWZ7kS48Av5B
qwglAVB8wPuC5F3R+xsx5V+PQP9OnNY47w1na91k4Vz19ytI/iHYtKd4xmhm5eQr
nq2PfkZRngheNAEZh5ry86dHXyNUWdPwtJBKfbB8XkD71a76lasGy4Yokl46swfj
zgWElrRdY7E3m1ci3N9BcpgXsDyQzsOs0eo10DnZlnaXtOR20TdS4uXPTj65RYib
Hp6w+gO6ic+scNuM2sCQ/XTLxORh7/EaUSMPGgSZaZiveUniuaDM56Vkh7y68l9o
2V3EoSvKV5tTUssWFnx4ZOdmjEPmYp75H2luJNpO/YVLCV0hIiX4LVCvpUcSNl1c
jhPudqd1CYU4M2h9C2jvV3wP7DGJRvQtmfRZHmHQuGzCR5Jusbmnm9VSsmkXP8gn
yg+GZJjRuQHVo/TL4tWXiRCeDM+dLPNnt36rlkBmVn/1uavXnASx51oir0ieY/CF
RfP3KXKYLElBpRNcZ/9MbDHgqnt16ufcTFS6AyFFkxJrmhgTK+B8c7k3rAmRZGua
74/XEWD5jAA2/7Ca/hnBN8JMXqP1gpIiLgM/rNH1Is45o6sYXYLjzf5bpyUdRpkl
nDMR7+tl+oGRcYvY8BNNNtLoLwRxEKryM5VnpVXo0dkW1ibiYmk9mgura6fu0HsY
jjRQqwq8adKs3/AYWZADdl2GcJjcyF4b2CzhFx8eJh+SU7ZTPDGw+c08SJzcRj2D
RrigllBF9RW/PAYB4TYqmJc8Dc2EdGwjGrT2woudkITeAdqEmEA6ZhwL++hKQvxn
CvdiTDUxtddKdFNDDockbnCu11ZLjbAwACtcHJ0eOaz+uVOUtIQPbRoQxuTf0PQr
9T0/gZA99cavuzbgz0QKuwmAau+3LEgB0Vvr/+d7/fRhpJcgxMe56n5rcfV3DqbX
`protect END_PROTECTED
