`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FvsmCOKveQlZD+gN6R7a/ncAzq6ngEzwX9k7hvEDDzX9SZJ/oKhutrIaPSPkur8t
y6yz8xY9EE3+OQp+BY+vwXdUK/dAX2bAi30s0fV8rAi67QVT3ZpL3w31Djv1E0zy
OGf2CNSUwek/1mrVWHV/3ckKp8ughmykgtYLKXT7edhJxmkaOj6ViCnAglaFN6lz
oI7VHt6RGShDrD/HKHzbTlBe+djxfzPiOlUKBmCRO1tQJ1XmHG6sI/lNQvH8ujy+
+JczXmuTljgPQyioUwjXNPNFx8X0nUQ8FRcdlB49+UWZTq1EJbzkQtxZPsnnAjLI
/FrL7ywpRTON/EzwyTIY5V0739tDTRdM92rtMYDKwHJhUG229DfMYcKZZEuFnjt4
VzwR1AT0xGXtIZ6XbL2IsZseDBVmZELG2O5Tul7DE0Khc8piHzSy7VbeIfN4i9lu
ATVwf9LsLHLc4h+FrhMHzOhstXS5G58HXy6a3/oByfqq0VdnNXao53CUOt5FiTPd
c/z/4Sqr3WbwDiblTjinofzcvn/AzWJYYecIWnSiXrVRLPoPhwXNBW0+CT7LGK35
sfmNAZZTCU6abw+0cWV7Aerx98F63y/GiimArCwtSPe40wsdIsQ0wZyHxALyPjiL
c2BeHXL9ILhUGW8w5Da8Nd2Zj/HOuDKb1PZ6cHO0+LwHW2vZadOfbD8IdMjfha5D
6bHteK9NpVhj+NODHy2ugPKde0Q+TAGWnhU34ZNZqERLG5HhCLOclcF2bG6oXTUz
RYgo7EVhtL022R3jsP6Ou9DY9Xa71PRb9AtobnoeXIYVreigkpZ899eQcg7QsQqq
tz7WyQe0/IEN8yZxpASiXeyVnRbf15hF9ugjXLKF5ZC1KOIeXXMijHU6paY+Z5ML
uHj+egXTLRcSBK3qHI5Ye43ej0T8ORKQd8cnp5sf5GLNSG0OqucAO2ZWtOF0nu7s
PF1iTMG56uPsFwiXJVRhuc0O2LJTGiY5JVj5wlZon9/WoYkiL5qx3QM6q0MVdaqN
Na39IDY5L8qymtOnaV3sUAwuEm298o8oNxpdmxQWopBY+py8KC7YXUAPgpce5et/
gwiv54iaywhPiInokmwN8D7WbudtgqO5scuuA4Lt5ap2tzr3uro2wP/O9AS5antE
G84O1szBUrBDFlvFnWllr2XrqSCKAMl+Cw98IEYtPZcbdwNCRowYL5lxeDRYzLfk
DzudmBAi7Lcun82lx2syWW+BCPav/DN1iB9FqSWy260XyMG5le/Jq6CvGX/LC/4z
HbqORXFdsYWZ/RMM1D4gcvsfDOHSzaF0mbPj/OCx25PXDPIiulzr6VyPJTHN59i2
v55ZJe6WUJM18UWM9uMsOF1niHPIPX4zQym0KDgNP2C14Ig9OX6hvOJHWEwnhwLb
VAJD3U6wy6cqq+SDTVNNmZ/9vP/iIgp4CymL5zKjtj267K4FfCW9iYIxV92PFrpU
8R5v5MSDQJ7Cwx2yxRMls2yoFgJsUw0kFQKJFzklTqDi8NJlx9hRWUdHX0LZfUJG
XFVlemx1qXNO4oCMjw229TtZYC8UO1JdYyXlyBzdO32jXBr3YpDDTgqdcsLCH5Tr
IgaWd44P+B5Tsde6/x+EhfBtFy3z5DgQN/XtSvmSno/5wHHMhJH5Pa/R6b0jlR6C
hx2dksWHlccGZdlEsqKpg9SIcMbYVkUApDg5w/7WTaHwCS9mnhsOWrfyV0mp3MFx
h5+dlDqvAPD0nx8O5EELN1phg46uRMi4NjJD+gWOCXpFx9aHZ4gCx3VQCM4Ypt88
TxPHUZhsNeZni8xMDgFmopG3Q/Z422EDSNYDkFybj7da63oMnJJSMwsHQNhdKZTx
9oZXxGn1d5wXqucF4gb6TJGziwod7DCDvE4eZ9B+1U0IbB/HfD/Kgz0E153eduB/
/YGnmRy1FdJpiY2NnZaV1s7QLiSkla43zvlG8ibQwzRKyvBymCRyxLtMHsV2exdz
sN2jFJXmnvNUBxjRGXwNq+Vpgb3/cv0I3WX1IREapG1WtJBs4s5PLUMOSCLx754c
EXnKJGz/D2TwuBmmOazzl+PWTfRuBuYeDItfU8D6SLby+1VrOgq2ba3gnN77sfQ9
6R8ZEKg9uE/tOXAT5bjOCoAcl9BVpw2i1yVNmGjgjkp+zgjSob7apAVTAiG4Z6SP
csIUFxUXpKmJ0IvFOiOOJEZBv1t9OZw/TksTuGCaCYAz/FlpKOgNLphNi5YjA9fi
TIFI+xNHTGKnonBGkGxGKzDU47GIhVAP0yL0Gu+GD1OBEYenLjyQqAQgQeEuZgl1
PQ92Y83bL2YEPWE8hEx2WsEI1MocWrCCuQJvhM4A9Mr/ucEcc8UHCW/Fd18/SoG9
a3DpX/S5wCyG+x90z3dPqGB/gAgCqyvt9upshGOQqk5RHfv5NpXdnDgRllbtDMiW
9TCGZGnZzF6iaoXqNYGJSqfp3CKYW2WaJjyzdHxGaKa8Ll6z606OjC7JZU0SNfjg
bV+flage3kIJy2IA5RZFOKYGzJHMXZBpzMctvkc5gJ+pVWie+Ns7VPJ9HKmY55Rx
xhW4y5XMWuMh90R3avwi0B86Qkyi9FNEjV3g+HsShLxAiUI+P2uM9pHq89QmwZbd
z+hH36ksBHnWKd0VvXpDvg==
`protect END_PROTECTED
