`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ILqAShc2HHmOObSfmR0g181mctld7zuUX/u/KSa9mTtieAU/YnbvyxEFljbWc0/d
aI4k8/u3b0nPceBe9VxeG+Qdao3dtOYMbLzqHwi9TeiQcEuapyYasmq4MH8uTnTN
0Jk8A0q97Kt9CnbKDUk7x+jYV8CWLHNbqJoT1FVXK7uSdmVv1cKrK9gV+VhduSbC
AIjuGiDPkmGOyZEvwDuyHu5BJLgmHiDcejL3OhWEIoFRiLaOQrfrnyrZJLFsAPCu
OSxu83Gp7DgbrBx+Du8fQ7t8DI1aNOBE1Vpnrw8/L47Z0KjBl2fgwwDpgtNOkKX6
KZzxKtP723Iw0mVYM3ZKcSGnC5nRzLbUhjLx1looL3kuWPn35+8ORxpUCrBt+idS
NIhJNfK6+4VlDLQJ+eTBkPyvhjXJrFPpHyNk4MI7MsIKx1ew215owux4RB96QJYL
CmkqT/bndkaT8xpk4HKsztBDskEf1a/fQQ6pWewkk953b3MNgMmshDkadfQojxp+
ZprXPglUCG/V/UTs5PEgLNYLTP6O5ezQZki3LPVxuUOogrRMKkXg2oqvOdvgAMvd
qkSuy6tkqIWN9OKtvoSGLjoVncChTKYizFmpRfGnZD/NtGqyEDlcZ0PRRT/G3zZn
eMywXipEcC5BCS5YZ1NnY2deegOf+bMJH2siwVvN7lvr1bGTraOf4ogEDj6rsYMy
jROyqF5+izgu+ruuQPnSxiywwRkSrX+nBacwZuyf/KSNJlVkf4ZD4wlIjxFOx+h2
DjTQWhcc3hRfgF42RK4F8kgwpjw2SXRcHA2DCAHZ5Cj5z8S8jqnfqljOdX8Q6fus
SpQ7SoOiozgY9zplhIU2VrUV7a2wK1qilBlqTsvpXf0KcEXrc4VpF+AX8BKYCGIL
ZD9BuvY/9qu9DOC6dFWg016iowPrdBEvKq99Osm/xBWVdAYi5ldT3resSCUnU2qp
sFML/XLQFRozmUjtpWC56G+Kx4xAO/Q/U2NgvAYgm40ocuvR2h4U55hWLLHKA+0Z
9C5xCHjA3lzEkaGa1Yt79YIPHFm3lBkBZQtPKivWXw+MPRlN2RB6IrBBGcC9fbnh
0QcIzIdAwN3Oj900cyeI18eGWwIE5Sv7tA2C9vJMlYl8HvjYHdja6ez4Sj/1nrNY
twYCyMJZKQpvG29B3paIfSCDUj7hNCLq2AKlgGLDX1WmmUEnaBhBHOgRZL4of4xm
n1ySMOGF8b9jZ4rQQ9KcMlrrYqsMpVMsikx8v+IsIUOwSi4sfMAeHLDN34+kwv7m
v4D1TvmZqRW9LjDpjorwglWJ/GTc0NXwDnM0tqhsJ7d4FdQ4iBu60j7e6NvfPstW
T3nBY9iZKyZO6mBdF9yrtdIghecn/YN4umsrafTV04e11Aw7H3iEQ0kBJZiNOKwh
QHYYXpQ5NkRHLldGCfQB3ic/25fjxPuLEThuDF7deJ30670t2bNvkCd9x4So5Pfk
zbnRZzzmBp4252xDxybBHFAcQ9vI++1CbEWFzbfcNBS0Fx+ZbMmKf2d3SHmZIlAd
NwE1Wre+q8uszGlXnsYe2Cz01VpaqgXURQc+zhew2L1Yop9YXDlQNCJhWgpJ+3KJ
6tZ3rjEvdbgAKKpMALLil7FR/k5QjKKZk4G2ABwolDk8o55V+/aRxzf4ixt9SZjr
1mWmKHKKVNiRAqbggWeejXZpXXb3uB5/3efOTWjAlHp43aUNu+F5e5qE7tSfFyD6
kAFHjVCNbMPH1INdHyB8PicLDjFWddbxf9HU0y7rHeRGivBpP2cIfz9l7A1+qGsd
1Fv7cBImdpInqCDmGzvhZNw72htyD46W3x2FjePDGt2SJa01FZjyT7AWsB/axOPF
fynrx3cglhlWD0XoY6YTo5mI1RSXbPycmxNBN6R0D0Q0smU0gaHCc6Gf0nIC0/KA
RCFA6b2+YOeS4YmuHkcwsvdCe/FkQ5PIGPc8rAIV8LqbiTqxihDvsugbGstPAkSI
/PWY9QPVJ1Q7hISWBU3kBEYHROowxnRebj/9s6V0ZLEB7wk3arCaPEWBlHq9FjUV
0PoEPC5U0K/RiS+YjtBJLnOyvBdLdfPX2ESBiOY/PwI5xOYWT2KW9SfNrZoQKqjA
157dEiyRawObSPfpgsbp/X8hBjmZdqd7VL9pveNyUqf/kDPZCQZ/Csiqbr7n+A04
TQFUqdYXLyl3faVCfdivHkkbe7Fq+RuH5kpbtXWbaxePI1ss5h/Vnn96n99Mq7T6
f76dqdl+3ATBpyb+BGjq59GD3KG9d8j/DQzSl+j7VAgJjkvGFBEjTfl04q4Ofn8S
3TNoUw42ZFP2eo9at09/BLkEw/zjzWKJKl+mo3g0UR/MA4+Wde2RRZOG4E7wFJJX
5Yn9fUulmIZBTrDuzqytnwO8YI9xk5bGwY+aRgWcryIB8Fw1WIRVU855DEhs0P8a
WbzsxZQckg+9P8WV+CzuMMugcrfuMdx5e3eyCD3VF1lTJ9Z2HJLkX7l09uClJiNC
7rvMxOrJqbFUCJzUAdNqPtNLw6oDy2qPMpVvhy3P/5wt6kjpFaEwfuNn3BT6UcRu
M24ei3eD53sRG3A4Yf51xYUP/dQ+MnxIF/1J/9pru4yPgbjNA3UQg8uJg3QkcIYW
QWZpALd2wgFytCQ+GInabagJVFrU+i6UiETNmA6NMJSNHTbb6ykoj7RriNdx7j4k
GZg9tyBJpyGcULzM9o3EjTSm0Q6K3D0hMUtbsahLLvULz1RQPWA1VEztnsibczm6
1j6G7rZx4WCmFHqEtgpPfYC3JplJwX/UzYBwrWgKy3q6TfDwKxEDHizbrPqNyKxj
J+FrbqMsVxxsqt2Xqoj2kecnh6/IaFpuAguTf1fsZufXE589th4kcaT49amYgq7W
CfNCkM6mJnXMA2Q/JKlvZQ1edvkbRJqBDFqsS+pd59OV2gbVutX51GMqSfsNvucb
FI1dTNz4cdaR93VU636McjVtmdfKfk1onr1H6/bJFgqraRbb1xnPcwPc6ac8L2HO
ExvVRpc/tFXWrF6QU5GVSXlSVwcFbsUF15IpX+Dzrm3sXLXGPmP2uEUIdVCCbW4I
4M9G0aR2C9VfuoSZSzg+RLFSAVAOjRdqJyDq7WrcEnyKU4mogmad87z6icROdliN
phPzLRGt/sqho9crlFLrBfAZwvUXed8uHKFdYVffiBbqzjeu6EL97xSz/YMB0XaG
nTcMCZpoHWyH4pe8oUWqvHc28MKWMJBhVTflJWBOT2nj3wwjilOyMdkVnnNKPWi5
DhjT9Evl7hHvecQgilrvF3qcixhEglmWLetb5f6HJo6t7l4pDBVi6SsuUrSFvNuv
As59HCMvVd5RzTXjsWFUpF0OSHH1v3ez1sYYHMiGE9pytOH7Z/kMdEOpmFm8x1y5
ONQ8hwuetpRUMuu4XFAgn5L7X64qd6cLVX3OSs17M0NZ3q0b2PX72wMThJV09o3A
Oh6ua8qseYXVmCN0xofbADBZG2bLs0n4LF8rnv9SF8kVe+k/TTDrU5JVgXoT65Ho
0EEzQPS8xO2tm5JCPtd7dnrN6L/hELuG/y7TrmXNEma4Wjbt7fmllKNsgHijcTG0
wpI21kSIfWzgguApZldYSNka8ZT+lT5gcHxUgeGArofABQTkqKiTbtql26GmCT4N
PNrynOW1gmZgFO6ZAoJCWPg3whqD2QAE/nuHogLUosvrzBK9GX784Kig0qRh79pC
Z76pyJFzeP1oDx7N5xjtaWcPXuMbCoF+K5lQozR8COnses2C9LqfjLKpGHk5mXMT
vUny0Wkvw8frEQIwsnefVZKWwWDGGjL+9puwmih6jHlLzTCla9uOfBPyXJXGRFcY
MxNrzakn3dpYUaF2oBoKNEQLkErPAZ1ZnIDKUbzQXBgJ9stSxTygvb3xBFGzMc8E
hhZyVcHgCej/toImSw5pmG3f9MOXPDvq+WO64zxqu/Au7u78dCLAZ9UbPHiSSfvv
Y8lclkv8fd7GgFkwSN52kcPSmbhQ+rkOUaT5tPjj0VQzZa9KZe9lIRRTMUqrCbT9
fJ67T/9+H6mXbASqP7wkb+tR7aZlNz1QvRfZDvt9iVEWszt/GtkGWCwWvaUDvukU
RkJGbfWYPlKNiRodSxCSRNRYuvUhrlwxykCFAxxjD9jGeEd+N+PESpNbk/tle2J9
4wSK650WRv3izyodsPXA9GDOErpq4YGrO/y1a4ebszL5orHYWr5kejEDh8Qi166S
jrqxIg1o29fcu0D98Bewd2YbqgnCXcSrtkUmCgxxdTXTyTSwN6keyHemApgmfIHX
/BZglpRjL2dAaZMuMLXKObhg/5d3fX5SORt3xljwROz26zK3IGvWLa7uk9KCr+iA
DkLBWXrbOQ3/cim1n/a6aMZCQjG9dhvlYWuMa/hD4gP0/lhyKjHOAZN8S25S/AaZ
QfgmKVPlcQm8v+IGrFS09SHq+sYoe7+liFnPIGbOYpTrwrt4uqLjcW3jMBmqaGyT
fJz5FrH5BnzXN0qYte3EsisveNr0ifwMDMAm1yQjcCoOGTTqfk5nyCyfJyjsUqs3
MHaSznf8xNG88j5p0jlSbWh403dwVkPGuWRsvumIsDX4fH8MJicbclD4ihwuvqip
N9BauQ0a+92dEg7h0Dka91SGt5fgFNJskoCEtH2bEeZwtYPZZ35YRelT0eyf5syo
lV0mxaVL8qevbCffZK2zFnmmaJta0SHNzGxgxYnprL365e4qSXrvevKWNBicRWq1
tToqU/hJwUHjuGPAdi2jqUdp+m+/Rqy0iwNhkeZ/6Y9P4y7jni6zfuch1sfJkXs1
Lx6OU6AfjijbCQBJ2JPctpj5g14axwEZEiuR1MkxD65uKmuJwqXK5Nht931rSmRh
PidzKFsE62zaXiEqFBuHNgatRiJ12+g0qMFUgDKCMzQliBzALNZHjhYjn/CBNPZ+
kOvk3mROK10kbDKVEeqOR2OhOi+h3Ndsfz577ywiDv+hkKOS6aT3ebSWT4issgGV
cbjBrdRkCKa/gXz6v3ZCR/tvsQJr0gV2+8u0geN/Xg0teGQIt8sRM1dLjE20JvUe
/RHHTFDvqmSEr24u3tkvOv5LOdh88144IUSQoJaAiFQaQ/ElfroWdQCJUl679GcR
pWUhf+9rvE9SCN4JXVX4lngq/mCPjJfDLJogdT1hqBmpwvnLevCLBTI3jBAs8PeF
fVSj7RATFjaQ6uP+JwWyTItQW0dE/eakijTeEOH/mHV9wTcm0RF150403s8cpG4R
U85BdibxaPzvxz2TOs5WDq0MsuXUV+kGAXUxiZpGszVPfCmR3ZLLGFKxgYDRQ/1k
D8MQLx8+mZUdtMQwGNkapXL7teHQV+EnB9vODiv5XcsLp/2i7pweSdCVgtbjEvHu
Hrcl6GWGK+o6Ri5/ShQTtdfdZMxobEepxlqBkE/t7CBUMDGmpi7SX2adcPtGN3ei
oWUn9KsFG0p59Py1a/FNfQ9v2CL4FgeKU2YNrmdU/BrdbEYLdYcd9Tmfy7krPdyC
jY38cHUj4frtyQDRJxKQEKsO7LD9D5rGBNbe5D3x2v9XC6bigBFeKI2cuVUa7ju7
r5AXgDjgRZynjsqLmV4pzEd9OYgU5o0yl2sQT/2ZDdY0Ro8uLVXM6+YRq0LxRy/y
w2ja7Qlw8fieiBj/do7XDoofvd5AFK+aienvZtUPCgcwGAP+1ZeD21poqlLl2fJ+
MKWsH0OrhbSu5uLFq6EOdXDdtGZQVh2hmUmbeFKkKIeZiV5pAiMteP5DNWsZr6qL
5bGbIGAEq9Mjf0dfrotP9W9Vnzq2p56NycY3G5uaAIiMT3dcJQ6oYiQALJFPfSHV
UalU6xHwSWfO12qEm2JtbQ6Jiyo9ZuRDpNWlyYU8QjZ6zUXPtHLHPoyUEsmwwHFE
8u4gsjI7ZM9zUWCOMO8l7bMW/4U5qTK0b4qJ+tlJSot9y+HViD+u6ZeVI3X6Te5j
BGjkdjr/7HkbMZreGVhZlycnrvS/iIM5XFJiPR5j/4QtMg7bCUNm958zns+0WqR/
S7FfNpWqQhzHdvX3Sn5vOpfLsy9Ub/agHadiSJ8itcUAhn1PFdfUYyHe36ufMmXX
QHyGM+zMOD6o3cdoB7fx9GhX8yJmeGo0eFN21J8LgSy9NrN8yguBUBrG2xQxsg4o
BFW3SdCTORBgPRh6j6+hqx1SJhJwXOo5+19ZPSBHlrnFAoCRIDV7Z0iE1f5s3Y74
wm+CgX1mGU6QC/CuYTWGwrdbidPFPqsQiP35oFmRNWnjba3Tndl5nEYopIv9lCDY
Rv8wGqtOZ3iQL2wQ7Vl75S/UGo6zwYkOaQl3ErsZ5by1u+ZwvpEQ6eXhFMxYfj5I
0Rw/mUcGTSvloxt1WAl8MkNDWSCRIBTOzzIH3cAiiA5T4vVzU5im+1IRCGfbjSQQ
2Xm+c3dadfEmcniqG6KL+y1y9lePycdb288XKTEErl2fEq5Znl88WtMjd7sZOXvO
9NpMIwXZE95I4AI90q+8AryqQpa2INRttOAho9B7y8dBQ5CqQxD1NsVqN5wWxERx
pO+06ENfxf6KPGXvl4aBBjB7UtorO/XmElP1YaaajEaj49P56xWJHKDQntWsqGVH
XWegyovaP0accLYHmX0yLa9dxfA4uaWpF0YDU0Ow0JpGlnxIwXZYDG5faSzW4q4f
p/3WmoAY6Ro8ZImgSr8fHq3YVUlO97wbn+1KGAmQYJFNthmGBBUvZDjVUSeztzh8
WYjYsH5FbG/jhkWph3LEZkiuI0eGQ2ffZDsopWDrvqB0VpqKrCpP4Eu+hJhJLS/N
Mqza5JAHqGHwb6bIptY6gRg8yVd5hdQJtPj1hyMBLfFjfwfPTglvhWZTW/3EDeV/
X66yWbTF9pS5nxKjYZi2Qm/uWvywq2RGARVO1junPtaJDMubd7m6Tue6RqvjpkQ/
fQU2KvyJVxgyWmulwuMMXWjoJIetVPXYxW8hxoEfGytJQZUeKysT6OScUaH72Igk
ht7WSkWK9eMPVAAkWcX3Gly1V3bowtdhU2R99xfFdmeOxwrSByeUR/XjraPvxthO
UB/5b/ivaShRglgxtMlza6Ps48KK8qP7x9HPLggRjNKtSTDT7XuTHDkdB37dK6zL
MnW1uXsmxgH6Fpo22lpUcN03xL5jRacCIAyh916lmLsagCRXpGAGSqBjqrEELuEy
cbxKn8cHMgHSbOqp9dvKVg5LhIxPPlZYYGhBva+P7JzdjcmXqLyeA2abFy8Rkubo
W2wDwnchb41CLs2vsO/wRARyovd8D9XBqlejpPlEKm2mDiy8C/8Uo4S+oqpGUTo/
1h+d0i0bHJnD4Knpp/LJu4NV+fagAuJgPFx5BibHTEBF3GiSts8MMXCbUYu0ecFN
CA+vWNUMXwDMMGq3dRnCNPADOzBHTszwTfpORrIDyh2B+8WCSPyD9f6Pryp9nIDr
XhgoGjOJHPN3LuU5fBP6c2z0rxLNhM2hBAw/3TAXMVDoCOIhe8DaFg4J/MrpYIuY
mEqsrqt/yiwbpvfNEvALpDON8j2bGyYGpwg0v3RAWWlOq1Fm3+Y/2JPvaPksnMyY
MWSSQLJW7FIDGWLzj96J1gn+XKmZwuVgNy/NeFYnJdg0H/UG+euLZo1DZ/jPHeep
a5B3DrMaddqpGz84QOkaSVzipNt6lDaTqjcDLcakn26ptVE456Bg5eQALexofEV9
kvtvGJHil5jNu2RaWetFU0CLyj8h01mHaHpU4YfRi60z03vpPbZ9R17ANT+JC2FX
cewSrzq0/eq72F8jfCHxwrYUdKnKPyyTJOti81f/Y9Ph7oX6E5fLbNMJhwJQB2NF
kSm5reDOU1oxe4L2j8ddvx9af4bnqNTjDv8UTpyDHy8kTlwIx/mtR8I2VwgT2CGL
kJMf5GDyDa1obMxfUnqvQKG1MJvuVk3HQgLfJzJskHO8NLMmTIAD23bECgB2cGVZ
owjK8Sb5KLDXjEerXcqT865rl8gzCIrLtXbD3l+CyyzH7/MUCDnc2JMjs0hp5UqZ
Se6oryIexUdhhd0aHhjPNbK5L826Lvfn8Aka89Poziu7CSPNVWlNSxbhUACaPVBN
VOceOkTGNsXOQSFff027RU1zSzUbd/63sIZE9GfkVknWBLbgzvirZY8NvRYCqvwO
rL1ieAG+txmQenByWPtM5lLhS5EwzDmTj5TMm/NICayIV4rSOc/CxwKqyyMum929
gA+/1/kmIRe+M1nyaZ1cl/IQHTlCG3Kap3vyXOBHSZ3A2vZ/CadOxIkVKK61XDqQ
tIo+y+FLg7yL3WoBWUbW/gdNdqaEToIFXe6OVPnE3ooXcoQc+2iDzKmN8FWeg1O9
cyos1QjpY0q3gEK0BjTWz3iaQ6g5V6E7r/j0cqCa8IeuAZ4+Rnty6FEy6o+e72jD
WdHv3NejsLqkLwZV3++0Be/KLraPxflhYMRbfJrXSt/Q1OSXRXbpj7tIIgK+stfN
ICIvcxwQdeQlI/TF9cM9MonwkqDT8XANUmWz+MkQKPqfIBgLucR2x9agl9JGHrzP
nwjR7jTdfCfwt4Q7+MkjUCW5YXxQGK8fakzdhEcw3R3NXJqCWU0l7irl5HhKMwsz
9q9/7kP5k8P2D0OJ+tXvdYnNlH1Q06L5C/SqCFW7nZ8so3DDkkSUIUC2F7KpQbnl
ft2qOm2c+JG3sB4icGR70kWW8FHjBrz85si4/eKf7iQT7t6q/UiGHe3fojfU0pcQ
M93T7JVIPmuNKoCmX6FzDkiv3YXVNoCNkeVhnjVAQ5CUSqEtNM/h+zy/r41TtqQx
p17B7gMU+eehnZnzgTlDtrJUmxADScPw+oFn+zTQ9bKWS3TtfQI3OG2eBqOYpQ5G
pmTs+XWSIqZK8DEeauJiMNKINN9B8on0Ts6hHaYEviI8t4sut2GENP/MNSzHCBLm
d3If3kTNX1ym4mNcptFvUU3h9UfbP6ya0pMiFkAC3D1kyBkqNnskmJSmly7psRZ9
x9x68rPf9FWoDJdCTCGGZuzcONFY4Y70T4Y7mSORkHv5XBecOlh0URGZBvQlQ2rh
jD2Rgb0joI/YMXnLy33+e5kYqVqKEo1ENzi2yNdVzmQMKthhze6jkMxOoFz76ch0
8mZB1MEe2S3eiVxq4W0iAGf+ZrfIadqOLdN4C4JODGYfxJDd0Yr6WGv4Qwecgav2
oBC3xrj4M6wz+xi4E3yk190gc7MvR1gp1ewNaA3vS1qRk5bvozvbcRMk57I+sLsy
pusxEHdZE5K9/43x8I7CAgWWWu3YXqZR0isNRbRUCsR4e1mOyXJQ2X687c6kWPdY
wAQq23oVbEawsOTSVNx8Lgr9InKx7uQ17Ysp+shDipxINXPN19X6Ozs5vQPnj24s
`protect END_PROTECTED
