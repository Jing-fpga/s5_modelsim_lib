`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mdJPEbnNAtojS4r3XI/c6tGWElZa55JXYBBFE9KVgarGv+f/FrzvupJ0+Phaz7V2
RFkFsKVHa2javgbvRr/kR7A/BJ0iA9eIhP9qqhrI53/Cb/UQ3Rw/N1I+W6vAyv9L
kQKGNboaHYI1NgK70Ev7F1lfGGqjowmfSm/ONm53jlFeopFpACbD2oQoIv576vmc
NJIxkPB+efnq2tFkCKJyqW90qOJumr2U99aADdn6vyteng0BJ2+yUnUcFKbEMjjR
BCKorRCokW49aS9gLefQYDNDifrSDG0rKM2dzQfpn9Zb/4bQ2bYOZ+f7oV9dRyqd
tnPh8vxTHpd3CSSUk1LqXZEbxJxcUOtSb0MSNA6iwApbHPw3Fornr48wUFPK27kz
eY/KV8JmGsdAXu0FgI1Ea1Dp2jMSWq+YSwARGgWjvz6QBgbONeuhX/IRJpyGLXWf
b/LsiRtCXyRSkLsG8PC+etqS5ITO04spxyOxKWaM4Tk=
`protect END_PROTECTED
