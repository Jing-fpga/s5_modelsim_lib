`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jJ1T5CJZyFpukJmkaOm882CPv1F9r5EqvTsZUycxZ9qHpTZFe9oxZBuY6lNKIBsy
Dv4OSKZHmCYeJ9f3Ym2Ox+SWMfDeLmKwlxKAbulj8oXt8+jfAbLN5s58U86z3Ct3
MLnZq0z7I2oMl9c3+0R/UTp+jB39m72XVU3arWgoDCFYrqawQibzmJE3wRvsK3rZ
9YAv2WxGN5cFRn/PXturovMYBqH6EtWY/DcRMjyx0bExjUSFBJEcNXpmqjC2PTMW
gWxSXF7oh/OUXvvPWywbGp76kWM+Sa4zErnPqikd5w6xCKEXR+sFOiK6cHqLxXZJ
LwRY69bNRvwFZ8h57S2eUehCZBAfYWIqLB3H2ZXBelCMrJ4j4+IAnMMCuQRF+K5j
kM7f3DnUGyfuaySaGK+vngatsIMYIBlXnVQannBichlv+g6bnt3z/MCEespMyD8g
ANv1vVGDspZGYR1ZjTTEmrx1FOhDNMs5x68M5HkKQWXSvmkFOFMdg40E9N0+3zPB
jN2JPFzl5mBaH0ndJagAo42ca7yrpdgzuhdn1qPD8jxeiFd1sOaLRNM60u7/OBy1
YwHNy1QQgOp1Xv/WE+5ZP56S3wfIb/2AqIWrcZsBos8aRQ8fyp20RHw2nBTB5nU5
0ROREo8ReESN3RDP5+ACeA3813mmxjTRLQXdMWleUSf6suU+Xf9/Em1+ZaXCUt2h
MpKLm7W0eozQsltKb1HZcGuN9eyfLzIojm6759PuDga5Fl1VWW4k8xknd+4MK1fk
CtNlaRWfKeV0ZwHxhxTO65V5Cjt8GXXeq+LZnivSRhZjzJrLBJ+A9tEaDVbYgYE6
ECVpLnJPzj5UUH9eRoUlNHOaIK76fRfIVv+i/NiUo2VcsZ0WcdayBekOf6GlIIUM
oNMLkFJFhNjb1/HIOZyWd+gwDWglmuOgbqBy6ykyhO6TjTWK8TR0Mp2szuw2dvPz
2OH6laZabOJVzSagKlxijxpqsTD+2iEllWebFchyZvspvUspQc3mDdiV8xw3QVOB
dagzrOx83ETc29siW5ZmD8TY5cVe6l4jwK+1Fqnq/vOgu7ql9lv5jTTlRYhJeTRe
SoyrukAMbWq2n7plwo9uowqPERFOwsuyn99zHwaQk+h49NUr93v6wlwcgdOM7MKi
tcxrdmCaW2HptS37b5foBJ9zE/hZLXlttgAkHCvwoR3GF6MJVwwd6m82fAbpL71/
FqEhpNPvxSpYdMfEqBMavPb8wm1MK8+S/U2PueojOo56uft14z3yI342ChZoiAhE
sSd+b5TAQtKuqylA3gdIVjj13zAqNgTkWwngcPzYEEQcee1Uy6z7eqzR4stOV+Mq
Vp5hB8XQ2BM+E5PPp59QzfHj8Q20TJ9ekJ2dYM57YXsBl2kbVBWVyhbpDBWCspfG
3DvOi1jjPzlb5iOIoR22HaDXBk5ztxXpMt7i6e8sbXOK1A1D+dXYfyeYYt9GGzul
xwPyg5/sjrytM7ePppQUJGhhsoroKS5nJ5Aq7j56J+0u0pOAcN/0UmoN/w2LUHJA
9glcZkxbkYsY60+t6RYwaIVqBEruRNcIV7oN0WgjIBZvYGrjZwm59aDygKgMP9XV
RFVqY/edOivuHIO1EGwdsLC8hYg4nthxlwKVSbyDPZiK1DJq0l6MkdxHO8D6xkVR
SgHeG20OPlVikyplZAy/nAwVbFRrqjAewqLoYazXkC4=
`protect END_PROTECTED
