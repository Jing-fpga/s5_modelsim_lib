`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lCXUUZoYqdyYxyW26qbbJBiyaCiSf6SJdjSKtdmCVpJjUX8fH45ywus7bdGOgEd6
pbcGevXt3FWvEyVJ6XNSRDJlgcq7Jo172cPHluSSgYzmqcLBjrFlj0AlFUj49kFd
qFvUrHZiFUajEYc4YyYnjMofMKQCj0ReXM8VgJ+EuguFHUzedFhJprLs/D09WvDI
jEKSSErdvq+dAT4j9s6/ebTp4JqTnLmUXB02mdmUUWbcpjpejoHlXsrtTb134Oz6
sPhnwwENYVPJSC5MAONhuATIK/Xe+Xylm28ah13ZbeDZANe+k14+A6o5j1tmzy6v
77t4/fHvIq9uwMc35mN6Z147tJlbUdTpsF2/zO04qeHdwwI0gNvjbyW2VFNmMLeB
GcE570fOjMA2S7jeqGLT92Mw9BFqx8Q0197cb2JPzDFRpg42g9EYhCV6gHwO9Ks0
7AGEXtqQH5KtxTP4ueBrZlFhDZixkHWKLc6y1RP5yi6N+6iBmEpESer2QlGm7gzO
EI0jC9tncCgqFGVDrNYyqF6kU4LNPl+nMC9+gwMKz+pshn/marrCFCwxtIBCTui0
rmOQyHwboFn/CCqOnAr7dyFSCAzkcohiKhQNqk3nBtKC5XoFCqvTPUxacUtTUgTm
ZgA52N6krOeHHdgD0Irmodth8P4AYrIr57nA74i2IX39XPEUtMhfQy6lXBf7TfN2
xZzInWvuVEMf7iB0B2RPaMeiSYTKeZ2FZOKS+Xmt2upjTFYanxkPqTs3O62M/4cz
rtZeRFsP740jMDnlUvBqWiSAMZymZKclK+ZyaluTkZYaY6zM2Z/GGbovDAbCBghp
BFVq8qTQ9MC17ACMrqr+ZnndEEtl/s6rY/IpXyFhV0xh6DX8jpFxoAedvbheq80d
3iNU6RpRPieq089nP2jsVzA59k1OxVUIMVBdpF7vCQfcSiJQakI6E9SGgMkG5Cw9
flmU3Ty/jMGXzFaN/s0SI6vsgSvugDNft1y5zkBNmjhA2URoYjakT3WvSM7vwxNZ
F8NcLPpAveyxOXWcuoxVwR5kCEAUZk9UIi3XXvrKI8DymnHn+S8yAGTecI+8J3n1
Ggspwp6Gf1ZRj6aBhPpOf6vLx1xiSPbbIjHk5j7zm4ZufYHPC01h+YV/ZsrZWzo1
EVEP7K/W/5r8INzDE5t3LDiM6+GtSGc5o5n7IFQ0gDTDFsE+MTyD2IT6nLuaR6jk
oF+bhTxeO/QBYyG7ntx2SuOic0gVDWmO07fc+OMBaa9yK6ZgMgvQpHnCMLqXJdNX
Hr9qo6HQGSDEwy6Gm1yqEqklO48dvT+5T3zhwSDfYKoFe4HjrMdFaKfFRwNGZAZn
yflsqq1qCl4qeuiniwWiiD1KMp95zc90v0d70OOwNI3xn0M7MTFfmIAPKtKrRP63
ykJ7+RhLApOLzhV+scjYXRUQtNYRs43vlOs5m+o6oRemq2wciqV2JpWa12UnenPI
btgL89GkvkE1maw6KYypmtMaPDwr0uqi+LwvIM6UvmlJkMAzVCERICZrHDlXBgub
TzLmqjdQqWU6Qtrvq1nUfX2V/CGp7cjeO9kSAe7sGocnngvwezqMykC2sKNjzgep
`protect END_PROTECTED
