`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nUvFQ1UZMHn3AeTGgiaMkdivtCdEKgcj1ixXc+Rp2juSt/xLOmvjlDoYob79gSZ6
wpK0Qcx7Np1GOsBn4dnh++57Q6cf1Ue5xIV6O8wcbasxXcPN5c2TJpRGBnQfr1JQ
e+FU6aB3vqjoRZoEeNjT5hJdC3y+XoLXhS/MnG0X3QkM0ZotjI+DDZgALYuJ7NCl
+ggtYuuXY3Q4QENNVPmPvNliEpebGtwLUqVJqWMfksb1fMPOE+jlX07aZ9EhplOB
or4mZ4gQm0yeuK0xwVU/X/VuDnZ+0Xd6bNiZjaTVNVWlBmUhfDb0kDFUG2j3udQc
qmi0UPXp8/tN5RAm6USGJKjyOm2lUeDltKmLFUgM+/jwvEgZszRR21K8NY1JNvwc
kYWzjK461VxpnKIjASuwwqsQ07ZM3CYry6fNO9U06ytMYeFfFT4hY8SGlqBgwHB6
ZFbidxj9u8jD6uvTpPVVLyhEJMx29TFaUq3ZwBxj92/lmp+NqJU3PYpDFFn8FP6n
uPW0QjS79MVjlTuhF/pPjepY77LgYv1eTwMcs4KGoDqD+EyRZiDhrgboSpnTjUqJ
aDTTT+dVIkNXhnWOo385kOmActziomxiopijDVy+0z8A6te7ReE21phKR3V5WctV
Xv9+wwbNVcC1LuWel+BVmK+q0s2Z+U3PPGSJP0gYQ4YKVeyOXfzK1Wp7/epp1GzM
E+oacnjCW1jyPkNBrjPhIcs2jbi5DvzkpcBASbOismPY9Q5F4SlUzuS+R2sXfAVw
CNnoEYnOiO9Wu4NPVsgUIYyXVBc534iM6GL7w0caiHzA8jV3XuMPyIZoZmG3lu09
YxNBbZENZxv7hkfVrqWjyF+ElksmNzPZC4RZa001zrcrBCmHfe932bSpa1PQjolb
rjxzb74K6CFzoivNZLwBepy8SrTZoMTtiAANrfvWruAlOFa1ihFzEbpYdrmUC7Ni
i1VOZUMTjQAz/Bmg5/n55DBWcJMhpJOtFmi+kavNCyZRBBQnBZw42/UFvF6vN4uN
bX3iErRrqFsBxtNKvBHk/baw31hmUrO2bR6JhKl2GPOSuO5n++Dn66nfqA6IzZkB
I7+TkeW1Sm/Q++XlzTdF4A==
`protect END_PROTECTED
