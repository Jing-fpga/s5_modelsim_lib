`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BxZjGSm5HjuaJWzdjmKTPmOsNf04FfUDIzDS+tc5ylVKKcZ19s+V0QbFY0pVanBN
zkTIWMTuYD8sD3UpwbQcyxUSYuf1jLTNgnOHv5tJTBT4kw51qIvw4qAE3agX3g4F
JrE5jQPKhOdM2u4kxr6KjTiBIQW9K6hv/9oUCuIjn1bRA5U5Yv8G/eNm++Xbzsh8
IJn7if8NN6TX4VZcNEGRaCOKL5Ow9TN8UuH6oXKLu65w2wsK96U6bvAofMf/um7r
O/9eD6g6uHahpBzMC5v2rcsVOR19GOTaQOdZBQW/z8SK3llaCovfJoJWCc+9S7Vu
597WI8ZlqU7ykSJcLjvnBVKjwSATq27PAqVpU1YkQ8P45+qFA/KOTagFeiEKYX3Y
G7g8HutbWFaGsZijkwKYui3rd6zL5pnJzM0W5BGTiYn9Djg33SvGFia17NNAmyEy
pe7TnEGfkvFr19DPCd/fUbA/l9vHuFKcFD6QfAuHROoDrkjLOSTbPSWK9IuWNo1f
iTT5wcRMcot6wQIl4ppwPWS+Rp6qD///+9sbhRJ0dln5sIcXijuCV0qa+Vm2a60Y
6VgCNSwa6Hm0IAo/mNOjsxf7VftFGJL+B8wG7xEIekZdWmZuQtX6S5rFDIpEMLaw
dXJF9JXV/Patk214pF5VeeHPjz7YHRszj4qt6nmOOjA46jlmvGO/t+DYmYfhVnow
u7v92zZC/4vchu51I+T6VnSxoI/qoujDmEuXamyQWuKU5aMHX9mD9u2MbCAUAo9Q
UWwLDX9XvM8+hypJ3ahpvqtUQta3rbshHmsxljn/i3uAVWBAnP1T1pHkh8bg2hA0
xLdTr/HLXcS4+0XQzDIxdH1GjHynS+rH+xxo07hgSEI28FB/97FagcR9Myg0CASh
cW7P9JUgGMo9grTteO4M8tMtqSt9HSo0KNlcMH00VbO8w23YUzQPXRTO2Dpl/1bl
yQFhi8BKhemzcwafvq9nkbGvnFai9BF8LjtHXS+Kw1hpRtwZnZS1W8lLYkDBgyP7
bgH7ntw/GgOZKX/9pRD+DGhMqCSyllflNnnt4xzzWpDlmqoWBmnBY4No+h8i1VFu
FdjFiPQNYnxvdNxvia9uN5fs6wBL7+N1oD3rltmsOteQua103nVspR4/sYWE9fVM
XZDGNqw10gJSEM/Ry/ZXWE5SU4qmA0ZPtfbw7UYE+TQL4QQ2uot8JfRRxeFthBT3
lGTVw9DqMlVeUsMvQV/8eN3++xeE1cr2fsxkHF/h4ktgUOtH/qvMKSdytTFVILrR
wP3TeeZ98RR4CnK7M1mgZ4aRzXJRaK4PRNUr/jIOkW4ICUCPufdlfOzEAYrx641W
QwI8CezX8pDNQ06Uu3XxphVB0mnXGv8emaCoEwL4F+6AppDUxUYimkAK0O2suknl
Uf4psA2w8u2BfTPyE6zyYTIXxI4l0VdzmV8/FTYNR1tcTU6SOuQACnzmdYDp98I4
FOw0f+BBYxQPue/r2hqqDjTdIfTQacNM7t6i8J4CcvauigIPW5VU14FfFcr1iToY
KuK1IfM3j6FuyuBGAFCiFEY4eu5yTAxmAbklXdcBBkNxe1DmqFWhaPhRh31Z4s0V
+UfBBqIBMy87e41kBCctpKKSabMAacZbI+5pDhfmPfgjfMZ3kHAdhPEPjK/gBckc
3lFnClA33Ot4MlID2Bx8FHQ9TAMtMy7wvO4mVnef4JKnYi5DVUtMGsvZiGmqBkqg
pQLYfFkmBn5dX+JINcS3BirI/6kV/UyrFSw+ILldI2wzrwp4HdtaZ+e4ufmWkbvb
yHt/MBp7HOpUmMVQunnp+lcAVmZhXE7rr5Gy3mLUlPcIuR4poGFfwfR0wA+nkxU1
xj1QYnun2IlGky0mdRwWDUtIeS8kcLEMoQLBbjf4RCvFGnMMkkfpizEMp5lhrwKX
wuXaGaAHDCDx5+wUXIoAsu4WJHaAG2S+pF+lkcysLnY=
`protect END_PROTECTED
