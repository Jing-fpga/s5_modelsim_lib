`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5YorolC3anHsGX8VYReEQLVt/M6+wwCTG0mLR+mpsNo4JD1pxUTd0nXPlT92iZRH
puZUVfaa98Xo1LUV58DimyxspZ6CPo1W5rYSLimYflqn++aryIcwtPnWZOvdjVuR
lsltpZRSb0FonCu9Al+Hrzf9aYbjY9L/NiyqTO/zQPZSGU6Mpt0KVcT8LTvG6rGC
YSstbttBFIwHgUmAgm5XUYepUda95w1UeeIqkihX1LxJEEbJx9IU3l3OqoqLDGli
VEgCFb9hC6U0eVST+h2nH7zzJJgYEaokw8pIkjgv0q5nEm08COq1HRWLCU2xRLfp
1euzd1mN9n5+GiysizHv668gMu381KkruHgjhjzlQnsh0Qw7HmzYzE4vRX/1s7WX
3Xm61gqSoHYHLK5FHjEdbSMbO3Xz0TW9Km4SOiS4pdqJYZK2M0MjFXFUuCQ/JDor
abhnxTd4QblQM53d3y3TGVhQXJAB3L2oYW9Au2ydBiZioXkA1smdDwcXGusMxSrA
O+sKIWaOLf/tc4aUQoLnvJlXCpEOEUlJNQe8SwXXr1VdqhDeOIDJzwR0tY7xhe1X
0AfE+awf472haWvq4Ei+MYwcR6iiPRis9JccVQl5lWXNDNDzL+mwthHMH8D5DKoN
Id+5BSh/pc2sahTM3a2RPogr0d0RjjChZNBIMWJoU1ch/c8+YrD8s+J2W4PL1zYF
StG0SQgEOoYJLCgdhOJB/8yX9910ofjOELLJMaqZB/DgzIHm5N2IB1N/eFRvwfi4
Z+VxqgJXMgdObVXYK1XFV/oKnkep3ca/tzBdBbfJdAvZmfHFwkSrqtf6hn07p/WF
P5FEGOeLZq/uhlHLaHwALexHOgC5paS8etS9SrwJKywOHkhX/ZDeT/vRQZ5SSi58
Gv7V0vw359xzUmDLr4PCGsEwKUZsvE4V9CaFNI0siln26xRYsvsubr/xy7ncksSx
rNBY4sFk+gXYGOH0rpLiSlhIDVuHTGnnafgz3RDynGtw81eN4g5CELIcNZk1aLiV
3XMnQwmrUUsG153C/Ws1F7NT+qmy3IPJ0R8k6dfBet5xBxi4SbPGQuYXEHbY19WT
fwE/rPtZmNQ6KKuAsU73oPIw41kkxE2nhdjdwSnQ91OoikhmBNbP3r6fiNKlnrpW
FLlezzc2dnp8XkCAz00oy3WGAb3B7kjxD23upvKhfphn7oDicSgBah2ju2JqZ+zE
9PrIWKc7GOO8R6jKAsEFvFN1qYl2F4RHLnEYtWXDJEk98CDiUWpkVJmjycR5NUDT
vVmWKLVKM57OkSEsVP0W0l0iDjIGEXWnrU2IVCJVxTEs7yPpk3KevdZvcAcVUxVY
R81Q5TGgLR0DlKEfi68HaBinuwKYoQrH2kN1C4p7kYSj1dqC8Z31uFqV3LOPQTXO
1tEuSvLl+qAGrWmCCTgOudvnwwaBnirbfDpt+QNuc4sy7ccuiNfHsh1f7uJxGE7j
cgWKB/LJXqP7oD15ECvCUlZ42G7PuoHyo0qp431r7kKvjouGeB5mYAthaYCNO/1t
OUVRxc1Gj9fwIS2A0frwDwde9G89VuD4+2MSs1XbUwU1rigJK1q2KkjOPK6Hyohh
SgCwY8fHOVMT2YGI2pLfWif0ol8F43bKCLcHVATczJE/HQ2KIys1WUORTnFPwkIO
/4oYCs184ZKpELsZgceGzquhr1UhtE4W00+BdGuYHvVVLacmgD4IY2tElqcRWRd1
RoJFp1sgWGb7oYZc3gW0rZpA1DfcFIfQuAam8QgCWQUEKqcw4H+YV+96r13O9XCX
Oa0Z+sEAStFzdOFa3qfW9EbWY4rfVgNt1M6EJnEzwes9EmhrIB599AsqCh8a2Euv
1CckyW7QoZ0uwoAIbbbFh8sxA2mrBLs/KNH3a+zTabR3Rmtwf0d2JYLf7FnaYq00
BNgNY2M65lmgeRn39B1R7MtJX/z2OZpzop55aTZXGe5D8LLKvJOhDH2x4dOOyZDm
zwsKZYyuICmuow+cfL9mSjscU2Jft5aYMbxkqjWEpBzCBvrvI8EKkApNMlWOK/Cd
YyconCAE1kMQ8yto2pbXjVBFGNHH/xzQpTE/C7tcWwxkyRyeT+eEh/rZIZEGxMhN
NKEY1VSYw+muJq+VhDbxszhX28Ou3F3YqX24GHnSyjSSFr1CcxcxdshNsUYOGxH3
AV/4Xyy/9Y2vn6uPc6LBeic5N+p4U06herz1dZ5L2Jcwv6JnF8Ip+8v7rIGx+yj8
ELwzyAvF5gW34FA+aVfS2GF9GdSfMpqYbh/vNzdPfQhnKkL1lNu+4VYdwl0s0Sxp
hHgxTbXaAiWOEKx9sBN4rIsZbzjyihDstuAxZDneqKbQM5kDis0YprIFumpwyz4T
hltNZrdjIpepYM5yQQtQ3ZAigWGtoUZuWirjhE1VWlbVeNzIucKwQ5u2x60onFDI
ctXxWNvYzHcmCYSUYyjy1ZgDjRzRT5Xrh1GhJ5p9kUWWYlhSq0ZU6uuCidUnGi4a
cRkbDn5nAKCQuZRG31X5c8pQtDdbcHoru8oV13WsfhGgK06iL56DO+uJMiGpMgT+
WbQUWbQtBqG3zaS1dR1xA/axfNz3pylSDZRcxiqjAd+mVVdO27wotpxG/9DIHzEv
pa2/sXN6MTk9Yx8SxrNFBq+/FL6XcsTXV+4hLoDg2MX5j0BiujwVfY9GauiLR1xk
`protect END_PROTECTED
