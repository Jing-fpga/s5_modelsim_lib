`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KRYETJgCadEk7uvfGGZxTUobngw+5yrdXcxAh7yKfeMo9ZK0FOgO3N1nNoQ8cSyH
UCrzjsoNJPXEXH1Boixp5NhCpXBfvhsRnDVFfLuNwa5WH8UmtU5N66HPqMkx2wrl
1i7eoyXwQ5dpN+tCigeLQdoPWXo7PvUvYjwutx9+2aTQtmtNFH3pAQsSLRbP76ky
xiKBBWdSjo6mKBaykB05JlQZ9P80tWRaIesJOyimVlkYmZxYLjWHN7UPHmSvLuYm
v+Y2r6dqhn1tlN+p8pztypWng+V5yd0L4lVd9brGMXthddtmazASDgim1Aa7iOc8
824PSntmUzuU7PLFnWvf/Z+iDizu5L3gBauAopMSAEiC7Drh9BSM/7PQ8tGCqoXp
ImH6uaRIYPzMJUgLDHvQJDx5vEo2u6whErnmzxv20NOXvdRHbuOi4rZzTj3shLRp
efg+sg8oOcfVWNzbezXQhCsN08+f6K2OAdpppTWhHCid0FCRR+ojXnyvrrxD15lH
K5IfQKIeYfwMLBavJis7t3JTuB6s26Um9SS6aPRYn9Qn4FBUo6qAZrOnGe7g4d09
zAJXRqD7oJjnEThZtj0GdkJF8aZWKYNzILLEscg9u5nR2zm0l3jx/OHO7H9XQ6Ej
RELl1HcNHgCN1TSuRdHTNBoAdzwO/q7JVocSNFwfogppSfplbXnUo7JxlmkGBTkt
TgQ3uZo0q3iA2qIu6XK3pKbdYqUEKB7yDiC4ilvxhPcXHhkb5b7yZZSLOhsCyGGz
NFN62zl1K4xTEt+zwSm79uiKxacxFEeUAzvaZZvEX6iKHOcK18QZxqYzymB65kh9
hKnP3/4xkDK5gHXP6K49jt4Pw+hGeMCxMpQTmIAjFy4QoXOmudxpUXprOfTXsbVW
fDZwMU0qYkskekuMeIxrLg1YHykPpXVwqCvU15B3KYR2gHrgiAnrXc26RmrSnaZF
/EnE8nxn4jlFDvm9igZfSH9Sre4XCfIAXCqbDPMkvD0XV753ou97GDFNrHaCPMpk
E7USOdtxX7R8XMj0xF6Wx+a5Sps9752DY/S6blKz949e6AGzSWfDTgCNSMdcapgY
t8qsv11qjGPhA9EcnviC9a/j8DviqTcPscOWGCXI/7iyPuHzTBHerfYHeLhJ0m6s
66/b/Q8zDCJDWMfdB9yHLi4apJcI72EE+2B21EaY5hN3RhWTkWONi+/zhYNtTMfv
l5SZZ+23QU5p9BcHLdS75Q==
`protect END_PROTECTED
