`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sCvnh5vvqiPtbRZ4BIhf0c+5ZXld++yRwaGluWULaU4ILn3IOObQ7uBp8f4l+tUM
TB5Fj8Q0pAB8Via9U0ZXMJd+Y0XOnNe4TMbNpEWhesM/AxJGty47mw3Hz/PC5qdd
PjAMYf8eJDydbDp7IxbzH6ueaDhuWnTHvtg2uROjC7myCO6RZ4zyg5RiA+2huiQU
bzIYpR5kQJggDB+ThoHpDZcwU0xd6g0conBeJofoDiioIb8JzvkBypx6i5A+Es/O
WLD2tZskJrqFsH8P3fU86cxH4/UojlK878V2y8JjfcDsEu5JdxLN+GPldK6YLlA5
hRqRAzDRqT8DTMXWoxtroVJt0ktm1ZxS1ZITOKOugMBlN7KE+JBLadTPS9UroZZK
pUgNxeCvrzB5US5NKYjzSPPQMJ0XuW/HehGYjsoVO/CN7JgCZDCqKcZ4oihbie9E
44h5qJP7wtnvRB3a0HkKXk+fLhHaqSGXvdtSivj5rnmj3EhHhosYb2ttTSrIEAEW
DAhLy8Cin8dwJcHma+KjrJX6j03TSkyD3A8RnK48w5cheqoSeyn8C//ZMCTJQyAP
dKLqLLK32eV0fTNHknVOFvPifFGIfiHR5P8dGNRdMUNsVYLixqq6ODaWOMHR1M4Z
Kyi5op9z2dlS+AsRHoNetSMeqkELGQdy3kyZE2jLLEWiHj75ZPVANoMUbLtfbliz
R5erpdU7gZ/ugCm1idUMN6UoDBxKh/C5VUQynb7M9L2veMU64+jhP6JXNhd8C6Mr
p0ynE2CoSVX2zoA3t1AVo3ROoOEVtNl6pMXzoS76FtovJctEseSCVXX94fXzUijs
KAy0roKPZ2R9N7gR2dbl0QpldPx8WTuLCr9ivGZ9PoiyomqWGhKERAwdt1xUiW1V
+z9PwxgEhzI0odolpNnWdRC9Lo0D0r0WzjVOKHvQyKblWfH1rrNhOCMPLZyusdpq
TAQvcZL4Sf/7HThzZWNIe3YuecXggrY7zXXzcBtugv6+hlPrDgyLnEPuKt62zD2h
JyCQuaP6CkrGz+Odn7n5lgkHpgIQhWqSAeHkJrzvhH50fUA8c9vUJ2nHXZ0Gtbg+
kDafG7qaIXcV9kupCham7rSi82tk2wWbjJu2yxOJsL3TEjLiK5UJkMv3BA6XvmMw
0OXkfojzR43dpqrwgb7wtT/WnhFKzRyf9kx5nfFXYyHwN3iYmaA/VcGvEdRZzNJ+
S2bxEsdDuoHzYvZ8QCT12nWe7O5AcC44Ol51OuvKf/7Z6oJbWJGD57Xb3wZPzMfD
cqD4tG6P0ssnum8SpqGTnvpM+6zMtO0fTpe/h8Q7aPPTxnVHZPHNrz4t8VKVgUrT
tVUPzjCk4ynxc8WEuwZq2wv0AL683vguXN8M0x3luDz0GjPgYy1TUjLWHC466VGJ
Cfjv81onz7Iov2iG90BDU/NmDUV/iSh+MfSUEMqXdCgro6vm4az5W+Sh1FF1UWKQ
8DVdSdYkHu/eo744v/TAVFmcfExtZm8jnwiopHWBfe0yxggr4nsXIv3e/CYGK68x
dzEsp6L2Aq/APXNSRPZkFzS4LhoZ5BGMhpEmn3HXONeswqElNCNSFRBnqQyojb9S
HY5JuzF542ScEYKFiDjLpKeweuJYuBuuyJPOeexR8khnpHQkuUG32VndKAfG5vh0
nEuPmUa5j4FPVw508T8m2waICutGDqZtf9NxEJVelU1DEXvPXEFQ1+NxOdZvGHUp
6Uyh5Y5XT0w6S/hl7FLcgw==
`protect END_PROTECTED
