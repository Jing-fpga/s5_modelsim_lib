`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sHgEetT5eUEMlivufnrs5F/6JEEoq+zM6G5//8C0auyqSCKFagfyzSl+aB2lO7Uq
3KoJn0OFmyDYY6N302gEzm0eE8Gyy8b2IJAkcOoih9w3dIviR/BfUVvVGjZBn1Vw
rykbcrq/KRLhuPBqLO5TOYireSVY3su06kAHkKsQ1ra1UBP5X20YNZnRr0u/dW8y
5xHcAKyPuj/BHHwW/7ak+JZ6mqUOgEJzr+y3kMsFbkemq8I+T1gczWsfXzSl8acc
lHkt6/5cLUA93id6cdbpozpBUhC6t2O4HUwWP5IN90NjU4/jKFhQOoh9uXgAYoso
UgQSTFnoYWRSqRC7+O1rdXH9vjNVXlUBw4hsEm3nPEgBc3HGLkBJ+I8i6LiqMfmk
iGVAPEcE46XYRzwFZ4yFnJ14HBZK/zi7iR/1NwHbiExgRvRWR0kcg3h9qjmVKWJ8
eRxsShR0gBy9EZj1w1jV26IOMQLX6nRdTJiirLPrU7J6lAJ1SORnRrxKauZWmWzY
tCcWXVMJc1y8h+elrDsmznf2q37hKFEl+6v7C8Es9eOBIE7aW6EV17bLZ+pLAvcM
VMOQ4/QEG4VZhzLSLh/XI+4w4Zg5n7Q7HZ/LYytU0UNgBlCDXZwzjZT56oloztQc
uktEVuo3gTJwk34pegcvQMqvSvkjP9J0tKW0s6LWa92GUoCYWlaHqFYCFky4gqkd
1lYvrcQ0BJkwFEKlIvMVlKBEX7iRwkzr356VybrhimGFYOD3QA6oDzeASVSvmcNB
XSwzX9BxHSaX72XoooFLsfQ3dk8hnSxRcqVmBB1eoo7vILEew3/WsM1PRTq2wpC9
QFczLRzcwuohWU3ELZX0uthsfsSwYd4vN8cZfdi6vTYNz7lgWuKKQO/IPMF0b+24
smfX3vPv/bX93+X28FMcXOrxDA225wL25eE0D2av2dus7vRoWh9Kcbr6gA0O4ROn
PpwjT8d0c83ZxpiVTlRPh9p2z3tYrSw68KVG6T2AHJh//sNR6gfA1c9+U7208YXc
PZ9s2v6TQE/E0l2aloTBGwJhXoe03uWPiPuSGiYepYNSU7XiEghMF+QlL6B+MJhu
vSeLHIq01hhT7JgGj+7UoumdKgexfQpgY0senoh2sZhxoQILzwT4Pc/Fau3PyQtO
Wivn4bc7Y/NAn6n627xEw6D2mVNAlUQ2ghgGHMAkgBTw1RQHxhu/OmthYGH28izs
K1PCnciE2gbvWrWhjLOWzXvB/pqGiBeagCpaZHDcd85PqvRFNe4vqgj198PAZ1TV
IHaxZlW2Oz0wD9ne47MYnwvca074YJasNsANLsAYR4neRDBxZZV7Tc01RmH+oi//
yP/Z1AscYL4psXavvPJVPyafZs6JKwXoYW8naRGTSYnvIAy0KviqmFzfVtN2zO2l
TvtdCUlCgA0MqbTWioQiaPKOzCCEIrtCrySGm1QamuIqeEX1lDNuNyKb9Ua7hjLc
/N476872qUoujfwua4qvZgs+VoXYByfiKeoDcc9AHDq+A4BF1qwHzL9fpuH3FgVN
/gVHGqHRltOLXspdrNS2mL/WvSNWHcU961l4U5YbT5N+7bdmlciRqew3aoplz8I1
tZ6lg9J4RSa37uoHk3QIUnMS3CWt/Y7H7+rFhzr2Ot1TN6YFz9wGJ/AR6ra5zRYL
`protect END_PROTECTED
