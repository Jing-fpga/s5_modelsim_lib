`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9mV9DltgKcuSx5XXSLGBukL26Kc+bKAsV56p61Q9k2unxpVUlb2O45dXl9Q1eTrj
v5wLtID75Bx5Tcf+2HJUmK2JsCThCuiKl1P7TmAaVWtzSD8Cp2KsWyqkBWO33ycO
2dDRNQCZcPRTAZcQKawJnQPL0fwuov9ICHbKL1fdZ9P1igzy91JhWPlrgTDpUq2B
YzKb3nMBADlgaKxITjc5ndZKYf3IyxkhUMeR2XCdSJ/jqXcRsL+peKP6RHfDGQtt
OmvKH55Trd8ofyjsOpJg/jEKCWPO298vof0E59KGysbrnZhqmkg5Z5jZ0JPyraDd
o+JeMjuSyOLx1q6qx8/vx49SiOTgEiEy7JQpfLaOqhe5CCMMN/V1Y7z0Af5qv6n0
TXnn9NewKSzwwxadw0v877iJONQ40XErbZfK6jTjBGTeEtMo00jCDcsq1xvtqyOE
XPZ73Vojds7Q94zvzKi4rJz1nu3f2DmC9JqdErKxVXprTH8eWdKCZuTvzRuGiNfF
13HZ3SQA5lRVA2auAqW1AV2YdmhafY63jQebkLyHjGQe5MMh5fIchsRTOIgiadG0
gVJCb3cvi4c3gI2+Yr1/3G3UovGsBVuOgkInlyzUpFpYEztrbsTeXmHvvWrV6DsA
+4vT14686qXxns+Uo/EmE/Qj8ZL0wpxqV7dbJhE7PMdW3W0gqifXR5hW5rFLHnEX
CUKBzeQ3fSlsWRrg+fcR/Gr5MMUT11fKbfyKO/QcExcMvDgsFFqxn4CUPlAE93WO
pL+3y9H1g9x2kkVBBoEtaiMEih1JzCg9MBGCazciM6yXWxwX/fq5nYzZ2fgYWD0x
4fSHgm8CET3GoY8xVm/EUrgJmc0Q/UkuQXPmnbodb6uQDhg/x4VNvIfjpRkMFfnJ
5/EKvehCIBw7DjfrbDfARH08yaYgy6G0C5EL9YU59dmxarblf+8rDsj7kZ5Lt53n
ulTMeWzt8q2QxqLvJladzD+yAO91tRqWD+XrEcgZYrSXYQmfBh1FA9JGGgeoM2WX
x1HeBxs8ah6oczVu4NJU0N7PIvKB9VPrwmUeLEYZVbV9ZGS/7/uUqpK4eqWW4qnO
TwHDE+6mtykXSjkdhcA/wIhmpyUO+EjzWOOjQxitHMIu3PmT/QNcKJFUe8ABnj6w
MXVJ54KCFIlS8Yecbjw3Qlj9A00nj1XYdnT6I8AFRBqW3SsMWae7d0nPB1jrjk3U
2aiYirMBBsHDSQf2QPAZytnNikDArd6qk92XEsZIAFoxsK99dQ9nkAEdxFS9zB4b
+CN4N2av5yNVCVyWnSQ/LoUzabYnIAjVrebKGcIqLOo6LZw1koa4tTwQxypvqZxY
7RVvsZ9swX6STaIypthrrnwnRlU68AZLNsSESg1UdVALt3OYweyrYTHG8paa2J5X
ZwnOQz7B8myReVqlO4+w6kPWGnr/cQHqcG5ljdSkAWoy1m2YDdBd/Cva1U1Q9E1s
Awou25Ba18xKQlWThS+f7g==
`protect END_PROTECTED
