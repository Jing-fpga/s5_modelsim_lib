`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nmnCuUgPtAjTTTzZCCHqtkLoX4dpShnsGjO4ViJTbHRLIZJM9aTKR/gnMZp3kLtn
OyojGNSOgYDodxfBsZkIMvzhJ9ZMYEM1LLXNbsJXanPa48esa/2cj87Yqheu/RsH
/l0nvBLplLpPkBhc7YU6gERB31NEpUpQ6fMvfWTA6VnrGVDtouaCgpLLi1yxBf5t
MNI43H/wWXOi0ZnEqxz3SnwVr81u4tjHgGT6gwiMh9UQuA3BbckYFkNo2KfT7VSd
krE9/TR3043062G868jOa3dvEWALdjGx7rYLE96h9TsReqgFpzmc3LpZfQuDzYdi
bhBJ5nmQRWLXMxwMejVfyQJ1ROOFz749jv27ICARy3HNQFxyr0WfAldzWBU252OP
HHKNZYR4y77ifpXdCvl7QK9C2tg7XtcylUg4Tu/7aD3NS8JxxAhXpdtbaMrRlmeo
uosATb842tYs5EQ/h+oCcgxwlQNS4dsSUm0sA4L9pFNpNUaY8XwBISHR+d1t/B0I
dv2GxcuykW/27jhpackJMkwoRHxOAoBWDhwfcxU3Dj0Ul/SX4TCBwMc5U04d/T8d
Bl/cDNTL6U+oFAufmdatTQUUqXsxK0JVbjSetnq1C884HSsLQwwF/SQG0WQnNv1/
G797eChUiz6UHaugrCec+sXpfCMtMrh3/kl43wYnoBGe0KCw2b6nC6XnJ0RcGDJ2
L4DYMV3RGuA2EiT3ZR4PX8oP/pNfYPcoYLalRSXqEHqAiiuzEJbK+LPa0GLeWZLI
MJ3ATtS3KI1AVQJbecvltDwr8TiXJabc8l2GCyvmMxgzlLSuayIjh7hOto/77ubp
QyujrBLkXSebddtys1ER/ow8IrnNUzZPuSX1bInxhKiC/wW6/2GpxmrZL/cJczz3
GEJs/JjeTA9jnPrewBSyhxR+IbPzelmtXBVcKUdWVY7L9i9aAU6ePr5GX4bwy7Tv
pB8oXgtncchnqkhYW3CxrCL4zCEpOkGAVdF5C1sBPjwlBUUMS+E8GsV+ixqlG1ZU
FD55EGt8HB7GUPJMkOTb4hY/aYYRpC6DK6HIgZ7ZpoyLlry4HkyiSm3RJLhAXViw
I4RfF2rECQKsHB88/TpT+vVR/dwLodJJIRH7Xw8dH84kAfYyaotFnoueO+WUGZTT
Ocq9Vwl/gDwuTdWbXc+taxKiQLtYcD0cOHQAjC0n8hs34i6P3w7H/Js0INsGCEep
OZiWpd8Z+yluP0OfOsFHswJVnXhvjZZyWmDiEtDgVRgXMfEjzXZIclqh/omyROST
`protect END_PROTECTED
