`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BdMrX8NjS52U9Oltckp4ozoD5GHcspNm3Ui3EVHy4ikao94Ddp+AFDO2aDknTkWZ
m9vCN2+5SmrrFIiMqjxfpGiAD008e0qOrMnAXsECGsx2us/5v9D6MDfdWSmYkS3F
jXIt6g3h6m4UNmgzy0+vB0G3G1coXbObOyVFAr1TGDzWFcQdYvGT0Lp4nelS9LSk
Z2rsw1yrqkqi6Ods4Y8Jfzt1U9UjJVCfgS93qlR5DfaMJiDGPu1aX0PeiC/iCzC7
E1nDFGCTy3h0HXkUztuY3oYzABD915NZwvNoz0bI2Mr7/3V2dF8CMUJ6xMkqxrVb
l3Wa8C/GN9F3JlobI8PkgT9MLZjzCFTo9djHl5NLo7ldGZxh01cw6qQU3B3Ya5of
hn33zA9Ilby/4e8IWZAHPyZq0CPJV+QWCWcU6H5xAb6QqLPm0d/TLK3miR+r+qZf
oMg7mzru6UdFxZHyG9GApJo10On7nxMtxetJH1V5C7KQrBF0Mt79y9M2NhWm6cI8
IJLcyfmVxStgG1mODlulzdCg5mPwYfdcbBq18Dpcz8IB/LrHgTMN+KEkIcVFk6ay
pnbt5YCO3+re9mw3pChe6FPvA7sN8NaUnTptlxb7pKqJ6pvvIZYTpi+M1jmN2gDG
maUnjzDJaRMPO+6fTWlVQvLjqm/I7STSjQK9m3BqoflQhkkw4XJRL5nMmJgwePqC
TGcljrRxtFKIB5+JFNmQlsQPjUt+kf4FSo4UZkdRL/ZfblhdqnjgbexW/yVrVU6V
Pm0X5koUL2P0mq+NYLngCdHVfZkA9zBWUttckVXRvfYIRAbo4c+/Ykba2kj1c0If
oClEh6FanZOaZO/g+u9JVtzAmyB5rycCFDZk2S9GVyNsiyg498pg2UTEC6fkT27L
wk06NmEb1cNVg951+lIbK7pjloBzd8Dccih+Zsy9aAdBYfqTM1ntyY0OjYaZgI4C
o4J4nDOAZKqmwe+becMHBadZBMTA0cId1opUmkhhmibGFnJk7ClHvEIUe/BvsL2V
fP8jzMw+FPDXd/s77I9cjHe5tITTyM8/vT3XI13tvgkE4nOB/xRR/n9x7atiYTBG
v8HGp1JnjcGsANGwVu2ixf+S4jgdjYCxFlajrEFiceDJZpPWzpwAXOpFxo8+gVxJ
iMSkMBmXFzf+UMtU+KvtAywAmgxUaJq2s8rCkJoBLUM8yFCoKJin4P1qS0idHjiV
SxPN6ZF3bEJUWWx0yYWP6NKGgVuUPX3ACnRKtp//ajVbWbKdFvRCZ19eVwIQEzSL
t1cHl1sEexunJuFmZZS6M/AubG6jeU9/WDKGBFgRUwAZOEL/lH9TsfLXGeF0kr8H
4em7ZzLl5utC1uFyJOtKnruofa2q0dNsJi5R0LmJHDaGxTJyR9q/t8o1NK9kwNzB
I2Fj32aokmk9bbLE9RAyDEObfxtSi4AXAuhH22raNeix+07X7jFWLz5m95vf9zWF
cMu71XfYs0coM3VJ71B1uKngL19i013TbzPnuWMqmWT1OiiEnZx24U/0RAVzjGzB
VUskpJnNFSTqfHf0cYjPdqnmiCavIGkty42lrV9pDJ0Tnf4eqLZsyXVXNNt5jpZq
WyRu3NYdEjPiI6l/buoXxnj+Z8sYHps0Mmqm3l0sOkAzJb5woBFbqpUdwidXnF6H
rnc7kYkKlTI413OxpMgXP2etrwQfU/x+ZOmVIK3Z/BtIiIGLzQ5n5vuiye3O1ctU
AfBpYoeG/DubvVQs32/V4PyasLj0cSFgwmsib/7gKgE+fqFVYy7jKpIYD6XpMmhW
bpB9gsRIwy+jAtDBbCFN920vnlfrMjstiUJHleSJBlo380b23nlkuySnU41uSE2d
7mVR5skeC1u/Ht0NyWMbYWWlpkIipgC7LM/60p3d9XocGOaysakZJRyLVwV0g8Mr
cLCMSnBSIANQjW6qSAlZ8SbCr/jWSJjs/D0lIFL1PAgvGvXMpKj+ucJGQ2D/YDuU
5aw2wPZ+Mf4cf6vfL6BiioTkN25A5xzK1ydDpltAqWP0swfceRx6qEperX3rUdXZ
RST2R+8n2ULsbYbGZ8C8vOMDMk74euKkIZ3Dpql2uMz6KJ3d06Khtwy0WLp35+mr
kxg72snOLjwq4FwQN9z/mi4R/DXgNQPgVu7Sw7/1dVGzKwroCS3KrQJ4fJInnj/3
grLE3Uq6yAij5EBWG0KzzdgdIpE7ag08qyIP7/Vzqig0XpxmRhFgQKIMkAqMf8Br
EL7w55Bpd++UbrL4Dq4Ow3Eeyw3SHeaA6KM6bFA9cy+6WvBTgkvF98bkc8B7v0B4
YC6Uxo4tt7TufCBeEzZwLcEHcGLpwuRkJyz85Nqe8CLnd5V5lNsbcXMiEo91QbCa
3rMM4cLzJISei0vE0VqE8IwXJFG12iBjESGWt3bF3W++qAUdPIFAhvdg5rFfJUf6
GlkgYbJnFN9gSG9WEjDaYRx7XcQAEIntjZ7IO/vcCOCbGIqxsetjkbJKInPXUdMx
80rLLzbupoJ8FQ4jqdSDPBQAY9ZuZlCgHRhPgd4R7f5sO29PCvsL6w+7L3hC6KGE
HNNGk1/tR2IXTi9p+6GxHSj0FhrlKDgAss2R+vJWxmeRfv3jc8lNZLIt8d3vsIL9
PfLZDeQEcMQ+XGrOj/Dsx6fo+SWdrJO3r/SXTSjWIfetzahL6kOdi9F20w2Lsf2G
hKkQw5m2i/ndY1iX1WqcgaKSkewiqLJpA896Uv2BjDKdn6Dxn2oYfxaOxH/F9jMf
k8xHrZzBXUU9hqOSWagDO6jY8d0WcqqO4bVhA8q/azShzkscFkUTKukwrIDsqIXN
WZNlhTDrK/PSZefNjeAeh/5PgJrfk7GF/aAidIiTWDXuNwNfmtDVYaGIsKy9gxS2
30m7SWSrG8gJgOdoQ9N5qC/7PrhDGiQzE8konFKcv8eQ7tBuW9fApLgjrYuo7UOg
RZBZIZ4QfwKQRyGj5bdouSUKkA7BWTXXayUsXE52+cKmJ68rQc3iiwyOfVtV5WKQ
YdlB8Bby6jtXWeBfePvSd5/jp6qCTQUyQ5+oPVZ4as1Fw3CZawHb8exUuVAPSzRs
QLhBd1Di+VURHXSeNHYAcTkpgJQ6Q4O1SDKtPEFi5NsE1PGfAbvJMQG61gwhn3Sb
jJ1n+PFLG8a7MeeBY5c/UloNuCl26MAXEFAUvfq6BNEdz9Qx1D/rzHIPjD5ps9oT
D95h9iXZNDsU+X4oMn+HxMGJkdFGhFW3j5OAru2HI+SAe7e/T1xBkwJYs4I9LNWM
ExXz87uV61+oyx7czdYe4MVOpFc1tU+PStmB5p0oKQ3XKncpsFeZhZqPo4meYma/
EA5OVvHos2ZkOPN4cuBVvwRv0HKpQi/8dcM4TECd8kJ9stzYeUNb+ZkIdtzuNXa7
66W+FQ2hImSVdV3f5TqSsqrBSLxwwMZPHDBmnCh+LOCEzA8zPY8zsvn4XClzaN0c
8IusS/sYByOguMytLh3kglHXm4lkrE9a732PobULNDLsXytPLfngZ8pCt0p5hNXT
DPtGRnnzoVO2ntJ8cyvx7l8u5xeu7DF330KyY3xp79Q7Wf1HR/NS863qqX8ToxJm
3CE2Z4ZXQdEh4I3XxUXFIkfnYS6b9TSMola0cSu9WdXh2xkFox93HFOYqs8u1qPo
Xa/x7s2cTCEW1HhlDz4I9qnma7KTxaveS1OjiwJQS2oxGq+V1x8tU+BmqzH3Ykkz
3Nm/B3SeM51Nw2XF5eoX3kYRNCoYT6bdrpPEQbZcnPFVTlfTQLwnV53um12lYFsO
R8g5kU0Wk5WpyHHbJIqyDV3sEFR2AfhJUnqjz3zXz9B7Rni2OBvn05QoosThF9aV
czQkEDyUmlIsEsN7GSP/1a8Et0hYCumxfffmU57KvEwBkLgKU/IjJD5fndaAZKp8
HdB/ySc3oANavW7LyZidvutROa5CmIWQ+Q94y/ES3Uwy5y8NnQTl0zioQCOqK18L
ikDyWToPNlbL0jZMWRnAb5t6HJtIyZyvyh48y4zdwlqvLev286OiWUTYFnesGkMM
Bc2DdIlSW7KOeDWFUpKa9L57hd6a4x/YZSfdoxNob4sQ8jasjKGcg6wR4rh7hFd2
18j5JluGT6hCpsdMmzBgSlYkF718bxzWfBzT/XdsUJgWDUciCncc5MSL74qWWNn6
EdNnZXsa55p1HeIQNatxAXSeKQpLqHd+2cLkZi7bmXhygirsdv9HZQIywU6zHetF
5z2PecNGDUmHcv0slsDoZv/wb90Jhbz2AahxXXHOdw7RQtqsYS9mqHQuKNKoS3Bs
2HdZI4Bps0jsTB9NO2mEXjCsrZZEeuRDgtcRevLa2+LwD5zH5tw6fDmssrt2Snt7
Wk2DSIzx7AnQMmn2vopOiY4Z67fB8lJhGFOGV5Vg2h8TVwPBTTTLyH4C6tts7yD+
OnlmT+g5UvDsP0QrjbzFoPtlz3y9yd0vKq5/JfdaVxU6OnRSzFLlCSv42s9cI4HH
Oac2DZzznZG1ValUxnr7Gz2eCheyXWCAp9MPWD1m8Jgimgs23H8qjIn6D5Rt4a0L
sLZAxybrgUUByMmIJfWjlodKOMqE08v+AHu9JYlN7Te+4ADgW5KIOIs475LS2HtE
4qdqOzfpc/G0+ZYrSFeturfv21vBTyuJexGPZM4f5ACZ6zEDDrRC8nHq7g2cT17/
jzRG9lFo34JrCQ+lGU74DKDK/r3Kf38s16G6ZEciTEcOI4F7ewy+G2ROc21jLlAe
44OqGSIWzJTPO8V96fAK6L9GvZymdmobuwiAfznfwBaUA4KgcsEokVJZrtQspZ9S
wqL9HuKJA0UL0PJFmrK/9ED9KTDHR2NhC5+IqlAJCpXXE4qPMhMCFbPmNwAKjQ1p
JO6f3yDZ8b9bAP1ch9cJN1ByM4SPmnOMIyGiYXDI2fhmmVBqcxpLzTXxKl2Jr9id
Ah+Veu3v0ATl/7lBkQQvWxaDpI4CHLYFqi7VToXmurXC77GKcYd5pJcE2XpH2H76
I0rt4e6oGHQwU3PccHbHri+TyWFbitlVmlAcWFuE6NDwM7HNidqO19GYZIodJcpE
s0q0Lecr9bO9bo7pPbuaiYuBlJcDyqqi6qd3JWuE6T2ilW2xP6DPtK4TIAgB46Cc
/wS80Atq+TxfyKjKzzEhLyvSt6GOKTyhYM//Wl4umQBIxResoARQEt9pQsMU2Ad5
BkV0iO1lb/zwlFbiZmfxU6ajirSzle6JpUsJ6odxUm+R04qiSQ9+Tck/AJs4rnmF
9J+ImM0tVBGHWXY6J+fAdaveORL5mVq353XA3DaD4MTSjhMz0lbUkrgMhpMMl7Rg
SiuSyaNak6v2GkDKQpUk/GI0vM4YtOFIelrYN/Tpi52kHS8gFu7sKsxC0UlZPKbI
nvfhKSEgU2fiwjyCjthXb8v3mleQVTGr+xbgFZLNWEyErSXJphiQb66HK2etNvG0
Ox4+7TD3505WqAkmmWBOktJkhQYBb4EzUMcd02hbwltIsUvOm5wlIlznbZgpWOzk
G+wvzZOdWEtWfBWVwn5koocbFx/r9dQGkZphn5f61Vxh5LlEsKqq5iTm4nsDhaut
/gc/3p9ryhPv82C5+aVmhQgEwYYVG9jzgLuvwWrwHME5130petxWIBnmMLj4HFv0
yz8vrtGDk3qHYD+gnIBQfpWpT11XtKGwRCoXlJGyrUCu69h3hxM5+eU0FFPvFUjj
BF/XiImX14SmSz8Il3l3WpkTMXiznars1p15D9q7BnBk3jUstLliqtKgFGOWQ7gQ
OrvlArGttlM4iIwZ4pnyagxI4SNKL7FZ9WPjMeHlXlkVf9kzjgzdyP5QgGiiGDQ3
CZbkq0eg8lo3CXHU9F3wRs1WfKUJXk3QxoMw2Ga3dfJds6iaK2rqCzq1cKQQwYwu
DcxfLKAZ0vLx2Nf9RxU5U3kwxHji9+E9q9T8VjLj6nZtcqXMEkAPqBv2XkJQhJ1t
KSJs/NOHciagjXK5VwU4PavAvEL0ezDUnv9XGB0fxAzP0ZK8k5ZYzSz/dIY8EzEZ
Yu0UjIsNDFdjYy0Pixg/7DSc0oiZaOVQ6xsmrw4dKGnKUAJ6TNKkekZh5nZr1mVF
J7zMslpxlt3a1XHIb0px1F/bZbQXquVYKU8jSgk05x036C8o3tt0jrQNom3kj8JB
BmBA4/XsyCa9SVbPIlX6D8PBdG1/cJy5xTW5LBuixM2FVb2Z9SMZyg8Oiu6mdZ53
DdUTx2d9tdYdKRbNHSIiy2D/V1eiQ9JqvfsF8ZtZcFepUqzRrVcyPARX/KyG3bQC
hWM3g0z8ylofL/eJsX0tBOVGd+dyxEy9mpVpEnI0h8ZsznFszc3R8LQyKxuNjOZs
rmo0xHbDt6LYMXAXKX3VCs8DxnazndugkbHX2VoCj81wlQe9hj2JUJcH5xlU/kwN
jZCY207G1oOScNHowYhRPx7xhhsvm6zUMUmpMYZDabyYj0nBkwINkzib/tQhdFqx
a9iYw8Qm1Sjh7Ufjl+5PWggMNgVQ2NJCTDRdn8MHyqDUEyO8n0mr/OKflEwa/HL7
EvWkifPqIQmL5F7CkQzvVRjRf1qg7jfZo9zOQVtV9lLMcgPHmBkwh3Xsk2ZtdK7w
Hch3EYHcMtlBKmlf1MyBdEgNdlS/MQSlpvsVKub875ZYdJNJyEyAqQUka06/Pyfm
MSSMsPTF1siLtKSGwd4w2uuNt76Iq+TSNxyVkJaE6e3BVHmCdWbMLZb+j1dSmYcc
DJHWFepoIKt8loms36bTjtVZnwdRhRVKn115KdH6dgKdurI7n6iI5tVzyQgZefwe
mdde7yO9KeJyCjBracjzOkdK5MnzNnl3rB2eLHWbIaBluMAT3RVQ7wBL3tjVejLF
U5FzculIA2FpgvGyAbbvwmvv5GagRL2OElG4S44Bq2q9/n9qSWXZmP6X3f69dlAF
uhv9Z0xxaWMO6faTGQkFfiOPNhYCr5/U0dKckbpVyHnuCS/aVu4tNzDjqaXoM4VH
BVVuhtg56szEkDG2YMS5HA==
`protect END_PROTECTED
