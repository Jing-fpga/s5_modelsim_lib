`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LaXxaD4TXaap5YyjKKE3jr0klIfLfG809NQn5kHPBpe/r/HpKEzemdtkPASPHygt
L3gzLkSQZI8vzPCuxRYxfAm5YBOrqExjR1gxAB4UNVDyY9BWyuvN36fyLGxfnjHg
GCkAggoAfYmNOsZTjg3Bdmmqbc+LsO5qeLP7KAdw3RHVlFNO2UYYPP+zSsX9tB8h
BRNWv4Lm8C9SvezA/nHCEfNVmAw4UyumHzzkehmkhBC9D1/StVLtAskqt/bP9fDS
KZ5tu+HKxgrieR1Gz9pzEniVk0ZFHOqUJyORaQGuCvDOn7dWv26TNIA1G3WFWpiq
ljQQmlbqKi0y121folUI15uFZD8+4S55lVKWMHx1aWAOePW3nZG2wqpvbk2qFymS
gARmBFe6O3YKVMR14DdRtrtbgldYqtk0rJhUyCtMYTtFl5ePERKWqhDU7pA8yX9w
8k6y/T4ac4WWqJ3ygpTSLQ==
`protect END_PROTECTED
