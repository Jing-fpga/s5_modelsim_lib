`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7MyPX4qycSBq3zxFl4P4PcvBfD7Pm3bo+nvnhYGCjEGW4r5mZbEe64y3sIClDRzH
0TDNGWeoTL2v+JvxFlpjd9x3DsxR33bQ+Ve6kn2TYSFmb/XXx1ZDquv2WQpeTlIg
N4d7tYSmBVwUqLdshmez3FeGC1IHlU8IP51kt5sltPLitn4hit2LdVgaj6G8kg0h
pm5epTvjml9iLfq6BrmqiqN/Wi1tk8n33A6/ngLD+xrMBY41voVM+L+2zBFlgk5M
b0C6hqUzqgE1eHYcmFgMt3iq04ob4KwaJfxhwZCcDZdY1LRBrm8N8bM7MsoE4yED
LU3yN6s/4oeOTdX0pkoqRdEYsfGQmXNxi0l2cZVb4iqvaE02cC2vR8eHmmfln1Qk
YeDOD8LhB3Suip7tt8jkJ+dr6lKl5bkqj71AOIWUc5vxAfPqbyqhFhIhc3tKcIn5
r5kdhbhgs6dlDzVqTmMZ69xO0bIHdcV61mE/pcj+xJxZ2KWUGnN7D2fligZvZ7CL
6W5ecfPcCX+HIk8NI5ApWCJBGEA14RQV7bneU+xqU3hcMjFz4x163HKUILV2BNcg
j/xZXhlXr72tlB3UCOjpfDeRpWmXv0knTrHUsPNCCucsFbbfRTh6i47Cd9DS3Vku
Uul29rPMNnAniiTEOTkd3/dmAjB63sD38cu6O0lgggdvInHlUQABEtFm4zxord/V
sB5naQtAZEQ4QS0mI5sF6Y3MtJO1H8lQZCiDTgizi7SWsUw3P979vjXh9l0F6Chb
sNzk1/8hVRSafZOK6EmRx/B27uH6Dus34HPRf6VGN9jGgp6clJjhbCFkRWx1RplA
K5CEIS/VxYcAllMseLvgyxLpNqJBdDpuBZco7sX/AqkswOZVvwuIEUxmvY6W2jRJ
MB4jXKxWNIZWg24J8rc3z+DzGww7KCNxHWjMM9/VI7WY0mNZyfEvehlE5L4xu4j0
NVx2/SBWK5wX68N6togYgiHWuBmXxNYNSk4kEpZ4QP+r0tk+81m/hDms1aNY6vM5
4I18qB3PIywidhkKHIbbMGflokS1MB9ZFNNwUpaflcoyqtgRe+sfW7fw1HwQZjzZ
EjmVELAcYAD8Y8j5ixVse38UtiKIuNvgBsP3+GixBLAoFRR9lhzBKUYOyXyB0SmO
0ibhgnxFjxhhAiVbF0vtpdXVd2sVqRH8qAPyritb8ZrTQN3WxnVGrjFd4MbraJLt
pHUp7Kfj4SiUbOohkExxiVglsyZdbTAG4kYpCuaGwC3bKcNga7LisSA5e2jNYoGv
FV8H3q1Vm3T52MtKQ9h59xY3p0++dF3MpQqXdgbZ1cDsp03JbXpsHRxlhT9CcYOO
SCASupenY5V6oemRAtM1ryu5dnGS1FF8gomG3ueV5Y198x6Jh/88vb52MZRboM7x
KNeW1pvZBLPlO/ptNXjc35bGKbIyTh2ELpJCNGE22Atjyq5DNLM4pI4E5uCCjVF/
kU3WqzA0tUN7RRxoGmFrIBoZaOjRmtHkc7td5vc2tKsxC0bxQ96CBAn1l9nwe9pv
mPbbjOL+W1KTzDAXEzqNCGZ6hWM38VlmT05yJKWKRPA=
`protect END_PROTECTED
