`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kUCBNJylxi7GSpJBqedzckb4wiROy1JKQ73LvEjZa4A2cP4OI3mQVtre6j0V37w1
t/wKWw8cP0ZgdY+hCK2/cnaxoT8c1uPdMc0g3JrdstuinkzanD3+qP/CIDifS0qt
ywGQWZHQ9loEkK2pKbiG7ug4/TQxkxV9ym8nN0Yg9CEWD57rW7sRd7K/PahG7osx
+4Wju/wuxy6XOPeepT7ZqcNAyxUqx7bANv7rUb3UCNsgx8nY/POZpMcF90Va398D
WTqeIpUdwc2qp5Mc2Fbr9T/RczvbTJGnffaZPef9YBJJkXCr9SFiv+8RKknTwp2S
a7EEimro+uRx7O1I9j0hPba3Ct1XLIrmTMTChT0Y2F/qLgk+Do2bOrORa474NoKF
o/tTdHAKCrXso19qzXxEfKD9EaU3hVPMm8lt6s2PxHEGmTEqbRIS0murna4Jtwhz
2wGV9zGVe2a+Z5cI88tUU+1/s7qZVEVfrPDPU0P+3IdGerjdFh9oMgH+nFVDHJiX
M8VDpIPOqtXdwsNTHXXStmcCIe8i8nqOU4+8kN0IRnpyUnmkIHvHlhX290e+aDtP
ODxPjt7Oz6vyF2TldUn7qHuhzJcqd+ACY/IY2B+5E7Hp3VTOEVZTh7GR/mbJ5JZG
lKUkPi5SClQikE4cSoRKaYTIh5BhPFTwhhEayT+9ks1KEfJG5R3JQ0HOB4iGWf/Z
gOqU3FIwbcHHIhLu4+VkCWCkthoG4gbjslBKFq0pd1xTbiqd/heUtdDqkQfKLq0F
7bzgV0iKRAURFfPBTRLmcIGjhBTQbnbJk7VkjTKHW7We1czYTAod5Jvi+QyB7cF5
1uBO4WH31up2zk3Cl6ThFk91ed0lwazmK6CNsMcQZUKxvNBPksFMk+dceTaX5LD6
O3Geo5AoUICcg+mFR6ezWJbxCdRiAIWHykJV7o1noXDsJnpHXyyhI1iAVxAXlWHe
3p7AhCdVZheh7cYF8p2R/xnhMGjJ+Zt/ZCApey9ZTMdrXwm51GUvu6YwB+HyDjtD
OE9sQKmHiJexpgw41/OPi3LyY/GvBp22zf+oY4S5aeGTmF16WGxNeYxPLZkdi5N3
MFqNplhZBrshtueY7LbN70JHfN2TozispMVRm/4zjr3zLBtf642Uz7wv2jo3H6ON
fECJhpCs0yXE2makwenglzfLU8r9UAEdEWzfWfQHIFI/9EqD0gyWFtyaPimjGFvm
UN9QbDuBK4sUw9xAyp/Zm+s4l1ihkIPR6l+BRwBz5R6LKNNqrWporV8y3DVIJK5s
0VWOMcfs/0WVfkeEVk35poF+z9kN8/2rFaG1jX65BM1jfxYWYVrfDmbydGhHQXHa
6eYmHyUHN/qTMzZewHg2YuIsgINl90iaW3/KkkHf31R52jnGiie0lX+csA7SJGDl
hg0ZRDYAgUgbwvZc6kHu/5g2nrCu6Ql00O0TRb602VrJdQu5zLhMx722fSU1LdS8
jLKcN7Y50y9EG5n17fNFzyVsJCJUW47sJkHWQns+RLA=
`protect END_PROTECTED
