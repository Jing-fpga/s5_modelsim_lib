`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vOdw/eLZeRA5FENMEpb8yI+eFzX5lSmAgkayjdneuElUG1/fKUf6+rMFOvbP74aU
lXAJkD7CIPJIZi8aj9Ed0IAJRhJEOkbkNFTdshYMcpGWAkX/YJ2QCXmcZp+RwWqo
dEnDFCuWsDu8xZKP+bxA9Q2VttrdxHyKmO3DRWrkk2YY2T/QHRVdPjKiIcQsWWmK
27uGU0EBLiG4BdAI8CW4AJwrqGnwnMJMIm53lyxCDs2OlGBZ0qIvkYxlzRnRPkGA
qzegrgDBIfD7zgzsR8SW2BLqBoCgzK4x/zftpfUUZFFUy5opIRspF4Y1LDSJfej4
JoLN2wWWijHBVDicm/H03pxJy+PVufVmnp7PRHhx9Sde4XReDrQm4Yp6s7ICznYb
YgwoffekSQrMl4ZtkL8E0ZU9Xe60Jh2oBMWU+59qnASCrqVKtExK8IAkY+7Yfgj8
Zv+UODnsld9++qI43TykDKx+XbrrCMqjh//gHARcPoWL2td7hOkDwQnmrl/qmX10
6oTBiw5G75TJHXz4VNzhm5xDVlwweq6A+NUy/D3jpAaUj8mkriXIOJyjkd5Mz/Ra
NqawWe9igakNrg1Q6ow1WdvgUiysEltacSiJWwAQ1nxX7sT8+1LWBYiSW0W9MaX1
DhOKC1ctJx+1izPT6w3PMUCxAv9tGuacsxTY01e8WfZm3aY4NL9iJz4eIHf3o3Aq
8Y37ANKldKC4uxFMbAcgD/UaM8LDeF8wM29t8gj+3wY=
`protect END_PROTECTED
