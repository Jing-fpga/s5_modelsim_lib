library verilog;
use verilog.vl_types.all;
entity stratixv_hssi_pma_rx_att is
    generic(
        enable_debug_info: string  := "false";
        var_bulk1       : string  := "eq1_var_bulk0";
        vcm_pdnb        : string  := "lsb_lo_vcm_current";
        offcomp_cmref   : string  := "off_comp_vcm0";
        var_gate2       : string  := "eq2_var_gate0";
        var_bulk0       : string  := "eq0_var_bulk0";
        eq_bias_adj     : string  := "i_eqbias_def";
        atb_sel         : string  := "atb_off";
        eq1_dc_gain     : string  := "eq1_gain_min";
        vcm_pup         : string  := "msb_lo_vcm_current";
        off_filter_cap  : string  := "off_filt_cap0";
        rx_pdb          : string  := "power_down_rx";
        var_gate1       : string  := "eq1_var_gate0";
        diag_rev_lpbk   : string  := "no_diag_rev_loopback";
        eqz3_pd         : string  := "eqz3shrt_dis";
        eq2_dc_gain     : string  := "eq2_gain_min";
        offcomp_igain   : string  := "off_comp_ig0";
        var_bulk2       : string  := "eq2_var_bulk0";
        offset_correct  : string  := "offcorr_dis";
        rload_shunt     : string  := "rld000";
        rxterm_ctl      : string  := "rxterm_dis";
        rx_vcm          : string  := "vtt_0p7v";
        off_filter_res  : string  := "off_filt_res0";
        eq0_dc_gain     : string  := "eq0_gain_min";
        rxterm_set      : string  := "def_rterm";
        rzero_shunt     : string  := "rz0";
        diag_loopbk_bias: string  := "dlb_bw0";
        var_gate0       : string  := "eq0_var_gate0";
        offset_cancellation_ctrl: string  := "volt_0mv";
        silicon_rev     : string  := "reve";
        eye_pdb_att     : string  := "power_down_eye";
        vert_threshold_att: string  := "vert_0mv";
        v_vert_threshold_scaling_att: string  := "scale_plus_1p0";
        phase_steps_sel_att: string  := "step20";
        bit_error_check_enable_att: string  := "bit_err_chk_disable"
    );
    port(
        avmmaddress     : in     vl_logic_vector(10 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        blockselect     : out    vl_logic_vector(0 downto 0);
        lpbkn           : in     vl_logic_vector(0 downto 0);
        lpbkp           : in     vl_logic_vector(0 downto 0);
        nonuserfrompmaux: in     vl_logic_vector(0 downto 0);
        ocden           : in     vl_logic_vector(0 downto 0);
        outnbidirout    : out    vl_logic_vector(0 downto 0);
        outpbidirout    : out    vl_logic_vector(0 downto 0);
        rdlpbkn         : out    vl_logic_vector(0 downto 0);
        rdlpbkp         : out    vl_logic_vector(0 downto 0);
        rxnbidirin      : in     vl_logic_vector(0 downto 0);
        rxpbidirin      : in     vl_logic_vector(0 downto 0);
        slpbk           : in     vl_logic_vector(0 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of var_bulk1 : constant is 1;
    attribute mti_svvh_generic_type of vcm_pdnb : constant is 1;
    attribute mti_svvh_generic_type of offcomp_cmref : constant is 1;
    attribute mti_svvh_generic_type of var_gate2 : constant is 1;
    attribute mti_svvh_generic_type of var_bulk0 : constant is 1;
    attribute mti_svvh_generic_type of eq_bias_adj : constant is 1;
    attribute mti_svvh_generic_type of atb_sel : constant is 1;
    attribute mti_svvh_generic_type of eq1_dc_gain : constant is 1;
    attribute mti_svvh_generic_type of vcm_pup : constant is 1;
    attribute mti_svvh_generic_type of off_filter_cap : constant is 1;
    attribute mti_svvh_generic_type of rx_pdb : constant is 1;
    attribute mti_svvh_generic_type of var_gate1 : constant is 1;
    attribute mti_svvh_generic_type of diag_rev_lpbk : constant is 1;
    attribute mti_svvh_generic_type of eqz3_pd : constant is 1;
    attribute mti_svvh_generic_type of eq2_dc_gain : constant is 1;
    attribute mti_svvh_generic_type of offcomp_igain : constant is 1;
    attribute mti_svvh_generic_type of var_bulk2 : constant is 1;
    attribute mti_svvh_generic_type of offset_correct : constant is 1;
    attribute mti_svvh_generic_type of rload_shunt : constant is 1;
    attribute mti_svvh_generic_type of rxterm_ctl : constant is 1;
    attribute mti_svvh_generic_type of rx_vcm : constant is 1;
    attribute mti_svvh_generic_type of off_filter_res : constant is 1;
    attribute mti_svvh_generic_type of eq0_dc_gain : constant is 1;
    attribute mti_svvh_generic_type of rxterm_set : constant is 1;
    attribute mti_svvh_generic_type of rzero_shunt : constant is 1;
    attribute mti_svvh_generic_type of diag_loopbk_bias : constant is 1;
    attribute mti_svvh_generic_type of var_gate0 : constant is 1;
    attribute mti_svvh_generic_type of offset_cancellation_ctrl : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of eye_pdb_att : constant is 1;
    attribute mti_svvh_generic_type of vert_threshold_att : constant is 1;
    attribute mti_svvh_generic_type of v_vert_threshold_scaling_att : constant is 1;
    attribute mti_svvh_generic_type of phase_steps_sel_att : constant is 1;
    attribute mti_svvh_generic_type of bit_error_check_enable_att : constant is 1;
end stratixv_hssi_pma_rx_att;
