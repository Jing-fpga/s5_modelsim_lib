`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P0oJ0UGtyAFbeQLwJRj22o/qvIkXgcfPi+Ls5SmZpMhU4dHm8cMO6L1e70gJn6YA
7nEKMx+nvQsKafsfmW39xISHALt0zG3w4x8/gEVJ1NofjUgLt7k/2R9lCNlNh4JI
sPWV4SdTX0JAaCAs9r//4uOKE9Zhyh6QH8M2+bw8ltiWaAJOzz2Jqq3wRrZ4oMFe
N+0N+u2BuEcDHNx3TycgeQtrNA4FDIZAyH1fLD83xeNzLElx6YTZd8Yz4KauD/xE
MFgBQtgnOfMp58cQODHAXNAxsq4kx1pBdFpw22k1DMCSR8tQdnuQazD1XgEjgnTw
JA6gCDR3Op5ipYd7fZPnEHrsliWKxkZznv1bl9Bmc4uGuHyRm+zaluNbq5ELc/Y3
HkzRy2O2/8ZGJpZhxStF40ouCyA5a030PuRCpS9NmyALYsUrtE0AZdWv4Pc0XxTD
KDihDP6C5TLyoSZMm3e3iG9Jzq6SzaiRwOUlVOXa6J4amkvL60JZJk5zrzmGjUR5
0cwobiwVQ9fwUVJoNVW1rZklolHjFZegXZRtTssNP0hGlDlwKpqmADlxgTbrxV8a
T0Kwm5D0KZszvwMxFISL7U6taoB7YvhGvm/VlKb62vfbia2aGd1BXKdA6vir5teF
vMYm9Mzh4GZGCXYgfwNAXhaOePBhcgB9684wmj8DW3hsYsO3GLnnxjffMWVDHy8E
yiJWcTXYOFek5YQMyf2cnc45Cbyjf9beEgjBzvQSjKhNJWJOUSBRQxdbZtKBCS+Q
5n6ViPl48YQdn5wgo3AjwrmYtkuG2wR566x6feXDtb6rE7GQpCoA1BjpkfWMzIw9
PTQo/rGPjuXmMfowqwQhARCSAsBD2521pLHAE68SbLE5NH2beaJ3JNw7tAL1WXdk
XXmvc9luraRKuLr93myrBBTa2dcIRSKoNKPIbnM9bqeFOrNhuhEkJJUm58kH5htf
rr2XihcMmTp4I9ajTFJYuH7dnYh8BjFO7j2adx/OwgYJABFSN7FL5X8h7dBHKaWd
cwUVli/MaT/XqUti+awt7cEY32dLBnoCVtCWX0i6wYvjJDbvaHdeM1Br6fHxTnqi
egx3e96hlshLEcdrVl1N8N72vhDN77bkFS+CV3ujypTqteghy/iI7pwTFu5pZG6f
5ZnS1WCMGTD2mkpwQPTuzjAUkY/9/bC7l6vf//hEPsCMIuU/S9HZHpWlc/HWhhg7
QF5T4qHdrdVS1ftI5n5ls0uW9oHOfjro4GLJwsVBI4BnMCdalN8QGiKy32tdDh3s
AyOrhhmFv/K+5r+GBI8BTz9DMWp9joFOWI90rWshbQbGwPTB7AWnb2zWIWO7sW5o
Q3m7GBbmBAxZJ1JXag/Kbf5z6VcpCPAQLRua38HjxSfJ6vOu5elS7ngVDpvhytam
mNeHP/Sm3MnaQpO60wXuwHrw+K9GPtY55zJ72RZr/Ct3986O1VxWUtKQV1rIDuWh
gVseFsNa2SE/CTxIzXtzGyH5bzbgHWLXXF/6dgoHqm9Ztso1DdORiciJ9WLhnObJ
6xuFbqxhNDp0G/lckP6ziwoL5f7KsWAyHLx9lVZhQOS58v+aQzLGr28Okr7NZQVc
QOwUHsAtbJQo0rXqiheFFanU0wrwtipI/ElKfoR2fRcVl5LWaDJ1D0Y7Tk4o6JGI
EHqY/P8/xxT9EXf71iTIQA==
`protect END_PROTECTED
