`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w12IHrTgVlqCffrK4qdc1FDDNIR2Yq7dkmjIlaSRiWu6BRwuruAMGPg+skjYPrVL
I9afN72wrWQKdcaTkv9+S4OR0miRmQgyEeFytEBpMqg9m6H2vksR//EXrFaWGakX
TSEi2HSPiWU4sgOL8FZwv+TJ4b4vV2OpGRy7v95Q2ytaWzWNO1ZaIYssB+pW4WR0
IMr8INxeEjy6D8cn498aXWO8lINHUVYi6yQ+FbaWfxt547pDF717ZICBK6q26iwk
+lSpinXrRlftvHN0xTTuXUyz+Gm5xpHRjjaIDT7WxC5y8PzzyUDsB7iJiWQA68YC
mW3b7u1bia7fJy31M0CYQqP24pMjpe91dOKJMqeiU69f8HVuIvKQ8WVOkvcfTFDy
5cZiB3bYHvg/hULkmgiywcinZbwVikcwcVE2weB8kxhoWds00fEY2kUQGql6E8Kf
yZF0PEjOiyAlqtDMtHpK4r36oZ0WQn9jR2tsJkni9UOw5YvzDe/rHwD0/5MnqboA
JfwUQNalxo+/qZiMuLTfCJoOP4hoi2v/sSl52y6SUyV7U3CPsNlgXAXiQ9EtFlrc
yiRFiBWJm/v83qPfY0EomDNZ5XprM5MFuUxMFHdUC7qa9D0Szv9spCKT7sqpP3B9
puzsSi/GgkURQ1rI3RmVvuWZzkhf1YsCXXQYZDBsmcuxk7VuNwhju5ZEWuoktj+1
Le74b1udVpK7QQHfsZvdvCRm7uvlXyqf3zgbCIPK4zGw7mx5ZMc+dJtBSytL3dwx
FOKtynJE2ol8o1ouhr5yBlv5SyLxSXPnBPY6tuT3dl3cE1janUnKK1616ICPUl1L
t8unHgSAAx//mXjxwRSQJcK6ZPGUN7Si/e/Pn+zbkB1JTh/k5nj54SUJ9aXgbeLm
x+DWHye2+XAgCbb+WP9O76RW9ecEK8WEo5Yd4CCd4Kk/xdV064ZLJWdMTJHtJvJp
B+lQSlDyUv1y85SBdxVyxBwEAhoypUaDEcHftsK6A1I5oFRTaDZuTYo/Xhx12ydn
cy3t49XJHkCxqY3ejWwOh8nD8NlElbC43vxYcTCdpblX4ocea5vIqM4EoK4LOMhu
L5SvFYsvDVXaW6hPzONRMxy3To3bUaaKjpEST8/NtN1sTA6Sjk2GPsD7Op0kK6z6
D1b7MOd8tLXE3BqPcd48Rc+CVNrBjqlIzz2utpFpYElj9aUHaD/KEVJU4MsJgMlK
k5cYRVDFud8aInYxGp0BluXbnPDvUhXlKEIXA8mDkdNRAun7M5IGp4FWrS7qOiEV
`protect END_PROTECTED
