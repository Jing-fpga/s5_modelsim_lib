`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AElghOkgBK8cFErOcWS8GuC11Id4tup3moF7SL75i1OlmfgGRo4yAp7lOsx/qb1g
soYJ3t9p0UQ4H9gFeTtPiaDc4rI1Oi7PD/dH1YdKuQnnnVRcrBpbSGVvEJodsflF
IGZlwpGXFb9jTAnLcwNdzwfZHh9JZqVPidT5lJMQ0azhSJ+TY8B2Kx3BqwTpIqej
7Xy2TBN8Zjhy0W/Yr42Y7nUdtoHaOO4+r9rRC4US69zJ0f90VlbOcNU+2iMCFRvO
RImFZu86wS1U0YmdkV0k2ifowoj3dwOwIHk78Uqu7xzX78wuUFX85D3i+Imx5LwG
noBEIcoQNEO0cl/2wg+p7EyKIdG8mRvpwly+/GA1J9nGfP+TO1rW0TZwHTnwNi/6
p/zCcUF7AvsiegfN8Od0uwJlzYF7e7QDUGe2DgjWR+NQu2tc6tJ0+Y+WL7TNyCPv
kYqzzrfLibTbeJ9Tgm8gVqD7EjT+yd/2nb36BE+uco8TpbbkpEj1iV0WvfdaxIb5
eCbWQXV99BFITgvCNvY4JCG5c9tSIUEvuCtm1AGDGxqaIZhsEbUBIWNQIVFfw9re
QzKpkFQBLg4zsgLnGn1K95vjlJrT7d87GVULqOOQZDiJ/lgJxLev/GJ6sbQ5naIE
bijdoGcmM6vIUF5kRdccG5dTaemDKl0p4p17qyBsrjlZJDhb6Hm4UdAl2kldjcRZ
Pr3G4tv9lABYOiX44DwpEBwMeXli9nV8dJ1IBZzZYhXujaMKUVKFQdAXBwv36Oxl
YvK2/i3hvRmkVHfCUEp3VQPDBkRIRrpaP0puxvT1mozdRmghY33JNwF1ABda1ErB
+uElocm75qXtr63asxVBp+kha14DpQ5Fpd9b6Kjg4GRPWiiwPbEBGw8EMtww9cpU
eg+Itw2ho+V8lcvJmSpAbXqCcGSIUH3XJeYw15u9G/JEguH009fGebyDiNX33tcE
oTfCiIMYD/c7AUrMtjBAKL+IJ6c5TBKXq5et2Syamj/7TVyd0ZJ4yEII5y++50W8
bW3JBCTWe2KXsfsYcM2JI0VBLTxUWEzOxCBaSaEFePKz8D3B5f2nxb6qcbmYWyqa
l3ugGK9NZwtPt9mrbvgle0XUUAtC45t8QZHA9fVj/p4951Rhs2s7B6L9+Fiqkq1J
5jnTh+qjnKhhmclMbK8IaPKnojomZ1j1yrOK6uSjn/5WrkPmsnnpbYTYU38Xgiep
mgZb0SftnQcPQ3Wv2x5z6i7RgZC+Qk0nFy/rDxlnKl/ZOtnOEn+ugdDmUCs7tbof
fHxDX8LAuyhHD/MxYD75pZiRrhHOK2dCc2uJefhHXbJl+wrWN00dueP2VsktL2Af
+6+7Aen4+jWstutXjZUvMB2gooU7vJjAcr1mNLvVAP35KS3Dg+C58gLx/gg1Gkh2
OA20uxV6apOtaVwyhT4h61hsuxYz0HZy31bkfYVS0G5pjYBDa3IHE+oejCRZpV9T
V4QjC/q+oILTRQkQR9JLH0o5HK479XjGXJtLuv5ixY5cFIierD2U89WorvCoux9L
QQCSum9p8/VQAvtvwB62+QcxpMde59CyeWpNa0BkKl4QJa8ZFcZ7c5lSGfZeDbMy
28S9iCGbhMHWyJAQpNusigplrq45JcB8Zfj3y3fuN5+Qcpa42z3noVnCBQ9G8yab
Xr5GzJS4N+1AtT1DR/LzwoUm1BUS4xtM1TUxFF5PekqlH+WcBZi1P7Fy7A2gfHz0
9OmqYudCR5AiAl5EtIQTnY7qmjlljcY+mVQOA166NsEw+JirZiiCrx9FyShU3gsF
OkQYaoSDKPmEIvBHy9TR0VrKfkZAFsQmF9ba4CUWv6IW0huxSFG59tUZ9DLY2x8n
ZPVROwdZ3XzAUeEZ+lXZfSnI/GefonHhCl2PgTUgiuvQIeJrWovrkx5JblKKXjhF
6LJfPW6lGZtYqvuPvsS4wQRlPZjuJIKVt7M2I31oPeFk+hznOLF4VvEqTSgWV5wP
7DBSRd0dPj7bLSNptwtiHbvV3n6CRF5isO3OpSeH7UBCulT5P+NDpen+02jZUO47
Dd69xy1qBcaK7B8M/FbxdgTzaMiAJpO3VIRmpHdx5b+VZbqH8y7qeXBApnp88tX/
n9I3BgyOZQ3P7fhXH8QyFmT3pre/kMGLlVZjZwrMDAaywy3fYKlQuLx+sLx3FVdB
ftdkP6+vq9varW8jW5thdqvVWCIUiKEiKxs0tYjSt30bdzxJV69cLTJI5J/bYCuP
hbnnEOfAwYQptV2mB31weCVY/daUQms3Br/rPqwxmpEC1OEfq0eXeuu7cvZ5kOg1
Yci45MN7fZmbF7XxHLrItgKMdKOappGPEhLXwKfl4i3KHwS8jq++KG6X8/5IUGCe
qmA9woOu7tXHvIg5KinCa72t4UBd+DitDqHnHiDCAbSDs3ZXC4TZ3I6YRo3LhCSM
udJDfWz486C8O/w32YZmYlCzbhzCXRb3Dv11274jDdrh7F6vlJvzN9WSGzgDLMWa
Nwfpw65qbjhhbm4yjGZzq2rLiw3CRw/O8It66Ril7oKwD8uasu6XqOJmWLzX3drk
WsQy7tJ6v8IJRi54pU5vj056zy5v/43Kgth4u669urkFQPjnrSg7XZjt417LevXs
J1G/8z12XABB+7+j5ivrRuz6Yam0NW3Z3z4ts6QoZClQiJ8eATTYezJStuSpS5QR
nZlLkFebHVs9oaQDzsEOVOws5g9s/adn0yuigIqL1rrxtjI1zg8HQO2Crj/acASe
fCgo9Yf9LUqZSihJlYLASTnI7L1FrxtReC5YTbVX6Nn+8O5f2BNaf75fSisQLjJe
`protect END_PROTECTED
