`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ec26hpIKn+Ey1KVsfZAtkMcyY/eoRWHXp1RBTZdQnBY1IWpC+mvyykfs5mDjwgCO
K0LbrlKW+QYS9iXojgD0EigkKdWG0S0SRnVjE8nZq7HqQo2udgfamKrzwycRza/P
E/a3ziPbF4QXNxtRNpxGhShAnho9jxxydoCUR90H3CJzXSB2G7DH8b6YS96ySjjf
Rj5Td6MdzCaNqETzRbR/ekj5KyRztQcvNxQ4yW/I9C+X1VtaEnhgtyVuGAl4Zbih
1C0eUf/r+AAJAsI1Jmxb4o+7IbUivCzULnlydAV/3fzrjgARe3T+V1ScNZlxKvJf
TsEBu2Dpmu5slqCloZjppiSHo6yyyXG1dDHvSKfMAAOUI6cdmmHA6BHGcpZy5A2b
/lpfPFVMxKCLrCU3PN0ALeN8oypPsBC5l2mMAC86nWfHk+83DaaxZU/xSYuiIUjQ
1au3k2tvmRtrbF+O+1cyf7zQjdK0VSVk4vQwnIy6A7LV6sA6XdQscMXOGS25mpOg
He1V2/adqmmANRPAdK0XIHmioGOXIKIeSs0wceKYdBl8OnaeI28OfPT6cxbeUYom
FixNNjRGwn726vBdDQGUOl1vSZaJpE2MXqi+543tzX5mjqxG5jvIAEiF695T4Ick
aDNrXgJUAAwlURwIJfil/X6KB7O9st1qLHG7C8c0TKZfOsK28DKTYZ31dlp7Zklx
8Sxu8mudQnPMilgx95ezbgpszMYWYvKazK56oBl7lK3gc/rzodcfQShr2TkDPmM0
QNbOcJooLXwWGb3nnqyysVUEeeaT1/F/LtgYSnlCSqaiu0ma63pZZEgQVQmH08zH
b+Hwc4Swu8N5lNRKYud7OnjelUcyQWHfZOpxVcvB/tKGLlrmgXQuB/x/qKxrFT0C
dzvIlCoUw0vEGabwp7swSkKbU5fEpdS53Byfxj8aijhHLmUiNTVt1uCpbXmwmqk0
TBv/ngf+VVxdr6+wV1+dkGTY/TCiJ/4c0ivKNjnCImNq4q1EaHOy4z09LF9ba5oN
8etpfNj0dAZCMMaG6lfZio44Rvcq028errqmiMi5Gmxm/ZGyVb971zhYlgpsj3ih
W9tWpBe3pAryeUn3YFhIKF4ZBuAy+C2Lu46t/kDQvHpWEYifsSoknQEme0a8TNNd
M+uIMO6+kcAecjZRzujnVE1+Jz2wkAcetGtPHhv2hXr5Wm8wbT+KiDRNw5DC3PrA
HQzZhXqexJi/BB1X5dge5S1vfIBHhAmUcyRTdSvl1fRoSBEzekGAddcUSddIjPgB
Bo1TXlDtBdF1Gjp/+O7Wtt8RW5CuJNTz9VAdHUoO6z2JRbxMv7ZaO+h/S3z7eKbm
8XgQgUHpKARQPy8Fldbe2Mu7SdBctwWauIeDahVmDwAOI81braC7V32jbBCcaaR5
HwkBSvGDZfM9xTK+vH8B5gKE8RPRxVAf4xQUwe56OAmYlEo+XGlbdzvVn2gmDywX
eA+Fe+NutN28K9DbBdBjUCjx24NrhjYpD/p6PXSllaGFLDHtLtKL6Ruj18GRYtJt
rfG1jhvtH8WdyLTl021+SqywynowAspC/YuIghKxhtItwZ8P6nFt/ZZadTQAaQxk
AwcQdBUApxoMNmv8JdptDvEXHeNv7Y9wxvMrpp2HlkL67k61L7MsuMR0EtvYZdZk
UOalR3coLRYpxbt/Pd8fRdF9fxD21XNTWG3hqHnvBWLrTVB1vU8+M2jpX0gG/XSc
Sqt0N9GIAzvJRKMMKPk13nInJ0a1vPnEvfdfxxhH9VyHE1xq5DeUAm/84QzkImah
6gWn76no9BNjs4gCkywH1z60stuMy4JkRbKhFq66gGxtFzT2JiRgYS5U/FbSIhr0
O2eD0z7EsRIGoTEFzVg9O8zm+FIcaFUFlOEB51AUhTu1p4/WVJFUjKx7oNb8/80E
p2fLrEg8dlvAGg/pf8YAn46vPH+vNdNDLTD+hLfol5f9jOTI2iTB/3pxEyCWs62x
mpnN1e/mPiu6sjV9tDWhCObC1kV9JXzzaVUrFA6yQADk1WWgwDH75ebe2e4isGaj
J/TJvVP4wD+me7j/saVkkZRczIbPo5h1iJbfPlOwkP4QqT3ADzdFUJ6aSgVf1YAs
aHdq/VUxF1/x6eX2uMOUkfAXRsjH7zkKJoTh6MFHxUX9bhb+yoe/NtvH4y+A9mt5
pDn/xhQPhFspl+50amBJ3dN19Ao8qPLolnYzE+KVlUOvNvsEcgYaEAZrFekBXq99
MHoaDHt87yFWVvuu9LIvfTO+T67qR1uW6CRJqIm9HlDvC9tdi+DMfaG3+ULTPdKX
DuCHNhtfCSgTPXPYEJSiV2cLWLMgDRko3YpGQrZdQMw3I3XI/sGlWMgR07bsXtam
EmHtvNcF85pNiRK+qXFE48D59qLOzXilXjKnPCmKE/uOSJprDCB6HyackYP2YRpQ
gugKJAdu4GmRZCzyOiQgsPWkKNY9DQPT/YpjDni4LucagjTlSsC/irCG/4gHsUdM
kqYp0J+uW7DXmQ8yEBf5EXYx7cRR/fqwIEa43v9HshI=
`protect END_PROTECTED
