`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UhaYs5B6FlXsouq3/j88lIkPIHgHgZqHWwOU+RgqIYjfheqgXXAjyViK3ixWg1WT
IYhkMHWdCNSM5w50I24ZdL+aFrgHKy8Svtiq8swZuZ9HFOMfBqGKANbwTsgbL8hq
rQ0ua7CiMsVHSD1Bmd8cMmOQV0pOcrIPohSci8t6pArhcb9cW1K7af5Cy5oKoyTj
QoVYNTBuM+0Mwu+9myy/LhzNMb8ONVVCRP4Lh4h4E5Xyh9xN2bXZLVF/TU9ZZ0pO
K7RMNwDwuWxupa6cMbk26LYerMtMUkH2obWl8RK36lM2aRMnjCCj6lz5hEupwslE
DvKh2O7iSjfQQEcIKWqm9VaJfg2mlCPFvYm+OfiwGWkN3OhsityCuSK/Qye/LL+J
GXMEzlSjTIsuahhQGl2q/Nx5DraYSgUSTpkSh7fBdUqCW/tHXotfYX1oiYp8ejZW
Gl34YBeghedtJAVbay3DLyMh9zZJluXKcdKrLnL7AT1xjxxVYYR2RferhtFOCEDY
D0yxxWQgDnwWhRiXp2sgLrglHXSdTzL1RvHdcEHgqwx6XeMjwEzj2d4SF9lY4GVq
dT1Nrj9jE6/pNRwhrLkX7F30n81e/nn6sT3GUTFTmwaXh6F1hjim/rgXgqembBQa
Nhxw6BAo7c+0zAoCJXFLngQi5rOopviL1Os+BVXMwz7T+AjFNmMAOH46DO1eZ6Cm
e2lkNgx6V1EAlip2BAORRrWwqhTNHe2J8xCoiiWPsXMHwJ8lpA6OyuwTZAgYd9Sx
`protect END_PROTECTED
