`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l1sy+6uadW1oI4oAn6xoTCn3dYNx/OzQetn/kYXE+bSAGUH/b6xpIHCFwAIV+lMx
i+qD3+K4i8XxVWyj/RAneGo2ew6zQvyewCygmX5a2exgCplZPjX0yWX1ynbqRT2P
VoXQaYZ5XvgUNmYbBuHVHPqG23kb2zLf1ssHZxDsiSsAC/qz1dY5tjHfjJCVMyzx
YQxw5HBEp83y1Rrbu8xBRuN3zjTG1gSYwfCGqQx7E5/ivJ8Oc/iBlc9LCSaVOwIQ
i0DV8GDgm0hyULVR5lK3R7WvICaTqqIvnQTVZ3mIKPeipkxJWq89ozlndguwwRBt
mHvDUMAlew8XBjXHFK+QUDnKztdu8tuKIqywX/XWpWBLDqsCFqn5WfjM6hPhA3ab
AvSJ7z4/dwIBSgTQHBqzC1bHlyJWimL0vQnpnJGyO2VLz2/4Lyb21yXAZjqA06b+
dwDX8dzMd3LFkJcaezeTB1GnKiwzq0RbgBr548ZyomDMMO/48JqnWwVXNAi3/Fo1
ydKlF+9TO2ajL52HxxWHU4GTR33RnbhKEstppHLGWCbZzTNO8HonWgwuY5jYWOZB
`protect END_PROTECTED
