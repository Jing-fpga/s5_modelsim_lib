`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VgfIis35NN3cm+DWuRTD7kDiN8+p5N7VZ/kEooIbPXBILpEcRWnnYbeX5vAOB5Lv
ay0HSEbjcBvRRxAo+wWm7iWvJWMLJz4l+zdiXR8t2LkoJokZi1Nlty+Gcs0aBQLv
bR7+K7K2I7JJNG5rQdrVCe8BlyeL13mA1S97ylEPXyJGsVu4dPI6T2rANyxfA15u
SOW1r+yM+eU3rh8uZVUCZ09Wqy6xchvQP/KHwsEAmBITfM3NWnU6xUdUykVtkqbw
u6CZa4PKzJfPULn9ikcx+s0p7J7EFEGUCNue78Sp75A6yJx3k+3W4bYB4qrHx/RE
zMZYRRZFcAsYiz1upgovMI97fDRBLGUMQrGY+Cootv5IEXS2iGybkIqz/Udz1hFm
DfN8AuOHl6wye/jR+cJOghRWOkN9ZHUJq+uDG2naK7W3UyL53tRT+gBwSb59PMc+
3NnmjDJ2ci0zIICH76Wq5WBm607S4Wg1r9zDCt/fpufa7PdqLpxceot3L45n7ij+
j7/DH7lNVztP7DkBc6fj22udDOEa4ypj9TcXbnq2VLKT9h4x7MOUXw/R8ukQhtjx
cczRFGkFAw9LvhOwzW+8De/d45ZH+2dkA6Zb6HDoaBSfYpaJ+8+0Nc99m+/5Bced
w6PruqbvhRuxrQZOBRELx/ps2XvoRr9n/xmoZCrdqaTL/FdmfmFCcbBQI68+7iDX
NExekwhHvRwsjycOdE7r3stiy3GwMF7GQ/Sg2AGGPZTUMi47OZY31T96jPi0L0DL
kqjcaZMSbPqpFBkElMg0LHdSHCM7IWwHSWlJn24OerFe0FHhBdmOVFJ6w2CxnaMJ
GypjnaJFOtwXOk/MTokRhA==
`protect END_PROTECTED
