`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZVe7rTV8iI/9uBI0BtKVyR810sceKLd+OobyW8AihW5M+Bh5DbpefQwDE74IMEWe
/0h0je3TTTA0mGefCk5Ep+3P84ENbNgdXl7Ewq4yfnWCIXAv2mEJH6oX+yAOFu0Y
QgTiTNplYUw58mpnAOkIn7v53VhK0WdaVgIlhaHQ0hZt4JFSOzUx75P6gboLcLyO
Q75RHtYsxJ11YnNcaYhw2+hLmP82/G5AtgDfsH37vE83Fnr8rcC1/LkAjmn2C1rW
BzrB35QlRSF/4X1Ql2q7p/SBKINEhtJgu/CzlTqbzhxejzFTaL6/xgWttVvrhLuT
HNRVjEaFQJWOh2W4dZ/TKJgKhoT9qqZSftv3bbb9EgH02KJ5PHImm+MD3kpYvlfV
PLELNF1uMOe7UxavmocsqqRvHN7gZ0HTvndCeBBWjWToVelzUbuRAx1qhi8u+hBm
e6q6r+NhsOeY5HWOU37On9yX+2toGlLxLjuITobkVVu1hv/0NxgK3oWlk2udw/rM
ZO3DzHGGNN7jqFV5DCxoE6ctogpUOinK4kisz2P0D5y/fGWldbAijHQe0Y2WsAS6
+d34L24G0o6HJPuc/9mI/RTVEcmPa+BGlBuvqpDGtl/NmzB27li+Dbz+hhwRFYVA
8Y98nG7RZw61yTWz1BaC8+RkA2uECrDGCBc5v4pNdq82T7DxBFF2HfshxlYsz/AR
utImbGkXxlYicUSGD8NlJ0X59Sqonideyv6JOYzRJApQgLTUIDkSVPVcdARfPnZv
1R1mvzl3Voz+FHx5n5NImGadmod55mQApONfwVB1+mBdlqc5GPfwpTs6J/Nu7qF8
ZXW/Bp8FQscxxSBfqFvbVOQbKTcUQ6/hnBX1Xwk0txiJKjywZTYRv67II4rGWawJ
dzBMVLZ4wI2SsGsI+7qYcjL/geYhF9Fhkwj6w7QwOidVQtrUIoepXjARoycQydFu
07d+J5H0gh0nIhgOd4MKvdUURzQXNLTEL4WMgscbtXwqgQPMTWx3DlIrQxTh8EHe
4JaKQxFGVYRt83iF7FiVN8+xkpbcUJAXmCvBvTwbJG0o0eXbIpBveRuoNAcJTnHA
x8R/8OPePFQajiLcK+K2TaEVDvpqzl0xbXCHCQqpx1tRd/ejKn9WyUl+6ceNDavL
UHHxhyeANHGS/K1NiPJuXSEpfUpZ/iGKmiaMIzqNYS3bogicWAxQU/EiwpKnsEHU
NuYpjwF1JDJzSz7lLvnF+NJLJtw9CEmMp8ntpRgQNNYj2t85ojF1CF63CW+GQqYB
L+eoWecxhsiNNCTEsd8HmMxZXXM62EUbzjdg9Yv/HGE6XtrGt/Kf1LwWCFxU225p
ftOIkRKxHhi5fSe7LfjUw0JVsypnBdC9qe0ToUTaebAY5hipXGRLt7kLG5nXRvXn
e4Ovb8t7Uotextj+EetDsn+V0bmEvQXsaul1rWsePtyP8J9mbR/pkLscOthW7k8/
eyTANZwA7LoMLqUC/jOyGJBrtY+skPi/gdRJAvGleU46Nbiy1EPJHlZkH+x4/qP9
dS5VR3A/3CctlZwvwfhY9GSU4ygEzgNxHj1471TpfuaXHI0EVGMvP+hpdormR2lB
i/oJK+0j6EqxjL+dYKlHulSW20hfY4dksZ+5YkJJV8Q+SLjhMpjf4PO7LMtSO3pG
WP9QeQIhLmXTCJX4KC/0UC2ACTFYAA2sftbOJvV74Mf9IXBH3UUjv+H2isybxNIs
MEyrLWBJ6yFg8Pgny1ptc8GxJjZSmU07TzSyiuz+sFLepvkK8gWhp+nHv1OK626n
/pGEwyjWdC2HaH+xvMfGc8L4wTxbI4RZqat9BhY+oXcJOB1jqA1IlWNYJg7+UH0Y
Yg/j1VF71iKvWYj5yKbZVPEPIVJWhWP4ODlQRxjUzHbCjw0nQ4uYYWm8jpz+hCJv
lffEqKDox0dfL2XR7fupk62AnIis4GZkL/Mz/ZLIdos9A/DkS7LYWAsN4WrVbcvz
NkKiNmWhBJumR0ATdku2K84C1ouL9kB1M9znrly43zKOqaCti2AEYY71gYt7FSbw
WcJjaTY1iMxuEiV+ifXjB/MSwnJMAx8FlE92jbUPQANB+FcB0WU43QXqvUFRMgVU
+M8nq2S1fgI+tTMMHTHtuI89+bMq4zgbdkKPfrv913Hx+ZoxOuE51ukyvA5aPyKQ
x4eoPjSOiDIN+N5BeOTmtm21OkxgTvGq/gcbyFeROaZEZqTSH0bvKFL1H80rZqyL
UQ4R3ota8i+PV5qySustxlHNVQeFgd6VbLqxQVc1hCw/4JJ6HfUpJWXuIpgQzX89
AUb7Le5FiUcP7926BgkdjcC3oFb2JxoLbedp5RtdY1GaJwPOGoa6eCphIKoT6pnX
VsQa0EL4T30O7wiXQjWTMw==
`protect END_PROTECTED
