`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hpiIWCj4e67MtClsG3L2gWMEnGh5hkhG2JU9FZG9D36Yu4ai9R6t/d0hueulDtyq
exHXZiMmsDkN6XUy2o9DowS2DgiWAfcPCCsnh/ch1ZiJWCnGz/2KmsWPgIRn3nKf
RLnSQjBW3wXzTcZ8y++jNSH2VMxuQS35L144GTbpuqjrbw2pFH/ezFjYiVFgH/ud
5banB7w+B5s81UmlXdBAvW1WRD2mez4AuUOHrGDO06414xxv2s5QZQNDI6L8fT7i
nbFmlUCIg2wjxdN2niESxIGicbQdoWBz/mvxlKOJ2lnqpIYiUxRtPSuO+x5tXv6E
2MmvRXJLEHcGwsclY3yadw0SKXUzweLWk0i6Z6bIdpF53otaX5U3CElRqk0ypgoD
/skMArwPuKgKtsIdKakzQWGa9uMfuJ4WiomknU7awOTaP7Qg9dg3bKIY9BIZNgHy
hHQg+fWnlMILlnvPiEC8UtB8DEZS9ucYm38EO1Q5DWdUGlxaKerpod1Ncdl1FJ9T
+/JLkr/zpiVqVcW9tkwOyMYHYij501tw0Ie8/ohUz1XO37+UPGqkDVVZeaC68W4L
X5zGeoxHRNRSuDBCf4JGdf/r39w7PhVZw3uSwIcIkC4d13ZG+bLMieot/q1XCXZ8
VkqxphtulCrWJqa3cu9ofPtVEcC5AYfpE3od5S4/Gog=
`protect END_PROTECTED
