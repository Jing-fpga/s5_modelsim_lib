`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YqDvKVRPxlfCohnF0C1Pcqmbzd9M9meIgU9cLG2nteiDGLLufqyxXFP12Ehhe2VG
V6D5boBu4+d1Zlool08VUv2ArFkbjPpY90kNpTxV/GWc1Ts9Kan/ApbADPt86kLP
BzC9IRXExbyyi2i/W59hqZ6Rb09lxIra9aGu1QsNlPreO2U/PTq+HaOQzssCP1Ud
pSn+yC82+UjpOlyC8PQbJIbuOUJFDYTnvdGqdVEmLWvyJYlWwrkjV/nppoLSf0NP
hYY39r9LuIkj/oMv6DCy0s5Xc6G7Vego82aaa5znxHQBJkIXgFJEJLWjbatQwVv+
nYNjWz9b3AViCuIk7Wti7HgOitFhCCqMek/KhDkbAy7wp93Ph/XIL+Q/VQap1QOk
wyoVIoZBbdjlv6Npo2gnPEBVjI/v92rL8zFkEiX18AfPX4IyBJkNXI7Kw6tjK/yq
701txlzQHHevJ2p6YcWvUKWndUi90xgTTN5ztfgr7KECjOC8qMbAxD7FkDlTqH3k
mUPgcLPg14TBVUBcEWf6RKMAVTjUfx3N5PCeoqY7gaOEHAqwGkDGlSVWFTmFCnvu
VK5KajqWudpW0zhauUHoc9QvHJOLDBMP9knE7XUKJocf+h9LsQ3j+MRcnfF6cxAe
5i6S811t99YQqvfmhs7Xrzzf7u1KpaorUbiKShAH7YJXWM8JtA696rjqWiZw6Ocr
avaKXGgnpSwmuH2a1Lj9/8Nv/Zb52cB1NNyv3DLtFQAcgjK2JdiO8zcQoRauMMQS
OkjgEOa9nlw2Pv34nIEBTraNO2YPaPs+RekDSgJzC4Fe2akGaR8nORyifaZS+Kvm
MVGjx1hZFdGpMR3X7s4Uy7n/anysVc4srQdFoXgzc8v3Q75zOFgeOx/jFYcDIp9u
qwG5IeexMset5Jr2DYwPQul982CfwDjZkdnCqJtEqZDcIW1aebUeLoCRk+a59qCf
+76p9/pEPZNwgNaEnykE9GfvcyUvI7NIvuD15S95P1LdJK9gCssjsOYhRdHHJyBT
0MiyN/MahFdUDqwt6HYHrSfzZeL5B9ZxJ8jP4a61WVGi75+F2qdtFFQTrNJa+BD9
CnK986RaTpi17be5gIZ1cGed4kcgpwgslHowO95yKJuCRIUPDQue2+QntWP5bgx6
XJVTfUl7regxRQYP3u4/Aq/5sSY17kR7tZHupCacbM/0vePoY4KQ6AjerVPFGXWH
cVq9jyHqYj9PcfIhGY55su1OjvzgNZYOEFmj7Ltq1ma98KRwb/X+3/2/gJ1nJfFY
XzCzQOAyAtluXTh2yUDX84oGqlE1VKhMcq9FSZ4UuMNFT4xdjncN+975woLBhXkD
ASg71Q+7aiyLekRa6ffdMZa2DkOA5gAdVYLobEN2hWfTL6nGPgeX/gEVhXjE6Xl7
ioGZjObp+b/VqV62WjOTl654nJIVgaUgTZIb3K/ehbQ=
`protect END_PROTECTED
