`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gZkBKwgvCFeFFcqUfjEmR5iRBvrzJtsyFge8N7ssXtQ72goCcDLRlQZpzaukx+82
T8xUUdDi01HfT2SNX++oBGOY+WAVRd3fcU4Wk69hXl6ozjLnBaKB7tFlsKpwxTuU
lCDYisskdcnmB5D6xkKxUw6Xh+sREEK3GhjP+gRfipWN38dIkU2q1P4CTi3BGWbQ
ZXwbJCYm/1KvxcatVd3UGxbdx66etNoVdyveLGjag9LvoHiDowQugQ0Nq5/s4SWC
//lvTia+o3OfnaVrcGmMzogP6+ma/PWPiojrjOYFIYft37I24Cp3UQ95x7ijHvNd
D4TjsMQHwGkSblQ8/1vlMZwuk+Jkjd5w0Gc4Y3K/pHmjQZD13hllMlX4eekzGs+Z
CGvSpWF8hm3rAdzchU6IiMihgABBz1qI4oG0KMZ9sISrS0h0LWoqyOAJHD7kAGb/
7SAY+fiHaDX+fUKi+ehA2gS9WkNTazckGISbD8xgq9llmUZF+vF8y1oqlx/w6H02
orlMvJbw8VNAPme4LhdXNXNrpOGCucY8LnbPKiyw27FQK7lB6Vi13MsIkAYf5Gwi
4RDIDz6lzN6XM+kic/vQaPWhMBF/ovzG8zI/my4e3ymqf1YQ1Y6qfUNLErNyzy0L
Dbhz6LVN+6bGMK/urFxAdrGNIKD884kDGz2DEu7ee1f283xwIUqVjVCGPaU58d9i
mzwDxWhCOVN466SudId9ZpqcQ+Z6EdpwaV2ayonOZCwPtJHip5ie3zRe0LgNN+g9
mdIUBPxFdcTOCxvmmwR32eFmumqhzqXgBrvNHm/I4bKhw3+JUoe5sj4aPd1Ws0xg
guNGyPPw5A7hoGQ1cgROl80yGwFESfBVxlO32/hrGclXGuoKx11GvSwqZZCTSAQR
le3S71bcFcOx90IQvVkgD3P4oEWsYjZoNNU8c0k1x4o8wCVdZ2ermDZ9QPgVFf6H
Ik30ZYAIQ4uWDQF4oyt1CkmXAsZR9auBTQjnbuOn2fo0XuEN832yk6MeaNaAwciP
90jhCO8JwIag9T0Lwo87tqy8xvizixzYPuP8IB2Yc2KRojrdP9CqRaer9O1Id002
tCHQJ38/DDY/vwMHnCnqnxBCIOm66s4zmaPRHPxC6AN/P8CD3/klZPedrKH2Qikx
NGNfHWGWVZZYtWnpRwgTacMUEUXuWvgv7qOsquTozWUA2kz0pTAyRD62li29UiPe
NzRUTIJmlVswsFSt5682ZVAkhFnnmrci1ZQzoTO+dA+TgaWMj0MieLP4/myd/Q6w
T4WgmvcvG1CcYTjY60KjjVhWPDWJRWpncDj6+eNlookCgb1U/6z7kpcsOiH9/oj4
xhoNEwnCcwC4C2FcONy59WjymN8gwDP3ig5zQtCqwn9dqHjYUKw4TjUOAmF5uHuX
TofPUHbZOYK3Ei86nBW0s4RvBGYYKRRDsp3SPFRNOrE=
`protect END_PROTECTED
