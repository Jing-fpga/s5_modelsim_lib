`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yLTP+6nNj8cH62u1YlJ6mw3rUdvU6Zwz0PHFNV+uSdN3a5xugzW4k74Q8nTik3Zv
/WKyhLNFm5IGxnOMUTgcGeF82iaSmw+bZ02Ji4mtosl+kBcGmthcPIgE0UMKXYSI
mwj9NXfD4nsEcjY+/2TGPMy/ZypGtj0y7N26VRilerICBiJHPPvXnRaB4KvGbm2Y
JyKt9Qk4HPS6buSzr0hTA94z8PNFBfuehwj1tnWN0aOfeAZ3ejS7u7ZuheqXUJE2
P5mL3Tnwz6pJBB/y1YKMbmLHPvKTncYZv6guFjM+q9ngovtJXjO55dTa0G4d2oNo
RFW0yKDnWQwaiXu/r/roGomNaYR7Tkr0Ie6XfcIIRDQi4ysCRfHxfc4NL/Zvo0b2
jSh9N13UM2FB0VcxGg0VvS+ABj69MBbbzBKP6Mn10+kQPtCjeH61BtT6FDGwuBqU
0zGAf0/aJd72GHvwDh8kArIkR1N0evemuRwRGVxQaBpErqvVRe6bY5OIQNTMIJdb
27F+1+B7kBAYXirnOAkDev8fkgT6u9RZYTkPQuPrKvSVvQDosbRBP2EAYxJqAIA2
IdK/ZV0dCfKWhZVuS5zSFoN0KePm+9C4dhcQ2lOTYowf/Q4fU3GIXEZ1htX2Q24I
E/m2Ra/A1QJdO/djNXUQxqLJvInTGDiHXdSwxu3TFBb5B6GssYuInP9tcgK/u5BQ
pxP124V0aMSArxdcF+H9rKCszo2aHpho9Ev+qgX8eFxq0jnM8qPj0meGrIKuZJFT
OCNlG7LDhrlJdkryJGyerShbEA374t35OHIVV/dFzv7bs6feyP+bUsoPXxHEZlk3
lsqETtSk2lkfisjOSp7J9A1k5TyQDzZCmZhCgPcN08CkxDaQzyZh+2D/wIyV1A28
b4OP13lXkhuZBbSFzqPeobJK1fM7n9m+R4v49e+SBJQYhZqwqkUU8r5U7UGI2lC/
q2raWQCkaRTWYcOoV0G8su9KsG+l9FthjghfTWWA5fnnuMF4G7a9Vj6R+0Kg/tGV
B8DkF2T9axIyVniYqoDeqhdLUa8KJOEM09PT1Djhx6nBdHtlklctIknzaviUCOQS
gI9lFGr39JsKkWrQlMyODkizIrMYk5oQDA4MqevScG5sAKWOMMA2h9cx8zvtTP6g
vyEGDWWC7Ny3r4MyJVDzS48hRNQ/Xf69YpGaXdRzAU+o/6se2Mwq1o+I+Y/+JbyB
3oNf7CUa7LnMY/X1L+mDEtN7Pdq+I1KoadFN256OPVAHXLdqVL5iPyoGcgZSGdcD
MVSfUudPJqYt4o+vsdospV45X/NV7GUf3zWDDX06VBLaOVfcKu2qyw9ahzpkN7hK
7fMK822OWbNXnE6Rkkg6bSFSJ3Iyo626BIy67s2mJcr6RuqsjKxn0fX0AgaYj0oK
VYeYhWuRYyD3AjgIimm1NeCHXUkf/lbmkDAhvx7yyLAPoFLG/vRDMp9aU1+BQx2A
xHK4kDRZS1zcs4azfdN/pavzNxJS9FW5SEqemzSeODegj6vomJd283NGoiFOcSPo
MLC25xbbOgxt7EryvBpduh+rXoJCOB582pxiKRruJdSNKbzlP76bxjWFny2X/9CS
7xEBgtdyaWghcTl/nRH3zNryx+rmbzzux5sgnchxRb+gC6+2IwgZLXow9VT3yr4T
YqH8XUUbdzqWOGnf386oW24Eb9pV2aqoVWQuN9hmUFXXjlRMR+f5f6PsiTqkGWKC
3wQLvJeygFAWnveDA6l7JYI6oaac0PiCPkdsuxFEXoYEqvCcrwt8VcxTm09NpOBQ
jZyzeEBlIx4IJjO83Ddc2AZlWyZeILdBrtEgEHxsk8+Y21XFPYnDHNOX8IvIcP/a
EPON2ysfAlNDYsSSTllEg2oQBbzngf925KPJQtRglWIXOXlU7Zb+8KkMmT4b8Rkm
vMBZIym9d73Ouw+C53Ncnx/MEuZVzpzBzsHER3iG/wfqHyl82jtEdteqB56MYLlB
laZqvCfacoHKyd9r9X4Fu+dZ3u2UJhYkHI/ahExf/o7ha7r/1iTUIBrf3yUjb9Jy
MPJS88KSPF2cjV8wU79Mi1JrDzkCZBOe9tTI/zIG6qg3zV2DQJuL0wWop6eye3El
QAw9coTFXlamrLxmpH7EE6RjPrenDni69LmY2mBlYiv7fGMylrSXzyplrSfKh2Zr
WTgnGZzi/KnlsFUYTkuh0Kg41YLE2a/iowAqPq+TJjkIGxDpx+Vw3ACSzjBdQZKy
4ytmIa4AKQCB7wRbHJKQf8xVv+LjyV7GPT0fTQxLK0rSqTsK0RVOIccv3hmER2ZK
P2DynS7gp2d+dzpqJbkryw==
`protect END_PROTECTED
