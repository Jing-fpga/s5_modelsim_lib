`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MjJDVH9Cd1ZfSfuQ5deGsezF1EbyjcrYcXDk+s+qE5DK3coWtxHZy0VJ9ECRQOtT
nDTH3FlwM5l06kFxKtmR/PcoaFbSQaNHxHRxImmbuWGciDkJNk1sq6iRM11sspY4
dTqTM85mSPPn2u1KybUYUHB1wNpoBUxZA3bmBFCZ0gNETdJaX3MTZ7uUw9taWlpA
Q9rykW3oNjrPWyHqTNCN29hB5I51o4jLmCg9E3F2FSZUtVJTnxleCcDGWCM1EHcs
0GPylUZKbQ2FEX0VMdvBMnxMDt7IDdBbLvI7INy+BjlyTFMA4oddp7O+NaZjAp3Y
5AZxtgHhAe+haAJWNaGR6IQNmZ1eldaMZdMvz3l1UlLRMtab3TjMFfRa02GtLMyW
IJo4cGB16j8/IBtryDEXs6JkAABOUKzMPO78zEBJU3yWCU+qIRU2N04psfThWyRg
AukdOvEOXj9GUi0P2PgJzmG5vuru3hqxehwtSLW4ZTP0PBjfgYsEI6P/+gEfcwNr
Magfpjd2f6QIYqpsMFgSJHgoPnzz5zvraB66U4RWhjwRVFk6uRFvmNV63OV7tJoF
5QTMAMWZOMeoIrid1/G/YOHRzkXcgWdDKZ+YozS17/EVGK+E4LVDNyNMQzTQ10Vm
afrOjPDBFD3vTMiyKWLr2JaMxr386JZVcclULh9c2831nJUHoK3bj/B2v/vf5kD6
mENctEZFkAFXOgu4WEpXspjsnmaEcffwfW9Kp29HFEcT1z1fATENiz/a6lhfASO4
TZeMA8vo8qocy9i7CRjYGUeoAr0Md5C/MPbkiqTyASnOf2mrijNP8xRrPHxDeFpN
EApWPNKoiFb0lZlJewWKy5o7JuBupTWMSxuWORsRkjfVeh5jFsB4BZsj7JB1JN27
+qCFz/YC+USd+Ywx7zsZj4gfnuhv6ESrupjIgeXXW8jbfVA+HiAqVsMTQxOTK8+6
flBpiPQ0/GDoW5mATw5/QxCEa4f0z8AmNj/EkX2dyz1X+kATUGQszb9xI9Am7wId
h6ZaWDv8+jOn4qQELlsAOgUz/bT/5wyCT9VhQ59Z0HQBTPbDSoCvse63/Botsc/b
qvRXegdAsE4M063reC53UTOeSQwOqTRoVhj5dcJLPNwgvVBjVm67UQRvG/svxizt
CYha2v3ioSmRszzgf4zfYxl0k1r8FN32lOA2zPa+oMB+A6sFqQ0aH66lYVP70BSN
kXe0BJjQvNMKus/VoRn13DthpRnNQ/UjoDZXITRt0/g+DUWCjnC22bcNuxNhZnTt
290nH5gU+kczoftqYkNFWuqMtnCzvGayz0LihiB5R1nJA0Pwy/SZSK1BLeoP2fdE
lQ2YCtMko7AsW2LnklskYluYzNq9pBnQ+BHU3LCdF91d8kBFcoEy2o4gp7TB91Rk
Bedxcyt9xEbswf1OOPr/Md25uffhCTJZB/wv+zE/gtpYpGJC1wXTOHpzzoGACbGQ
33udCr57NM6eEUiCWBpaedpUBWOvYz2V5uaasKrUXaFcgIL/MwB/op/JAvioZx3j
84CJFJxlZUjULGLAzAovfwMvtYeYtW1zRDAl2Ol7I29iwx8qc7NUXZun2UiPANII
bu4ebtu9IVBGbMjJOdOMFi4HrAhUA1IQdiV/wdvuzF3fuOcdhUqLxQED0xv3DndT
oF87e5oxLln4YSD5STvNiKurqw7pTNJ3IZzNnNR1Gxe9YI9DbtCuNXcm2J330Ye7
gfFusUWAQcmHw4ikN4p20+jIkbWJ7XmcgRTcVF8XxGCmSYicQVpKUGqbn/W3A67f
JbiawjuC8m3qeIUUnA/e9ZY6kbwNJLYrbTe6NswcOI4VRZC0vgTFP5NDhih+WrUt
Wo+xKkVzL4ddlichzADAlssgpVLA6YGDMekC55KYCRMVnDE6VKHAF8EkwwUgaTNz
xVNA/4a/LhQJWjprHqmpmN4zwX3FCm9KSUsTx7tFCYtm0YFxu73hkiiAnLoIMSpZ
x4TVG6wf4mnKWIp0DkRzFMmAILO53fJJvu7KqqoYSjVHlu3YNHVYlY4OADEil/9S
VZyys8ibrs3Z57Laeph+9gcmqspFXpoKfNK9v1zmAmb25GYyqkWyxMAFACvo9PKX
s1DGGvKYgyICPZx+v4SrOIm2CCBPgzfljtcIcOom+L2q++8IBj4SeEYwDRp+E443
pI+yFu+6LVCJD3Gnmf4mW6PYk5+NJxjJakqYXibCzsS0r+vAsmIKL8y8G4IQhlKr
QltXdzJYceQ4A6yhzDlxe0UlSmQxx64snWYpoV07VuCUm0Csb6EFOi8HC653YLHg
WnzjUXeLYsTeKtJhOBJGjmraeibi2V91TndqX2PIyYVCgMmIuqbN3pgbru8HhFqc
PGTyLpuKm6oC08377+PErvNjorEDtx3gYyT8HtmxHPrhNCu8ibrRhLiuRZIkX4ti
gj9enjWRzMMF3SSAOSlNuAnxxf5aaY8BpI6uBrKpCzjHwBcpgIDdijAtdTuM/Ako
MxxoIM9a3N0ipJrTq8+CjsJjow+x4MKwX3y2JWAdo+59LJBBQbpVD2hZRGa2ylhN
QTFBLBoe53bTV0dbc/NuBnwUNyjPbXc6HZlY6Op3x3GWNSYPMuz4TcvfFIpHjYkE
ioAE9K0qAMWWanx5ykSiEw==
`protect END_PROTECTED
