`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
btaIGxOXFuzPXY1kVwZuV+SqP05HTSVykX2rd21DXw1OcwpLhL1IOkEZl3ixc623
zaQ45JDGF6ny0NMY3aJXZIssjpm9/DuYXQRZOBuS0+HTVCfwvW/woAaj3x/yHvY3
1dyGkUSm4J0oetpnGQXOAfS3mI2ICA+WB2v8tMxtg4DkgfpLqKVljtilumfwwqma
7nofSd8ypThmdyUfpBmvwQV6mQsDBWcm5ODDIVamaGRok6iaJEb0h014cZguL5sD
+l3+zrTZeRLgeYe9BrmBJS6OABJhOgohFgOLQr++0JtRKnUtPnVJNTKR5UZfGfqT
JfQ0ZvnPiXKecXlnK8mtroDOTJQQ9/ESd1ORD4ENGABnjUpVH8/1Wf3xGLJ2YQWn
T3sp3Bs+wLOi7hIL1CGaO48FlzsvF7p2mFXDeGe2ObZI1QoOnqq4OcXGPOguT/xl
XKkl1hSG3dilm2ks+6W8R/C+KYekcoNRyn/avTDm5EcG36fXFg7yY0sLOfQ6oVAx
IjcJkPwFwEuXPoZY4DC196myZbPJKrU+OqFyd3YMgF7E9728FTeTGic15GKt5mjW
AdhbLS76Ng70SziYfvK6CE68BH0azgGe8+PB9L1+r3f8SxOZ2RuMPm/9+wGpdMvf
`protect END_PROTECTED
