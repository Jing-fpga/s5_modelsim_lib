`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mkGf8MJayqxKGL6VCH5Sl1vAJ4R/lf9k9OfTiqaljX9035THTuFn7aetymkfouUb
jai8h0JCTFzMaVaA5guc1Po0Drdygx28BMH07jfp9dGpxB7ehMSHYYJcN1ubu9/d
YDw1F2yAYxjmqGMH7GU7KyMLXCqRAiGGgZxF2RailS4vCIcBMpxH8UTksxsRpGIR
fezw6F4U1gsu8KRREXAqv2jHSeBfyy2d/vohai/ADYxploEyujrwZj5UobNCq6Eu
C659RJfRx29m8SlXJKToO0LELMtBwkDUeGfTnpJJtrBMS3NzRwJcYYop7iREvKiZ
FTgSLh3ziCOpqzV9S9Bvg2YRphPLTWiiI3MRAWboHnOpVWc7X+xZYxCFCDJenZIv
/h4l0Yp5D/tTEWQOuaDq1Abd9l6vOcagEsj11XtG/W4oltsCi8Buv84/D7Wfn0Yl
3XfnktK5p/971qsXE2eQ9tilozFCSJ3muJCAaEg+euWNKD9XROuqaWmifpHY2ArS
xu0HcHdByv7jMnGUBLW1kZWaY2Q+2JO8jU714H5P5RqgtRFrtt8h3BsT6AybSkzJ
ao2Tzj0aQ5aBuisXQbMcoZFQUjfZwT2Tkf92ssUPQ2jj0cP50h1KpNglEB2iR4/o
fnf9CAXmdEbXwN3BY/ghtgpl0BKnUO+RBhhsq8oaZs/l2nZ+Apzm+O4sHai0reBY
RYbXVQRpefeoW5pLRyoP2RQejroVDAtZEJ7xVP2jiNFOau/qerWA6ViPPruXhQqL
WBZzp17CexLgpkNqkSG4Hw==
`protect END_PROTECTED
