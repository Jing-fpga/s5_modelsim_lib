`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
18ry+f9Aik1jNkNkWKN1fQRYAzqlFUmXzWYDumGTAfuicf1icrlvsfbNAnAxouoT
m9Z0XDk8GKBVzdlQQMyJ5G6Da5cTZtPZ87bFIlSsg6mlziyan+D30dkZnhh/WWMw
T1x74oCpw4QjXe/JeqbUBML83gz94S4xPFvyxWkQmwaJvotCX0ZH8jFl/H3K9GoD
Awwq5KiEyqYNYBEvGQLFBx2KNQzL2KK+QK+AC8r922Asepk21kQ+rWH3Fwid7xP3
HDNgYZKY8+Cm6811siEu/SFuYonhWHWW4vUwun7+87LBgmiG7jb3F7W39hhnLYsn
EyWHEuGBpfcZsIgik8BmRE4DnMhUXk+EDpl57CZKVDFar767Lkts1Kt4wjNzIS+u
etaHU1fLr/BpONc2rCsSFtTHO3F/+558MTHvJj/cHPdRP/innq0QOnOmy80Z4Dbc
Q8MasHGJDZTRtU/dTTF1HGswKUwNTIKoYf7TLhUwyatFRn4kDAp0soua/ZubbBTC
KaB2ozawPTorfpSrT8ZavgVl3qb01MjW0aDyVDs5iY+KegP7ilXFczYOX6lhbXIM
xMXCgD9rZTSr6OD9ZnUVbxwISYJU8xAuKGuRCMNmK5mrjkq+jiZc5qqZCeCF5Etb
tV5K0cNApv8YDa18Xoz/0HoTovDoxnL0d3oLXaDLm/8Te77C7CQikiDA2GQNMxzs
mGAVOtMzQW6fFLFnyYqGkWUdLE2651XwqYpvP13Eqt7qKFuC7b5jwhGJOt8KkXaH
WtTbRZ09mOQDgUcZ7bhXsuwt6TE8mq/NXligB0YgPTUtCQqP5vYWKliBlQzDtJ2h
MKad/4t7LE0qqs+GkwEM+po+MlpgxNPFmk4C9QN9xRW2XAUaYGRF65Xjo4Br8kF4
dohIcZLGt2A0GZEnpSyQLSklJBGIg/6+u12wkMujj2PBe/1X0VSlkCE+6bDxVSIZ
xlm+G69O8nvtyNXviAOd9G6jggmvwO4BoriRS3fUyUACRDs0mMt0QEVXJ4ttRKEY
q2gRaJC+nr3mFyMI3WKy7dG0kQ5mfhPu8soSLmc78uNrBsBq36MBRLCZZzfQU+bL
9o3jOh8fXjnJGazVtVLBtPlYELZCY38WXvAGOtp0Cw9DmavJDehkYQeOJ2m9OZfB
7LresfpCStrere/bsDzvp1rg4l36hp+nrFUGGP46qbo=
`protect END_PROTECTED
