`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S4mhQem7YkLZ1Cyzb/iTyfYpxA3Y3J23K0E34PG5pEfq/1kBq8DzTPFVIgNNlAIF
waaGzEipKek6KOmPtE5RgixfmjNUpq22YjhwHkAGEG1c0cqjna1KspCe8wbqrgsG
tcILHCHg0HsaauVoeLtBMIlLuCijcurW9skwdFPb48miIgVA6HVXxAYZeQQkq+j0
hOdBrSjIWZDftWg91GDQJDEKtv+lyBrOEmLuR1DVd5qWuR/Oi7o+U7Igoloclp55
GRUtIYjaKz1lvH6cT5JXBozt/uZML20Nhm21F3RHucRQDQKPRIaRrXo9breSJGjR
tTe6GF5Q4agNeYLQWbjmWv+NSUYUiTxuMGBI6YWyvz1w/ivErMjW3nbMe5DzXN5L
PXJIRSp7x11lshDnnvPhh7xjZ44RrhjBhxMKlrDquJkeAtz17kPViTeVITvh45VM
V7AXUu7Jjr+QOC1yyp1ZuRQG/mF8driUzpCCNGhGDseX9gmlaWtu038QypuVXGRh
SrZEGNmeJrRJqjpABKqw54ZXrK4RraE7bKxks4sPs3rP9WUd1/v5OEaF+v9ymrvR
QU0whI10PjS8hDczbQ8VfFe3T94yjHjG7tRGlnjT7Y0awyl/RbLlcw0NdLHAgOam
0RLXB8JB7wpsIMpyxbL7xcOWcouK+pCX0TG4DmQskj95Ajm9m5AP5STf9j1/dTlD
Wfven6O4CwfBf3xoBlv3BCN63a2KClwNDUc2mMwtiKznzM8OQXRvXSIzRC3yEVyr
Ttv77ZyLmmtcJfEfmNzPpFg90YXrwiO6PVBk3LrnK1ylnAl4w+oCsSFAsNW53L6k
jSY/wcEx/yQtWcApkIrSp9WCyFyi1h0aSf1ANznegPNbpw1V6bOXmX3uVxlgDwH0
UksV1nHzw4FN5E5U0vmQ61JHkssODMtAhqekMa7vUe9zYYb9TWGTOAz9RwH/alpF
7MM5zxjAmeCcN1Mckpp5vInxsuKdg91glsVwJ12vbHZyqPauRaq/wPyoyY/qY3tE
Y+Oh/+5tS6b2s9Euo8Di4pjYkaqaKprh7m5RLsOs3+6Z7BVxSP8qETYATQDyRUKA
1/rfh9jIJ/OhzDXHFjoA0rpRnLRDFSeAQOoh6HaIR15G/mN0l1Ioboo1LPN0gZ17
Y+lFHUp2eP2xpKEAxJGGYb8L3GFs1ll2ZvPfuXka0RRjUsFQmLmRdqg3fGJm40xL
H3dLeouTsEU9ru0NU2nHrlRSwCcy0pOFMBxKNKNzsD6e+Lyf8AFDYxZK4fOwPlGr
XGGjAFNmejwM72Bj+TPz+m4/2DdPBYikR4lwZO/BgwNNeUND05Xzy1+UG+dnsp3o
5W6LalNEPqt/lxnRThTo1mjlMfbl2DXzMp+6nWUP5DUoz9sLKFz0E8YXnQVh8pSJ
LcrrQ5sIhwW2iAgE2paF98Jfiam+KovJdedHJ6F5vJYGBUtgjTU5AURbhsyCMfz1
zJ0gkxyFgk9VfrFMW+5ZhtiyM7+4CF5fulTPO1nPrFPsPWu4U5Q6k5/uXsM23DV/
89J60vpWDeBf0HeRmD4JrsaMY4JtHRz49G3cCDp3K6xJF6euj/lR6z/LamPpGBLE
gxmsey7mnjb05aDeC+Fxm1mInLpkV6WkHUOHSpNMSsOKq5z4pNu8zNwXxw8FSmD0
+ei90YDGUJbJnUwhmqd11tQFSsYCanaMXCJArR83e3Int/PTqYvbTYNxfleGTx++
/k4i7jPISANo2U+qKMpomlO830coUmt7L3WbkH8POy7lxUaTT8c5VNsyFxMsPY4F
z54pDogjPcoEH6tfIYjIzAG1gRaGuzisdwn/1tpHrTM4U5TEu/pTaHJBn8tLAgDA
C0+ubujX4AKTt5T89AbPVFLXYXvoW+iMuepFlVlBstWWYfbNKfJ5zLexDhX2lPLz
O2SY5Pa1omcR+6CHG69qMzOAXHG02urhBROJe10P8gXbA3PXUZd5U+yjCdA+jJZ+
/XjnXCy6/A92jaSMoOA/9bcPhsV+ioyJK+/lHpuwyLImyeWGsK61opo14DTKl/Wd
SBQT89YsH3SQesAvXht4RGbJaiZXQYncHHRMrFhAbU7qPBkEXZjMTQ07hEpUKKSJ
LOeOVSOj0kJHaLXWtFuAt5loV8cOLfchqIOGTGyZWPSRrO6aJUHQp2o8NutTSLDr
tdWoZH6zhEEIcuMNSoDHyydEYikXhImmdMaCfFZEnIg9ZhWmSq9iFfOCsclMohtF
jGqKLXInBJlRnF0MB4RrQys9wu+s9UoG5pRdhIyvVsYmi0/bjfkta4GW9k30O08H
1/Q8KvU4G0M1HzKUsPASnRidqUhMAYzHNWOG0KMM2J2w5IK3RU/nJvjxdkGBVuZ5
g/oMutJWr1Zx9BbfSveeckVtlOWaS21Je8EvSuzLtNH6BZ6TwqmLlk2/TThycAma
vG99HHdw+YdzO9kqqPs2SYZju1U050i3axd8xYAXjndLLSxlvPGM9GwgWWQ7j90C
Cz3f6BFY2NKIoO2peqH+HmsFM8l1z89rxmo8jHXtpmvnAy5U76sv2Rk9xvVzJCEN
bzfPYpWSAOKP7FqMVlsO5i0fL4LS+a+blg9qFdZtSiylJWo/USmUsoeSBI+iGp7b
InEU+4+7TYIdXY9vKrLGy8f/H7ZbY9b1oBGILPsESTZFipObO2MnUi7VA2X6yVDA
SfRPfDRrL+1y3+kTBHfgI32LfnX9sKY/O7+sdzYtfIyl2yT+2Vi1k644zV4LDRu3
VzjrfIatsmZUTu9lAltwjZGCOEKhgxTDuNtok1nkFPYfbr5PvyEw4S0Lutyax002
B0LX2fHDsigvLaa0ckngHjd+d2fBCW9wFgu4YcDkDSjdZTPkv6p4PZOPR82f0QBu
r32c355uIdpni6wfFEzpaj4ijGS/ydUSEDFixuL8Q72d8hyhp3VJHMNbOGlXpi3C
PDWEplUM6FoN1Cbi5jEDT8YVZO8IYHI8ZsEj/frgpD+utPjTXsjWZAKqPrbLjSLv
9SPl16bRI+jRy5PGknqyxwC/IUdisvJvo4jOcAN8FCm+USPc4hj1prN0Nplyelb0
ZNop40Q0B3DzR7ppr+JznC5QvCrQ9p6anfLgzvM/vvvp34qbAJVnG83PgeoM90K6
ivi3R7NZLSYwnFPTNUQD1/OZ9Jngd4Pw1Mc+04xQSGJT2pNr8JBTiEuNB8XqVY+g
1leW5hYsWqfM+iQJlUy4TMBKB1yXNlMH9sbX5jFYPuYSQhGeHAhADn2Z64FRx0fz
KDLLMPHhTRScAaqGqowrtwU79N1Yq46s0VbtR6VVfpXhQToJ2xrYDmrxZ42fUWmN
nc/ORMCdCAzfQTW2MALGNZjyPRguAWLwZK8Airi3zfAetU4p0ynXhjaMiWyHG3pr
fA6usNQWZF2kcSnso6j4ZSAqRLP9zcFNZvVMivYE67KQuNbSe2s6LHoYrTvYKGSn
h/CSumyDkS8ox53C2uE0e94EU14iFAvB8JZ6qNRA9+j6Sj3UAMC0zMugCBIDFEm7
HNWQIUunCiIq02la5I57F475L/5rtkxfIhFCTLixslR47oCH266fVSD91jDcSoP1
HAxCI/Cq5RSuvlKHmAJ8BPbMwGjzg9ngMwaCnbzfv+FB9eFJXZe/towImY+vEDll
FSBUmwvikaIV35jIUeIR8uCv9uZE6Igbia9KGvRZMqi8JVJGRCdeyzAT46DDuNXe
TWOKxeL1woMcfpIVQMFbURTbqQuN4XJvktjIDC1lgrUKBEqyoJD11fh+0z/hlOvV
SnJtCrvB7kvWPKEqaWxTKJdNcozldWOHzzMCkCoe2TlWOGcb0pBYyTjm8QMejnS8
WJk2gb47M4sJzJ9UHB//FGArqmuB1VqbvaL3OLyVI6vt7Kx5s3LAo+Q5VhGR81nF
G4Npv9Lv9PLKl2/EJ44KUIPxHxS1KWq+yEzgSUJR+COSYS2XMXvzWWAluHISvism
lqv9lcLUnyMExQC+x55WG4dqlgdyk0jbTIVntnRG4B0p7lwY0yKxs51c89eFRZx1
r5PbM7G/aHtMGlahbNUMQZf748iWFXFxGunaCq4SmUBIHhSJapI4dVnDG2or9Wdg
Seq3ZIDszQ/YRn0wbC66/H5128Be+eFL8jehKSB+bqyIkrDFx1pwUIWhGjJu048K
wIIP98+1/jABXznb7sqcaN+kcvsj1ISNd9UZ/el0mPpwwd1y6Jsy9oJq6Ep3xMKv
1llXq7GM1NoKzPPqldpq4BudXj7Pfa2LX459da0Hc3GbdxA31eD6AGT+6I3oor2b
hXghBrGxFeF0dONNeWrskqCm4r7yxFxj7pxp0AR0C0USheCgxFjPrKA+xjTHz8vT
5flVsjLh0Va7WzQfXtZRWe5bdhbNHOqNJzQ/NzlEiBCQTRFBBaonK9c3vBZxzBbS
lL6QA3EEg/2e0B/924Clc/w+cWqwVHT44WA9iVUQ5hYtLcFhUGGjdjSjILqT6lcW
GD7f7ByigzAPZJVw49nBCtvoIPFw3hDooCBzOOm32meVggkdJAgIfuy1z2ZdqQ5o
wf2nCNCp4R/K6OEmf2DHJMPiFOGuzHfU4LJ1If4BOoiqsAEnahZn3bYeIstM4GLU
8z0yTGyIFXvqvLKBI2Eav7rRvLafJu4MIjyGwlB5ejhFaLjaqD084BbvytVJZH31
sK4lZCIkbEqa65Jjh66y5JPWctF6fFiGSCqiG0KEaotDmPnTf2AlU6R44HaU9bNG
oxQ3UGZebYbCxbuGEydO3+KabrLAMLJdIK/WPi7G9GclhfeP5OGTHjgLMDOHIX2n
mYLP2h4M1AlIa9QJ6QqHuigGOCsMIRga9/GehmfqPYmxqIflK3YGWf2Y+S5OiNeg
IpJ99NUacfua4EIIgjfJVXNa2kdQ4/bzHgabi9+GNqPKvtccNQdbb8Oj6C91t0Aw
rYvLw6k+CF5TDMa6krEBbU2i9taMdihSQV1KqTYMvcQ=
`protect END_PROTECTED
