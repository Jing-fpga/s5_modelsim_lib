`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NQPZq6jcTP8ULSAQpzzFDaTWxrs7uTvG1l3HP8/1jjBKFEBdvKuN+uMr39xcGDsu
dsHQfiQBSTPnt5WolVaSSpPRdslzU11n3SqL1CcQ/I9ZFLi51xL5AIGGEk25sRj7
UnM8GoVxg7mOjhJrxqiNUGcxRBQvfd1i9N/WrIIBTkeMz2krwY0zKgYufu3Avtd6
VxmYgrYlEL77WTVRVGEZT3rByxn0emMN3BG+shptw8WFed+C/H5lDcQLTL0ydEQB
+Unq3Y96lbMB44NZQvkbnQi5/4idEoHHrvXDBERnpWk0I9rqGYE60nLgCB2jUD2r
t68mdkj3y5pSvb8Bxap5l14Rl+xBQ1GIFGWOiT86AIlmHmln6mXy7bMmGiQwrkf8
/9jebDXK0R3xyBtKzZ0xWT++hZVkZtObd3uIbaufO3VsTW6n4z/VCO/HctFqkfNa
BK4C8sLXx8bVZUdU6thNIi0QskFJO0EWLgziReAIBU4wfZm6ovhAm5fwvM8NrIJ0
Henu5Vg1VV36ODfa89EFKa61YRd3fuouinBm817AzGhI6cmYa8+uDTYtxJXu/5bZ
ZweSUYQts2FLFOeYwWd6g093M9bXvKPOXjs0HmQEn19H6BBcVVQcahwfuBivVJP5
tqU4TyPSu31GQTMdtKxVceMqhRnATFKwNAyoHrFkkxP3E1locUjyANSqiyWjMEQL
dwO8lnet6EJEae2Q6BWdGDZdyAxT0eqWd6oWLn8aQxMLgh1zddLYNgZXaaW7rUTe
K1dPRkeLlh6ZMfuPytsAFnyAbMmC7XchTP6jcJXwrrhYiOfbCxqlVNdpY2nOSka4
E36DEOXnalXsD/JWCQ3HYbsJjp2kbvOxNHKc7LZHmDdojInw/Kl9AiAa+neX3wzB
rLvD1uCgT4oOGSQ7B29qqs7l9rynDzCpOT5L3M8cAK8KK5rIp3ltixLBvtl4e6pu
QHyiEzqHE36jw18LM8M1HXRHar9Jm39hJLLHvenOkQNZMNCJ6eWFD4veP43dEMLm
dPPgmXv5dvPj1u8iH87BpFTG/kDMHgs98KzN/t5BLaOmEvzUcZ+/UIaffEQDkpRq
mi6qsJ3LzChYhQ/Demv751ydavmjp65gxk77hc3BUo1lJWW5zTrSix6yycKKVLUR
D6CqqJZw+tLzQ85xXHn/M4lcgRRihGapBDWW0q/xa+gKk2gYDPOi1q7j+wPk9URJ
qf/Yr3x79QfmBugDKQFU5eYYjlBDnI1VFGYJHU3fPSHoeDsOOgDMr+KLT7241DJd
EM2BI/jaW/XrYLRK02YpKqLBMyyijjY5D/NBQ1m+KlqSjB8F+AIhm8EJ6MWG05OI
RbLadd9gMwYxsfdLyGi5AJ56N+W0QeuOoVODHkSuQ7HKBshAOBU9Plbl30J84NHc
Q9FuB0liMOKSt/d6XXWZvhcD9rNhB6hyA9vkG+Z/G74rI3wflmDZ1cocJHwojd0j
KHY+Rt6eqsbcnugUF/uOSln3Pl5/GgLJiYlEZibG92C+8VNhmb1jyYz1UqDI6rcw
PJgbujOOOgLoFhpBQimm5btwb/DUoCVL+1WbGPbyZhfDa0cZ6L+EQAOKEh5h9GG5
zmNjM8vZkFpLJsI04GIVdzsIHZ9+NS3Gs6GuFqEv6Ur0vnFb7pqcsY5UYpK0U/ZG
wQh4k2532ctgy+T7CfzzqcG8u49El5BlGTxwFwooI9fBnQr24z5T2EmeyUdM9LKI
+o/Svm0mWERuw8zaGt3bQrshY1OI3wg3DaTK0Vnwj3NLOyHjUCP9CtRYnMDHq0wL
gxXRGEOB1jZ1G1MpgzrsT/Ycw5u+s7hyEGJ74OJUib+YXI6fihM+uaYfHNabWYQ9
Es7zANYaD8/PXkp3iIZrcydtb9b4wkaJKVZuJEGZrt2w7MSal7AU+TR36A/aKdCK
W80/G+bK/jPyMUV91mk5QivwQaQcI4obKd4USEcTv3ckKgejhkrcIWuCjiFenoLB
rA86wPZj15QGD4es1qpORulHTy32GqVvtIWTrD5RVhbPtybVB51avXAGy6bZwmSb
OsYMW12SqKwj0+UrK+xeGCWs3DXt8tH1T1t+l3LyVVw3guSbVJpGJfOC+MP+0JAi
8VlCv2YbLP2jnJLmCkeo5Mo4pDKquhh8MqP0/obA90CDevM/HrQISaAK5dd/Z3T6
SdtO8q8ZxHnTB8ndJxcVzfhD0BJb+zldrJkxsi+IZV+2DQuOFAX8MgfacJcOrG+l
v2cxjJMytc7B7GLtba+Cbq2MgFvWoxeHMdbLE3P7qGi+xy68d9FUzOvehpcnfMW4
TFA5qRsno8kfzM3KCLIkqCtptPp8g/0EWnYYtP/+X1gM0yIS/UYu29ET6xO1Ycuk
Q02Ae8e8B/GAStc1a53u7kJAh+XbFPSw8KvXuvx8ZZ6OyaFx0S/GqUjPiVOtV0JK
Vli2HYobxzS7fHG4Rvh6b9VaacWsVT5KTGMplRoT0l6EVyM+75W5v62Xm97uxNdv
3WDms6TWm7SuJ6W1eSuWr82/ECnrFFmExhx7aygeEzQSy8kjko64nSPnHCJIOwRZ
Kuo0rG2zGH+j0qwpyp3+TcHebOVtHjwXmF5qBZUaa41A98ABXCtD5VjUzPxCBBpE
OmBEZiocaymJAS2HpV3CFUndaCu7oG0rN70hTdvb0OU=
`protect END_PROTECTED
