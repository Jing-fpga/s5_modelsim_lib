`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lCLJwc4p3AkXhIjJ21I9umjO0EbxwzPH48me32CyeJMKCZqPDZxJmBME83Ej5tfD
Y1FLWlr7Ol6dQLIwJOtateWqVHYmmXbE4cSRJxCTQ8NFeDyrf8up15sWz463OyOB
WTNtwqdDMQn/frr8ysFUbDsJcwg8b6MGjNAhEk2EsZMUGa0pYIbP73Ct9QHa6oMv
fl4gb0vvt4Wc33f515TapQ0RPQtvQyTDirX/86DnixvQ+U759r0ClAIT+9Zj4yDG
brS8KIgbG/Kdhx8qdzdcn1bCU/D7aCAaFIdVAj+RiHYITQrnzBU4iT/L7HZ5o8rO
YG7K5m3gBBzb+Z+CPNplIG8NL6Ri4SEPHUY0Mf/J9k1nn8h+e3HNZZFuQ+PXlR2G
OO5a/oFYKkeHQHcNqt0R/40wWwIS3ufScjV2nLW+mtsLsTd9KFtMTMuZfcXehC4k
HqWJkt8iIfMcLHD8AmzsUPO3DE35dmmzWsogOfUXMtynrHBYWGlFy1+/JShI4bWd
nuZ82h2qXA4oTIRHVfmEXQjwyFDUfAA/83TkaeNbo3m0MVENU7yEzlKQ876ydreU
htbKSHWRv2hLouIk2RuHLKnjutTHTCiQgfUyiWq/a69K7GhdAJ3t6KEt3xj0HmrW
EAjIzeuiMNe/j9ggGva5HIR/rW0BpPbVL7pPcNiJ82LjiWo8AKa77chNvMuGDoIR
gsa6Q5KWgrW5VJspw0PYJuJxgBsA4T0X9NmEOBYyoulFBbZh4xlf4vQsPpi14r+q
CGwIrKs8I4wBhnJng5GYRoYhjuZtYZQvEFNuO4n/kiY/82YL4KHVluinIqUsodAy
VENeYiJYkE+Y8Q1kYMS0Gz0lu9fOapvcVByEtxGmd3DDgsnHLaSRTL4Tt3zumOKs
PJwf5Rb/TNZUd0eF4P/TBFWK6/hL/TKbhhX8yu2oIlx2YD60JchIABFj7+UFrkwZ
UNWAXhTuKxZ1ZS/au3i0hNChTab5Rp0ZlhwNvAs07h4pblcOpeLrwLYr3XPMDurw
mFUGnKlWBVcl8+/HLVZZWbUjuNHR/UZlsAfb6ooAFYST08jU8wSC8lCrVTfecpD6
8l96naJWZZFQisuT/vqhfduzjeKPEJ95fSH7btadgGCcMTDfgKKhlJmAJoaoVK50
UeVquXsQGQ/po7O06Hz4V/pj1HyAFWcO4EWgQk7PS/xtGXmxPNbUcflgSQ7S3lDo
cWxA7bBtosE2Y5W5Hm9Fjvb9N28oMLCLSi09I7X6oEVJZfqzQJFeZNGbwnumBhyy
yvJINKgqoIb4KSNcMHlFx7EYN+mmYDRw2mLwDZ0azRfhisDJQgUnAR7FkPwT88hk
PlslBUbTNCOzhr5YaLUnOpwk67Sd2vewv2f6pxyI4iFA0iRbtKXbFQMuz9LuyFdz
K8qpGxSnz2D14mXv1dpOh3KUfuzstz+rpqzLXkDzDMkegH02wJoe5h9HfHiH1Z8y
kHjIYGfSrcoBK5qwzrF9QjFuoihwOz4GSUK99B3outvprzgxjYQDpwHQeH2XIy+9
Kq06baEkJU/RXqrkUwoeC86fw9ddDGykElcxLH/Wf55lVVQvc3vT7phbB43ZzJcS
vMmfmFUxC+gxwvWMPLtN7wtT9GVCUvaZrBKt53yyUJnhfriFhJoLya9hFivBArYq
AfJDs7todnBrfeBKhO3hOPCnqIc1Y1JgFRIFUaMNDptxJ6QbwxtJWvyPEKTl/+9o
8xhe1hqtuLHuUFDEkZ3sL7NyeGl3GOwZsVPlTDL+UtrfwwCI7inQsas7xYz9cn8I
iLeq/ZSMkRjljOlUnMwRLLkGLnMcySEV8Ou5K96NWurvbpMHFgN1Tjak6fVBZT96
QxCXC1Gk8glOoseUBie+5cQAb2f9lB+Qq/qg0zN+POtzE2j9crkj5XR2KJ9Fsum1
ARUt6NpShAD53RMK7Sict6Taigj/eHnfwXejRWbSqYOog4jwo604LLGSV4T+f/lG
oRgTAukQn/IsxG/IV1Ja2wetmY9BrMNo6Sd2wVW8FveL3b2J+Oz5BrVoypBqPIu2
EGBqIq5Qdfm6jy1YH0/6mT7Ma+nGbRzzagTsWmh4Gsk7oMvtgK+HzJwpC7Z65UFZ
Y/NgyLYL/+/0MGwcr3Y/NAzF4aFMaG0X139r9PvcBlbaRk0NIdpU1pdS8PaxjS0J
R9Y58M8eZToqrGj+tMJZwFL7cY2U+JpyTFUapapF02gVL5p/KaaX9+CXGxEfPUV2
mjMR5sjw5hYjER+uElxQ66QwRdmJaE2T2P5Cgr8z6nrG0uVolXYuv4jzDf5nBw60
aucegsdlw8whtKoQM5h6lYFP7H3LRRLe+TRf67K4eCi5s7y4acAwrq/MbTtZLCvX
/2aAyWV0kS9BP95fn6jNhtGcO2O3LLT/X+hCX+R1vpJTPnskzP//Kze6naDBRmym
pMV0fUrBdBiVQWqIXUEFMad9C4R71cExdawYlyS5cUCWrXmeTi3P53oLt2EseFND
64RcUAwF/wNmG9ime9KSCnrqwefCbx23mh2r8Z29aNiVm4Nl60o1aikSptwhYmDr
Z59FiAlnmrvhUQRLthfUWUKNI2UXq9c+i8t5pImPfjyI4oB796/cDHVSkCpIlVrV
qgEYTIUamyOyCjudstSi2RfeE2Vfl1qI9u62Kcn3UCyMPt5+4EPeX+Z8my8dpl6u
QQV7TWohGpNz7TEld1811MqUrGi9gl/o6UODJFKIa2ish9lWXpHV9uy4Z8+wqKln
aTi8RxthU5/yCfP4BcqQxr4a3A+pxw3LMuiq6Cc43Wt6Dt+YpXAJDz/72qJ4HKRV
+5q2maVnBWqYrPgDKKGzooxATBn4kJTtACi1luQrAS6DUU6VjQzXKqk2zuaPiH0s
xdPSIXs/3S3mHolT5OtPZZKJ0Fob6lT+JZTfL9zrAzYs+O2DixIzpIYAbF2V0sh9
rS+jHVVYfoAW2q4a9iFyHFc82hVhdyRTiN+2AneCRrcly41azkH3FLJvPbDFb20U
rqBE02VwNtLZsw+pdg1XbTg70XHuZe4IsaD4twTg4vnmQnnx9RxswEa6tjt7PiXo
K/abBkpEmmgzO04U8AWCAIFO5poNmBtdkuW749bby8l8Ha8eV0SWqqSi8zXV5h93
vvFgVx8RitjgcFFoIkovqs+tvekXAd+pCrb5nbNrodTzmZWdsMFzadV55nNDuX+n
f4UnbGdrxpnbyB16sMs856O1dIvkM484RUZ2QLRcm4bIRwbkI1/HaKM73M3fiQdE
trko4gYRTc7wPoVkgPjspI/vuY3k0OD3J+bBlCaJPp3xSb3ZYW/5fZH4Z1HFh/o1
tV+aC35DNb6uTbqEvt9Rz7SY8Z4WnRniu9BOgHnxh9GSCQwFGjTcvwt76WsxXYg0
fcNDXjfTp9uwEc0SmmJYcWI8+6wihjq7YOmWAtGYvdPr9/NPQHh4F76K6TIIBI4d
Y6e8hDAfYT5M13SVGUQVAEx++VtU9wJlu5t67yHneGMKNXDHBj9UpczlCR9CiqLk
ObPeu+wFM0eguuAofomTCNzyf9ZFpA/fC0DJId1UjXVr5Jf+S1H+4FOALZimJD54
glP8cl3SMaW3T64rTHCbCbNG9kceuE6cYLkroinKblIDgDFsvrpjbnlqhPqyhAyw
TL1w5ejKxbi2N4YBneC9XU8HBkohaoZBCaMH3BUIJPpyfylGIlGusNv/SDOQHhTk
lM/Pu5XrprcI9Iy/DMZ6qhI7wrXYUoARh8VQRXv8hBF4pMsQrJbNLcUNjwUCdm1f
T+FEseFh19InJWkAZYE7hyyUzro+RW530TW5n4yat3DjlBwtGzYbBgmk7nUqfmSG
ewILufcq0C133NBi3SB2oHGYlGTGukbjjGrd/kVpjz26LoWE4+UDT6qFdbX/K9F1
POfiZtVhYpCaYGm+izuX9Pzc0HY4RGSjdcsbkhdFxQ4=
`protect END_PROTECTED
