`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UGLkq1xa7x9jiO1UIsLAr/qjAFpnMlSr6hGBLxdJTdIWi8RmqtIOO+f3Fuuvj6dm
Ijj4ViI80DtqmYZkgXQgncvqMaY6t73+sa0Ric1mkm/Yvvwgwo8NtRTOgSq7ejwL
NOImeWeq1x1XPcxv9KJKGFff9SweTsANDa/VrNO9M8Pp9sNj2bBpmjo74APrhlFa
TqRLcOin65xJ35/tdl3MCyx6CtCaESODd1XCDY5We4kk6svpkX/hbGhQnEGWuMLV
w8yqouDPmn9BHcbnWjEn0gHRJEflypJEf32avWFBCldYZgq7VNRZkiUJmL0+WOsl
+iM8q9wpJmdKZVHesoa66NwW0raLbWoE63FQiGw5xmSiwtDxn749Ihgch+SXJMbz
V4OgkyTAWLp0cEOqRsyHQ93dDIsNtUkMacYR7zX/N2GtCUL3327R28zoGYxcJa6S
hSwSeu2omc/ruJMR6DpqU/P3jafjvwCS5maaeF3J/5pQSXQHAvD5+hVBKGm/NEHz
CTszofFBEHqwe23UEg+IniatXkkLVM3QKu0NXoG6EY0=
`protect END_PROTECTED
