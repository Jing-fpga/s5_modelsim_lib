`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cETxgs30tPx0ZpVQTYASNXv20NvUpUhRKFCGbrH0TnvpoQ0yjY2kdqsoJlbP707e
3KI2Vgqtbn0NM6L+r6/4pjCKaWw1yLBxB18FakErLx7jmto2/TzNVpUWCUVJyeIL
83R69IuZTTIE4wpczZXPSYWkXoQp5ETxiCeO9XxgfYELwCrinoO2bNWXiaqFzP6y
nhJmOwOWFEFBnH8C0iR+3eOEuD8VjWVyMRoGV/XjSGxiejKOgS7FYstYtD57mtC1
mB1rnDy+s0UQok9sJNXuPO0XSUhtDVU0CiukwK0fn2Jg/15DQ+kQt6OuMsKijy5P
Zelc0XkbAI/+VSJT3gcko88t/vPkM1kyEj/JPOmduMjI1avvYl5QQOwfRnlEWoEl
OmVQURYmWnJlfoj98jBJuLLUVQ86d/jx1hYKabxOyOt+s8oKgoi4PzVXApSWIp2T
1lYriMpZ1l4bwRJkCUnxwQAMMK6EoaQgTZfSYKrPHw8=
`protect END_PROTECTED
