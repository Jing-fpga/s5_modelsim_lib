`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5eOGT9IaZyO078C08wgUhMcdbPocTA+HK0davu5tYvvGYMEdO7qtFhV24pRlx53u
eBTRn2do/+mYzhTJ6xVlrLn24E7IUiKUVBa0x7nAOAvBXalq1R9DvB6jxq8Vl/QT
Iap1Q2BmBS1SDCWEzheAH1wCjn8aopFzk0G75xFuCc3dDaBNPgr/lsY2hj6sUqmu
A/UpLtRgNs7vZGov8K7/h+PYPioNCloiMXNdYjNBMJ9cW3skKE913yEn/OsaYQLP
BAiAXPP9mErK0twKUklAse30EV9tY5tMY0IJ9ReLMf0ep1wA1PSFbQbtvdAxk9V9
fBN+YvlCgKy6S31QtjSCknU1N2yrhQvWrSmwlo+eUPQR7eMwXWEnS5o1JGa/2F2t
AC8pPbkXT0QLmLOTQlPpgLMOOZpBkKFP6MhHsY9Gmrgd5yftx6i/wBFV9WxYf8xS
0SNiqonHH8AA3VA7YGQHbh2NATHDVWfmF78vA8XqlSKHtO+OnaJYZE8on/f9/rbj
VjCbz/v6MWpFVxs3FnQTg2iqxcBlQG9GR5FL35H5qY3XeuxPJFO6pKjE6rha5yJ5
RG2Mikl6nZRFvM5/zGAi/tIL72PGTYF30+hqXIAoItClaBUWm2jQoklEle4zOBfQ
dvXL0FHwJxJBzGE9oNmhVlyH/RP8tmXIHWpThHurXHCVJi8MrW9Pfvof2LR3AzTV
QuKPc+8/2Qmm0UB241RIgckNOEgj429SakaQ0LWaJ6nnI9CkDA44HYc0cFzrBb/3
7Mn29oXOk8QH9koJISTmZ9GVfYNyFfuAHn/wCRu10dUX5TNWFhW/V3oSSYiwtCog
ziqDodkPQwuH5VyHyU0RcPfPmRrnNfP4XdKec66WT4E3gtHkhso6pfJL7z47GZLk
NzcRhBjwjjspKkKFGPcjPvca3sVV0M73slyh1NGdQCxMEYblqzyDZW/l/UfZhQzk
OhYrmNbR7vI1z29gonT8Q5+o3finAYnADTJyOV8QWbqXtMBwWURaHlXhbal19Gh4
bFurodzxBF8DqoP8Di3fX3g8CNwoyI6StaERTV1n+trXgsjmz1CJ9ELycZz79Uao
sZKikl0Lptva0El7FkNjT8PrbBTzB8+5cgohrOuhmAA=
`protect END_PROTECTED
