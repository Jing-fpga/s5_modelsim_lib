`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZlZPzxpLCXcq6JnrRAzKqAWA5U5S8ktnGpSPiL6OLSnwRoUQVC8EM08B/bnYtoux
iDZ5vLJN+Q/9Ny8EA6fQyUx663a5sV2ciC67aUgd3B/Dju6m2Kf4RupdrSEqg2zN
9RpBfS5xmLN87PY4jo9eMB2BHrUEkTa5CqyteL20Enj+8wtDswLH5RX9YP50I4bv
hngq9SIrzttREHCuDuHjbs4/tk4rFU8K1vt9hB3HBkHbDo5oLqlgi6YVXA2C3mG6
Su9lRJZ/+uMQ4SmrXCvc1+VGl7/go2NiyJMWMjQb7GxaBXYI7juPFLIIfvVU5GLF
opeqiozT8dHooKJc0t2XxpTmVjpR/MTkUKNQ2eNWWvtKHGGIGAxpvMNJLKPw3Ftr
6cuywMxRc+j8Q1J8DyrSzRTDNthgmo4R1lCupmXF8T4raowEc9/q1IQmHJZfjFYb
6gk6rrnJFqwhSDkXaOqgnf9E6MYAxxPibIQGevfjBNoJn6kWCsWd5RO7QrpsnUsi
0FIHf8dgYUF64kNCfjRvfDTApDLZMsyYfCt/zwpUoTY=
`protect END_PROTECTED
