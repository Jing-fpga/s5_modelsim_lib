`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0kNblJ/ZMRvB8Dz6cQjQhPA9plOEXWQOAxfvghx2e4Qprwb7phxIlS3+kPaEg0J+
PLGhImYMV3FAAeaJ+vyWOs3MdhrgUSX3JAy+mrgtIRzIUZyoCeXmoI3tBzQDmDv/
Nh4LLB2haRC4bE5nQoSNdE8yWG0z/ySUT2RO9eqtYj/fHj20EqaH8aBG2Gx59uRn
RNWJWVEdrSzhmxK6EIRn0A/wyr0dx1i5B4cnUsZRebByQKfY7eNztQDXXn5pwPiG
ts3SE8IqRwsX2tlXhs7wIlLIhYTs4xZi0ly1kMrhXdbhByuLQ3jtF2A53M+KJizI
befGRtdBdegDXXyDa2fu0FvJlFIANiVfIX0AfeD35s07Td86snZqJLWgih8sJ5Do
X08HM5rCJcju3tqvIlskTxCwwbOOqN5aeLUR4Mnoctjq0Xqq51Z5b5VIbKn7pH6k
rxi4jFbzSE7OWKN17p5T6TYrR5D6eCWB7bw9o0/P49S9ZcAp4uLYpCNKRLfDbEyw
ybi5WJBqESlLsAB2S8fcH7yBSKvgy9Fr4G8MoiPdeGaS/h1SGbkkuxzAosiKcSOf
aOnV5y73DTzAcaYpCpKHGl/WblMus1fk1ucRLd6pQ4sS5m9pYaNufG6z/mYRMfxD
QzoMtFkTISjLHjDIqXTwtw==
`protect END_PROTECTED
