`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
na7xQhC8pqEffK3PdEcYH2+R30RcPc34GnqP3Xir1p2S6dAofPsqkOrj1DbJEzO5
0LKNybw/L9YCW70eBdlx0qQmI8pRWHMcXWB7owtGklnLkPgD/2DMOW8td7TMhQgy
O3SNQv9jjsu0E1bKz5Yh2qSK+oHLTyndFvDI1uZThqApgyI3RPu5Sp1GbRSwSx0T
3PCwUO1WCbl1JwfSlntuep96vgP8uqY9rhDA6wSs+XL0gcHr5+yKaX+6So2ipHoW
oYTpNJa6lLKwl9JayGtJahKZ/RlilCEegGhLfZT6g5tKwiB4lXqywftgeHz7+tvb
JEGppZ/VN6b5q0fQHqnmGmEta2fd2xRU/fVpNtYo8OnQkT9bAP6EV2Hx/Tl4jUPY
KqcvMm3cWh5D5cNgTYr+D+QhPdjfJjZV2fYXS4ezOs7ZoJj4DRUMedU2dzsMNU9N
BYpxfyvNGHTZ2pmxX1PuJlbyFeP36byWS9LKWrciwd4K4Uc8smQhvJhd19UPgcpH
lAf2Ie7+ubj30tClU2Do2GlaoXSdR+OZ4cxLTp73ibQ=
`protect END_PROTECTED
