`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Im3xvhztYU9ORe9A9rsqXDzX6SHkoRs8jSYNTmQ/I3g9TE/a7/inn700wQ6uCEJ6
6sHT+5Ocx4k1JT8CQ9GpShXGlRSs7A2NGd5i8YXoT/VDT991vjo8BxHdxoCjofkz
NCaE+SL9GE6CDQ+4FkqIURCZWDOSlg/Y6IzsB38YFyPJO+8vCbYXJrGLjNtPbSvV
mXX1icgfOuxtyPyjNoZ9xzo64YNOPkE/l+Bv0qpkjd+YI6iTbRbDmXPpIX18UKUx
KtEIZhy7CA1OcG8PeEiF8NlFduGYuITK9uD7jyVwTVYYD5wNXwdnQ9ZhQusA3VNI
9y5CSMgO5INC9wPkGmMCpEgQWFgukfu+8eSnrQz1JK2tZVww8Gc5wE4VdPeKY5aH
4BccnD1OlX/PB4FT3oKaHSdEj+LRjB3gEnYuCsKP6gmhLbyOXuVA1zN/Lv9KlwO+
pPRjHFswSGsrpWg6doYtRk+ZmtoSfrrHGUlYYGr0c+yFiALLc9lAj5/ZZM5r+OAU
uRYT7Lgyf6x9Fap5DidcCoA9G2cZY6hrvG95tmGHM9aQH8y3wQoT0jhNo2vdeQ+B
6OBQSU/WiJhhMP+v/3Nz6KmaLKmz5z+C4C2O5hF6YoNYmYks1ya/Srk5R2BQ331t
wD7zUZ6dHkP0D12jntblm+h168mEgYwyKyb+P56M1AtX5tTZ76oLgZYh7Ln++r8e
L9Rxo/WVHSi7MesJ1XpLqw==
`protect END_PROTECTED
