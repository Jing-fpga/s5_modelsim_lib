`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uYoT0f5rcIbNhuWbWnx3Vb9yOeDvwKiNFHOTclxLh53B+SSHdbBXPiuy+D6ubfDY
hgrUPHRomRvZMmOk3q9o5rqq1dkZNNFvLKm8IXLZytbCRxVbZv/UN2Rjpx2ex4qh
LTRhIv8clsZ0SHiBW2TjOZBqZL71Gd7NfOxp//8+D3QKb3T9b+H7aqUsHK52Sahi
fIXj00no/33hcLgvjW5nflP/VrBAAaxxnJA2KnpjK67xjAxbEud8wF2mLjtX6gFU
e+Gr79dBDLrRiIaVaqXiVt/Ldh5/JctUDfzaX8ubLq1HyJCpi8I81VzRdOYD6C/f
I9w9MiTweD4yqbpC35MRzm7UmTZxGEi85N3nc/dTR84h0uLa5x4ikF+FVcCIQeyN
hfmoqizCp06FAPCTjkNqHY80D7WVL5O3F2xuHGYx3xRGvE+Jx9QHDrrUW4+xcttE
2fkEdUaYwoIaR9y2sgyQc99AK3UfyV3Yw7IuP/beJEMUqk8mAQYPj18IhFotKGXj
c/mKMoct0l9COMSAa7qPE+EiPmQr9dT22Fd/fLURR9gZLdylFc4LNHIUf5Mtp7N9
7YtA0QkXZpHmREz4zF+bi53PF1qdD/m02KL0nytha1INRayOS8Yr/L6HyE/EVT1q
Ou4WsgiUxSLSOK1EnRDc/Z+fM+0/v8tuA7vfrG4egSbjBce6ZLfgZvvTg6WZ/E83
6a/PPZ2do2m194TT8MjnDs8rItT7odcsArXF3oqaiopt2R+FQQvSYFLZTkGrEhVR
+Bg2DOlDVh3cNbx5LXVqMuhWd6uuooYKBj5L4uBFCWnztRpIho0N61cB0eg3UoL4
m5k63VqGNXtkosgGDJhmhQ7vlPLRassjxC+aPHuQI7YJ0JB86Q37XuC2yf14Rr4N
nQoQVlXGS3L+0zJv1d1VMTJ1PJDvYZ5nGSb3SB5RBA1cyFjADxab7OJuUxPr8P2/
8Sjlu8W0mSAdQF8s/GfiiV0kROfTXsVOrNTY+ymldJPB1DkDskYC/QR2qEbDSoVC
18bTm2sjDT84nPMBuCKVcfsCiPOtz5VtLQOmG0yibXSBSonXf0+HNimTogRuV1T0
SkOvLX267yOHXxT9T2Vd3os8lsOpXAADXvhiaz7v2UZXnrN8DL9dgGo1wr1pip6W
PkH8sWGZv7ICDPDoiKNcW+IuJCRBCxMVcETofazQdGQnXbWoNnXuUm3LYHqQqcKK
fqq92kqHgTTHJH+VXTiPsFzGFcYXDGe+4xCcz2IMs9zZq0kmYQe0HwAqQRyIGaFJ
nudzMR8Sqne7Ao3atpYd65cK0tzT7kIFN4JaG1YHBFglxFsqTTWv67rnS9TDeBZC
qRzSmR1mFK6dsR8he9E/NMXNL21JhBhnqtMS10GGpm6OfQYrPkH+P1QukU3exeEA
ZHaSR0vUpnFwkIcQzVo6cLr9dIGfX/VZ0QXOsqWXmXOa0KB58TaqtQLjTfVAOVGZ
36tlenaYaiH2TNDRu8VTveOqs0ycyMpKF3AaWUPVB4tlSqdw3wJXHFAsS4aSwYb8
pwht21Mr2Ox8QOz9dFSS5Fwoxzfvax/0Ku7eSCBKvShL9w6DCAbZJYu24nKK+/5N
9X5ell8TVngbawVuTsBx6/mOl0qXj1eym3sbsuhQHu0TGgHMnlpNGhA2/qRi4e/4
JdG2GnyIgJ7gEmY5pTmfTMKbj++AQIU13HPy5L/lBIQ5hitJyUTB7RCakMvnxDwi
JcUqeEPYR+XL1BgdU/VodS6WVHVhs3JL6eTAOQmrlncAr8q89Fb72KG3DIet66ms
QKv+8mXR7wStMdnf9QtvJ4iRsZv446EBlviXFNWeYVP4rMZiSNa5wHa4sQLVT2Ki
fGPgGQswqYUVMcJoCluIDJVMgOr+9uCZlDGTKv7USrbLq4nhIn1S265hpuU8T051
KwB35pA6J76SF5YuSaqI3hLIBpM0Ir5gZ/BenmNx6K5zk8ohz5xwcMoxg3XCVeVZ
5SeHwcC8Dt1Pzu65ySaruK3rtO3wOghUB3inxO4Auv6XrLrYwWsHIa4jSUeEsE9M
TrhoZUZez4cIxwqtFKz/vMxapCczOVJK2cTvNOtP2tmNrb8xgjCncPrsUj6gEQkO
kbYPs8Q68QSuRfJusDmE52NX+U6swfh8umOzvAcYEGY=
`protect END_PROTECTED
