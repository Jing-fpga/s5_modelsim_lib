`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fUwkh0jCqijOujxre9Rh8bcLgMpSdopGfFN95lbpUfp2Ewo8h4OGGk6etybm/utd
Bx8f0+sUHaUHy4aNshgIuWHOZiJTMw246PaS1nZXEizUiFH6R8ff5NlRGfZI+WhZ
zF+bDKIgcW6032qweiofJmwQHt5B2FKanhXnRt/UOR3lnd+I5eT/2XwpqY4DpOOr
a/kbbsZhQoAmiQHSS1jE2j5VZ7UxqY/rzLpT8pDjATzvv8iaX92el3VigWcHtasZ
47K5SPsMDrUCnIw521MkitLj9FQq3FyXykeVmdblQ9w5QadW1V42C6HIA1weidpr
dCZhtDiETWsxq57+n7l1rgbTIXQxn39NKfkX0VR5nYoKJBOWWjvENx2LWe9KA7vL
yCTFTfn2lafiXiU9leygsIrEMJp9KVu+tMfE8f81O5CjhhGDZgNEdxmCHQ6Eri/M
8unwmCPT4+kqF4KO1PtsD9kC5pXP77pRSOHo1xKXTSEgo1prw/2a3CPv4+T3uOM1
imfIN/twTGJrlTaKwlDcY+1103g+9UBUi9xRhHIvTn68NMpbZj/C+gUyI0GtZhKC
LHo4xd7hxbVt35gwuu3puREhNpyIt0o6GQ0mqCxMDlw=
`protect END_PROTECTED
