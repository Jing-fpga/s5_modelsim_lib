`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aOhBmx3kXf6n8T3krXun2S/IRydkkvAuFaa6sKxP2QpzITI5REHIO81yfpauSEr5
7lwuI0XSR99tHkZJzcvkSppcGuAe30youARNlcEMcemj96wRCklAbqEa2YaSb80q
7BDSCe0dokh2K141pL2WlZXG0KPqgX+TxhR9fbmsA6d8cxgoL4uzXR3C6HAD5L+c
mSStKaA8jyavWBJxdakBN+vCrRqqKLuqTNzIIcM2RUVxAVnRVgrBzjA75hwnhDvP
0/uOynvWYEVFsYBCVPBO+ATu2DCRpxsISrACOdCkqoW8bsB8yEMMdCTCYfYVY28k
I32TC8rGLJ26mfe13jVcT6VIqerXBxt0H91MrehLBC2j2NeXWrlCSNui/utELWJf
OBTnSKThrL5nF4p0ANivCn/FNeMW/MDamTNqLpZWweD+dH2s8TAed1zERROLbpmO
ktEj4g4hKGYaj+/8R///MGSq2xJuWmJ3OnhU3eyHwvtHKraAydJ2lz7sNpBxtMY2
gG6mDmPeHbtXf8Q+/wwmI4iYKp6idb1hoAfnTaTiSmLMJHzw3OqjS5Hp3JbMoKmz
v/6TaYPVVQWSthSAkx1l4Zhr3LfIV1B3olOlPSnKYzpwX4wOIz2hKp+eSyBHLys0
bp1edSaAFKlkLJYumW02Uqe2PsolM8keizudEpc0a4uFuSoyfuYRh0/mOsBv52VD
T5vZftl2tF0qt3/01MjhS8wj/pJf/5AjsQsAk+2mlZfl9Plhkk3Fv2z6UepsjF5X
lodtq0OnP6m29Cq3UjwZxCenyKb/pegqjiyVPks3uuCPqiErd9e5iEUW7aL2fxAM
twmcayBiDt8c+ItOBowU1+ZnOSD8oBrnEV35QeZNn4+1jOHH/fZ0qG6eS6cDIlXs
Z3qRrBTCLjxJU4MfMhEllnE3q45+JWPb8s9MqhJvHxxq3g1vwXD4w4QTdqZ+HnCU
+j+TSEEhGodBGdwOcPYH6PbOi5HBb+A9tynNYHczzsDphDN/RU2+DEBNsfVUrDiP
jmW858fIxsvlXHl5HXbeAmyJ9VX301VmavP2gv+HRnRGPl05psI+YOih3u/vQIUA
N8tudCQxxUkUnWFsT/vDOud9QYSw87LNH40xdPoaeUUGQqyL/k0tU6WGCa4xk9X8
/xcKHqlMQNUXKw5MoqX9/IxHJAU3Ud2g8XDCTcMTBoNLg+V3NUY+1DK2RTM+IcYR
siJ3K61REubYC1IkiaAHJITJmRBSpWjziWgoH4buqauIgJsPjupstMvKnofse5P7
JGMYIDHBacPP4V1YshxEOsnjANfz8HPXcul1sEYSzK27hF3KNCEIfNjNmp+PZFtG
Kwm0aZP0axKZSlS4spQwVsTsMCprnYBGru3EdKmOYQ0B6v9ei04YhnMfI7ZaPOjY
zB1ofCctVNUogRGXXs4cjWWBhsBcc2vulqZH3iLVCRvT0anzOxK1WpYGLXU6lrqL
31l2F6AEF2Sxw2/oyMAiLLGaQvEQie9p3BQ87scvPpD4KmOfblcwcxVcmiUrIdME
DvHF7A0zlZCJquh+T5sCAtE6HUImr0xvyLROxJn/bt2EdjTeWyOolu5YxLJ9WCJU
hJWEumDlpDweSF+wVYnb/C6Y+BnzUoTlDlSF5/2r+vv9FezHhO4h0IKdXr8GKGTl
ljZYzYmgt7z4lxpHawJE5MoMTFyGcLOxkkvP7Oz/vmH1lSNApPyl06FqFgMGDzLX
MtZVUSoopAAA3MKm4TvKm+b77TS4PtLMsZcuj9/9/LohHU0DY1vJlY64tzcJJlJP
2l+DDnbnUaupYA1arx8mIB4OBqTUW/1jDeaAFfJALS52HdKUIPAMLwvDrrXTemXu
un78WkYuHxsrn1EAVKU/gFSUxk5QA1ewJLfH8OCUENBZFiSi7Idy6tJY74V/lxru
3kzcrq1X0kU3nLlNvgLbdc4P7NP/oPlUGSQwHAddP854+art7kkmiGVP3x3pfT7d
7dm08RxgAnLmAJsb9WZBfK00gUxVpjr28LiWL+obrorYwDDdkhiGXJU8lWAOlnmL
XdNqU3Sf+Je85ibZceUE7lRDE3E/Re1rGAf5NeIKukDFgXyYthnSd1ZnC+rxJIft
cKPcvf2b9DrZmSZHTgH/4InU6B+YCKo8938G98vlycTf5gmJ8Xc3yh3G6rHzhAAg
i0Tnx+eOecPD2+3DEFDp7++Ut+h2Ac2prccxEFv/XxDjzVf2t5YznGnJaoWMklB7
NPOYo9u3DeyxnduQFIFN8z+g173yCYLs12pK2DHN+UKiVQpze/Oo24eqKBobJqng
WmCEsOR86K0r4sIqXLeJTtGjlQhvR0x2/7y4lC96A1B9HjFPfFSSEwoR9YlrqHmU
OIetY652UyAl3ln69tOihXEyPSivEyikAbQFeGS4miF0m9Ktiw/YdUcVy2vs1cHJ
j8r6YCxGecOo+528aqtiQUClmD77rvmPcxN+fTUhHqk7xoXsIKDj2qWUG+QFa/mk
C+kGz0l3Cb3MPcvMZO6y1TXlCjfrRM1wEvYtjSmisDEBbPqY2alKYpUFTU3jerBl
tBf9W6uYv+7tykoaXLbHJz7s4w6ZhpQRsFG3aNUt3Pq24vi4ZB3vwdBhY5yohCL+
XFBCw9eelZ+U2HLwUOPw7t9AtNs1LZbxmN10YMxIMgpoyzRuYfaA3al9O5m2CGUk
2ak41B9Xleef5Lz4w19RrcTAAIx3O/EUwYEZl/lp26IJ4DVFr3oqyO9ohGtBhNOX
UQ7WCY0MWliwJV/KwzPOrkX10T4XLLv6EbBn8duy3TpDqmoL4/8U6axwhPcBdZcC
pNvuXuH+YhcJAVaH8jIpNH/HbIZW29uZ8Kqc6ZFXJHQK/D8zADT9bTGm64ca46m0
GzDMYG8vty4qXvDRwx43Oy910IGvujvStTYu7lsduQkWhwn07kajccwg34lSDb7p
hTRVMS07gdWz0DzVwjnkR2yE9xKtL+PdyUIgmFvIDXraldt5qur1K2J8U1ortm70
KtCDa24QiqiPbDBqM1f8FZY/zWD/nrDIShJcGoKgm14rQv35awX5UxbNt/9f15gV
0APykgsJm8Qbf6LwRCYuatpICni1KzFTeAjUdWuYBKgQd36GVR8IPYAUF5Nw3jBG
BmCXbB3ZlQIoFuisJdya5NcfXUjLiL/D2rYVH+DL+oYqwuXNskBI9pWuGeQmYLeJ
JsG9zwi66QAy7jNxEPX/z/3c003iIqK9VLTQ8h8UbeQj34rg0JrGPXrotEOgdx8T
7aI2lfrFb4+S+EveKDOqS0Ip44hL+BypaiGPO31u+prjKbo5xOjMaYwaTiSWWEo9
dw+lAy1EKxjV9lVEiyuxxsBFubPzvPGWGo/oZDNW2+nayB+ZErU0FuFL7CIEObhx
vLeuuVQcX4KIdx6RlT4PPc3NZEc9pZNSlE5waCZ7+mnlf2o1XQVVawLSsjPVeoZJ
8S6ADMNEDrR+drACcBNLqsVowRmVDJHdXw5ylKbxIvw=
`protect END_PROTECTED
