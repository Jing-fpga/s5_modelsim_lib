`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qfkm2g/bLmJsImxvmQBcrJY+dmM6YaZsUq8bFqw/rHhkWCd7Hz+r/rMt5745brhG
zGPsmXlExmTqqU7VhD5EOJW99FFoKdNobEoeilfnX2fq2ft2XVL1rqjwrE1H2IiB
Ep9djnZkun6xOI4ZKXl0xYENBuloLJl2zb3+40XKN+tRKyhUwebAwwGi9WYYqk1r
oYXI+fGmjWipY/lrDkUkLniCrHsNHzZb3rt11/qwSOMLdsxMls2wvwmd0WjEplGg
Fir4evqiQhGPkexHx0+K08xeVteajREHIS/zEgDSGCxuco71vSbao0O5WhBYcfRu
xav3CdOAW8rksR1xb3JRgiHl8fFxRybJ6kz5R/mGjZzrQ/O5Exxh8QvNZpgVKYSI
TE+05nFGqZ6b+2YuVhHtfqIBHYwzmWfr4JF/me0X9D5knAE4M5D7yqDReSam9T1T
tYmQTyOKGvbuaPqnDXl5+Exnre0sovBN53OyIiGT5IP7I5BhfoDwxXvC3auJjki4
RaM8VMGiwY6hGHv3+s36WNmMP4BiI7yqzMc2/4kd2gWTMJTcd9xuxgRpCbdkcaXX
9u97gmoQMrKRmPIh4DwzvO3WZIT1sz8RdvZ/qhSnBmdAid7F9iFQ+QJVXuJEY7lb
TaWQB0u/5qpAEOYEuMZ421u9G7eorZkhQfab5y7RaF+oIhWU4yRBtWTHHXXFg/HP
WXgtZSQ6GH+dC3EhP1D0wkVUpst8IbeZhVYcOdF3P+SLeMJMx2UC/rHFFNex2mhq
Sc4n0LClEI/8z/yTk4a+PHEep1D+Y0YrFhTmxj8hHz5RonT+055AfUkCEd8JB1i4
6/wzfVU6hqtV1OlY2EzTkqU+wdrsxhbO8HPT+N+a/wI7Q8jnP4ijSjPqfixQU7FW
mZEXJjJmZczVYTvtzr4i1RtXGlUb4xVmtwXhLJPJPJjB8Mvn48jPSV0Bdr0WT1jb
uFv36+evKmgRQNipxVMbdnJ2tzhts3nY0sxSWIuFbb/4bHtRNIdqsunT/cu2bSgZ
dw/RykbH2yVFe2ecy3Hk+ayqQFXpTyw8eRtKydPKZQawpacqR7CE4Au+56F3RDZP
JszI73frz+hBJbT8qN0+hDFFLn6eUU+hdzeoFRzG0wTrpt/Hx+UO2H0FFwemlfZA
qo4MeQtyLH/NUyY73NLIdbudSN1s2oxqZ/eYGzXuhF+DKgaWn+EtopgIVrH6p17d
Kdnak/M8G7C+mAxz1EyAveT4KbeOKJ5kkmawYY0hJm9kkcjMx9B9kWCGabZDYH+R
zNVoUFB4j82FYEC2O3ARaYz9zHqpHB7J8XjlUAcGjmARyms1tFQGuS9mT/u9i4+r
0CjJsnEHOTmW66Zj3768pTabwsLAoGH5PWdarOosCbJdmZkjY7UE2LsLt4TVdYia
0Ilt0WtxVnLAGjVoGokhCBrWT429N+lXN2UW3wtDyVbvyBEsq2cQIH2LYUvrwX0F
XKfXTOv0POxaYyMTiB1Z5FUH+eGhb1Bqg8S9kbJDZmOwj6/XTnnULUVLKIoGppQS
IK1oYq3rGzGCP5nUltlz/ziGRwok9qMzg2tCfxfVJI4FUgdxotMXp5/M9LzITZLZ
K1BzLYaWG0xLVRGNLfAqB7P7bxpmp9W4GaL150m907uiYRshanMF0fGmsz3PZT9N
DE3BEy1dlxrPfuDStiZGOJxyTYQOL5BEYK4+syl5TqDgkvMjNKDLsiD4SkO0oQ2l
kNMvfZ+ZCzG0B4oREmgl0Q/dqEQYYj85QIe+6PJl3Dlp3UGpXWCb1H6/T91WynBy
RIqtHjRL+vwYpaDxyrx06uWwqs6r1r3GsRnbJBNyaQuivxTjnYeAv+HF+ruFHwHw
uzX4XohYBP0kdCEklSxxRBfacsYu20jMdJVBGvVG8lilJsC1WwHKsSufdBx704KR
H9nIwqsmk7LLq8WGK3iKsER+BFrA+MGwp24YBmP2DBj7mEo43W3KDrKmMgmDI/JH
spEOhRUaOWkBXFe7o+bsOf3XrFIBEIBjsZHjVYd90+jxbWhnvrCmKe8hbxBbfnWg
+yX1A12CmOg7AH6HsCajhNIriRz+nuocGAOAe1ZZLHt44ZxhmVw+LQEYw7pjAMid
RldkDB3e9zvccegGsfGEU/N3o4wqWlRkHIe4vyU27uk3bWB5IM4hJCYHraOsvLaD
+IFy4DRlcecABJdOKEqy8wKgHJnw0yIqoMo8v4XCmvHQRuygmkvGyoeksyMi8cgQ
L3kESiNILJpI4wPFulhlvOCIbRuvsE5eibgsFglIu6bcm5Xwd4uqBxjKm+FyrjT3
MEeLLs7dJvybFFtD887Gl/hZaHx9v3QjR/AW5KfsvOgUmStz3LmrPoqjm17I1q/c
qMRBdaa7qe79Q1d5GwqA4Fm3fLHU5M6e1r/5vb5w9fCYAh+SKYKEHEgYGietJIkW
iCq+RyswCKRJw8re4dvzRWgvlmp/cOEYwmU1LBBY7xlI/h3hSTZZDehqPLg/vKYm
UJOsp0BW8O8x2tXdWvU7JhA15H6mfEPh/hHeZHcckj/XhbUSp6aX0cZOJj1J4PBt
YN6vr9AkUTk5efUdXFz9wHmbn82K+IBlwRVVrUxpS38S8/OOHSkQqwaMnA4d8eUJ
VHGXqTO9HPQWlE+jJhMlw3ZSyCgn4eZeeq7xP0kZlEaplzNw0lM6Ke0FGRPFoBB/
/K0Kj0bSGScLvNGQFjOyS0aGl26Nrf/AsKE4VtDtMWVfP12VG+lrMRpw6W6r76/d
y2PR9zQOWWxdhptwe7Fw6KljLQ5ou/ddCUdvfxc1AI8Gfs2oSOJ2U371Hz8QmWDl
kSmR/owbA7SMGrZg6Q9nJDKFzTUbMT+iuG9y5J9yZCDVwIYOdVbPXe4lyzvPDEcD
4MzlzBrZEZeWyJpif6m8t5XzWTSmXYQhyUoEHhJknviY9NE56cISHBDEXJyijduC
W2/GjKGizeCxhgqZsbojzVtd9XBsTxPMvHmd79+JVYbENRmG+rKmNV3QtBvZ1kqD
mgMQ/Oja5EYLRh57kHmEOtl3guiCaxNzQfSdy4Hg16fzKvpyqermve82xoscham/
4PGH3QyPzsrumUQie8EBvAe6yoo+cfTV+WDXAS142r1usWDR0c9lv0iJnLxZl0uD
xGoVkSOu2a/KjbV4gtkCJ6VkNbpSBbLlfT4C4HO0BaHlNlaVhsILThx9g2ayMSsZ
qXip2YnIkAffzx4v+dBjHN9kBwj2SGc1bc2ulx075c0s9/KGeUc4pmro7/ogREuC
le4JsFEWNkHIcsFSYg2OF+8/CuVmCKT2nLywptp1rKVR0SSulZe/HYShA5rO2wtt
sNVMsaJqzfWeexAe8gDx9ZR41ZxZjpwe/tifwpOAX8uR5LTW0ZKOLVrCkqYeL796
Ch0y1JLmHgQsRnorsLbThPMYudHcxSY6z9fcg25DndxVyL4AEH1V/lyhTyq9ARAf
eFjBtxZvhwzSOv2bGg0SWRfcfOnhyPBX87ukXX+XO5GJhrd44e3OmF94m8OtUyEd
CznB69xR50Fpb/fX8vKhNl7P4I/p1XfjZBz4OdqZhJkYnl+epv4ciio8BW6DF1aF
u1+Q6kF2Toi06fGaqW037GUnd/m247mKoHJ2Ye3xSvfdAVQQ9scqwMgyNUx5vHHH
PeYep/PYQY91GRms0PzQWG/c8YSkSAMtmfg2kleCrS1ehfw7TpZBR2FpBHnTgZVB
Qf1L1QSogMPine++hFZA5jPrd/8slGcjVj+40FlNMQjvdKaRnBkSwGLP+i447hs2
/iRUPIXMljCBkEs0VImXxZ1Ym90YEvYeBB1bOHYTijCvPJXh0Mu4gLJc7rxd2ZMJ
Lk/pkkvxdFgtu3IY6o5LG33ZId/JZtaEYKsWP4bzWOcnUn7PNOl8q9QRjYflz8tj
9IGLz/56VgCAsfbA8scIFv2Qlpbfz9zkJEr25gRvGb8ibyS8cXiYtmK1RCWMZfUk
WxdC63Ul9Fuxav3pUVOo/c5NhmOd5+G6v2Nd1vfzwwLgdHFoRvap3qzG/5tFIcOO
Bwlps2BUIM444r1jivekDrbQIu4FFXo457A++Xu8vxI4p7X8GygSZgKspt/hfkq5
WqJSqSBR3W7+VhpQWMLAg8puj4m6rCCxDL58YU1z21SPL6vB9iQ3KPFlznc2X4is
d7gHtza5s0IfWnCbxspnE6DShttqgxcvt3aRE+PR2d1qXLkwxKI4SonQUteyC/pZ
qwgLbl3kViVhpjlde0Pz2naMQbPTZOTN4uhvzfkucfKBYdzHvrgKF5Ry9ekYqtvM
9812GpX7vy9+7SsJo650dG/MexeeP9WBeYdhOU41JRmmMXprntqMzXYjJd5yILp7
nBVLxn9h38Kny+2RVwzmrweniowDds4T8ikg+COLDs9ISH/RW7hhI1av3IKphD9e
ywUjb2Rakgp3AXLphPHVFtIRFovCYKb7jFgBmC+0N5upbIB326Q19q2Hc/2ltd00
5MNymOkmldwC2tekaQKJF2Zvkkv0jhU+1PupQ7Trk8psV2Vj5VNXPHok3KkplhCY
RVaGghgh5GytfKIDMw+vzjWFZozC5UtyiKzUTTl8Rr61/rvN5a8fj9BLM1dtTwiv
PslVFaFaOTa6d63uMmqk2E6gFHIuvVzSSPj7le9omJhAIR5H8G67h7iLtD6b5ECb
OMjziD18fqsCFEGAnR06eXjTFW/mhDeee7m78+mqrUUsfWf/Q70mwkigQ7Zn6szK
LG7o5xkapoAXI4L7nfQUMDcp4miY0n6ge3keOm8/MlAUVuLNlgnJurwR9ccgddoD
R3IZCzSX8yg8dacDIRNV4dtF7o8nBifeBV6AWEVImoSo9VKeBT8gjSSnIpgfbCIZ
ZnrnLSDoDkI4+gB3HzwplS0Cu4kDHcb7STl1uvjrf4D9tlImrdCyx0qcIxf3/Oiw
yERUQclfZAqGUfJ3i6hr9W5dmtUN9kTfcxhLc2lLbNWCdypIiACBX1V6ze5kzqOS
LPzzwODpJEIrTgK6qa3XC4h10v433oS02Tk5Ai/9/IrBjcO/DkspcBIKizMV74as
qGJu7S5Q9FIHf/SWxxEtmAizFrBHBbCDx7thZm6tcEbLxUL7O3HavTE0AYEF6nkV
j3yce0cO51CrFIr9bc9x6IGmHHwMSvXgy3VHZaVnVln6cVAr2wNEApZT6h7jmSl8
ylaSV2r6aSk5F2lpvm1F3huOTddHyibJvvUa823qsg20JZQik6hbywe8fNmrLlLO
V4BrduKgFQBypXFFGoOoRFAZeQnYAHiBrTgBEne+dGgslAszB0CT7JEg9sX3ABzX
unosmHIuKKsOhp8wSDbNakUxsWLprbDEMNJ6EO7kA6QPY/eWf4wCFIXitoZGlvum
cr5t9PHseTpG8mDzmTf7DwYjzSMEIz95kd8IjTFJScfKjW4q4ic7xqQiwBveSwrx
NLNWnzLIVldw5k9QTKEYWr8jPhl6jPHioiTrpYEKVxWMUWB53PJvkQx65CngyzOx
3QeeEMqdd6iHTkqNhqBj9GA4zbRTLYP6/zFSnIKNtbJNZ9W3wbPMSJ1xWp6NzDdB
qlMjOh5zitDx/6qu4Hc5CM5jYMBvGv6B5n6Nx9iyrBofWg6vd45vzxXRuaxgiGn0
oU94gxA40CYQUwLF24dhVP6CWNcDBXNNaSCUqw9/gHLJl4AKhMY+EZ/EuOoWfBQk
sTjcTcE2oFnFPU+5RAdOG/OZImpeCoMUPAckKt9IyCKW9tkBu5Bw3anLGWiieXMK
Xjom2dxgUZRTXo0QAVP7BpA2PjLmtCbkcsrpXECBlLKDXRiWAe7pbmryW0jnOg98
GKB7nyHauLlWYBV9ypUXSKd2s7hDdcTzE4XJsRMIv4eUXVNHlfmgUXNPH7q/Dwuk
wq7W9w2eXPx1pXu+LO33uulMwQwmqGHtm4HDo9qbuBvIJbmUw39ytBS2yFmNYgC8
/hoGYZutGwSEN3l+E/yzMbhfqjEriuIgH591i+hk/QsjJhYXP1GekBQZwP38wQYu
aG72P0TP55TBEiQF/cErXqj0n3PtxWMFz8onCeV9xkV0frfNuhmo0oIBmtOkZiE5
Qc2+avA7jaXR4lOeqjOCiTcodp1cqqLB5wrdDlKmyjciEzqy6HqTNjce6mxUZmK4
Lv141Bj5fTbgfWYfdzDRXwJExY2pNqhQiNTpj/P0+ksvYWh+hpikxFEH3ROyaKOQ
HGptjrpn2ms6yBHOIcUnauOAsBOD23YaMpaBl401DJ1LwYpwCGKLxpTySSB8qRUN
NG3xufnBd85HqaYm3yzcItd/yAwMX8YOCGqlWuJw5hw+mtjuxcak/A+BtkAgwASl
/J4rtgVOMEeP56aGgTEcDa3ioclGy66pHy35b1dNROHkCZoz35To4UjCkUSJ9sXC
zgHj2IPI5q40gL7VgmvvFisrROBG/zKfW28BaHGa9+6M9psNTtsDvgSxb0osAKB2
bZTrkcFBPCiyWGkuNquOdRKizSZovlU4whOrIYEhyXY4a80ZFME2SHPhGvmIoatD
9GRPh2vbCchKQmvVO+JEZKzHsq4XpjUBIh+/tRVaTGixwOjtaGoG4Y7fib32KJf9
8cLOhNa6zDcieyQp3Yz7zLjwnx21daR//KMzzlk8RNNmifIDyCy8xni3o5AK1p3J
8LpmyGMZ9woxg9rek1odqHbzxpe4CuR58a1R4FqUz9J5LJ85PdGAUvqD3L24xpEY
bO25mf4vcoiTCDN/EjMT+KtF7X1RPMT/BaNU1Qfk90VtcIl6/FXjdEXtuSic4gs2
AoDBV3Q1Mm7U3XFYlQqIB8idp/MG0tpwQxHh6x0+6poTIy1HgAnN1H01/u3i55yS
ZklfQ396Sf2UGfOf40ZKH86sma4ybMb5DtI9GXaTYw4KEUTNyeJ0W24Js4gzQAoE
WDrUBFSNirf3ZLlHy7Zs8ZE3adC/xy2KjSiiBTCSlTlO+uri5+0ZsE/W4jeqGfQM
LNsADhPMXQEWGb1NOmnIAlm6aZx7L2l6jmHXDFYRDY8VOlcfGVF6jphMe0BioQ6N
Axx/ARKk/btgO74EqFydZdpNtQV72QaHHksiUn/q0/OdvCn/4op5hWIZa81kGj6a
RVgzt3ZZqgLn2vUGTIDAcGpeUt3perlrVuuESzoiZFQcit8UPzbP/wDbIe2k3/Sz
yNMUyru5tNkvrHtrjLM4rph3NhAg4KdXt1m3WPFcHUpIcTequEY3Tgx/KKanJrVa
aSy9NbBU3s0qhKi898b6C9Cf+9KB8XCmsdB5waNwf9oLQsdWxKcH0Y8ysiq2ek4X
Y5GYcYgzDaxv+RYenjs/JZ8KqFjlkclwARC+WtDSr2Hcxgxl5fXgQp0bSg4A4RGY
OqUvDuEboXeciRxXbkax4kJTvHkZSyYyZLtfHtFWd6YwifV4Vc2FTo25+79EjvuT
lNE4Ow1hXRozV4Wx59FwlQ7pLxYi1XhPnbrBV79HTWNVWsafotwGzvLBTT/k2V0n
OqY0Uehj9hDwlFw0m2klQbjKPwHeoP5PDz2NYcyy9/t47yHr/tF14/z2H+Jqzo2p
4O9qOkoY6ux0LtHRrs/3VyDLFKhECDc+h64md29x69YUUPnzOZ5fGH5CmMZ9LLIn
Z3tByolgCxeEQndx7odYRtITh0RQILzXG88htBsR8ruOpL3EAJsGXiMz3GCIxFwQ
+43HZB/cr16Necbahqa4zBOme2yi50zv2SsS/tGobx4XyHecF1iNTP/sKrhbDDHz
H65bdWTpMRxRTFgX6lfjAn8UOdlHMwoKTMgwqVRjI9B/Eh8rzIVD06KoIJEe7zF9
n1PcTqvhs3x0zV/rJVGcarDxOQAaMfq8M3PXvSx8d2+2M2/gC0OPR7eZkIUXhE3R
XrLGCxPtxYIhPdXBNjmGqEj2sL/zwZDjnuwIP9iCXYcLJDZ+u125MTZLIhUieGXt
6Kewh0pF/KO4IH3j5S9c1TT+2ocYt/IuXN+nk3a2hQQFnIG/UmqjgAmWXm1F7ObC
DCqi1gBU04nNLyb2RWI6Q9pDFlmJZ7rBfjVjllPP9kOtsMW8ijcDnWHD3zCFfnGw
gsrFRmOhQaobIijlt5Yp/GS4bQY9c4U97q+QuUbt9wOrPeb2uflKp9RnHcx5QNZ8
ClABXxyKX0OVCrKI3Qd3VM6JbV05pFL4WQTTguXJ1//PwJMhLthATELviSVaHRn1
wEzLin4rESW3kXyRVbkV8LevGI4vMuOi8EmNYdjWpFFgH1tzCfUfj/mY+g0K2daD
gb7teRHZ0cvSdMRmRuwOGplEUZIw5lTalHToU+QWZDz/SZDGINfI1Eztzsq2/XDd
ClyaL5ECHDKUTsp+/ePYBZNe01mN4FQj1dFfFqZSQWBjjGQ3m46jGtgeTuI+0mMM
n2tRVu22bi6kyE82AjN4lF4djt/fgw5nCcqavbd6tkht99kno6IVXSpRjUCkd4FV
31DHYEgsqI1s6N75/Ueg0AONKFn8CVl+5ZVpm13DkBEQkoypAng6K1k5FEcfhM6D
maI3hZ9KO7VLODWXgbbPJFh/nZPko8q7nKOpidpVgsU6pMcrhf8Bzdgk3PCsuZ+s
wKJFByRj65sjgK3t92NkYdLiSCH/xksq2hGOusmaEaQGafLFekxi8cyXBc3rGzsr
RnREGQJlTMeYtOxzzgspwViB8QYrLgSBfvT6yyUaZ3ot/FIRsYXRJIEIOAPLCE3R
4KtPk7st42YIDUEBT/XTSC5JvX97cHrlCpHrPSUajOTXOz3sQSPQFHoRHtCIEq9p
Z3BSfNeOznf52wIdcAN5ghxc6tgmYsc/FH/gc/0ihHBsHpkW7nZP4PMFq/sslKgx
dLU2IL2Es5pNhmtL1Ksmnur/fZf/fy4IJxW7U8nauZUEplyciOqqeIuKyhykXA/3
o6SraVpfxXQoJYwb6Aul576vhlMr/IiznY0zaREJ2NC5Bvsvall/tkSu8PDuVTde
pt2MbOqN6zzfC4bWxKVzyz8+Hml3uqGSrgBiE4uW4Y0jdxYquisoy7tk3rhFdZPY
lTa4b5jjaDEgQWyZbeP4vgNevWj4Ci8Sm3mdU+wJoJHdU3N7moDcUgKpZ7tfmd8J
SeyO1M9SfYmjh7A9ubDxWIN4U4D8UFTIE2bNFAVusU8oi8Yog9OPKge62ODCwJwq
ZqBF1dW0bR3f4HPYsOpEA4a5CTejnKNEkkAPv3hErHwwfCX/NAYiDiD2s9I0F3r+
MP4nZpK8iqx0E2JorxlnRLqS1CcYe+v2GcRODKcRGbY2A4W30nq2papE63+Fn5vf
0uW6lRQsZ3qxCdCdRqg7aEajlQJ9og1iSeYmk04JTskqcPmOKzFPN9t7gEOqjcbZ
7NV1zc/pdAwPtlqVS2SbPtZLbhe+Vru+zy7AXfCH6agSrbuyYyCsoVJPL1htSPHN
4tv3lwgT6uE2oyhiilV3I/6iITmKd5iUGc+KdF1gR8Lt7C2gSleyNg2aaMORqdVv
6LaZVXEm2av6iHBsP/hJ72kT2wlvLR/orQSW0FPi9+4hoOmozQIgHmNeCW2ZWqiy
jGLR8IpnzCrHAhM6e3hm7lp3O3oz8863EHt1CmkNpWKEmu6BmE/9SfuczwNqx4T0
Pe5TFjVlWHVlrK/EwGnqOJqDMjPsEZkwUtMNMJq1lETR5EC3gGhmhb3UWnR1ZYYv
1Njd+ivscMlw1QFjoQznUisA5q3y1NFBFWOXfaQhZodSNv4IEQeoRPPm7HGQZVur
ERtdj1RNzCRhUxQgfa+aiO73FyxoDCB2xqAemyWsFPkDnXernOfNSko9+naL0BYH
VsKALwpXoD/LD+g9QFytUpvpha56fmQmlrRG2kj8xTKc9T/8mPQPRYEJR6wWU/db
mn8XlxDF/jW/CA3Ovsdc1TsTIO8vFmXwp5lkJlxjYYRrK3IK2RL0SF8l+71tLa7y
96KysDP2DdBXncnJcO/MOyz2d54nDjQUUQGvjYuS4w0L0mJQZVmZg+Hv4MtD2dzW
Ggbcb4+yvChsWJW6A3ai+LBoQNwBvC/nuiw5tvNNn5wqvi7vQiWWiPnYgHy0FKUm
Urc3qpqLBBx93X/Gqi7a9ZC72NGezV9G2k+JOV6FetS60irR89UStOFzlvcDVMBr
ozLz/9wdoS9b8c+r8rregLMsPDIvFIDeyV36LMtV0hFP4wmLd4B49KpLTrCSRCgH
dAzIYTGcZcoKxax3UL4dW6kGBQtk8drKOKAqrTaNS7knbLlg4CNqLws5TrGj3HOa
1YdJZeWYUWHd8mrL2akbB0p3KkG0fuRB4LG/4M44lSK3qoGk1TMKhf9P2zQQDV2u
UTsInHfdtIv009qHYpLaUp58ohmX+QYxTWLi6w7BojtOJy8SMTD7U/iUmvKcqf7j
Q4QVKfOU1j+GsV1l9D0inMf0Qor17TH2UWDpxsVJ7/04BiE+R6ixulb/iiQKxopq
XpnKczb/jK6elBzulupImvta/vA9XpPc08H8on/y2Ncv6zqEg2qcgz43h4yOj6mn
Fh+zv1Yp/GX+BEWU7T/bJQAXXdlMNTTXaSR+Wfp+EdRmBv+jHyc2iqz4TlGKeLQd
K4Fsmh9eTudFe67HrIiSv8fAwGpX62hHwHgyQtW9UuCqSHMs6Z837XB47ZxLoTjk
AdZJmchDapKtB8RZ7dochjZnUGZO+xP7rJ+oNT7sigAZ0QsLYeR2EsUZ1WBKkKp5
JQvahMfPN+mMcf0rHmVbQNBDw54An+FCufaEBpc5fClCF71jbmeTxfhwwgbUHFRd
8ovhsV1OIHfGM2lek0I3h86SkBvFuAIzMH+4xQURAG5J3OJwSTyH7NpXCu5mrdUa
6FAaawVt3dmmPuKpxr4+xKVCjFnyX25JOp87DUxUNr2SModFqhED6T0bk/A4HJ10
bc9lWBVcncnlQOmMnv9F5zXlUnpWhV/jupHWvYPeuPWsMrx7XUEATabKM4YnWRBW
fGCEts9PDgnSTrcfKNrca3Bx0hREreuHG6VGsWlh/Ue40+8NG9v93U9znqwz1jo3
aaud77IvybGnsjymS1FX21vd4u4fY6UBsL+lVB62mBytX5Xm9NDV+6g1HUN4uOvy
RVGeQx81u6Toe340oC8sI6J6PhJfdwB9kwFCRgs+cHcLcR2r0z0sNDv2rnqEcfOb
yCMwK7BrO0nMYuirMKiPQPH/h6V24Mbd2THaYMX48EDOjUIQ+p6SE07w4oEE682r
B80jFc11cOHx9d8XPouhLUBXMRulg9bM3xoKYgHW8xw=
`protect END_PROTECTED
