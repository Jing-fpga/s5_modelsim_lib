`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uRmWSls2F6OsIxgM7bPaBt3YOMy9lxfOHhHfK04XBuNHUWoDet/msnxG1cggK3tT
iHW9+5/HtiU0//FVJCIK3139sx/LlvusFjqYLfUO2LjVwAgcUDioyWHCMAMy8ZUo
qlCG6vwihG2/SyvmRP0F8tysb3LukvjeOmn21SyFQjGOGIe7yhk0j0nJDr9zHH2Z
SpD/l82yMz0TY6llzFnfJUNChnMMpBN8WL3DeNCVSokpneDLbScxKOeV/diIKw7G
0JT79vO4nToDeLHNpYUJdcdKgloycCcmiU8vA7BvaZmOJCu+uCgZEd2zYCnfMa8b
T/+WBrBU3ZQ2FGgEtSTEkpEe8IgdwAGYV7GFA0FLxyItWTZs0GpPtIm4h9CgPg5n
OlTbE+AQRMwbhTBU9fuClvjmAQZ6phOvTTxcyS64MqJRnjkV5noOXG/VrYdDviom
795jhkJqml1nvRhCruizQ7RKCdb2K33BZnzIQII2R5Vg8vG5zR30s+0fb6arvKmV
Cyh/DdMZ2LRuHoBK6jyGeSYOvzGHe/mZnat+iVFKLz5/lXcAaWu3YcqUD8MKZq2V
1tnlDSSwdkGo8BijkY3RyjL+wbii4PnmmHVjNejLOmHZHhI9xhiaVUkLiecSEsOF
el+VeZLrcLcsD0T/ySETyXqHAJe3F7eeX1sSLPdBmhKdc/FqXDhoucU7mbKSUVfK
TQ5bttT8XzLBPB/WHuAGIg3uI94jOttMBYOgJkNiuQLvkNTdju47lbnMcy6E9J2S
+OHfaQuYuPuH6dlxkLWDOdq6rBENIyhrkkGedszrOSwWO3FlBH6mzToTjO27hpm3
XP5aAzi1Ly7YjqIzZUM9jPLbwnK0VCDXlaMVWgHjY4117Js6Q8H5D2+jh2v3dhep
otZWciO4wIq4RE7Xp2Ih+Urri5QSoEFO2sxm0twWRi/91z7gziB6iA4doiudM0ah
C7FxgWsGb7X3zT9A1FchlA78KUXRmSxOr9oQGHLwbtjIWg6aLJcpqpDqkEcKb0er
MXBhK5By8ejx0XioLxPkscIrEgrQ8sA6YfY6LuuYENCkUbOM3hDh+BqMhkVprswa
10GJXAikJIPOjQFWFa4rdH0rQBLyluha81nb4TTxXH55dUZ1pxC4pQH3NxkKlaCw
szXXZKN2lSIuN4QEFmBgfIiuYYgkohZvNcOqBUmBFUYm+LMQiXms7HwX4fARLSLe
756YaG0M7KSwlEVvNSGQra0/9c8Cb0sbwQAPRHBOjJYI/82xkzh+wGVvsqxwr9lM
NHp3jz1d7uFhHOJfrv/Tq+ocZw2I6igmb8HKPbN6DPWKltKRTHttR9xHYrAvRT4d
Yl+yza0PWTopRsUUzWFCrV3JGNPg0FYBnxGWCrZVg2jv4x0N28qm+tgA3R/KVtVV
5EW8Q/IMNYeKK8eSQ4K5OBIUnjkuvlvXJc5himb7axT3CK/fW6sl0kwlkeKzWI9g
lqn6T7RNrxBw+KFvKutNnlizz8/tf4n0uMhYnFrCgyBbU/ewCOrAA7rNX7lN9g79
RuXHxubrxNpPXUCFaUjfwhHB28RLxUPv20xr+v2Hh/MCubPOJ7tXtf+52w9x7/Ef
dEeYYljDn2+3Ar4ppE5DG6PxAt5DoLEwZWk9gtZiV/LfReKPE79R4tGaXI1GMMxV
zFeztLfdxgCYoHTWyjxrLEzQUUe4yin8EYytRqv7HFysoDycpAGVDNpT7snbtA7A
Ae90+82tz6/3qSMZqSCohYdW63aLVkX2csyw2zOf4Kmmy3aO0SXyYLrMCwicAyhn
xxrn695ARUxJr1L7ArMIsMcarN+TB5n0FEJHpM+TBpRb9Hokb1nrlly2kF+F7zEA
efzA4UwH/BKIE03pQSCMHsO+ConhI0N01PYcdjzEpJ/g2xQ9PXcDyRepeGNUbWR4
t8YjaNIKa5yMPA+97yPytBOsr1ZqqQt8xbGDKKHOm2v3Wm54MVLDgGEuAX4r6H5a
LrW7fjLKwOgXVHDDjH1Su8c+Dvk0tHfHFAvgcpnkFWgMMZ5IKVywt1ohIPzISifi
UxumPKgmv7Z6t0OKEKakEPogpf6POlFjjfXJiN1BFCk4dcIEIUzTHpygjVPdRshr
IsA6YqnvBUzUXlx45cBGJF/UW3fdLl3G+KsZNVtn4d2ZZT08kQfIQvaJH8GgLppw
FX1fhpb28Yl1n5joDY+pZ67lg2+wKjVRIUvJknqDiHqttditsKhRplp1VAToUD3b
8Mq+Oja0dBbB2oFUbqJWwZbZe7L5iu/cloXTlU2uocSkbW5HboknmAO6WCx6xjRU
2j+c19FxhXDqG1sEhGAz9WCdFJyOk/N+gbhdB3yWgAUXAlF2OtP0x4z/H/JQJiMc
u+KBz7gENl0cNJxfs78PTeuirVKJEdg0vl2pp7kDhxdnZ4FyLDZ4EvKXXIONuvfX
S8rtxaBEVjZ5erSbtQ9fKcbNKBUQwNL8GVXH4MpjqIo2lF3/iQFYjiyZt0XWjvC5
9joHRS+4QNRK6S30VpBpoBRF3kyJ4IyulE2w8nd9/IcPksBGGTdXsl/PB6A+KzQx
hiF5Y6gOpHqPKUxEqS9Z+ZnWgMPWWIIdhdblzOxxYQyk34FZTpDHJsoJwLc/hCRz
RdwhOcLfM7/5R7GRtIYmXxxQoKgO4WS9SvaFUVL2cMif3AXmFN5TmLW+g4O8qaFH
Csit2hmtc/5QwzEa+Uxg9205NP2HifLm64RMwNBS3hdAT1WuV6xFR/NyzYxKK0VV
MC8/K6CoWj1txEDkgj0x5lfjOUnV3Mcu8oAaDXnQczT1AfkvQ6HlOdP9osBeVPRI
heJDbqzD2mmceqMcwwWdsTa+MjFqbdjlK7BVlUZLbqPhIyBllgZGGpDCyKI2Gyd2
nIcIBB1Z5Q34UdmuLuWmnoBQe36f1lQY0z7OUBwtzAXsc7Qyez2wkm42x7ZE39ax
Ky2xswtRD1NdtdF77kUYtmfML8bxSJS4X7oKED9uCn+JSWf1A5hKguiU7AXbLhnF
g1Xy/jVCY89P3RgpFRQuxpvhyXO6qfXBWLm5QOfpfpnkCmHe2CvzEb1ziY454nnm
+XVGnrGZALp9pdagFvyoYhxfQJRx192SDTWWxs3ZZOyV84bkwWLLLIOlmte/nNH/
r7TWaXUCvDHLZmF2gPygfo6YaUbwECZDemjIap2o8/yxcI40yZKcQzFnRpKvcbJ+
ihbVKRvkF/vViEHKCBtieKP7+A+FT7sYB11WG3g+W0aKgkTSP9SE3dZEpwjmRsQI
mh8pxRa3eOW8aQtUyEhJtXwPHBGSfjd3IF+mp/BiDCb5EfzYS3UpoS/OY7j5ZQOt
lDotpOh04uyz8PMwI2IBTd02Vf3Bbii8G5UIavYIgeRal35xbLswWGLekghmVjHt
ksx/Bw4EUTRS9DCSj+5wrA==
`protect END_PROTECTED
