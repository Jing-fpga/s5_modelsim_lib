`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TzPYNFJNgubE7rlMS6Z1AaoztC9ETZKKq/PJdk0CDtLpha2vQAvqffVsClkjcNCv
pMCHu15ySoZFhvybn9nwURdNr6pw0MU/Hp3Esz+Z+yBJ76P5CPrS53YBL2bH443c
kmdHlZI8Hic/QlhQRhDlH+NaSSNLoHdL7yk7ZO1F3upWoeQzP6kVNLK8ZtX4+m2/
pQoMTNUmTO92nIY7F7OpyRFLgrWUtQld554+WNl08NF6IU5QMIPXSjiXBz6k2ciD
7jxOXqDYBSGQpeBdbYy3y47jSsLoM9LbFcbmY1ylzGCF+IJlxDAa2KbXI63iCUSP
j7TQmPgWm9PZepcBeHuncVU2bNMUE9iT48iFFp9tsG0Q+Q/yy56HtWeeyffDE1VC
IhMvgrNXPbzJK1kn19rfSG904IJpOs8CsCM7VYlZQpDaIZnGd4L8KdziqccdcUCJ
blHic2ePzC5bJ/gQ/XmciFCjuhkGl4rhstLdxJza6GMXIMzAzDDEutKdeaeIyGMp
V9htgbd5cybrmPc95gk32AbJTqyJfo1Yg47usvkvAw4PZUq443Buv8BvnJioRhIS
Uha4wWNtqvUmjTU5H+JXPIWpt2qBg5LAGV059kCV4P7jvt/Uuial+yVd7RcpXbvR
hnsGSDShKzc7lpxfTCkHIFfk8qDlbjA0ZfuhTugISbIzzmLS8NLzh4MG47TZ2/HM
0TsLa9riGvrtUA9lGi5miMAlwQ81378dGNSMVXgRdcKFFTttxLZYsYbepwdulzCC
gmqsmJLhyYo2shMz/Du378tDALxLnGKEtRq7ud2omIM2DLKZFm0hqj5y5z4kakcM
nP2zdoWIHosMMrSX4A25ghlBEr3KjUoYe7QT/EiT6vG6urUVOIdgmKoL+XPw1gOs
oqyV+hMJmQvzlXSuUxg05rXGUn+7KlwePpVWc6TXpNQVz+J/+NVNDUbirIwcCmo8
Nujo1UhrYHQLhf6+9ZCfGooUq9DKnxgaK6n+Dvvmu102Wj2gdp0aJSm4bCUI8u6E
I4xFqeE9Sa/dJP5s8sqLYx20m8yGxnTN3s1B08l2sZncCYVXClb5VH9EFDGZpEyk
g0OR7S4oZ9bMMFBFCGW6qIWRyDENfjBek9fR019tv6JgiU7Bf9izpVJ7URPBGjfq
eGpSTkVrIL0Y1l8Qp7SyVXf6m0PdJxI/V8Qvouq2r7U32/XF4RPQqywj+KDLt6nd
gVIApNdZZ1RLLhk0ZLiDohO1jMavxnsvAALTrSgn80K06P/h/8x9McgABuXNTBpW
LpMTXeRQBHK65+UamGFBunMMCTYvwIDebOXLfsqoG1e8Hm8Os3K/T1g5cbOhOtNC
p1blqf8kAKHHgLhwWf3Q+Zlf9PG9/sIQL7lnMKjQI4xxg5akoaBycdnBPRNsg8qB
l/mcOvaBC5LGVPwJ9TxmemCxUM6Rcjf5VI4PCWO5R6qewvsrNzbRdWi4F923wU60
pUrLiUQ14vtHu+p0EYco549gMyK6iKMMKOM5THCcQrrvgjc+peMYC/hh7YWC2Rxh
/BeUftwRHCiYEGkndr3RfnSLr5W7mG+d4KSozmG7xArfwtr0tWmfmXyCX6eEzBnz
Mb57gtCwAPUdaD30rnCvqRCn3bKwETEhCy3th+sLcUBTyKm426Yi/s4r0bPakRXE
hc5rmFRjHqOHfj1Ty42qa+dRnWRebmp0zvLM1fmdXntypZPkNWKH3PnpIPo/xKxM
ciMNcX8ZuIEGfqAya1hdBtBvAqFZJmCTciNYSzCbn97Kk0Joe3+z1wdpeZ54zBNx
mMGfGC3RWflDktR9LH+z6cen5WfgFHgXDbwmyo3erYVb2JITbvEJHazBTi1ah2Ai
bWTvpryIsk6NXs771Dsalz/OpsAvXYttKukv8n9eOv5GpyCEcJcyARi1hMq0hvTc
kIRMapDWgRraCf6hSUPxJXBDaaANX6AQzky3age3cnJwMkuqAu0TwOPqwQxBT9Ym
Grqy6CDdLDQmGBUfuTg4RAnZj2b0CvtZk7VUvY3+FcsG1xMAVm3L4wChJpLfNRSk
fJcU3n1smR+MjIkVLGBn40bpJNudWHD0uw0pgugzWIe3jRat3QRWxgUoEm/ZqpEF
4PVdtXzkoqoM7ofsODambPUV3gAqd2txUydoabeKvdm3eL0G5BInhL5/iAdWZN9K
r7MMdnLUMJEWopiIIFMt1mJhuWyA+xz1hPErTVhlM0dDJjuIIDu4eZhvSubCQEmC
6jzJtT61igBdfQxpkyP3YWYYkyjcz2q+kZp/zKhK8pdbxdkQcMiM/kE9cmglwDLl
j4WtOmpxbKcfs44tMGrSeiymg6AYURnNdVANvbbdgzN5d/jbtKdXxCqrOKwAFNnO
f5fDEt2pfkB7L2nm5Qqh2JsrtiTIAuNU6hVCEjW9ccnEda8xU/ZEk4az+9e5GsID
dfBYqH3D9SycjQosJHJE3hyevflNOXT4FsAx41PyI4hTQ+aB2UZrbtTlXDDC8uqw
apEkWXQ7eyWEkdZerIEMlTnjFJuE3b99E3goCgZmWFlO4Rj5qZjwEPiWuJ5egpF8
VPKjBPugKGKsBohNh08r6FArXFPT00KqeWj4/OVPsU3RfBjDNmVVHWjqGpJ6BbD2
PtFf9J0zp+PBGnptLqMI6Lp87DqpxXkcD2pDnjh2gUHjI8vgbqC7bjlO6imXI/Ur
IEsD1zYRxTQyMSAf9Baj66PqKj+KSyNR8T6xGmMPZGHoRWfMXjZeVW56xvA74wj0
1DkKpMHPjCNxORhSQ8qhnq1A6Ug2qpPoGHINV8g14nzUg0jWKq9wwvnXWhvTS0hr
EbGlwYcPCYIy5EiVntysN8TcF83f6mNmi3Qayj+xkcB7PwfDvyE+873X6aYoZ5zI
VV1MN+srS6otMOzMTVcM986GEbvE3nhec49SdFh7x4YSRGsuG+ZKN2yf6O7uPa6a
82B2FTapLnsviKPbgm0eHeIMSPvqnSWLIbXEUj8BXRWZlBWhlr274i7IQN8rVHZM
1QZoR4Sd9qyRO5KqlBR8xrlNkjwzJjjI+SkDY/JX8WMgGqwO86W5AwlkwoeLnI02
g7ed29iS03Crj8CNangPZY7ce3X/FssBpzs5L+f/qWoZiGm4UXh21gncPrcMsxGh
3QXr0G4LkPmgm7GvYKRRT3A/6s0+nPsjqYMjXO+aaWQ0sTzuAg/Z/dm+rRTcuQ9L
9s0thO57mRToELkezEuApeV7T7l90FRd7lLB8ZH76rdTy65034NO4jhmElz/UNvr
DhmfZt/v0BQveCJbqzTiFzDFp2IW+pWrLxp1djkAQMW+RLVaJFI2DFiZP73QXhPO
kfipIv7+xiqZ7Oybf4xSw3p3441o55fk88dvNPLQJeJZ8r2LS148WVJMQTY5/6pX
rMIR3l5BUnLR7A6WjV2lFDiN59JsjjhSORYUzyV0DkdQP4UaIjWTicfHCyj7pXG3
11yRUSXvpvGKsGCUFLS4rw==
`protect END_PROTECTED
