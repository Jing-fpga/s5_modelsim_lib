`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tb6BhLQO/YsRvKBKgCkJ26gds88GQNriXzxpAhlPBTWNUr/4KiC8UvDqzwP4D5AU
iW8WRnmTRZj9T8+rimvh2lhqZoQaQ5EbnF/uwvnUT71Pz+1e1Ow8Oh6VOChkOW/6
f8lhX9gYIijB80Csh5eZ+YXdLqtI2tGGHTGUky9YLxl4ap0z0l1/rpCfK3bOWWP4
biXXRcWtgEvYEMoxMgXszExbCzOedn/FCWyKHXxTcBNo7TGA9dkT5UOUsgHhNyPT
yBUww2/vneUcjd1GrCT+6CG1/HXI0XZBu4WdALUHt+bA8pjSj/8RsQpPkVWcrwVu
SCPLHINtL01mDf1fGQ5zJCz2ckfgrvzNf0N01OrZVPGyza9hcAk/qBht5nm+6U+3
cAb4DiPqpE5Cbm1FxVV+L349mjCpnFZDnGEmchUdTBqbyEoSQoQFPqvu5vLP7tUO
XMdQnQV1MJBTMGLt7zCjrF/0Gp4ld3kjVmnXteq+SKFFdCOjQXMXlh7e+6cH2vyP
8qBgBi6t1gVrTntKmn1TVn0yKVKesu2WKhNRJ9ZjlXPXf99vlKVJtTyi/oZWtqW1
tzUhizdcqHTVc/Fcqm7K6fmyLw7knxVLIZPw0QZzK8nhs/2pWSxEFlOLOnSuElk7
mDA1mr3am3392w7nRjsFAaSa/U9XQc0mkBy40F+iFyJocaWF/NRvgEkfPDhDSTvO
kRx1+iPLrs7Gt0H1kUJNgYgn2NozKnFBsw5QjAjbXAYmJ4DJ2blY5fXBLLgwnrYb
MEkTq51v35nNweddqrKd7ml9gMEAhQ7a8M3qjo5BZia0o4eLtL5nTWn8wrl8D/er
TjlewS2KGzakfwnfOsj5d5TEVxqslF4WpW/dnDZu7AotZT51FStdRyEpmdj5CmSm
tCVZkAkif7kuo1kELasOBcilsvycy5lhLui6Z0SS07HEjxN+cIdIId8VZbJCru70
t19B5Yfhw+i3VKVkLyJ4nwX53bxv/nbiFt/in7zoeFA38MefDGBxNd3xllif/YI7
04yQGWqCtF/ZY6Heel3nWPZabt6CAbuXYU1v7WS+slf0EIhNqdDdiTjbg9x3yiQA
ByPEA5iTZoIycc1oSu0GiuO3GB1TO0d6xWe8qN6Pom9ZiW7w8gXEnaU9UD6d6EMY
tjZTy/34wchoxtyZVPu7iKGQ8YOB0BAexcYRdyuzZfp8JbtA/bI7sxz4NHoCixjs
q6Rcg3d0qsdTa5OUPpgosAT5R5hdjnClE4nLrncse+rMIA6hiQ0/tX1w1Cw8NIlj
FAA6lPe8ZXsDKPOTbIm6iqnUqV7cSp6a6HkhPFKCu+qTltEpMz7kDw8SYG1LwtbF
9/Ogn59NPRXRx6vfyuFAV/Z/MYifxU4tpOJQhkzOMWEVvfO5X+psnl3pxKH//RH4
joPkIA4XXJ2j2ZGsfGfIkFeZ86mORsbrEWzBz+5FywE2Hk8N/wLP/Q/6ID4bfON/
ugKExRlqB7PFzvxBYrm0Pw==
`protect END_PROTECTED
