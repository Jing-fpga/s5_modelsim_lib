`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VTVElqSwBGsGRKXQQjak/JMTSc3hpDSohhnS9NAawNDdSqtXAPygutzYStDD3q6p
pTgRrrg8PnfV+1As9BoKJVuzN+Pd7GXeCuAhxbUF73ltjS5XF1niX22FBI6TXyyw
Da15AT5BRFAOa0Evh+0ml87lDOo0vkLBS5K+r1CgKQUSNh7cHRQE40s1ejULyAPA
wkNyHAkrPbvYA5WoemUeZYK4s+Z0YnHd+NC+CvGCL2j7+aKcZbBkCx+3Eq7ShuaB
mncgxSgPOYBmUPSoPZmJtX4TAyvrRYvgkWf5HF4imrnyjLN+z0seh2FmdmJjBxGT
CINE0Z7TKyVwwhrRTRh09XzcRxrnqc6iwoMrESTN1ZNnvKDrMJbpp+N9GrQxL1hn
DinLkM2VXHcm7R9pkKQAllQTcbRmNnwH4UeTRmCsixlkYs4YbN6XC4qkJOc5tAK7
KWAzo87Nx2jcyOvQ49u46HqhyeXQ2VxcXCTHSrprbmDvwp13j5QPtYLjG+ThQL0h
f3qJFgK4G/bsgelB01Yj3tEotGySMqT5PfLW6asjeya+4EpryKt9QgU+9LapClfQ
Ze10VTuHO7OvMZwhAkHgxZ4g/V2pKSdUVVMnr4lNbJgtImzyXqciAubKj+9wroBZ
YmDnwVgrptJRTl2zidqserKX9Nnmz7o7AcUi7vpP/EkkNUlKq2IWOf8J/RP/rSTZ
1QLSLnlWwcfQOpGUGpoR5nFAtoTnviofv2f+7+PrrZIEwgrNnt6rVxaZV+6d4P4H
4Lrfx0GK4UESrM0QT2b82D55wC65dVESVl1kvEWMrmX/xfchbgjloLNE71VsjUdK
mzgAQ1ZQlgbYOpQcOPWu/O9p8M9nMHoJPcpm3l/fh66/prAqRkzGfbdgvdh92i2f
k5G4t56aLBT8eftjtIVJljxNiWDChjXZUUyQ3SmNLJAnWMlhN/kVHqxJxYTIrmQy
WMHqFE0CAX6V/mOArKhSyTfrPiEog/AltKzkRYgbg60CAptPAwVTD5rY5FGuXws0
TnPQAAowwAdT1jKh0SoqnLL+akM3RqlcXiCJhYW4Dxt9Wod+DLp6YxkIrcFPCdxQ
7J7UUFsbj0DDETmwbams7CL198Fj7BiFxHBr2qsupm/h+svWbHdYCjntvzon02kw
pOlYQNCd3xhSj9KsI6EAZhHCpIsmGEhJeqb5ED9F4sCqo0nS+TZM0HEkhtkowBuP
1LWE7tuHSKiDWF5PU51OuQlsO67A4mDxdn6EJ9mT/sPNVI7LhxrtWkafMQBi2f1V
/+K/+8TB5YcaKwHkeyvTfAmN2p7qrGcETWYtjDDOvngwm3jKdY7dzHUE1rrN1/wA
DUOcZTbQpeMHDaWaOEjrgHAPu3MuwNbNFgPQAZhyOedn8kzI5WCci+XMPn/+lmhn
VFhIVgRs3O/XUFLy0ASCocxZWyXeWN9iZbfOe4aXJFeOc2HiO6eGQuBJ4ZFGup+v
ron6udwHa7kcIuJvBZ9jYW+wZ5F7ZPlE3nIKWI8AKo+NL+UYfrMirUSiMbWVXAcD
BPaP1Md+9XgrApSpXvYZMDDZHRXlvkN0uCsakyU8SRr90pXn3kVJ+HjLTY7oCXR+
rQ5/vrDZc1jkUR5meSuywdADYeAxPwcIGuK/aOqFyRyLQgO5uDBxp7gCalC38R1j
YeoAAQs/Fo9KTPQr+dYRqfYjRsZJ05CAm9wMVAGqMBNsSCTYUgd+Cw/d3Zaqxk48
rgvScpfmGQtkgaN3g2aHH/CExZXPkGz3ugPRnT6hveylnqMHTQRjl/Vv0kSNsHnK
gHhuJDJUm6wrh1d7l5jEG7jSOJAg3MpliXImZHDwGGH7UwW+hH5R0x37Mm4aollw
7gkafDUnUpolk78p+hLa9J7Xvt+INcd+kAmKAoy2x4XvKrq+LYC48pj19T11Q1Ec
5mBRMhRePZJ0Of7DBoTAgLi0lZiIu/km1YhzQKlpdYeFvaFVBPitVheRQ1Heonah
YzpR2/rCbWvyRf8gOXFCtLd/irqZQNDPPdIrW7/5cmMMvssnkkW4vIGMuOOP63q6
`protect END_PROTECTED
