`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
STs4gDj8iMy4ULd5NY7js89/V7Ot/mAOvxIDdqHEMDhmLwRPyMlLbjW5r1zFw/RO
S7DJoDkkOif2jJev8kITNDj9J2+w/t/95spWVmaOsck7t4Z+IRteMfux9Ph+3+dH
KYdhlePrYCR+fCi7sx3ViICTXBfI7tX9HE4J7F7Q+khltDxvvtoPqeGCr6mGI6wj
8w1gB1LvCi78/TMv4aFQbMZNjZQhs6P78qCQzqrrapkzvVjvKl4c+SxbFZd8eakf
PFD28pfyeIqWr+9X2LHZmd1M5997FKVpx0uBhDZ5DXJJlXBQAQvKs/mvvFgtb/aA
P3vj1SK8I06XzUelyN7S9LsaTXYwqD2rvsPqwkrUBL5mRTKaDxT4giGILTl5sxNy
1f7l72wTpnBIeiLmnYer8l1o3goUSjmKFh/JL5cwoAfqeRd/sVvkAwySCdYmEUSe
Uz8zYIFYIufJNT+PgIqtzo4P0mVqZCFghjzS/e1XrBu/Lsk0wgVBWmSSlRfbVMGs
LTJ7RgDoXnAdBbku6ZMnoJ5orj4rJToVdiD9C+gc5bJqXqzEZCe47qpGAlpgBpRz
EBwyRqmpeLftN1sTCLP0dedyzJoXlPIBNiAJePqvAJqqzKoie99USrowikQwubX4
Qv64B3cHQREClRfc3mE0a/dx9N/Hi3jyOw0YsGm4hkElaXUMeznrszQKW1OQAeSx
+AsFxV3ZxdM+fkKLqGWeCgVv0NE7INLbTlc3ysUJaR9eg+8+PREMJqp0Os/9yui0
mHk5rJGYTGXHr94YiuIJir2yPVKf1K8pmE32zDNj2dWYx2lbCkSQ8+0oh+Az0sk5
EUvYitFykVMIji0v45Bs22zI4YaJZnvkYlaWQWY71R0EVDlyFObNKhks6neLcpHA
YXL332Bp8U0Ph8n1JEFAnxkg5SVkyZUuToy+ERNwM/sTp6AzDawFDLaRahRQI7Ha
CyNyDiZYO4UgFq4AmTGHSOxnj/UOcrHlIaifWlo117Dw+0Zz9Ne+bksNq4toHSCP
jwcLSQdc8IklPt7Sz7oXAZelrpuEYm2fPyp+DnZqhIWbEuD9sRvtNU/nGOPkass/
PNl4H5pdPj6x6G4H2f16Xeh+9ytISnOVGlX/3Ahkq6iB5bouQV1CwPV5Tuqo1f8D
5rv96A2eRSf9zT4S/VsabvKHy9c5Ie64svcQcPtffyvhnZWx/kfHpubzxPwCD4yT
EzrG0a7b/kX0kT7GWyVlvLDm+/gDZeKWmKpjrXn7Twx7coCIdskqBQxujdlOvOnS
mU50UB5JLyHf5mHb2jQKPbKuysSNF/GdpDTj+zIF7mLGmJ1GYH+eIC3cWV0kgaLp
JZdAG7OiVV1PuayypiWuS5uyjYiNBE3wt3A61ZeIAv/6P0/H3z+yvAk7gMPVbYAP
FZPSXJ4C5rh/q2eOGyzZ4eVglfxzpXSddGwxxIkvaKmi/5NU1267TOTehhmPH826
VRtI5ZB4EdM1A/A22PIUH1DrlSbA6RHPhYbPBXU7WyQahEGq85Pc94MHLkDJiKSD
Z/KIEMgPtrR0aQYcMwueKq8QO/OIkfWW2qK2tLdEw0/Y2B9LFftoHUNDAJG4mLm9
fAcycaNM9NHns+7d1Z1InGljNPwmF14uCYaIkhmGZt+QDj2CxW/Mn0ABg53sstEl
8kuhSZkcIViBRcLqGLUoxyLOXt71wjwK64pVA9DMJGbgDBWB+4tCFH9wO/N9MEUD
gmToyprUBx/+kcHiuLY540m7ntPfiT8UQsNaWzvL3Re20idyakyapWlxF3sJ0plB
xfif5rvWZ0YqYtO05U9EvQ==
`protect END_PROTECTED
