library verilog;
use verilog.vl_types.all;
entity stratixv_hssi_gen3_pcie_hip is
    generic(
        func_mode       : string  := "disable";
        in_cvp_mode     : string  := "not_cvp_mode";
        bonding_mode    : string  := "bond_disable";
        prot_mode       : string  := "disabled_prot_mode";
        pcie_spec_1p0_compliance: string  := "spec_1p1";
        vc_enable       : string  := "single_vc";
        enable_slot_register: string  := "false";
        pcie_mode       : string  := "shared_mode";
        bypass_cdc      : string  := "false";
        enable_rx_reordering: string  := "true";
        enable_rx_buffer_checking: string  := "false";
        single_rx_detect_data: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        single_rx_detect: string  := "single_rx_detect";
        use_crc_forwarding: string  := "false";
        bypass_tl       : string  := "false";
        gen123_lane_rate_mode: string  := "gen1";
        lane_mask       : string  := "x4";
        disable_link_x2_support: string  := "false";
        national_inst_thru_enhance: string  := "true";
        hip_hard_reset  : string  := "enable";
        dis_paritychk   : string  := "enable";
        wrong_device_id : string  := "disable";
        data_pack_rx    : string  := "disable";
        ast_width       : string  := "rx_tx_64";
        ast_width_tx    : string  := "tx_64";
        ast_width_rx    : string  := "rx_64";
        tx_sop_ctrl     : string  := "boundary_64";
        rx_sop_ctrl     : string  := "boundary_64";
        rx_ast_parity   : string  := "disable";
        tx_ast_parity   : string  := "disable";
        ltssm_1ms_timeout: string  := "disable";
        ltssm_freqlocked_check: string  := "disable";
        deskew_comma    : string  := "com_deskw";
        dl_tx_check_parity_edb: string  := "disable";
        tl_tx_check_parity_msg: string  := "disable";
        port_link_number_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        port_link_number: string  := "port_link_number";
        device_number_data: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        device_number   : string  := "device_number";
        bypass_clk_switch: string  := "false";
        core_clk_out_sel: string  := "div_1";
        core_clk_divider: string  := "div_1";
        core_clk_source : string  := "pll_fixed_clk";
        core_clk_sel    : string  := "pld_clk";
        enable_ch0_pclk_out: string  := "pclk_ch01";
        enable_ch01_pclk_out: string  := "pclk_ch0";
        pipex1_debug_sel: string  := "disable";
        pclk_out_sel    : string  := "pclk";
        vendor_id_data  : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        vendor_id       : string  := "vendor_id";
        device_id_data  : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        device_id       : string  := "device_id";
        revision_id_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        revision_id     : string  := "revision_id";
        class_code_data : vl_logic_vector(0 to 23) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        class_code      : string  := "class_code";
        subsystem_vendor_id_data: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        subsystem_vendor_id: string  := "subsystem_vendor_id";
        subsystem_device_id_data: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        subsystem_device_id: string  := "subsystem_device_id";
        no_soft_reset   : string  := "false";
        maximum_current_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        maximum_current : string  := "maximum_current";
        d1_support      : string  := "false";
        d2_support      : string  := "false";
        d0_pme          : string  := "false";
        d1_pme          : string  := "false";
        d2_pme          : string  := "false";
        d3_hot_pme      : string  := "false";
        d3_cold_pme     : string  := "false";
        use_aer         : string  := "false";
        low_priority_vc : string  := "single_vc";
        vc_arbitration  : string  := "single_vc";
        disable_snoop_packet: string  := "false";
        max_payload_size: string  := "payload_512";
        surprise_down_error_support: string  := "false";
        dll_active_report_support: string  := "false";
        extend_tag_field: string  := "false";
        endpoint_l0_latency_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l0_latency: string  := "endpoint_l0_latency";
        endpoint_l1_latency_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l1_latency: string  := "endpoint_l1_latency";
        indicator_data  : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        indicator       : string  := "indicator";
        role_based_error_reporting: string  := "false";
        gen3_ltssm_debug: string  := "false";
        slot_power_scale_data: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        slot_power_scale: string  := "slot_power_scale";
        max_link_width  : string  := "x4";
        enable_l1_aspm  : string  := "false";
        enable_l0s_aspm : string  := "false";
        l1_exit_latency_sameclock_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_sameclock: string  := "l1_exit_latency_sameclock";
        l1_exit_latency_diffclock_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_diffclock: string  := "l1_exit_latency_diffclock";
        hot_plug_support_data: vl_logic_vector(0 to 6) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hot_plug_support: string  := "hot_plug_support";
        slot_power_limit_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_power_limit: string  := "slot_power_limit";
        slot_number_data: vl_logic_vector(0 to 12) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_number     : string  := "slot_number";
        diffclock_nfts_count_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        diffclock_nfts_count: string  := "diffclock_nfts_count";
        sameclock_nfts_count_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sameclock_nfts_count: string  := "sameclock_nfts_count";
        completion_timeout: string  := "abcd";
        enable_completion_timeout_disable: string  := "true";
        extended_tag_reset: string  := "false";
        ecrc_check_capable: string  := "true";
        ecrc_gen_capable: string  := "true";
        no_command_completed: string  := "true";
        msi_multi_message_capable: string  := "count_4";
        msi_64bit_addressing_capable: string  := "true";
        msi_masking_capable: string  := "false";
        msi_support     : string  := "true";
        interrupt_pin   : string  := "inta";
        ena_ido_req     : string  := "false";
        ena_ido_cpl     : string  := "false";
        enable_function_msix_support: string  := "true";
        msix_table_size_data: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_size : string  := "msix_table_size";
        msix_table_bir_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_table_bir  : string  := "msix_table_bir";
        msix_table_offset_data: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_offset: string  := "msix_table_offset";
        msix_pba_bir_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_pba_bir    : string  := "msix_pba_bir";
        msix_pba_offset_data: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_pba_offset : string  := "msix_pba_offset";
        bridge_port_vga_enable: string  := "false";
        bridge_port_ssid_support: string  := "false";
        ssvid_data      : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssvid           : string  := "ssvid";
        ssid_data       : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssid            : string  := "ssid";
        eie_before_nfts_count_data: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        eie_before_nfts_count: string  := "eie_before_nfts_count";
        gen2_diffclock_nfts_count_data: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_diffclock_nfts_count: string  := "gen2_diffclock_nfts_count";
        gen2_sameclock_nfts_count_data: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_sameclock_nfts_count: string  := "gen2_sameclock_nfts_count";
        deemphasis_enable: string  := "false";
        pcie_spec_version: string  := "v2";
        l0_exit_latency_sameclock_data: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_sameclock: string  := "l0_exit_latency_sameclock";
        l0_exit_latency_diffclock_data: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_diffclock: string  := "l0_exit_latency_diffclock";
        rx_ei_l0s       : string  := "disable";
        l2_async_logic  : string  := "enable";
        aspm_config_management: string  := "true";
        atomic_op_routing: string  := "false";
        atomic_op_completer_32bit: string  := "false";
        atomic_op_completer_64bit: string  := "false";
        cas_completer_128bit: string  := "false";
        ltr_mechanism   : string  := "false";
        tph_completer   : string  := "false";
        extended_format_field: string  := "false";
        atomic_malformed: string  := "false";
        flr_capability  : string  := "true";
        enable_adapter_half_rate_mode: string  := "false";
        vc0_clk_enable  : string  := "true";
        vc1_clk_enable  : string  := "false";
        register_pipe_signals: string  := "false";
        bar0_io_space   : string  := "false";
        bar0_64bit_mem_space: string  := "true";
        bar0_prefetchable: string  := "true";
        bar0_size_mask_data: vl_logic_vector(0 to 27) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        bar0_size_mask  : string  := "bar0_size_mask";
        bar1_io_space   : string  := "false";
        bar1_64bit_mem_space: string  := "false";
        bar1_prefetchable: string  := "false";
        bar1_size_mask_data: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar1_size_mask  : string  := "bar1_size_mask";
        bar2_io_space   : string  := "false";
        bar2_64bit_mem_space: string  := "false";
        bar2_prefetchable: string  := "false";
        bar2_size_mask_data: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar2_size_mask  : string  := "bar2_size_mask";
        bar3_io_space   : string  := "false";
        bar3_64bit_mem_space: string  := "false";
        bar3_prefetchable: string  := "false";
        bar3_size_mask_data: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar3_size_mask  : string  := "bar3_size_mask";
        bar4_io_space   : string  := "false";
        bar4_64bit_mem_space: string  := "false";
        bar4_prefetchable: string  := "false";
        bar4_size_mask_data: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar4_size_mask  : string  := "bar4_size_mask";
        bar5_io_space   : string  := "false";
        bar5_64bit_mem_space: string  := "false";
        bar5_prefetchable: string  := "false";
        bar5_size_mask_data: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar5_size_mask  : string  := "bar5_size_mask";
        expansion_base_address_register_data: integer := 0;
        expansion_base_address_register: string  := "expansion_base_address_register";
        io_window_addr_width: string  := "window_32_bit";
        prefetchable_mem_window_addr_width: string  := "prefetch_32";
        skp_os_gen3_count_data: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        skp_os_gen3_count: string  := "skp_os_gen3_count";
        rx_cdc_almost_empty_data: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        rx_cdc_almost_empty: string  := "rx_cdc_almost_empty";
        tx_cdc_almost_empty_data: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        tx_cdc_almost_empty: string  := "tx_cdc_almost_empty";
        rx_cdc_almost_full_data: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        rx_cdc_almost_full: string  := "rx_cdc_almost_full";
        tx_cdc_almost_full_data: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        tx_cdc_almost_full: string  := "tx_cdc_almost_full";
        rx_l0s_count_idl_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_l0s_count_idl: string  := "rx_l0s_count_idl";
        cdc_dummy_insert_limit_data: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        cdc_dummy_insert_limit: string  := "cdc_dummy_insert_limit";
        ei_delay_powerdown_count_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        ei_delay_powerdown_count: string  := "ei_delay_powerdown_count";
        millisecond_cycle_count_data: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        millisecond_cycle_count: string  := "millisecond_cycle_count";
        skp_os_schedule_count_data: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        skp_os_schedule_count: string  := "skp_os_schedule_count";
        fc_init_timer_data: vl_logic_vector(0 to 10) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        fc_init_timer   : string  := "fc_init_timer";
        l01_entry_latency_data: vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi1, Hi1, Hi1);
        l01_entry_latency: string  := "l01_entry_latency";
        flow_control_update_count_data: vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi1, Hi1, Hi0);
        flow_control_update_count: string  := "flow_control_update_count";
        flow_control_timeout_count_data: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        flow_control_timeout_count: string  := "flow_control_timeout_count";
        vc0_rx_flow_ctrl_posted_header_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        vc0_rx_flow_ctrl_posted_header: string  := "vc0_rx_flow_ctrl_posted_header";
        vc0_rx_flow_ctrl_posted_data_data: vl_logic_vector(0 to 11) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        vc0_rx_flow_ctrl_posted_data: string  := "vc0_rx_flow_ctrl_posted_data";
        vc0_rx_flow_ctrl_nonposted_header_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0);
        vc0_rx_flow_ctrl_nonposted_header: string  := "vc0_rx_flow_ctrl_nonposted_header";
        vc0_rx_flow_ctrl_nonposted_data_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        vc0_rx_flow_ctrl_nonposted_data: string  := "vc0_rx_flow_ctrl_nonposted_data";
        vc0_rx_flow_ctrl_compl_header_data: vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        vc0_rx_flow_ctrl_compl_header: string  := "vc0_rx_flow_ctrl_compl_header";
        vc0_rx_flow_ctrl_compl_data_data: vl_logic_vector(0 to 11) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        vc0_rx_flow_ctrl_compl_data: string  := "vc0_rx_flow_ctrl_compl_data";
        rx_ptr0_posted_dpram_min_data: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_ptr0_posted_dpram_min: string  := "rx_ptr0_posted_dpram_min";
        rx_ptr0_posted_dpram_max_data: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_ptr0_posted_dpram_max: string  := "rx_ptr0_posted_dpram_max";
        rx_ptr0_nonposted_dpram_min_data: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_ptr0_nonposted_dpram_min: string  := "rx_ptr0_nonposted_dpram_min";
        rx_ptr0_nonposted_dpram_max_data: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_ptr0_nonposted_dpram_max: string  := "rx_ptr0_nonposted_dpram_max";
        retry_buffer_last_active_address_data: vl_logic_vector(0 to 9) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        retry_buffer_last_active_address: string  := "retry_buffer_last_active_address";
        retry_buffer_memory_settings_data: vl_logic_vector(0 to 52) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        retry_buffer_memory_settings: string  := "retry_buffer_memory_settings";
        vc0_rx_buffer_memory_settings_data: vl_logic_vector(0 to 52) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        vc0_rx_buffer_memory_settings: string  := "vc0_rx_buffer_memory_settings";
        bist_memory_settings_data: vl_logic_vector(0 to 74) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bist_memory_settings: string  := "bist_memory_settings";
        credit_buffer_allocation_aux: string  := "balanced";
        iei_enable_settings: string  := "gen2_infei_infsd_gen1_infei_sd";
        vsec_id_data    : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        vsec_id         : string  := "vsec_id";
        cvp_rate_sel    : string  := "full_rate";
        hard_reset_bypass: string  := "false";
        cvp_data_compressed: string  := "false";
        cvp_data_encrypted: string  := "false";
        cvp_mode_reset  : string  := "false";
        cvp_clk_reset   : string  := "false";
        vsec_rev_data   : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        vsec_rev        : string  := "vsec_rev";
        jtag_id_data    : vl_logic_vector(0 to 127) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        jtag_id         : string  := "jtag_id";
        user_id_data    : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        user_id         : string  := "user_id";
        cseb_extend_pci : string  := "false";
        cseb_extend_pcie: string  := "false";
        cseb_cpl_status_during_cvp: string  := "config_retry_status";
        cseb_route_to_avl_rx_st: string  := "cseb";
        cseb_config_bypass: string  := "disable";
        cseb_cpl_tag_checking: string  := "enable";
        cseb_bar_match_checking: string  := "enable";
        cseb_min_error_checking: string  := "false";
        cseb_temp_busy_crs: string  := "completer_abort";
        cseb_disable_auto_crs: string  := "false";
        gen3_diffclock_nfts_count_data: vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_diffclock_nfts_count: string  := "g3_diffclock_nfts_count";
        gen3_sameclock_nfts_count_data: vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_sameclock_nfts_count: string  := "g3_sameclock_nfts_count";
        gen3_coeff_errchk: string  := "enable";
        gen3_paritychk  : string  := "enable";
        gen3_coeff_delay_count_data: vl_logic_vector(0 to 6) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1);
        gen3_coeff_delay_count: string  := "g3_coeff_dly_count";
        gen3_coeff_1_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_1    : string  := "g3_coeff_1";
        gen3_coeff_1_sel: string  := "coeff_1";
        gen3_coeff_1_preset_hint_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_1_preset_hint: string  := "g3_coeff_1_prst_hint";
        gen3_coeff_1_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi0);
        gen3_coeff_1_nxtber_more: string  := "g3_coeff_1_nxtber_more";
        gen3_coeff_1_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi0);
        gen3_coeff_1_nxtber_less: string  := "g3_coeff_1_nxtber_less";
        gen3_coeff_1_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_1_reqber: string  := "g3_coeff_1_reqber";
        gen3_coeff_1_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_1_ber_meas: string  := "g3_coeff_1_ber_meas";
        gen3_coeff_2_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_2    : string  := "g3_coeff_2";
        gen3_coeff_2_sel: string  := "coeff_2";
        gen3_coeff_2_preset_hint_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        gen3_coeff_2_preset_hint: string  := "g3_coeff_2_prst_hint";
        gen3_coeff_2_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_2_nxtber_more: string  := "g3_coeff_2_nxtber_more";
        gen3_coeff_2_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_2_nxtber_less: string  := "g3_coeff_2_nxtber_less";
        gen3_coeff_2_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_2_reqber: string  := "g3_coeff_2_reqber";
        gen3_coeff_2_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_2_ber_meas: string  := "g3_coeff_1_ber_meas";
        gen3_coeff_3_data: vl_logic_vector(0 to 17) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_3    : string  := "g3_coeff_3";
        gen3_coeff_3_sel: string  := "coeff_3";
        gen3_coeff_3_preset_hint_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_3_preset_hint: string  := "g3_coeff_3_prst_hint";
        gen3_coeff_3_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        gen3_coeff_3_nxtber_more: string  := "g3_coeff_3_nxtber_more";
        gen3_coeff_3_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_3_nxtber_less: string  := "g3_coeff_3_nxtber_less";
        gen3_coeff_3_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_3_reqber: string  := "g3_coeff_3_reqber";
        gen3_coeff_3_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_3_ber_meas: string  := "g3_coeff_3_ber_meas";
        gen3_coeff_4_data: vl_logic_vector(0 to 17) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_4    : string  := "g3_coeff_4";
        gen3_coeff_4_sel: string  := "coeff_4";
        gen3_coeff_4_preset_hint_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_4_preset_hint: string  := "g3_coeff_4_prst_hint";
        gen3_coeff_4_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_4_nxtber_more: string  := "g3_coeff_4_nxtber_more";
        gen3_coeff_4_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_4_nxtber_less: string  := "g3_coeff_4_nxtber_less";
        gen3_coeff_4_reqber_data: vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi0, Hi1);
        gen3_coeff_4_reqber: string  := "g3_coeff_4_reqber";
        gen3_coeff_4_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_4_ber_meas: string  := "g3_coeff_4_ber_meas";
        gen3_coeff_5_data: vl_logic_vector(0 to 17) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_5    : string  := "g3_coeff_5";
        gen3_coeff_5_sel: string  := "coeff_5";
        gen3_coeff_5_preset_hint_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        gen3_coeff_5_preset_hint: string  := "g3_coeff_5_prst_hint";
        gen3_coeff_5_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        gen3_coeff_5_nxtber_more: string  := "g3_coeff_5_nxtber_more";
        gen3_coeff_5_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_5_nxtber_less: string  := "g3_coeff_5_nxtber_less";
        gen3_coeff_5_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_5_reqber: string  := "g3_coeff_5_reqber";
        gen3_coeff_5_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_5_ber_meas: string  := "g3_coeff_5_ber_meas";
        gen3_coeff_6_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_6    : string  := "g3_coeff_6";
        gen3_coeff_6_sel: string  := "coeff_6";
        gen3_coeff_6_preset_hint_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        gen3_coeff_6_preset_hint: string  := "g3_coeff_6_prst_hint";
        gen3_coeff_6_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi0);
        gen3_coeff_6_nxtber_more: string  := "g3_coeff_6_nxtber_more";
        gen3_coeff_6_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_6_nxtber_less: string  := "g3_coeff_6_nxtber_less";
        gen3_coeff_6_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_6_reqber: string  := "g3_coeff_6_reqber";
        gen3_coeff_6_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_6_ber_meas: string  := "g3_coeff_6_ber_meas";
        gen3_coeff_7_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_7    : string  := "g3_coeff_7";
        gen3_coeff_7_sel: string  := "coeff_7";
        gen3_coeff_7_preset_hint_data: vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        gen3_coeff_7_preset_hint: string  := "g3_coeff_7_prst_hint";
        gen3_coeff_7_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_7_nxtber_more: string  := "g3_coeff_7_nxtber_more";
        gen3_coeff_7_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_7_nxtber_less: string  := "g3_coeff_7_nxtber_less";
        gen3_coeff_7_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_7_reqber: string  := "g3_coeff_7_reqber";
        gen3_coeff_7_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_7_ber_meas: string  := "g3_coeff_7_ber_meas";
        gen3_coeff_8_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_8    : string  := "g3_coeff_8";
        gen3_coeff_8_sel: string  := "coeff_8";
        gen3_coeff_8_preset_hint_data: vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        gen3_coeff_8_preset_hint: string  := "g3_coeff_8_prst_hint";
        gen3_coeff_8_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi0);
        gen3_coeff_8_nxtber_more: string  := "g3_coeff_8_nxtber_more";
        gen3_coeff_8_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_8_nxtber_less: string  := "g3_coeff_8_nxtber_less";
        gen3_coeff_8_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_8_reqber: string  := "g3_coeff_8_reqber";
        gen3_coeff_8_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_8_ber_meas: string  := "g3_coeff_8_ber_meas";
        gen3_coeff_9_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_9    : string  := "g3_coeff_9";
        gen3_coeff_9_sel: string  := "coeff_9";
        gen3_coeff_9_preset_hint_data: vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        gen3_coeff_9_preset_hint: string  := "g3_coeff_9_prst_hint";
        gen3_coeff_9_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi1);
        gen3_coeff_9_nxtber_more: string  := "g3_coeff_9_nxtber_more";
        gen3_coeff_9_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi1);
        gen3_coeff_9_nxtber_less: string  := "g3_coeff_9_nxtber_less";
        gen3_coeff_9_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_9_reqber: string  := "g3_coeff_9_reqber";
        gen3_coeff_9_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_9_ber_meas: string  := "g3_coeff_9_ber_meas";
        gen3_coeff_10_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_10   : string  := "g3_coeff_10";
        gen3_coeff_10_sel: string  := "coeff_10";
        gen3_coeff_10_preset_hint_data: vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        gen3_coeff_10_preset_hint: string  := "g3_coeff_10_prst_hint";
        gen3_coeff_10_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi0);
        gen3_coeff_10_nxtber_more: string  := "g3_coeff_10_nxtber_more";
        gen3_coeff_10_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_10_nxtber_less: string  := "g3_coeff_10_nxtber_less";
        gen3_coeff_10_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_10_reqber: string  := "g3_coeff_10_reqber";
        gen3_coeff_10_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_10_ber_meas: string  := "g3_coeff_10_ber_meas";
        gen3_coeff_11_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_11   : string  := "g3_coeff_11";
        gen3_coeff_11_sel: string  := "coeff_11";
        gen3_coeff_11_preset_hint_data: vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        gen3_coeff_11_preset_hint: string  := "g3_coeff_11_prst_hint";
        gen3_coeff_11_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_11_nxtber_more: string  := "g3_coeff_11_nxtber_more";
        gen3_coeff_11_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_11_nxtber_less: string  := "g3_coeff_11_nxtber_less";
        gen3_coeff_11_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_11_reqber: string  := "g3_coeff_11_reqber";
        gen3_coeff_11_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_11_ber_meas: string  := "g3_coeff_11_ber_meas";
        gen3_coeff_12_data: vl_logic_vector(0 to 17) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_12   : string  := "g3_coeff_12";
        gen3_coeff_12_sel: string  := "coeff_12";
        gen3_coeff_12_preset_hint_data: vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        gen3_coeff_12_preset_hint: string  := "g3_coeff_12_prst_hint";
        gen3_coeff_12_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_12_nxtber_more: string  := "g3_coeff_12_nxtber_more";
        gen3_coeff_12_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_12_nxtber_less: string  := "g3_coeff_12_nxtber_less";
        gen3_coeff_12_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_12_reqber: string  := "g3_coeff_12_reqber";
        gen3_coeff_12_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_12_ber_meas: string  := "g3_coeff_12_ber_meas";
        gen3_coeff_13_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_13   : string  := "g3_coeff_13";
        gen3_coeff_13_sel: string  := "coeff_13";
        gen3_coeff_13_preset_hint_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        gen3_coeff_13_preset_hint: string  := "g3_coeff_13_prst_hint";
        gen3_coeff_13_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_13_nxtber_more: string  := "g3_coeff_13_nxtber_more";
        gen3_coeff_13_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi1);
        gen3_coeff_13_nxtber_less: string  := "g3_coeff_13_nxtber_less";
        gen3_coeff_13_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_13_reqber: string  := "g3_coeff_13_reqber";
        gen3_coeff_13_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_13_ber_meas: string  := "g3_coeff_13_ber_meas";
        gen3_coeff_14_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_14   : string  := "g3_coeff_14";
        gen3_coeff_14_sel: string  := "coeff_14";
        gen3_coeff_14_preset_hint_data: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_14_preset_hint: string  := "g3_coeff_14_prst_hint";
        gen3_coeff_14_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_14_nxtber_more: string  := "g3_coeff_14_nxtber_more";
        gen3_coeff_14_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi0);
        gen3_coeff_14_nxtber_less: string  := "g3_coeff_14_nxtber_less";
        gen3_coeff_14_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_14_reqber: string  := "g3_coeff_14_reqber";
        gen3_coeff_14_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_14_ber_meas: string  := "g3_coeff_14_ber_meas";
        gen3_coeff_15_data: vl_logic_vector(0 to 17) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_15   : string  := "g3_coeff_15";
        gen3_coeff_15_sel: string  := "coeff_15";
        gen3_coeff_15_preset_hint_data: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        gen3_coeff_15_preset_hint: string  := "g3_coeff_15_prst_hint";
        gen3_coeff_15_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_15_nxtber_more: string  := "g3_coeff_15_nxtber_more";
        gen3_coeff_15_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_15_nxtber_less: string  := "g3_coeff_15_nxtber_less";
        gen3_coeff_15_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_15_reqber: string  := "g3_coeff_15_reqber";
        gen3_coeff_15_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_15_ber_meas: string  := "g3_coeff_15_ber_meas";
        gen3_coeff_16_data: vl_logic_vector(0 to 17) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_16   : string  := "g3_coeff_16";
        gen3_coeff_16_sel: string  := "coeff_16";
        gen3_coeff_16_preset_hint_data: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        gen3_coeff_16_preset_hint: string  := "g3_coeff_16_prst_hint";
        gen3_coeff_16_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_16_nxtber_more: string  := "g3_coeff_16_nxtber_more";
        gen3_coeff_16_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_16_nxtber_less: string  := "g3_coeff_16_nxtber_less";
        gen3_coeff_16_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_16_reqber: string  := "g3_coeff_16_reqber";
        gen3_coeff_16_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_16_ber_meas: string  := "g3_coeff_16_ber_meas";
        gen3_coeff_17_data: vl_logic_vector(0 to 17) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_17   : string  := "g3_coeff_17";
        gen3_coeff_17_sel: string  := "coeff_17";
        gen3_coeff_17_preset_hint_data: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        gen3_coeff_17_preset_hint: string  := "g3_coeff_17_prst_hint";
        gen3_coeff_17_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_17_nxtber_more: string  := "g3_coeff_17_nxtber_more";
        gen3_coeff_17_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_17_nxtber_less: string  := "g3_coeff_17_nxtber_less";
        gen3_coeff_17_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_17_reqber: string  := "g3_coeff_17_reqber";
        gen3_coeff_17_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_17_ber_meas: string  := "g3_coeff_17_ber_meas";
        gen3_coeff_18_data: vl_logic_vector(0 to 17) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_18   : string  := "g3_coeff_18";
        gen3_coeff_18_sel: string  := "coeff_18";
        gen3_coeff_18_preset_hint_data: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        gen3_coeff_18_preset_hint: string  := "g3_coeff_18_prst_hint";
        gen3_coeff_18_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_18_nxtber_more: string  := "g3_coeff_18_nxtber_more";
        gen3_coeff_18_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_18_nxtber_less: string  := "g3_coeff_18_nxtber_less";
        gen3_coeff_18_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_18_reqber: string  := "g3_coeff_18_reqber";
        gen3_coeff_18_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_18_ber_meas: string  := "g3_coeff_18_ber_meas";
        gen3_coeff_19_data: vl_logic_vector(0 to 17) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_19   : string  := "g3_coeff_19";
        gen3_coeff_19_sel: string  := "coeff_19";
        gen3_coeff_19_preset_hint_data: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        gen3_coeff_19_preset_hint: string  := "g3_coeff_19_prst_hint";
        gen3_coeff_19_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_19_nxtber_more: string  := "g3_coeff_19_nxtber_more";
        gen3_coeff_19_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_19_nxtber_less: string  := "g3_coeff_19_nxtber_less";
        gen3_coeff_19_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_19_reqber: string  := "g3_coeff_19_reqber";
        gen3_coeff_19_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_19_ber_meas: string  := "g3_coeff_19_ber_meas";
        gen3_coeff_20_data: vl_logic_vector(0 to 17) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_20   : string  := "g3_coeff_20";
        gen3_coeff_20_sel: string  := "coeff_20";
        gen3_coeff_20_preset_hint_data: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        gen3_coeff_20_preset_hint: string  := "g3_coeff_20_prst_hint";
        gen3_coeff_20_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_20_nxtber_more: string  := "g3_coeff_20_nxtber_more";
        gen3_coeff_20_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_20_nxtber_less: string  := "g3_coeff_20_nxtber_less";
        gen3_coeff_20_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_20_reqber: string  := "g3_coeff_20_reqber";
        gen3_coeff_20_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_20_ber_meas: string  := "g3_coeff_20_ber_meas";
        gen3_coeff_21_data: vl_logic_vector(0 to 17) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_21   : string  := "g3_coeff_21";
        gen3_coeff_21_sel: string  := "coeff_21";
        gen3_coeff_21_preset_hint_data: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        gen3_coeff_21_preset_hint: string  := "g3_coeff_21_prst_hint";
        gen3_coeff_21_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_21_nxtber_more: string  := "g3_coeff_21_nxtber_more";
        gen3_coeff_21_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_21_nxtber_less: string  := "g3_coeff_21_nxtber_less";
        gen3_coeff_21_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_21_reqber: string  := "g3_coeff_21_reqber";
        gen3_coeff_21_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_21_ber_meas: string  := "g3_coeff_21_ber_meas";
        gen3_coeff_22_data: vl_logic_vector(0 to 17) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_22   : string  := "g3_coeff_22";
        gen3_coeff_22_sel: string  := "coeff_22";
        gen3_coeff_22_preset_hint_data: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        gen3_coeff_22_preset_hint: string  := "g3_coeff_22_prst_hint";
        gen3_coeff_22_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_22_nxtber_more: string  := "g3_coeff_22_nxtber_more";
        gen3_coeff_22_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_22_nxtber_less: string  := "g3_coeff_22_nxtber_less";
        gen3_coeff_22_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_22_reqber: string  := "g3_coeff_22_reqber";
        gen3_coeff_22_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_22_ber_meas: string  := "g3_coeff_22_ber_meas";
        gen3_coeff_23_data: vl_logic_vector(0 to 17) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_23   : string  := "g3_coeff_23";
        gen3_coeff_23_sel: string  := "coeff_23";
        gen3_coeff_23_preset_hint_data: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        gen3_coeff_23_preset_hint: string  := "g3_coeff_23_prst_hint";
        gen3_coeff_23_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_23_nxtber_more: string  := "g3_coeff_23_nxtber_more";
        gen3_coeff_23_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_23_nxtber_less: string  := "g3_coeff_23_nxtber_less";
        gen3_coeff_23_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_23_reqber: string  := "g3_coeff_23_reqber";
        gen3_coeff_23_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_23_ber_meas: string  := "g3_coeff_23_ber_meas";
        gen3_coeff_24_data: vl_logic_vector(0 to 17) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_24   : string  := "g3_coeff_24";
        gen3_coeff_24_sel: string  := "coeff_24";
        gen3_coeff_24_preset_hint_data: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        gen3_coeff_24_preset_hint: string  := "g3_coeff_24_prst_hint";
        gen3_coeff_24_nxtber_more_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_24_nxtber_more: string  := "g3_coeff_24_nxtber_more";
        gen3_coeff_24_nxtber_less_ptr: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_24_nxtber_less: string  := "g3_coeff_24_nxtber_less";
        gen3_coeff_24_reqber_data: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_24_reqber: string  := "g3_coeff_24_reqber";
        gen3_coeff_24_ber_meas_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_24_ber_meas: string  := "g3_coeff_24_ber_meas";
        gen3_preset_coeff_1_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_preset_coeff_1: string  := "g3_prst_coeff_1";
        gen3_preset_coeff_2_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_preset_coeff_2: string  := "g3_prst_coeff_2";
        gen3_preset_coeff_3_data: vl_logic_vector(0 to 17) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_preset_coeff_3: string  := "g3_prst_coeff_3";
        gen3_preset_coeff_4_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        gen3_preset_coeff_4: string  := "g3_prst_coeff_4";
        gen3_preset_coeff_5_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        gen3_preset_coeff_5: string  := "g3_prst_coeff_5";
        gen3_preset_coeff_6_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        gen3_preset_coeff_6: string  := "g3_prst_coeff_6";
        gen3_preset_coeff_7_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        gen3_preset_coeff_7: string  := "g3_prst_coeff_7";
        gen3_preset_coeff_8_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        gen3_preset_coeff_8: string  := "g3_prst_coeff_8";
        gen3_preset_coeff_9_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_preset_coeff_9: string  := "g3_prst_coeff_9";
        gen3_preset_coeff_10_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_preset_coeff_10: string  := "g3_prst_coeff_10";
        gen3_preset_coeff_11_data: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_preset_coeff_11: string  := "g3_prst_coeff_11";
        gen3_rxfreqlock_counter_data: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_rxfreqlock_counter: string  := "g3_rxfreqlock_count";
        gen3_low_freq_data: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1);
        gen3_low_freq   : string  := "g3_low_freq";
        gen3_full_swing_data: vl_logic_vector(0 to 5) := (Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        gen3_full_swing : string  := "g3_full_swing";
        pld_in_use_reg  : string  := "false";
        k_cfg_parchk_ena: string  := "disable";
        k_dis_cplovf    : string  := "disable";
        rpltim_set      : string  := "false";
        rpltim_base_data: vl_logic_vector(0 to 12) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        acknak_set      : string  := "false";
        acknak_base_data: vl_logic_vector(0 to 12) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_use_prst     : string  := "false";
        rx_use_prst_ep  : string  := "false";
        rstctrl_pld_clr : string  := "false";
        rstctrl_debug_en: string  := "false";
        rstctrl_force_inactive_rst: string  := "false";
        rstctrl_perst_enable: string  := "level";
        hrdrstctrl_en   : string  := "hrdrstctrl_dis";
        rstctrl_hip_ep  : string  := "hip_ep";
        rstctrl_hard_block_enable: string  := "hard_rst_ctl";
        rstctrl_rx_pma_rstb_inv: string  := "false";
        rstctrl_tx_pma_rstb_inv: string  := "false";
        rstctrl_rx_pcs_rst_n_inv: string  := "false";
        rstctrl_tx_pcs_rst_n_inv: string  := "false";
        rstctrl_altpe3_crst_n_inv: string  := "false";
        rstctrl_altpe3_srst_n_inv: string  := "false";
        rstctrl_altpe3_rst_n_inv: string  := "false";
        rstctrl_tx_pma_syncp_inv: string  := "false";
        rstctrl_1us_count_fref_clk: string  := "rstctrl_1us_cnt";
        rstctrl_1us_count_fref_clk_value: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        rstctrl_1ms_count_fref_clk: string  := "rstctrl_1ms_cnt";
        rstctrl_1ms_count_fref_clk_value: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        rstctrl_off_cal_done_select: string  := "not_active";
        rstctrl_rx_pma_rstb_select: string  := "not_active";
        rstctrl_rx_pma_rstb_cmu_select: string  := "not_active";
        rstctrl_rx_pll_freq_lock_select: string  := "not_active";
        rstctrl_mask_tx_pll_lock_select: string  := "not_active";
        rstctrl_rx_pll_lock_select: string  := "not_active";
        rstctrl_perstn_select: string  := "perstn_pin";
        rstctrl_tx_lc_pll_rstb_select: string  := "not_active";
        rstctrl_fref_clk_select: string  := "ch0_sel";
        rstctrl_off_cal_en_select: string  := "not_active";
        rstctrl_tx_pma_syncp_select: string  := "not_active";
        rstctrl_rx_pcs_rst_n_select: string  := "not_active";
        rstctrl_tx_cmu_pll_lock_select: string  := "not_active";
        rstctrl_tx_pcs_rst_n_select: string  := "not_active";
        rstctrl_tx_lc_pll_lock_select: string  := "not_active";
        rstctrl_timer_a : string  := "rstctrl_timer_a";
        rstctrl_timer_a_type: string  := "milli_secs";
        rstctrl_timer_a_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        rstctrl_timer_b : string  := "rstctrl_timer_b";
        rstctrl_timer_b_type: string  := "milli_secs";
        rstctrl_timer_b_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        rstctrl_timer_c : string  := "rstctrl_timer_c";
        rstctrl_timer_c_type: string  := "milli_secs";
        rstctrl_timer_c_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        rstctrl_timer_d : string  := "rstctrl_timer_d";
        rstctrl_timer_d_type: string  := "milli_secs";
        rstctrl_timer_d_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        rstctrl_timer_e : string  := "rstctrl_timer_e";
        rstctrl_timer_e_type: string  := "milli_secs";
        rstctrl_timer_e_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        rstctrl_timer_f : string  := "rstctrl_timer_f";
        rstctrl_timer_f_type: string  := "milli_secs";
        rstctrl_timer_f_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        rstctrl_timer_g : string  := "rstctrl_timer_g";
        rstctrl_timer_g_type: string  := "milli_secs";
        rstctrl_timer_g_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        rstctrl_timer_h : string  := "rstctrl_timer_h";
        rstctrl_timer_h_type: string  := "milli_secs";
        rstctrl_timer_h_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        rstctrl_timer_i : string  := "rstctrl_timer_i";
        rstctrl_timer_i_type: string  := "milli_secs";
        rstctrl_timer_i_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        rstctrl_timer_j : string  := "rstctrl_timer_j";
        rstctrl_timer_j_type: string  := "milli_secs";
        rstctrl_timer_j_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        g3_redo_equlz_dis: string  := "false";
        g3_quiesce_guarant: string  := "false";
        en_lane_errchk  : string  := "false";
        g3_force_ber_max: string  := "false";
        en_phystatus_dly: string  := "false";
        rstctl_ltssm_dis: string  := "false";
        force_dis_to_det: string  := "false";
        g3_redo_equlz_en: string  := "false";
        tl_cfg_div      : string  := "cfg_clk_div_7";
        g3_dis_be_frm_err: string  := "false";
        g3_ltssm_eq_dbg : string  := "false";
        g3_lnk_trn_rx_ts: string  := "false";
        g3_force_ber_min: string  := "false";
        force_gen1_dis  : string  := "false";
        g3_bypass_equlz : string  := "false";
        gen3_skip_ph2_ph3: string  := "true";
        gen3_dcbal_en   : string  := "true";
        early_dl_up     : string  := "true"
    );
    port(
        dpriostatus     : out    vl_logic_vector(15 downto 0);
        lmidout         : out    vl_logic_vector(31 downto 0);
        lmiack          : out    vl_logic_vector(0 downto 0);
        lmirden         : in     vl_logic_vector(0 downto 0);
        lmiwren         : in     vl_logic_vector(0 downto 0);
        lmiaddr         : in     vl_logic_vector(11 downto 0);
        lmidin          : in     vl_logic_vector(31 downto 0);
        flrreset        : in     vl_logic_vector(0 downto 0);
        flrsts          : out    vl_logic_vector(0 downto 0);
        resetstatus     : out    vl_logic_vector(0 downto 0);
        l2exit          : out    vl_logic_vector(0 downto 0);
        hotrstexit      : out    vl_logic_vector(0 downto 0);
        dlupexit        : out    vl_logic_vector(0 downto 0);
        coreclkout      : out    vl_logic_vector(0 downto 0);
        pldclk          : in     vl_logic_vector(0 downto 0);
        pldsrst         : in     vl_logic_vector(0 downto 0);
        pldrst          : in     vl_logic_vector(0 downto 0);
        pclkch0         : in     vl_logic_vector(0 downto 0);
        pclkch1         : in     vl_logic_vector(0 downto 0);
        pclkcentral     : in     vl_logic_vector(0 downto 0);
        pllfixedclkch0  : in     vl_logic_vector(0 downto 0);
        pllfixedclkch1  : in     vl_logic_vector(0 downto 0);
        pllfixedclkcentral: in     vl_logic_vector(0 downto 0);
        phyrst          : in     vl_logic_vector(0 downto 0);
        physrst         : in     vl_logic_vector(0 downto 0);
        coreclkin       : in     vl_logic_vector(0 downto 0);
        corerst         : in     vl_logic_vector(0 downto 0);
        corepor         : in     vl_logic_vector(0 downto 0);
        corecrst        : in     vl_logic_vector(0 downto 0);
        coresrst        : in     vl_logic_vector(0 downto 0);
        swdnout         : out    vl_logic_vector(6 downto 0);
        swupout         : out    vl_logic_vector(2 downto 0);
        swdnin          : in     vl_logic_vector(2 downto 0);
        swupin          : in     vl_logic_vector(6 downto 0);
        swctmod         : in     vl_logic_vector(1 downto 0);
        rxstdata        : out    vl_logic_vector(255 downto 0);
        rxstparity      : out    vl_logic_vector(31 downto 0);
        rxstbe          : out    vl_logic_vector(31 downto 0);
        rxsterr         : out    vl_logic_vector(3 downto 0);
        rxstsop         : out    vl_logic_vector(3 downto 0);
        rxsteop         : out    vl_logic_vector(3 downto 0);
        rxstempty       : out    vl_logic_vector(1 downto 0);
        rxstvalid       : out    vl_logic_vector(3 downto 0);
        rxstbardec1     : out    vl_logic_vector(7 downto 0);
        rxstbardec2     : out    vl_logic_vector(7 downto 0);
        rxstmask        : in     vl_logic_vector(0 downto 0);
        rxstready       : in     vl_logic_vector(0 downto 0);
        txstready       : out    vl_logic_vector(0 downto 0);
        txcredfchipcons : out    vl_logic_vector(5 downto 0);
        txcredfcinfinite: out    vl_logic_vector(5 downto 0);
        txcredhdrfcp    : out    vl_logic_vector(7 downto 0);
        txcreddatafcp   : out    vl_logic_vector(11 downto 0);
        txcredhdrfcnp   : out    vl_logic_vector(7 downto 0);
        txcreddatafcnp  : out    vl_logic_vector(11 downto 0);
        txcredhdrfccp   : out    vl_logic_vector(7 downto 0);
        txcreddatafccp  : out    vl_logic_vector(11 downto 0);
        txstdata        : in     vl_logic_vector(255 downto 0);
        txstparity      : in     vl_logic_vector(31 downto 0);
        txsterr         : in     vl_logic_vector(3 downto 0);
        txstsop         : in     vl_logic_vector(3 downto 0);
        txsteop         : in     vl_logic_vector(3 downto 0);
        txstempty       : in     vl_logic_vector(1 downto 0);
        txstvalid       : in     vl_logic_vector(0 downto 0);
        r2cuncecc       : out    vl_logic_vector(0 downto 0);
        rxcorrecc       : out    vl_logic_vector(0 downto 0);
        retryuncecc     : out    vl_logic_vector(0 downto 0);
        retrycorrecc    : out    vl_logic_vector(0 downto 0);
        rxparerr        : out    vl_logic_vector(0 downto 0);
        txparerr        : out    vl_logic_vector(1 downto 0);
        r2cparerr       : out    vl_logic_vector(0 downto 0);
        pmetosr         : out    vl_logic_vector(0 downto 0);
        pmetocr         : in     vl_logic_vector(0 downto 0);
        pmevent         : in     vl_logic_vector(0 downto 0);
        pmdata          : in     vl_logic_vector(9 downto 0);
        pmauxpwr        : in     vl_logic_vector(0 downto 0);
        tlcfgsts        : out    vl_logic_vector(52 downto 0);
        tlcfgctl        : out    vl_logic_vector(31 downto 0);
        tlcfgadd        : out    vl_logic_vector(3 downto 0);
        appintaack      : out    vl_logic_vector(0 downto 0);
        appintasts      : in     vl_logic_vector(0 downto 0);
        intstatus       : out    vl_logic_vector(3 downto 0);
        appmsiack       : out    vl_logic_vector(0 downto 0);
        appmsireq       : in     vl_logic_vector(0 downto 0);
        appmsitc        : in     vl_logic_vector(2 downto 0);
        appmsinum       : in     vl_logic_vector(4 downto 0);
        aermsinum       : in     vl_logic_vector(4 downto 0);
        pexmsinum       : in     vl_logic_vector(4 downto 0);
        hpgctrler       : in     vl_logic_vector(4 downto 0);
        cfglink2csrpld  : in     vl_logic_vector(12 downto 0);
        cfgprmbuspld    : in     vl_logic_vector(7 downto 0);
        csebisshadow    : out    vl_logic_vector(0 downto 0);
        csebwrdata      : out    vl_logic_vector(31 downto 0);
        csebwrdataparity: out    vl_logic_vector(3 downto 0);
        csebbe          : out    vl_logic_vector(3 downto 0);
        csebaddr        : out    vl_logic_vector(32 downto 0);
        csebaddrparity  : out    vl_logic_vector(4 downto 0);
        csebwren        : out    vl_logic_vector(0 downto 0);
        csebrden        : out    vl_logic_vector(0 downto 0);
        csebwrrespreq   : out    vl_logic_vector(0 downto 0);
        csebrddata      : in     vl_logic_vector(31 downto 0);
        csebrddataparity: in     vl_logic_vector(3 downto 0);
        csebwaitrequest : in     vl_logic_vector(0 downto 0);
        csebwrrespvalid : in     vl_logic_vector(0 downto 0);
        csebwrresponse  : in     vl_logic_vector(4 downto 0);
        csebrdresponse  : in     vl_logic_vector(4 downto 0);
        dlup            : out    vl_logic_vector(0 downto 0);
        testouthip      : out    vl_logic_vector(255 downto 0);
        testout1hip     : out    vl_logic_vector(63 downto 0);
        ev1us           : out    vl_logic_vector(0 downto 0);
        ev128ns         : out    vl_logic_vector(0 downto 0);
        wakeoen         : out    vl_logic_vector(0 downto 0);
        serrout         : out    vl_logic_vector(0 downto 0);
        ltssmstate      : out    vl_logic_vector(4 downto 0);
        laneact         : out    vl_logic_vector(3 downto 0);
        currentspeed    : out    vl_logic_vector(1 downto 0);
        slotclkcfg      : in     vl_logic_vector(0 downto 0);
        mode            : in     vl_logic_vector(1 downto 0);
        testinhip       : in     vl_logic_vector(31 downto 0);
        testin1hip      : in     vl_logic_vector(31 downto 0);
        cplpending      : in     vl_logic_vector(0 downto 0);
        cplerr          : in     vl_logic_vector(6 downto 0);
        appinterr       : in     vl_logic_vector(1 downto 0);
        egressblkerr    : in     vl_logic_vector(0 downto 0);
        pmexitd0ack     : in     vl_logic_vector(0 downto 0);
        pmexitd0req     : out    vl_logic_vector(0 downto 0);
        currentcoeff0   : out    vl_logic_vector(17 downto 0);
        currentcoeff1   : out    vl_logic_vector(17 downto 0);
        currentcoeff2   : out    vl_logic_vector(17 downto 0);
        currentcoeff3   : out    vl_logic_vector(17 downto 0);
        currentcoeff4   : out    vl_logic_vector(17 downto 0);
        currentcoeff5   : out    vl_logic_vector(17 downto 0);
        currentcoeff6   : out    vl_logic_vector(17 downto 0);
        currentcoeff7   : out    vl_logic_vector(17 downto 0);
        currentrxpreset0: out    vl_logic_vector(2 downto 0);
        currentrxpreset1: out    vl_logic_vector(2 downto 0);
        currentrxpreset2: out    vl_logic_vector(2 downto 0);
        currentrxpreset3: out    vl_logic_vector(2 downto 0);
        currentrxpreset4: out    vl_logic_vector(2 downto 0);
        currentrxpreset5: out    vl_logic_vector(2 downto 0);
        currentrxpreset6: out    vl_logic_vector(2 downto 0);
        currentrxpreset7: out    vl_logic_vector(2 downto 0);
        rate0           : out    vl_logic_vector(1 downto 0);
        rate1           : out    vl_logic_vector(1 downto 0);
        rate2           : out    vl_logic_vector(1 downto 0);
        rate3           : out    vl_logic_vector(1 downto 0);
        rate4           : out    vl_logic_vector(1 downto 0);
        rate5           : out    vl_logic_vector(1 downto 0);
        rate6           : out    vl_logic_vector(1 downto 0);
        rate7           : out    vl_logic_vector(1 downto 0);
        ratectrl        : out    vl_logic_vector(1 downto 0);
        ratetiedtognd   : out    vl_logic_vector(0 downto 0);
        eidleinfersel0  : out    vl_logic_vector(2 downto 0);
        eidleinfersel1  : out    vl_logic_vector(2 downto 0);
        eidleinfersel2  : out    vl_logic_vector(2 downto 0);
        eidleinfersel3  : out    vl_logic_vector(2 downto 0);
        eidleinfersel4  : out    vl_logic_vector(2 downto 0);
        eidleinfersel5  : out    vl_logic_vector(2 downto 0);
        eidleinfersel6  : out    vl_logic_vector(2 downto 0);
        eidleinfersel7  : out    vl_logic_vector(2 downto 0);
        txdata0         : out    vl_logic_vector(31 downto 0);
        txdatak0        : out    vl_logic_vector(3 downto 0);
        txdetectrx0     : out    vl_logic_vector(0 downto 0);
        txelecidle0     : out    vl_logic_vector(0 downto 0);
        txcompl0        : out    vl_logic_vector(0 downto 0);
        rxpolarity0     : out    vl_logic_vector(0 downto 0);
        powerdown0      : out    vl_logic_vector(1 downto 0);
        txdataskip0     : out    vl_logic_vector(0 downto 0);
        txblkst0        : out    vl_logic_vector(0 downto 0);
        txsynchd0       : out    vl_logic_vector(1 downto 0);
        txdeemph0       : out    vl_logic_vector(0 downto 0);
        txswing0        : out    vl_logic_vector(0 downto 0);
        txmargin0       : out    vl_logic_vector(2 downto 0);
        rxdata0         : in     vl_logic_vector(31 downto 0);
        rxdatak0        : in     vl_logic_vector(3 downto 0);
        rxvalid0        : in     vl_logic_vector(0 downto 0);
        phystatus0      : in     vl_logic_vector(0 downto 0);
        rxelecidle0     : in     vl_logic_vector(0 downto 0);
        rxstatus0       : in     vl_logic_vector(2 downto 0);
        rxdataskip0     : in     vl_logic_vector(0 downto 0);
        rxblkst0        : in     vl_logic_vector(0 downto 0);
        rxsynchd0       : in     vl_logic_vector(1 downto 0);
        rxfreqlocked0   : in     vl_logic_vector(0 downto 0);
        txdata1         : out    vl_logic_vector(31 downto 0);
        txdatak1        : out    vl_logic_vector(3 downto 0);
        txdetectrx1     : out    vl_logic_vector(0 downto 0);
        txelecidle1     : out    vl_logic_vector(0 downto 0);
        txcompl1        : out    vl_logic_vector(0 downto 0);
        rxpolarity1     : out    vl_logic_vector(0 downto 0);
        powerdown1      : out    vl_logic_vector(1 downto 0);
        txdataskip1     : out    vl_logic_vector(0 downto 0);
        txblkst1        : out    vl_logic_vector(0 downto 0);
        txsynchd1       : out    vl_logic_vector(1 downto 0);
        txdeemph1       : out    vl_logic_vector(0 downto 0);
        txswing1        : out    vl_logic_vector(0 downto 0);
        txmargin1       : out    vl_logic_vector(2 downto 0);
        rxdata1         : in     vl_logic_vector(31 downto 0);
        rxdatak1        : in     vl_logic_vector(3 downto 0);
        rxvalid1        : in     vl_logic_vector(0 downto 0);
        phystatus1      : in     vl_logic_vector(0 downto 0);
        rxelecidle1     : in     vl_logic_vector(0 downto 0);
        rxstatus1       : in     vl_logic_vector(2 downto 0);
        rxdataskip1     : in     vl_logic_vector(0 downto 0);
        rxblkst1        : in     vl_logic_vector(0 downto 0);
        rxsynchd1       : in     vl_logic_vector(1 downto 0);
        rxfreqlocked1   : in     vl_logic_vector(0 downto 0);
        txdata2         : out    vl_logic_vector(31 downto 0);
        txdatak2        : out    vl_logic_vector(3 downto 0);
        txdetectrx2     : out    vl_logic_vector(0 downto 0);
        txelecidle2     : out    vl_logic_vector(0 downto 0);
        txcompl2        : out    vl_logic_vector(0 downto 0);
        rxpolarity2     : out    vl_logic_vector(0 downto 0);
        powerdown2      : out    vl_logic_vector(1 downto 0);
        txdataskip2     : out    vl_logic_vector(0 downto 0);
        txblkst2        : out    vl_logic_vector(0 downto 0);
        txsynchd2       : out    vl_logic_vector(1 downto 0);
        txdeemph2       : out    vl_logic_vector(0 downto 0);
        txswing2        : out    vl_logic_vector(0 downto 0);
        txmargin2       : out    vl_logic_vector(2 downto 0);
        rxdata2         : in     vl_logic_vector(31 downto 0);
        rxdatak2        : in     vl_logic_vector(3 downto 0);
        rxvalid2        : in     vl_logic_vector(0 downto 0);
        phystatus2      : in     vl_logic_vector(0 downto 0);
        rxelecidle2     : in     vl_logic_vector(0 downto 0);
        rxstatus2       : in     vl_logic_vector(2 downto 0);
        rxdataskip2     : in     vl_logic_vector(0 downto 0);
        rxblkst2        : in     vl_logic_vector(0 downto 0);
        rxsynchd2       : in     vl_logic_vector(1 downto 0);
        rxfreqlocked2   : in     vl_logic_vector(0 downto 0);
        txdata3         : out    vl_logic_vector(31 downto 0);
        txdatak3        : out    vl_logic_vector(3 downto 0);
        txdetectrx3     : out    vl_logic_vector(0 downto 0);
        txelecidle3     : out    vl_logic_vector(0 downto 0);
        txcompl3        : out    vl_logic_vector(0 downto 0);
        rxpolarity3     : out    vl_logic_vector(0 downto 0);
        powerdown3      : out    vl_logic_vector(1 downto 0);
        txdataskip3     : out    vl_logic_vector(0 downto 0);
        txblkst3        : out    vl_logic_vector(0 downto 0);
        txsynchd3       : out    vl_logic_vector(1 downto 0);
        txdeemph3       : out    vl_logic_vector(0 downto 0);
        txswing3        : out    vl_logic_vector(0 downto 0);
        txmargin3       : out    vl_logic_vector(2 downto 0);
        rxdata3         : in     vl_logic_vector(31 downto 0);
        rxdatak3        : in     vl_logic_vector(3 downto 0);
        rxvalid3        : in     vl_logic_vector(0 downto 0);
        phystatus3      : in     vl_logic_vector(0 downto 0);
        rxelecidle3     : in     vl_logic_vector(0 downto 0);
        rxstatus3       : in     vl_logic_vector(2 downto 0);
        rxdataskip3     : in     vl_logic_vector(0 downto 0);
        rxblkst3        : in     vl_logic_vector(0 downto 0);
        rxsynchd3       : in     vl_logic_vector(1 downto 0);
        rxfreqlocked3   : in     vl_logic_vector(0 downto 0);
        txdata4         : out    vl_logic_vector(31 downto 0);
        txdatak4        : out    vl_logic_vector(3 downto 0);
        txdetectrx4     : out    vl_logic_vector(0 downto 0);
        txelecidle4     : out    vl_logic_vector(0 downto 0);
        txcompl4        : out    vl_logic_vector(0 downto 0);
        rxpolarity4     : out    vl_logic_vector(0 downto 0);
        powerdown4      : out    vl_logic_vector(1 downto 0);
        txdataskip4     : out    vl_logic_vector(0 downto 0);
        txblkst4        : out    vl_logic_vector(0 downto 0);
        txsynchd4       : out    vl_logic_vector(1 downto 0);
        txdeemph4       : out    vl_logic_vector(0 downto 0);
        txswing4        : out    vl_logic_vector(0 downto 0);
        txmargin4       : out    vl_logic_vector(2 downto 0);
        rxdata4         : in     vl_logic_vector(31 downto 0);
        rxdatak4        : in     vl_logic_vector(3 downto 0);
        rxvalid4        : in     vl_logic_vector(0 downto 0);
        phystatus4      : in     vl_logic_vector(0 downto 0);
        rxelecidle4     : in     vl_logic_vector(0 downto 0);
        rxstatus4       : in     vl_logic_vector(2 downto 0);
        rxdataskip4     : in     vl_logic_vector(0 downto 0);
        rxblkst4        : in     vl_logic_vector(0 downto 0);
        rxsynchd4       : in     vl_logic_vector(1 downto 0);
        rxfreqlocked4   : in     vl_logic_vector(0 downto 0);
        txdata5         : out    vl_logic_vector(31 downto 0);
        txdatak5        : out    vl_logic_vector(3 downto 0);
        txdetectrx5     : out    vl_logic_vector(0 downto 0);
        txelecidle5     : out    vl_logic_vector(0 downto 0);
        txcompl5        : out    vl_logic_vector(0 downto 0);
        rxpolarity5     : out    vl_logic_vector(0 downto 0);
        powerdown5      : out    vl_logic_vector(1 downto 0);
        txdataskip5     : out    vl_logic_vector(0 downto 0);
        txblkst5        : out    vl_logic_vector(0 downto 0);
        txsynchd5       : out    vl_logic_vector(1 downto 0);
        txdeemph5       : out    vl_logic_vector(0 downto 0);
        txswing5        : out    vl_logic_vector(0 downto 0);
        txmargin5       : out    vl_logic_vector(2 downto 0);
        rxdata5         : in     vl_logic_vector(31 downto 0);
        rxdatak5        : in     vl_logic_vector(3 downto 0);
        rxvalid5        : in     vl_logic_vector(0 downto 0);
        phystatus5      : in     vl_logic_vector(0 downto 0);
        rxelecidle5     : in     vl_logic_vector(0 downto 0);
        rxstatus5       : in     vl_logic_vector(2 downto 0);
        rxdataskip5     : in     vl_logic_vector(0 downto 0);
        rxblkst5        : in     vl_logic_vector(0 downto 0);
        rxsynchd5       : in     vl_logic_vector(1 downto 0);
        rxfreqlocked5   : in     vl_logic_vector(0 downto 0);
        txdata6         : out    vl_logic_vector(31 downto 0);
        txdatak6        : out    vl_logic_vector(3 downto 0);
        txdetectrx6     : out    vl_logic_vector(0 downto 0);
        txelecidle6     : out    vl_logic_vector(0 downto 0);
        txcompl6        : out    vl_logic_vector(0 downto 0);
        rxpolarity6     : out    vl_logic_vector(0 downto 0);
        powerdown6      : out    vl_logic_vector(1 downto 0);
        txdataskip6     : out    vl_logic_vector(0 downto 0);
        txblkst6        : out    vl_logic_vector(0 downto 0);
        txsynchd6       : out    vl_logic_vector(1 downto 0);
        txdeemph6       : out    vl_logic_vector(0 downto 0);
        txswing6        : out    vl_logic_vector(0 downto 0);
        txmargin6       : out    vl_logic_vector(2 downto 0);
        rxdata6         : in     vl_logic_vector(31 downto 0);
        rxdatak6        : in     vl_logic_vector(3 downto 0);
        rxvalid6        : in     vl_logic_vector(0 downto 0);
        phystatus6      : in     vl_logic_vector(0 downto 0);
        rxelecidle6     : in     vl_logic_vector(0 downto 0);
        rxstatus6       : in     vl_logic_vector(2 downto 0);
        rxdataskip6     : in     vl_logic_vector(0 downto 0);
        rxblkst6        : in     vl_logic_vector(0 downto 0);
        rxsynchd6       : in     vl_logic_vector(1 downto 0);
        rxfreqlocked6   : in     vl_logic_vector(0 downto 0);
        txdata7         : out    vl_logic_vector(31 downto 0);
        txdatak7        : out    vl_logic_vector(3 downto 0);
        txdetectrx7     : out    vl_logic_vector(0 downto 0);
        txelecidle7     : out    vl_logic_vector(0 downto 0);
        txcompl7        : out    vl_logic_vector(0 downto 0);
        rxpolarity7     : out    vl_logic_vector(0 downto 0);
        powerdown7      : out    vl_logic_vector(1 downto 0);
        txdataskip7     : out    vl_logic_vector(0 downto 0);
        txblkst7        : out    vl_logic_vector(0 downto 0);
        txsynchd7       : out    vl_logic_vector(1 downto 0);
        txdeemph7       : out    vl_logic_vector(0 downto 0);
        txswing7        : out    vl_logic_vector(0 downto 0);
        txmargin7       : out    vl_logic_vector(2 downto 0);
        rxdata7         : in     vl_logic_vector(31 downto 0);
        rxdatak7        : in     vl_logic_vector(3 downto 0);
        rxvalid7        : in     vl_logic_vector(0 downto 0);
        phystatus7      : in     vl_logic_vector(0 downto 0);
        rxelecidle7     : in     vl_logic_vector(0 downto 0);
        rxstatus7       : in     vl_logic_vector(2 downto 0);
        rxdataskip7     : in     vl_logic_vector(0 downto 0);
        rxblkst7        : in     vl_logic_vector(0 downto 0);
        rxsynchd7       : in     vl_logic_vector(1 downto 0);
        rxfreqlocked7   : in     vl_logic_vector(0 downto 0);
        dbgpipex1rx     : in     vl_logic_vector(43 downto 0);
        memredsclk      : in     vl_logic_vector(0 downto 0);
        memredenscan    : in     vl_logic_vector(0 downto 0);
        memredscen      : in     vl_logic_vector(0 downto 0);
        memredscin      : in     vl_logic_vector(0 downto 0);
        memredscsel     : in     vl_logic_vector(0 downto 0);
        memredscrst     : in     vl_logic_vector(0 downto 0);
        memredscout     : out    vl_logic_vector(0 downto 0);
        memregscanen    : in     vl_logic_vector(0 downto 0);
        memregscanin    : in     vl_logic_vector(0 downto 0);
        memhiptestenable: in     vl_logic_vector(0 downto 0);
        memregscanout   : out    vl_logic_vector(0 downto 0);
        bisttesten      : in     vl_logic_vector(0 downto 0);
        bistenrpl       : in     vl_logic_vector(0 downto 0);
        bistscanin      : in     vl_logic_vector(0 downto 0);
        bistscanen      : in     vl_logic_vector(0 downto 0);
        bistenrcv       : in     vl_logic_vector(0 downto 0);
        bistscanoutrpl  : out    vl_logic_vector(0 downto 0);
        bistdonearpl    : out    vl_logic_vector(0 downto 0);
        bistdonebrpl    : out    vl_logic_vector(0 downto 0);
        bistpassrpl     : out    vl_logic_vector(0 downto 0);
        derrrpl         : out    vl_logic_vector(0 downto 0);
        derrcorextrpl   : out    vl_logic_vector(0 downto 0);
        bistscanoutrcv  : out    vl_logic_vector(0 downto 0);
        bistdonearcv    : out    vl_logic_vector(0 downto 0);
        bistdonebrcv    : out    vl_logic_vector(0 downto 0);
        bistpassrcv     : out    vl_logic_vector(0 downto 0);
        derrcorextrcv   : out    vl_logic_vector(0 downto 0);
        bistscanoutrcv1 : out    vl_logic_vector(0 downto 0);
        bistdonearcv1   : out    vl_logic_vector(0 downto 0);
        bistdonebrcv1   : out    vl_logic_vector(0 downto 0);
        bistpassrcv1    : out    vl_logic_vector(0 downto 0);
        derrcorextrcv1  : out    vl_logic_vector(0 downto 0);
        scanmoden       : in     vl_logic_vector(0 downto 0);
        scanshiftn      : in     vl_logic_vector(0 downto 0);
        nfrzdrv         : in     vl_logic_vector(0 downto 0);
        frzreg          : in     vl_logic_vector(0 downto 0);
        frzlogic        : in     vl_logic_vector(0 downto 0);
        idrpl           : in     vl_logic_vector(7 downto 0);
        idrcv           : in     vl_logic_vector(7 downto 0);
        plniotri        : in     vl_logic_vector(0 downto 0);
        entest          : in     vl_logic_vector(0 downto 0);
        usermode        : in     vl_logic_vector(0 downto 0);
        cvpclk          : out    vl_logic_vector(0 downto 0);
        cvpdata         : out    vl_logic_vector(31 downto 0);
        cvpstartxfer    : out    vl_logic_vector(0 downto 0);
        cvpconfig       : out    vl_logic_vector(0 downto 0);
        cvpfullconfig   : out    vl_logic_vector(0 downto 0);
        cvpconfigready  : in     vl_logic_vector(0 downto 0);
        cvpen           : in     vl_logic_vector(0 downto 0);
        cvpconfigerror  : in     vl_logic_vector(0 downto 0);
        cvpconfigdone   : in     vl_logic_vector(0 downto 0);
        pinperstn       : in     vl_logic_vector(0 downto 0);
        pldperstn       : in     vl_logic_vector(0 downto 0);
        iocsrrdydly     : in     vl_logic_vector(0 downto 0);
        softaltpe3rstn  : in     vl_logic_vector(0 downto 0);
        softaltpe3srstn : in     vl_logic_vector(0 downto 0);
        softaltpe3crstn : in     vl_logic_vector(0 downto 0);
        pldclrpmapcshipn: in     vl_logic_vector(0 downto 0);
        pldclrpcshipn   : in     vl_logic_vector(0 downto 0);
        pldclrhipn      : in     vl_logic_vector(0 downto 0);
        s0ch0emsiptieoff: out    vl_logic_vector(100 downto 0);
        s0ch1emsiptieoff: out    vl_logic_vector(100 downto 0);
        s0ch2emsiptieoff: out    vl_logic_vector(100 downto 0);
        s1ch0emsiptieoff: out    vl_logic_vector(100 downto 0);
        s1ch1emsiptieoff: out    vl_logic_vector(188 downto 0);
        s1ch2emsiptieoff: out    vl_logic_vector(100 downto 0);
        s2ch0emsiptieoff: out    vl_logic_vector(100 downto 0);
        s2ch1emsiptieoff: out    vl_logic_vector(100 downto 0);
        s2ch2emsiptieoff: out    vl_logic_vector(100 downto 0);
        s3ch0emsiptieoff: out    vl_logic_vector(188 downto 0);
        s3ch1emsiptieoff: out    vl_logic_vector(188 downto 0);
        s3ch2emsiptieoff: out    vl_logic_vector(188 downto 0);
        emsiptieofftop  : out    vl_logic_vector(299 downto 0);
        emsiptieoffbot  : out    vl_logic_vector(299 downto 0);
        txpcsrstn0      : out    vl_logic_vector(0 downto 0);
        rxpcsrstn0      : out    vl_logic_vector(0 downto 0);
        g3txpcsrstn0    : out    vl_logic_vector(0 downto 0);
        g3rxpcsrstn0    : out    vl_logic_vector(0 downto 0);
        txpmasyncp0     : out    vl_logic_vector(0 downto 0);
        rxpmarstb0      : out    vl_logic_vector(0 downto 0);
        txlcpllrstb0    : out    vl_logic_vector(0 downto 0);
        offcalen0       : out    vl_logic_vector(0 downto 0);
        frefclk0        : in     vl_logic_vector(0 downto 0);
        offcaldone0     : in     vl_logic_vector(0 downto 0);
        txlcplllock0    : in     vl_logic_vector(0 downto 0);
        rxfreqtxcmuplllock0: in     vl_logic_vector(0 downto 0);
        rxpllphaselock0 : in     vl_logic_vector(0 downto 0);
        masktxplllock0  : in     vl_logic_vector(0 downto 0);
        txpcsrstn1      : out    vl_logic_vector(0 downto 0);
        rxpcsrstn1      : out    vl_logic_vector(0 downto 0);
        g3txpcsrstn1    : out    vl_logic_vector(0 downto 0);
        g3rxpcsrstn1    : out    vl_logic_vector(0 downto 0);
        txpmasyncp1     : out    vl_logic_vector(0 downto 0);
        rxpmarstb1      : out    vl_logic_vector(0 downto 0);
        txlcpllrstb1    : out    vl_logic_vector(0 downto 0);
        offcalen1       : out    vl_logic_vector(0 downto 0);
        frefclk1        : in     vl_logic_vector(0 downto 0);
        offcaldone1     : in     vl_logic_vector(0 downto 0);
        txlcplllock1    : in     vl_logic_vector(0 downto 0);
        rxfreqtxcmuplllock1: in     vl_logic_vector(0 downto 0);
        rxpllphaselock1 : in     vl_logic_vector(0 downto 0);
        masktxplllock1  : in     vl_logic_vector(0 downto 0);
        txpcsrstn2      : out    vl_logic_vector(0 downto 0);
        rxpcsrstn2      : out    vl_logic_vector(0 downto 0);
        g3txpcsrstn2    : out    vl_logic_vector(0 downto 0);
        g3rxpcsrstn2    : out    vl_logic_vector(0 downto 0);
        txpmasyncp2     : out    vl_logic_vector(0 downto 0);
        rxpmarstb2      : out    vl_logic_vector(0 downto 0);
        txlcpllrstb2    : out    vl_logic_vector(0 downto 0);
        offcalen2       : out    vl_logic_vector(0 downto 0);
        frefclk2        : in     vl_logic_vector(0 downto 0);
        offcaldone2     : in     vl_logic_vector(0 downto 0);
        txlcplllock2    : in     vl_logic_vector(0 downto 0);
        rxfreqtxcmuplllock2: in     vl_logic_vector(0 downto 0);
        rxpllphaselock2 : in     vl_logic_vector(0 downto 0);
        masktxplllock2  : in     vl_logic_vector(0 downto 0);
        txpcsrstn3      : out    vl_logic_vector(0 downto 0);
        rxpcsrstn3      : out    vl_logic_vector(0 downto 0);
        g3txpcsrstn3    : out    vl_logic_vector(0 downto 0);
        g3rxpcsrstn3    : out    vl_logic_vector(0 downto 0);
        txpmasyncp3     : out    vl_logic_vector(0 downto 0);
        rxpmarstb3      : out    vl_logic_vector(0 downto 0);
        txlcpllrstb3    : out    vl_logic_vector(0 downto 0);
        offcalen3       : out    vl_logic_vector(0 downto 0);
        frefclk3        : in     vl_logic_vector(0 downto 0);
        offcaldone3     : in     vl_logic_vector(0 downto 0);
        txlcplllock3    : in     vl_logic_vector(0 downto 0);
        rxfreqtxcmuplllock3: in     vl_logic_vector(0 downto 0);
        rxpllphaselock3 : in     vl_logic_vector(0 downto 0);
        masktxplllock3  : in     vl_logic_vector(0 downto 0);
        txpcsrstn4      : out    vl_logic_vector(0 downto 0);
        rxpcsrstn4      : out    vl_logic_vector(0 downto 0);
        g3txpcsrstn4    : out    vl_logic_vector(0 downto 0);
        g3rxpcsrstn4    : out    vl_logic_vector(0 downto 0);
        txpmasyncp4     : out    vl_logic_vector(0 downto 0);
        rxpmarstb4      : out    vl_logic_vector(0 downto 0);
        txlcpllrstb4    : out    vl_logic_vector(0 downto 0);
        offcalen4       : out    vl_logic_vector(0 downto 0);
        frefclk4        : in     vl_logic_vector(0 downto 0);
        offcaldone4     : in     vl_logic_vector(0 downto 0);
        txlcplllock4    : in     vl_logic_vector(0 downto 0);
        rxfreqtxcmuplllock4: in     vl_logic_vector(0 downto 0);
        rxpllphaselock4 : in     vl_logic_vector(0 downto 0);
        masktxplllock4  : in     vl_logic_vector(0 downto 0);
        txpcsrstn5      : out    vl_logic_vector(0 downto 0);
        rxpcsrstn5      : out    vl_logic_vector(0 downto 0);
        g3txpcsrstn5    : out    vl_logic_vector(0 downto 0);
        g3rxpcsrstn5    : out    vl_logic_vector(0 downto 0);
        txpmasyncp5     : out    vl_logic_vector(0 downto 0);
        rxpmarstb5      : out    vl_logic_vector(0 downto 0);
        txlcpllrstb5    : out    vl_logic_vector(0 downto 0);
        offcalen5       : out    vl_logic_vector(0 downto 0);
        frefclk5        : in     vl_logic_vector(0 downto 0);
        offcaldone5     : in     vl_logic_vector(0 downto 0);
        txlcplllock5    : in     vl_logic_vector(0 downto 0);
        rxfreqtxcmuplllock5: in     vl_logic_vector(0 downto 0);
        rxpllphaselock5 : in     vl_logic_vector(0 downto 0);
        masktxplllock5  : in     vl_logic_vector(0 downto 0);
        txpcsrstn6      : out    vl_logic_vector(0 downto 0);
        rxpcsrstn6      : out    vl_logic_vector(0 downto 0);
        g3txpcsrstn6    : out    vl_logic_vector(0 downto 0);
        g3rxpcsrstn6    : out    vl_logic_vector(0 downto 0);
        txpmasyncp6     : out    vl_logic_vector(0 downto 0);
        rxpmarstb6      : out    vl_logic_vector(0 downto 0);
        txlcpllrstb6    : out    vl_logic_vector(0 downto 0);
        offcalen6       : out    vl_logic_vector(0 downto 0);
        frefclk6        : in     vl_logic_vector(0 downto 0);
        offcaldone6     : in     vl_logic_vector(0 downto 0);
        txlcplllock6    : in     vl_logic_vector(0 downto 0);
        rxfreqtxcmuplllock6: in     vl_logic_vector(0 downto 0);
        rxpllphaselock6 : in     vl_logic_vector(0 downto 0);
        masktxplllock6  : in     vl_logic_vector(0 downto 0);
        txpcsrstn7      : out    vl_logic_vector(0 downto 0);
        rxpcsrstn7      : out    vl_logic_vector(0 downto 0);
        g3txpcsrstn7    : out    vl_logic_vector(0 downto 0);
        g3rxpcsrstn7    : out    vl_logic_vector(0 downto 0);
        txpmasyncp7     : out    vl_logic_vector(0 downto 0);
        rxpmarstb7      : out    vl_logic_vector(0 downto 0);
        txlcpllrstb7    : out    vl_logic_vector(0 downto 0);
        offcalen7       : out    vl_logic_vector(0 downto 0);
        frefclk7        : in     vl_logic_vector(0 downto 0);
        offcaldone7     : in     vl_logic_vector(0 downto 0);
        txlcplllock7    : in     vl_logic_vector(0 downto 0);
        rxfreqtxcmuplllock7: in     vl_logic_vector(0 downto 0);
        rxpllphaselock7 : in     vl_logic_vector(0 downto 0);
        masktxplllock7  : in     vl_logic_vector(0 downto 0);
        txpcsrstn8      : out    vl_logic_vector(0 downto 0);
        rxpcsrstn8      : out    vl_logic_vector(0 downto 0);
        g3txpcsrstn8    : out    vl_logic_vector(0 downto 0);
        g3rxpcsrstn8    : out    vl_logic_vector(0 downto 0);
        txpmasyncp8     : out    vl_logic_vector(0 downto 0);
        rxpmarstb8      : out    vl_logic_vector(0 downto 0);
        txlcpllrstb8    : out    vl_logic_vector(0 downto 0);
        offcalen8       : out    vl_logic_vector(0 downto 0);
        frefclk8        : in     vl_logic_vector(0 downto 0);
        offcaldone8     : in     vl_logic_vector(0 downto 0);
        txlcplllock8    : in     vl_logic_vector(0 downto 0);
        rxfreqtxcmuplllock8: in     vl_logic_vector(0 downto 0);
        rxpllphaselock8 : in     vl_logic_vector(0 downto 0);
        masktxplllock8  : in     vl_logic_vector(0 downto 0);
        txpcsrstn9      : out    vl_logic_vector(0 downto 0);
        rxpcsrstn9      : out    vl_logic_vector(0 downto 0);
        g3txpcsrstn9    : out    vl_logic_vector(0 downto 0);
        g3rxpcsrstn9    : out    vl_logic_vector(0 downto 0);
        txpmasyncp9     : out    vl_logic_vector(0 downto 0);
        rxpmarstb9      : out    vl_logic_vector(0 downto 0);
        txlcpllrstb9    : out    vl_logic_vector(0 downto 0);
        offcalen9       : out    vl_logic_vector(0 downto 0);
        frefclk9        : in     vl_logic_vector(0 downto 0);
        offcaldone9     : in     vl_logic_vector(0 downto 0);
        txlcplllock9    : in     vl_logic_vector(0 downto 0);
        rxfreqtxcmuplllock9: in     vl_logic_vector(0 downto 0);
        rxpllphaselock9 : in     vl_logic_vector(0 downto 0);
        masktxplllock9  : in     vl_logic_vector(0 downto 0);
        txpcsrstn10     : out    vl_logic_vector(0 downto 0);
        rxpcsrstn10     : out    vl_logic_vector(0 downto 0);
        g3txpcsrstn10   : out    vl_logic_vector(0 downto 0);
        g3rxpcsrstn10   : out    vl_logic_vector(0 downto 0);
        txpmasyncp10    : out    vl_logic_vector(0 downto 0);
        rxpmarstb10     : out    vl_logic_vector(0 downto 0);
        txlcpllrstb10   : out    vl_logic_vector(0 downto 0);
        offcalen10      : out    vl_logic_vector(0 downto 0);
        frefclk10       : in     vl_logic_vector(0 downto 0);
        offcaldone10    : in     vl_logic_vector(0 downto 0);
        txlcplllock10   : in     vl_logic_vector(0 downto 0);
        rxfreqtxcmuplllock10: in     vl_logic_vector(0 downto 0);
        rxpllphaselock10: in     vl_logic_vector(0 downto 0);
        masktxplllock10 : in     vl_logic_vector(0 downto 0);
        txpcsrstn11     : out    vl_logic_vector(0 downto 0);
        rxpcsrstn11     : out    vl_logic_vector(0 downto 0);
        g3txpcsrstn11   : out    vl_logic_vector(0 downto 0);
        g3rxpcsrstn11   : out    vl_logic_vector(0 downto 0);
        txpmasyncp11    : out    vl_logic_vector(0 downto 0);
        rxpmarstb11     : out    vl_logic_vector(0 downto 0);
        txlcpllrstb11   : out    vl_logic_vector(0 downto 0);
        offcalen11      : out    vl_logic_vector(0 downto 0);
        frefclk11       : in     vl_logic_vector(0 downto 0);
        offcaldone11    : in     vl_logic_vector(0 downto 0);
        txlcplllock11   : in     vl_logic_vector(0 downto 0);
        rxfreqtxcmuplllock11: in     vl_logic_vector(0 downto 0);
        rxpllphaselock11: in     vl_logic_vector(0 downto 0);
        masktxplllock11 : in     vl_logic_vector(0 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmaddress     : in     vl_logic_vector(9 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        sershiftload    : in     vl_logic_vector(0 downto 0);
        interfacesel    : in     vl_logic_vector(0 downto 0);
        holdltssmrec    : in     vl_logic_vector(0 downto 0);
        forcetxeidle    : in     vl_logic_vector(0 downto 0);
        reservedin      : in     vl_logic_vector(31 downto 0);
        reservedclkin   : in     vl_logic_vector(0 downto 0);
        reservedout     : out    vl_logic_vector(31 downto 0);
        reservedclkout  : out    vl_logic_vector(0 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of func_mode : constant is 1;
    attribute mti_svvh_generic_type of in_cvp_mode : constant is 1;
    attribute mti_svvh_generic_type of bonding_mode : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of pcie_spec_1p0_compliance : constant is 1;
    attribute mti_svvh_generic_type of vc_enable : constant is 1;
    attribute mti_svvh_generic_type of enable_slot_register : constant is 1;
    attribute mti_svvh_generic_type of pcie_mode : constant is 1;
    attribute mti_svvh_generic_type of bypass_cdc : constant is 1;
    attribute mti_svvh_generic_type of enable_rx_reordering : constant is 1;
    attribute mti_svvh_generic_type of enable_rx_buffer_checking : constant is 1;
    attribute mti_svvh_generic_type of single_rx_detect_data : constant is 1;
    attribute mti_svvh_generic_type of single_rx_detect : constant is 1;
    attribute mti_svvh_generic_type of use_crc_forwarding : constant is 1;
    attribute mti_svvh_generic_type of bypass_tl : constant is 1;
    attribute mti_svvh_generic_type of gen123_lane_rate_mode : constant is 1;
    attribute mti_svvh_generic_type of lane_mask : constant is 1;
    attribute mti_svvh_generic_type of disable_link_x2_support : constant is 1;
    attribute mti_svvh_generic_type of national_inst_thru_enhance : constant is 1;
    attribute mti_svvh_generic_type of hip_hard_reset : constant is 1;
    attribute mti_svvh_generic_type of dis_paritychk : constant is 1;
    attribute mti_svvh_generic_type of wrong_device_id : constant is 1;
    attribute mti_svvh_generic_type of data_pack_rx : constant is 1;
    attribute mti_svvh_generic_type of ast_width : constant is 1;
    attribute mti_svvh_generic_type of ast_width_tx : constant is 1;
    attribute mti_svvh_generic_type of ast_width_rx : constant is 1;
    attribute mti_svvh_generic_type of tx_sop_ctrl : constant is 1;
    attribute mti_svvh_generic_type of rx_sop_ctrl : constant is 1;
    attribute mti_svvh_generic_type of rx_ast_parity : constant is 1;
    attribute mti_svvh_generic_type of tx_ast_parity : constant is 1;
    attribute mti_svvh_generic_type of ltssm_1ms_timeout : constant is 1;
    attribute mti_svvh_generic_type of ltssm_freqlocked_check : constant is 1;
    attribute mti_svvh_generic_type of deskew_comma : constant is 1;
    attribute mti_svvh_generic_type of dl_tx_check_parity_edb : constant is 1;
    attribute mti_svvh_generic_type of tl_tx_check_parity_msg : constant is 1;
    attribute mti_svvh_generic_type of port_link_number_data : constant is 1;
    attribute mti_svvh_generic_type of port_link_number : constant is 1;
    attribute mti_svvh_generic_type of device_number_data : constant is 1;
    attribute mti_svvh_generic_type of device_number : constant is 1;
    attribute mti_svvh_generic_type of bypass_clk_switch : constant is 1;
    attribute mti_svvh_generic_type of core_clk_out_sel : constant is 1;
    attribute mti_svvh_generic_type of core_clk_divider : constant is 1;
    attribute mti_svvh_generic_type of core_clk_source : constant is 1;
    attribute mti_svvh_generic_type of core_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of enable_ch0_pclk_out : constant is 1;
    attribute mti_svvh_generic_type of enable_ch01_pclk_out : constant is 1;
    attribute mti_svvh_generic_type of pipex1_debug_sel : constant is 1;
    attribute mti_svvh_generic_type of pclk_out_sel : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_data : constant is 1;
    attribute mti_svvh_generic_type of vendor_id : constant is 1;
    attribute mti_svvh_generic_type of device_id_data : constant is 1;
    attribute mti_svvh_generic_type of device_id : constant is 1;
    attribute mti_svvh_generic_type of revision_id_data : constant is 1;
    attribute mti_svvh_generic_type of revision_id : constant is 1;
    attribute mti_svvh_generic_type of class_code_data : constant is 1;
    attribute mti_svvh_generic_type of class_code : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_data : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_data : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id : constant is 1;
    attribute mti_svvh_generic_type of no_soft_reset : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_data : constant is 1;
    attribute mti_svvh_generic_type of maximum_current : constant is 1;
    attribute mti_svvh_generic_type of d1_support : constant is 1;
    attribute mti_svvh_generic_type of d2_support : constant is 1;
    attribute mti_svvh_generic_type of d0_pme : constant is 1;
    attribute mti_svvh_generic_type of d1_pme : constant is 1;
    attribute mti_svvh_generic_type of d2_pme : constant is 1;
    attribute mti_svvh_generic_type of d3_hot_pme : constant is 1;
    attribute mti_svvh_generic_type of d3_cold_pme : constant is 1;
    attribute mti_svvh_generic_type of use_aer : constant is 1;
    attribute mti_svvh_generic_type of low_priority_vc : constant is 1;
    attribute mti_svvh_generic_type of vc_arbitration : constant is 1;
    attribute mti_svvh_generic_type of disable_snoop_packet : constant is 1;
    attribute mti_svvh_generic_type of max_payload_size : constant is 1;
    attribute mti_svvh_generic_type of surprise_down_error_support : constant is 1;
    attribute mti_svvh_generic_type of dll_active_report_support : constant is 1;
    attribute mti_svvh_generic_type of extend_tag_field : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_data : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_data : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency : constant is 1;
    attribute mti_svvh_generic_type of indicator_data : constant is 1;
    attribute mti_svvh_generic_type of indicator : constant is 1;
    attribute mti_svvh_generic_type of role_based_error_reporting : constant is 1;
    attribute mti_svvh_generic_type of gen3_ltssm_debug : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_data : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale : constant is 1;
    attribute mti_svvh_generic_type of max_link_width : constant is 1;
    attribute mti_svvh_generic_type of enable_l1_aspm : constant is 1;
    attribute mti_svvh_generic_type of enable_l0s_aspm : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_data : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_data : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_data : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_data : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit : constant is 1;
    attribute mti_svvh_generic_type of slot_number_data : constant is 1;
    attribute mti_svvh_generic_type of slot_number : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_data : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_data : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of completion_timeout : constant is 1;
    attribute mti_svvh_generic_type of enable_completion_timeout_disable : constant is 1;
    attribute mti_svvh_generic_type of extended_tag_reset : constant is 1;
    attribute mti_svvh_generic_type of ecrc_check_capable : constant is 1;
    attribute mti_svvh_generic_type of ecrc_gen_capable : constant is 1;
    attribute mti_svvh_generic_type of no_command_completed : constant is 1;
    attribute mti_svvh_generic_type of msi_multi_message_capable : constant is 1;
    attribute mti_svvh_generic_type of msi_64bit_addressing_capable : constant is 1;
    attribute mti_svvh_generic_type of msi_masking_capable : constant is 1;
    attribute mti_svvh_generic_type of msi_support : constant is 1;
    attribute mti_svvh_generic_type of interrupt_pin : constant is 1;
    attribute mti_svvh_generic_type of ena_ido_req : constant is 1;
    attribute mti_svvh_generic_type of ena_ido_cpl : constant is 1;
    attribute mti_svvh_generic_type of enable_function_msix_support : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_data : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_data : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_data : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_data : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_data : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_vga_enable : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_ssid_support : constant is 1;
    attribute mti_svvh_generic_type of ssvid_data : constant is 1;
    attribute mti_svvh_generic_type of ssvid : constant is 1;
    attribute mti_svvh_generic_type of ssid_data : constant is 1;
    attribute mti_svvh_generic_type of ssid : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_data : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_data : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_data : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of deemphasis_enable : constant is 1;
    attribute mti_svvh_generic_type of pcie_spec_version : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_data : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_data : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock : constant is 1;
    attribute mti_svvh_generic_type of rx_ei_l0s : constant is 1;
    attribute mti_svvh_generic_type of l2_async_logic : constant is 1;
    attribute mti_svvh_generic_type of aspm_config_management : constant is 1;
    attribute mti_svvh_generic_type of atomic_op_routing : constant is 1;
    attribute mti_svvh_generic_type of atomic_op_completer_32bit : constant is 1;
    attribute mti_svvh_generic_type of atomic_op_completer_64bit : constant is 1;
    attribute mti_svvh_generic_type of cas_completer_128bit : constant is 1;
    attribute mti_svvh_generic_type of ltr_mechanism : constant is 1;
    attribute mti_svvh_generic_type of tph_completer : constant is 1;
    attribute mti_svvh_generic_type of extended_format_field : constant is 1;
    attribute mti_svvh_generic_type of atomic_malformed : constant is 1;
    attribute mti_svvh_generic_type of flr_capability : constant is 1;
    attribute mti_svvh_generic_type of enable_adapter_half_rate_mode : constant is 1;
    attribute mti_svvh_generic_type of vc0_clk_enable : constant is 1;
    attribute mti_svvh_generic_type of vc1_clk_enable : constant is 1;
    attribute mti_svvh_generic_type of register_pipe_signals : constant is 1;
    attribute mti_svvh_generic_type of bar0_io_space : constant is 1;
    attribute mti_svvh_generic_type of bar0_64bit_mem_space : constant is 1;
    attribute mti_svvh_generic_type of bar0_prefetchable : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_data : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar1_io_space : constant is 1;
    attribute mti_svvh_generic_type of bar1_64bit_mem_space : constant is 1;
    attribute mti_svvh_generic_type of bar1_prefetchable : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_data : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar2_io_space : constant is 1;
    attribute mti_svvh_generic_type of bar2_64bit_mem_space : constant is 1;
    attribute mti_svvh_generic_type of bar2_prefetchable : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_data : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar3_io_space : constant is 1;
    attribute mti_svvh_generic_type of bar3_64bit_mem_space : constant is 1;
    attribute mti_svvh_generic_type of bar3_prefetchable : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_data : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar4_io_space : constant is 1;
    attribute mti_svvh_generic_type of bar4_64bit_mem_space : constant is 1;
    attribute mti_svvh_generic_type of bar4_prefetchable : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_data : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar5_io_space : constant is 1;
    attribute mti_svvh_generic_type of bar5_64bit_mem_space : constant is 1;
    attribute mti_svvh_generic_type of bar5_prefetchable : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_data : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_data : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register : constant is 1;
    attribute mti_svvh_generic_type of io_window_addr_width : constant is 1;
    attribute mti_svvh_generic_type of prefetchable_mem_window_addr_width : constant is 1;
    attribute mti_svvh_generic_type of skp_os_gen3_count_data : constant is 1;
    attribute mti_svvh_generic_type of skp_os_gen3_count : constant is 1;
    attribute mti_svvh_generic_type of rx_cdc_almost_empty_data : constant is 1;
    attribute mti_svvh_generic_type of rx_cdc_almost_empty : constant is 1;
    attribute mti_svvh_generic_type of tx_cdc_almost_empty_data : constant is 1;
    attribute mti_svvh_generic_type of tx_cdc_almost_empty : constant is 1;
    attribute mti_svvh_generic_type of rx_cdc_almost_full_data : constant is 1;
    attribute mti_svvh_generic_type of rx_cdc_almost_full : constant is 1;
    attribute mti_svvh_generic_type of tx_cdc_almost_full_data : constant is 1;
    attribute mti_svvh_generic_type of tx_cdc_almost_full : constant is 1;
    attribute mti_svvh_generic_type of rx_l0s_count_idl_data : constant is 1;
    attribute mti_svvh_generic_type of rx_l0s_count_idl : constant is 1;
    attribute mti_svvh_generic_type of cdc_dummy_insert_limit_data : constant is 1;
    attribute mti_svvh_generic_type of cdc_dummy_insert_limit : constant is 1;
    attribute mti_svvh_generic_type of ei_delay_powerdown_count_data : constant is 1;
    attribute mti_svvh_generic_type of ei_delay_powerdown_count : constant is 1;
    attribute mti_svvh_generic_type of millisecond_cycle_count_data : constant is 1;
    attribute mti_svvh_generic_type of millisecond_cycle_count : constant is 1;
    attribute mti_svvh_generic_type of skp_os_schedule_count_data : constant is 1;
    attribute mti_svvh_generic_type of skp_os_schedule_count : constant is 1;
    attribute mti_svvh_generic_type of fc_init_timer_data : constant is 1;
    attribute mti_svvh_generic_type of fc_init_timer : constant is 1;
    attribute mti_svvh_generic_type of l01_entry_latency_data : constant is 1;
    attribute mti_svvh_generic_type of l01_entry_latency : constant is 1;
    attribute mti_svvh_generic_type of flow_control_update_count_data : constant is 1;
    attribute mti_svvh_generic_type of flow_control_update_count : constant is 1;
    attribute mti_svvh_generic_type of flow_control_timeout_count_data : constant is 1;
    attribute mti_svvh_generic_type of flow_control_timeout_count : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_posted_header_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_posted_header : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_posted_data_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_posted_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_nonposted_header_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_nonposted_header : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_nonposted_data_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_nonposted_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_compl_header_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_compl_header : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_compl_data_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_compl_data : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_posted_dpram_min_data : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_posted_dpram_min : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_posted_dpram_max_data : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_posted_dpram_max : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_nonposted_dpram_min_data : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_nonposted_dpram_min : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_nonposted_dpram_max_data : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_nonposted_dpram_max : constant is 1;
    attribute mti_svvh_generic_type of retry_buffer_last_active_address_data : constant is 1;
    attribute mti_svvh_generic_type of retry_buffer_last_active_address : constant is 1;
    attribute mti_svvh_generic_type of retry_buffer_memory_settings_data : constant is 1;
    attribute mti_svvh_generic_type of retry_buffer_memory_settings : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_buffer_memory_settings_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_buffer_memory_settings : constant is 1;
    attribute mti_svvh_generic_type of bist_memory_settings_data : constant is 1;
    attribute mti_svvh_generic_type of bist_memory_settings : constant is 1;
    attribute mti_svvh_generic_type of credit_buffer_allocation_aux : constant is 1;
    attribute mti_svvh_generic_type of iei_enable_settings : constant is 1;
    attribute mti_svvh_generic_type of vsec_id_data : constant is 1;
    attribute mti_svvh_generic_type of vsec_id : constant is 1;
    attribute mti_svvh_generic_type of cvp_rate_sel : constant is 1;
    attribute mti_svvh_generic_type of hard_reset_bypass : constant is 1;
    attribute mti_svvh_generic_type of cvp_data_compressed : constant is 1;
    attribute mti_svvh_generic_type of cvp_data_encrypted : constant is 1;
    attribute mti_svvh_generic_type of cvp_mode_reset : constant is 1;
    attribute mti_svvh_generic_type of cvp_clk_reset : constant is 1;
    attribute mti_svvh_generic_type of vsec_rev_data : constant is 1;
    attribute mti_svvh_generic_type of vsec_rev : constant is 1;
    attribute mti_svvh_generic_type of jtag_id_data : constant is 1;
    attribute mti_svvh_generic_type of jtag_id : constant is 1;
    attribute mti_svvh_generic_type of user_id_data : constant is 1;
    attribute mti_svvh_generic_type of user_id : constant is 1;
    attribute mti_svvh_generic_type of cseb_extend_pci : constant is 1;
    attribute mti_svvh_generic_type of cseb_extend_pcie : constant is 1;
    attribute mti_svvh_generic_type of cseb_cpl_status_during_cvp : constant is 1;
    attribute mti_svvh_generic_type of cseb_route_to_avl_rx_st : constant is 1;
    attribute mti_svvh_generic_type of cseb_config_bypass : constant is 1;
    attribute mti_svvh_generic_type of cseb_cpl_tag_checking : constant is 1;
    attribute mti_svvh_generic_type of cseb_bar_match_checking : constant is 1;
    attribute mti_svvh_generic_type of cseb_min_error_checking : constant is 1;
    attribute mti_svvh_generic_type of cseb_temp_busy_crs : constant is 1;
    attribute mti_svvh_generic_type of cseb_disable_auto_crs : constant is 1;
    attribute mti_svvh_generic_type of gen3_diffclock_nfts_count_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_diffclock_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of gen3_sameclock_nfts_count_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_sameclock_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_errchk : constant is 1;
    attribute mti_svvh_generic_type of gen3_paritychk : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_delay_count_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_delay_count : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_preset_hint_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_nxtber_more_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_nxtber_less_ptr : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_reqber_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_ber_meas_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_1_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_1 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_2_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_2 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_3_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_3 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_4_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_4 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_5_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_5 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_6_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_6 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_7_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_7 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_8_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_8 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_9_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_9 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_10_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_10 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_11_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_11 : constant is 1;
    attribute mti_svvh_generic_type of gen3_rxfreqlock_counter_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_rxfreqlock_counter : constant is 1;
    attribute mti_svvh_generic_type of gen3_low_freq_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_low_freq : constant is 1;
    attribute mti_svvh_generic_type of gen3_full_swing_data : constant is 1;
    attribute mti_svvh_generic_type of gen3_full_swing : constant is 1;
    attribute mti_svvh_generic_type of pld_in_use_reg : constant is 1;
    attribute mti_svvh_generic_type of k_cfg_parchk_ena : constant is 1;
    attribute mti_svvh_generic_type of k_dis_cplovf : constant is 1;
    attribute mti_svvh_generic_type of rpltim_set : constant is 1;
    attribute mti_svvh_generic_type of rpltim_base_data : constant is 1;
    attribute mti_svvh_generic_type of acknak_set : constant is 1;
    attribute mti_svvh_generic_type of acknak_base_data : constant is 1;
    attribute mti_svvh_generic_type of rx_use_prst : constant is 1;
    attribute mti_svvh_generic_type of rx_use_prst_ep : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_pld_clr : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_debug_en : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_force_inactive_rst : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_perst_enable : constant is 1;
    attribute mti_svvh_generic_type of hrdrstctrl_en : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_hip_ep : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_hard_block_enable : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pma_rstb_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_pma_rstb_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pcs_rst_n_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_pcs_rst_n_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_altpe3_crst_n_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_altpe3_srst_n_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_altpe3_rst_n_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_pma_syncp_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_1us_count_fref_clk : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_1us_count_fref_clk_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_1ms_count_fref_clk : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_1ms_count_fref_clk_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_off_cal_done_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pma_rstb_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pma_rstb_cmu_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pll_freq_lock_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_mask_tx_pll_lock_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pll_lock_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_perstn_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_lc_pll_rstb_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_fref_clk_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_off_cal_en_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_pma_syncp_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pcs_rst_n_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_cmu_pll_lock_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_pcs_rst_n_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_lc_pll_lock_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_a : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_a_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_a_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_b : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_b_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_b_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_c : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_c_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_c_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_d : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_d_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_d_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_e : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_e_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_e_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_f : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_f_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_f_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_g : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_g_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_g_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_h : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_h_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_h_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_i : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_i_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_i_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_j : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_j_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_j_value : constant is 1;
    attribute mti_svvh_generic_type of g3_redo_equlz_dis : constant is 1;
    attribute mti_svvh_generic_type of g3_quiesce_guarant : constant is 1;
    attribute mti_svvh_generic_type of en_lane_errchk : constant is 1;
    attribute mti_svvh_generic_type of g3_force_ber_max : constant is 1;
    attribute mti_svvh_generic_type of en_phystatus_dly : constant is 1;
    attribute mti_svvh_generic_type of rstctl_ltssm_dis : constant is 1;
    attribute mti_svvh_generic_type of force_dis_to_det : constant is 1;
    attribute mti_svvh_generic_type of g3_redo_equlz_en : constant is 1;
    attribute mti_svvh_generic_type of tl_cfg_div : constant is 1;
    attribute mti_svvh_generic_type of g3_dis_be_frm_err : constant is 1;
    attribute mti_svvh_generic_type of g3_ltssm_eq_dbg : constant is 1;
    attribute mti_svvh_generic_type of g3_lnk_trn_rx_ts : constant is 1;
    attribute mti_svvh_generic_type of g3_force_ber_min : constant is 1;
    attribute mti_svvh_generic_type of force_gen1_dis : constant is 1;
    attribute mti_svvh_generic_type of g3_bypass_equlz : constant is 1;
    attribute mti_svvh_generic_type of gen3_skip_ph2_ph3 : constant is 1;
    attribute mti_svvh_generic_type of gen3_dcbal_en : constant is 1;
    attribute mti_svvh_generic_type of early_dl_up : constant is 1;
end stratixv_hssi_gen3_pcie_hip;
