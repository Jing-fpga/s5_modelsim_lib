`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LqEhMrcDRo9edD+6rva7hsEvko9E9S80wsGS4uFCnCxrlgeeEv1IeMB/ISIwTUCd
wc3kVva/nGwsviK4AfjaOfX3n9XHP8EnxY98kos+HN2bysLa7h3bEBiFOyCmV902
MWPY2wV4YeXzXoH43jO/mvHSdcJ0juGH6+F3nJQt/V5dwiufGeUitHpXw3Ujujtq
cPj+cCsH7tcSdky4rE4hHS8QvN2lzKqByK5oWXU8hqsYVxkE6JzmVRXkfvGtpvFP
s88n+mILPzEqIuZl0BVGKfd0gj3It+JWU47LcyPplSpmwxYtDgY675WFs8ILhgWk
3k6skcK0oFc8RLKLWepk2sCeFHlQHLHjmgh26zX1b1drkmIUGOMSvQ73BEwxyT23
LOerm5rl/Ov2nndGH6ffvrFx2Vy+bVvISRGpwodyU4a/g/Xmge3V8rhTg9pyNoZO
K49rIZnaIspYkrtvumLFAJAFrLRwheMeiqT++UhVjXGtKYZ4N4gUsAVspe/VhLnq
uWKkaD4ax5cq/aFHieqj/BfmXUokseoz9MtwhYQV8OGTzKMuZFegMJUf2HIzo4CA
VmjK9X0Pr2Fu4B5+fSsbAHXvlGrleEYu3N/QV7rmzZ1wba/sUJac3dVxPDzoX/+3
5NkgEqI/G9mmmCmkwNFDi0ok+bh4oF0upLv1Sezl5XIMuMjfEiHGer1Up0vxXEMH
9zBRHQvqq7dthr5EgekX4FY9PLR+T/t7H1ib1/fd7U9x5fA2yGxBks1tPKLvauJZ
1ySIOfKOqOiWXEzu4rI8tAs/KVzVa6WROAVZSfotqbU4vXOmeEkIJUKgBygl1kgs
9qPTBtnGmXYk6X72rWjRF6bDc88nBUY/R6/YkzBOIIRaWAXSHaALdxzrNCHC4jWE
B6omvi792IacpKtTJDjPM/pqZuT1Z8MDRDcEqkFnuLzV4QABjMmTeeWNPGWooDDT
algvQcOjmVTvbYKjg5HRJs1xRQAaYgczK9mhRhC4I94oozJTUhmGl2wkzmVWbxNc
Nhhm6uthVqrnGpWzSbwbhunOtVJ0VDhlSlkT6uJc84h4UKP+jQktL5OSixnM+GRh
hrBtQEybsV5RKblBUEydnNEWWUTTbZe2W1zfK0HzKiYrwt8kvZE74/WVfymGHZrZ
KzHcIyQct3ZlWjH3AoRbICAbKFF+njYTHP0QLJBpCB0AloSgWgYLgkZBgrPBT7/0
3HQVe5nsGkEOaNr/KiOMjefQ3b0ThrFdqRHQR2AM/C1QXuznddvlddYyRpRpW5JI
2rVFJa9qX/rK4+Clqrr8aAE+G2Ztdbs9Yz/I9/hJC52DWAd0TZdrvtKh59t2s0FU
9un2oJnUEuq0GkqSvOZgghi5qScchsr2OZnMgYmkCA82Bmqd+nLmH906M99bcK61
ZwCjrT+EIZwOtP0Rm0u3l4EJo+77+c8UQ5OOyKM+DEhoIHFDS+lonXVhRhYP/08u
g9m+EwKn7qBx6V5vaSLe7JZxJl48FHE+P6lnjJ725mQUs7yuJpl115ayc5xAmeg6
mVIMS+G2uMossDFn4/JhJw==
`protect END_PROTECTED
