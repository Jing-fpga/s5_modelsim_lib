`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VkYGM2CCu2w/7x+cDqu6GRaI0zET9h/HNbX7kNv3PMNY3sQTHPpnUxy7SfWOoo7Y
KCuBck4/xj1HojrJPFbAkA8lAyNJWAgESJJV2POi0ViU0d40ChqEtQCa3vl1KPbE
a7ZTzBcFoDVX+aDCN2FCJ3O85XTxFosGUPxBhvLLVQDNgaUS6DvIEiImCDwmbGOm
VPbDbFSma3KpPCtfoKB9e4lai99um5OcaKCh0//SN3oo8F8VBEP2khKnaxSyUl7h
CbT1RBMakjtzWqnGpaCcCyzw4+a+nHkQN6cLnp6/ZNKj0cFEUqN6WDTv2rP50eU3
h0W2sFX7rPEZpmDvzWXME6ef8SS2dHJU7UFnFIyLJ8M4UNz/d8iPCsKgxvyhroaB
i+VUHc2jY4Pc8RxSWyQ3N7LPI1U5POjYkj/19Z9npfeu+APwQkmeq6MYW1GK6nkD
B2Ikwr4TiU/W0dtPI03tLNXobeH1Y8WAQ6bVqiJ8aZ18IiixZXFU5bFAGb+BTwIs
bMuQoza95+i5vPzV/2xoljHYbiL0BlLPXRFz7TVqDc/AIlG/a4t2WpK14fjEHgrN
BrkYPokpLfoFTTSQFWauS10CRWjdGxfFKtbNT4Cng6flP2YRs3QRrtYaKL78zG0Z
lY7u995eFTl3yY9jFTkzy2eR4LXlfmgMvLor9MSdlrToLV9B8mHIyKLYAJJ4CWI+
GVTDmnGfzWDMcBH+AzEXFa1OmxJgn679Ry7gII1jNb7egsJ/lI8u3kIv8vBf6ifJ
QlchLxhUvqUNbGCHSulbWsZq47WQO9oZG9w+F6mF6UDDZo+L+XXhWaM7AHOiiJK4
s1/pPHD5TWI7K5fCgpo8oeeOmx3f1OCO++9dlGuj32Ma6OcWF6LgTVTzujPpLUNX
gi7pUs13RlCGKAIaSZLqirgbQryodkWWVTvq6MrQonG6T9FR1RPv7OAw2+F4wXCc
0GcF4t5HpQLl5h2+IndAvM5cmk3Lqonf9IkqE5W0SJA+YIv+zniqSLIto3zehy6X
2rj/fkpnzoNcx3X/aTGDZSFaEgNJkZgFLFcfaHGCmRuwLiDxAvLZ4y6paem3KTg8
Ll41zNamwkDv7taakkw9GEmsESvghp/nZYfDJkV25Ucq2+r9xpJ308ruEzzg6q9z
ZxZOoMK0AYlhb3qeBQignMCTPXhWKc6TTDFDYp9npBxjCJnECanUpFpiUtDU+SwS
2RevJAxc39e+hm20zTi5u/Q0cTSdGM6VP4XVkYc42HU60tNT9WBAYwQ/KQFFJSjJ
o+y1wDaQA/+M89Y59Gr1v6cJyZNlMneZ5mqKMzdE6vpEaAZQP+zHBiyaCdgKsxLS
bjQ6sDhE5koUFkff26aCgToLcHTzFprvPHJM8vUIFp2HpCRYxZHzGFwMBdsfya8R
ZfY+EAOVT3OpTXIACSVG4T5NWcPdBIG/QN3ZXs8l0a6Nntpt8b8LQaBjE3dkQeU3
r7g1Peq4y08DeuD1A+2ioypuJGVb8XavgamMpMs4f8QF5bFI2umg8jxefa21Yflx
5okauN752ARSccm6OZlVmF0mawpVjX3a3lUEZM027Yzqapf11iecp4V+IyqJm1Ad
r5m6HCbZavPUmp+Mzwue0I+nqVBNX1DL7nt4jRoKGk130wyD2PUEjX1qt9MINxVu
gW3fY2kgmcnl3lRBiiaWq7xZvw0uQKtRyMq/WvSNyu4n+e+G3w+2jSlLqHKeBXW/
8sCFqsSjMFh9N+vTw+RP+7S1q2xhVJDsteCwXovJGRXwJeZT1xUnW3M/fCqqw/IX
SPM+lzL0yMTIgbX8CIdzN65NFp/ts57CSkpr0zXk2EuKiTKUI9BFzvR3uwL+a2Ky
uXMpKi6bZNdMP3ZWFTIOjEGBExRkVj4cuYNX7esEGUTXwKQgKBJj9HRudFpu3ZAj
Nzks6bTsm0k9Sx8Qr7aJtnxqtCgj7yJojEjvMoK2P8G2Y0mdN+kp9b8fVRQF8ByX
TQPxeoMTGyfUwM/3MinvyVc/3FGE/QNpchTO4sFGX63p/lug2EKLlFOP35nzNuGE
93hmgwuKQQu+QBS2UxwABQfTn7eNUEiD+dc6vwLvrETCyRpy0pptwPQYlTOAcsap
OkfIZ08kOyOABSlqHUzQ0DALGVe8T4MbHUf80xTD2V3rGad71k8tsabM4JYt/Z5M
NH4/jBxfaDZSxCHMZ3O0JE9KZ4dce41IUB1pha148VSJ1RMojCTRdvdDhq+YIkri
qIQP2NmdBkT9XdtKWyZo3qkdHME4s5ylkId6ZLLhx79atq73g5dmOZriLnc83bei
7Vx9v9uotVHq/fGqXeDAfIq5q4rE/SvPY55X8WC10l2AT7J4KnSsUR5I6hYG5Kq1
Q1TqLNoS1Q/8JdUYD+kJY1OwTw3UuQQS5iY8saaQN9+UWgOjDkVpuB8s/Ga5jQUY
+7r+6Ti0HOggAY5zmjvTgfnttpejF4Wxzt5sGMU+VjzWY7jFa4ij942kB+ItTFbR
ZdaQC6QuV854lBVyVUPUCmzu9e2OtBtEtfCfY41iy2UatpIlbjyqIlmR6wK+nIOz
2PqfvfOvkBun1LAJT4kS7X5mnezrYdzg/9OT7YKF6fgkkKQ+QnWNzNGr84oXwaPQ
sTfV8oPWE4IhoOUs5CNPD45FXF+b+eDC9OYGIvWc0AqrmkdYambxJVqupC8wZtcE
bUvwb5Lw+6xQx2makhIDZcTxwISaVnG57gV4ziXHZvFWfBGWv7FSkSyRkZPNDuU2
GpWuh4qadFJjFSAs5brX7aCJkJd9PNyIYGcnjKxp4w9eMNqCu5kUtfOwgTENlD4j
q4QqTpigmLa0GQOWm2U74Ua4nWsJqtvcNkgYylrlCia3bgcqelJIIau0/OVHKx00
w6kMWm42XOXpdLy2TofDOFH/8359AJ62huOSXm3ewFdPFvJk68MLc756uy53geVu
2NsDvq03G6T0vQD9OHxRXga/Z0PT/WjCrfOZ85nHK/gKfX6Hna73CRBp1o3J871U
aQ/ckrr68u1mQhamT4cL51jfFG5LMzlm+CciFh21qCmljZy4IL5QDdrdh718yCPS
QMwzURKjELI+Ie8RpSt3VHXEvYVh7dzRZyiQiSe4M5CZk8eghRm4ofz4NocnHvHE
RJmOa8ahzxLXWckACvTeaVgZmuFCM56xEVHbizGiLXetNPO7hRVtEqGaGgoWVoj1
1BMfrd41Lqoz7NYFBNsrbYnMIDkWON7ZP8UpF1Weu7psUyY1jvl7BRaGo3iPtftH
Mc12Xfdr3zF5rDLZ6V5zYzIg54gV5q3Pzh5KNycO6ufWOBWQr+QJLs3C3J90adt8
yAhp+WV+nEGJmyMQpEnKlB5Yt6iZjU20R+dibsIqA7ESqI8QmheTRYOSWV/nWLY0
LP1YryZqEuJcBskAHD8sjGLNGkb8Po0ietrQII6GwPdwG6KKTlVj6YJ35OfcGN56
O2iI72mOG7XmIJUjTO9ynD4WHSX6/EH3+Xz0eikj0jglIeOrFC8DNeISNc1SPIG8
lNwcEbUB6SGN83nSldGeeYgoqH4wK6VbXiFjV7pcTLoVE5gPIGRjCndvS0ihp6QF
v+y1q9Rg/oGLr0NID1h592l7a8dTxPCbQYmvzJc0SdOzoKq2/E5g/ED3eXr8ieGe
BGd9/c35kaQmvC0o/p0ZjkGQrdlqyFzb2o6CnBmwkMk0f6FJ7NbcdHtDVy3ou1LT
tCvWO9xA7yfhZ1BbilzjyErERIbZjpjCPmMPtG3OqTY6h6vegXA5XG9HDvFEFhzb
K0hQphNtU9huQegh+P1soOVKGZuagbbQdaERG1A+wlYJ8S57IKKxziV1xfCCY3ve
Jl0HlvFrDUTRBVZoGypyucvTPkIqRY4Rn4I1HXnl/orkHqu7xhS07TOJqMjvUFfP
MPEjm2JFItLt/s/i46bQnkENJTv+botbOBLDqE+fID+XarRMWxa5wRDVjui6vJLa
w/l39TZ0qH0S5FMQEkI3ZJwCmERRf+yXK/3EB+lgzcBO7ilqbgmohsierHsf7JZ4
7fpO/qWsiqadqNegCiFbDFsroMaPmp3IoXS79Scx3UOyLTUkBrDwUfTKnxC2E1/R
v8Wu+jDdxrEEjUhRw+bOfV4UW8ZHX35J9+FnBdzCDz+w1izP8M2o7HmTrDNf9FnE
X+zIowi1vTfxeB/eFX0mm+Da1R3pHOQUs+br+uZKHBvWX75VLfcpFOgVjsC3nZzt
sXaJ4dSOARqh1vr+Ys6xYCucNJ7qftXR2VSv/KpS0KHD+VQ4l/ainUs41zG7dbM/
vbKef/uKXtbUb6kvpIq/9NacL75ezaoJqpVyySfgE3PeW7wOG+1PQvkWS7d2Lv8D
HONtHQCFCr8rVwpHwgK1DaSjzcyn25HT0K9m3H0iE3dSsO/ybsfDtMg7t9XX3pbk
ebDbT58n5GB/9nzajrRGKvI7CdrGfg6iuu6aElELLxrP84hmH+/9jaR6PLRgjGfx
akNz/lbYZhiUDIyOxsk8+YS5f65Y+MPq5uziFLXKq0m8pW1UMALZKnDOqmJFRZZC
+QtDwG3LVF6VUf2pt4boPOXBnecd8oUzZB0asCS+Y0HZt7G7kQ/gG+AgN8eY6mg4
j2+UWbnu64tJ1GKW4nS84pLv/kLP7p8aYg9ofrXgTkhgPA2Xd+2voPT5NYfK2HJ0
VMPNnTnM9xLQH/9kRNtJj/UjfAp6wdYtMTTvc7uxAlAv1rONhs2CxE8RDN4nqP4Y
61rRgtLwPT2xIJgjecZK4L0QfUplY1/xqXespgoTeWuB+y64oaEU7KIvpvLFOHlz
vg961nXagXVfXzw/1p7m2JyAjxc9wnIUykA2JJTjGCSrh2WeUtpBJp4If9FbeXXw
UX0wVRQjjo8x2EdlatuJ5QA7gnIK5iOok76pyQ4W8mXm1/VOfQSu6FK6m7ujPdNS
vN4yaNzsCWhGV16Z7GeqRjis4QocuZo6Uz0F/wf7ISMnXr9+UDK/Fx5zVECS65Wd
MCBSUpeYKBWrFOVM5ks3UMvC9u9/HXJbXmDu+EL0CyzayE+PdoeIFK+XCsnWefC+
mjctHtAW0hcLeULmxfDXxO+zA/IpLSeu+Ig07iXX1J0tdWwmD4ruXnhVgx8t5xZy
TvyuItjyFFh6BQEJkYGhNKd3RjYYCy162E3du7ppspDl5XXWGMcNsbqVHpePQqiU
7tISK0M0uWYLC8a6PZEZ3ZbaN/Yx3V0iFKvDs9DUK3Tvh8rEB61RvTxzxFp0cU3h
8ILWPFSiJu0Cc6jTttaoDxSNvbdpDRLYZmqbQHjfZ1iNpJaQVaTkg+8ndul5iDKx
XdDjiIQPrml0CFAlm6CKnASZ/fYL2KFrXIDfFOUfmf0LL+G0Pw4PM4yrr6Hp1x1l
cvenk6D57lrMYjB6s/2Zx6XihjUPUGmE+/jvPf5AQMgPHbG0BZg0h6vkSeNGb99a
6hHr7A4lzgPudxKjxvB4Dk/NZggE3kTj9fPW8NMuZztQPDR/goAd2AfihFcdYcXi
jy7COil/6wj7teOOOJ4ckHQpXNbXx5R69jR1wYsHT+y3l6FhdHiXu4eeUbGgxbi7
hP8116CqGoTSJbH4IJsFU+BI9uGJPhEKxYz76DtXPt5g0IHsbbwZNV5MNgkZ90wK
tk64wCF9MJ2Qjjc6lh3Pq5OxZkxaScSOioHX8Xtv2oyGEfxVppbmmexs4VG6LUD9
W4JJH3L4gLNKrNAS7EAU+njeSch5UDRICmyJOxT0fr8iYxEZafPd/KO4ZhPYFW1D
ppk+NXvFos6ichrLk3DZh+Iatrmhk4Fc4XYCbW23CwdJdoRQOSTilG2vp09Y6jLA
w9h8B5WJYCnvDEZuZb/zsTA/d6+UtbjDAcAva95IfUGgwF+mgb6nWyjEOU7/2Qpf
FnzJJJL0Gsfwd0wcJISxR8q2/9DQvuvgj0BYyxeQ5ApDvjmTha85KNMGES8cs0Lf
KonDfKhC98xYe5vDmNUYNq3LghGe7lDran3JicsVYf3KswCmFjvpiWuC/7fJSfpS
ECzbrXlFZvPaWalSudZJjtssqpJfGrPlhsjkkD3ktI47XvcWYVTq9S6O0u6u24vn
kcl/6vZaltEPUlU8dCL4viLt1/F4JvrL7/0G07NG6SdmsXNE1goO3mYAs66oY0Yy
NFqW4vh/PoSreyrLj4/Utrc6G9PzSoD9IscGdL8Z2iTrgBPl3kwd3ef5GVailR5G
5Z5IOIFxc0yxKbrfAYcPl669A2ZDKz6LO2jfQHAlRj0YTbxQMS5Iy3etU0w9IQ7L
s3DzILmSQO3nESw9wSieb1eL5DaAVISW29aI5PE7NJWQQfwkHrvjBtFFwJ27GiGt
e4zbsBMAMnnOGfrUmeKcgE7Ktnjg17Z5Gl3uB184dABwJ1eSdkdTQ/NZLZh53G5N
eQkUW67dPtJR4sDwyCTXZ2WH7zAlWqC2DyN2KeyEtBWCayuG5Xn40ABIRqCq1lFr
15RoDoeHDqlGoZ1BS3ywFpXJbT10FCHF3jUTET4aoV2wEkIC6vk38F0eSH12ACws
szttdo40OFhUztGZh/AuWelUMK5bPxbCMdgsKJWgo/YpQ2Z/XWcLl9rsGIteCSee
361JGfbONDUw6sPonlExZ2k/AGr0n8c6Km2KAy79qXQJz6pEIOI22Ocq5wvhPmp1
BZTv77nIfc8SqxfyXcNUr1ClsYG6hBUCBft4Ol7C47UPa8yoA+QXo8Ws4C3J2hfC
g8G3VJu60Bgm5eqlQ44RrWECjgdrOXeSHfVbVe2HRHbNkW3jdD5s9tUiLO0YrqE0
zS21CqagR4IInIpimyTV6eM0ZQ83XavkIKjzAtRIl7dhjxfuC7rMAfJD/Ib5qL0h
xXX8GhEOcj44gTGH5rNRhGzVA7O0zswbPHQpv90L65BczeE3Xj2K0EswZmQGDMbG
OlowlwsLqdnFDz40ngh31rA6EAIajV5NPKkq7JqvE/s27azwcQPp5IbOXK5D5xUZ
EX2Oit97h7WdVBl5ua1jX6XJjX+tu31i4MxkUex2680BhxOWrOeq46IxYbugjNa0
ZFF9jAcnk7cTgzrDX+rY2HlnkDSpIEBv678Klg7AFs4fvNWtQ+L14nSqWFde0vCL
ekGmSyySHLesJCJjxlQaVUm8inJhxlu5W4IBGW5PaNMoNwsQ2Riu3UP1vjc55SRa
RhFA0vUPFWTeQ7er7o61f9ioqNgf2aWdFLoh0b2hX/ton13sFH52Joex/DsxJttL
9e/mmYy65Ult6KZu+ntyPsJzZaEQE7hHzZYIvwhcjJ1CR2lMMVzBpzL6C5u5ySBk
26hxJmegVOnfd/xppYZ2xCLjhZeLcjnchdL8t/9j8H0imPqaupFZ99nSaQhdEtfg
C+zt35qpqT45mOzEFUxe/45bDSs/6Y+EzgVWTFdK1zkRvXm3egCgRvq8c1ONzyRu
kg0uePBMA7MlQIMPSsrda1E34LuEkJDrZsV29MSbKGK1bFubOyi04hO80TDB+aOI
16B1hZpN6pE1T4cB7QowT3wswGUP7s078+c302fqcbEzBRMHAeBE4Bxu6WbbuTjP
cnQOt63j0A+r9o6f7GJQ9/Uv4sIbUMFRE/VyjfgQ9H9/Bo0rJDNZXLc6nRFQjhXP
nDENuudXSZeC+uSM+/84NqkOyqEbs/sd1r5I3r30XCzZjYZvEQB887ezWP/VQty6
Wvs0Kznk40rQUPlzF0AkwByzCqeNb7J3h1WBqgyQXTbwCf3fYN73Z1/yIdzpfQ09
NTATdh0LDQVorMszK49xyr+Pe5hBWZ56RvNlRN0T+75EyYtMA/N8cRqPcxUY/338
49W5xhceUhFVfgZxRdvZxKbH7fNR9tj6izweHmZrEx7KjtldCliLmP9eCtTnbqX4
LP+e17gS4J6CQw/Q066RNJ1nxYGtC+behuEqdt4j+59/8nS4a8YJkY/yfgKM7xEL
5qNkZ4fAR7a2HX+Z+ibZI6e5G0moAdfMrneufGB69tsQD4jcXKm5u/9Zv+OYHOtL
q7tw3Tc0OcSUqYZy3Zgz+hBIxHeP9jTRJLcPvXciaZfQLGjy3NgXW+8wQpitkWIb
MQCrzqR+bsgIM+IaSRH/E1r057ZX1A4Ii5DT5/i8GFH2bLyHNeFRmO93qzXp3GpS
97IwIFy8Cq0gCyi5lVzGTj1AbRs4Fli5SV+zFsDfmw+1ZZUXwjsCZLP42xmUm57v
4n0krNulhHP4Q3UmURCugHoSZ+nD8N9yMmfcFOZqtlxP40uXUPauLA3rpH+Hc8TA
aTUvMU0IOfd9cY6N0g9+QMb1ZpLSUbuDsMVRb2F88g53QjVoOnzlhj3RiFX4tsBV
HHt7CnEQot7MCOsUt3U2KULq9Kzoz3jJhTsxOFqvcTK9W2FermZvHKFafOx0DLkW
rbUAKnB2m5XupC/fh+PuJRSagJl+DfiyTE8+06nf4Z9sEoDOJOpzMNzhAU1ZIJ7e
dJKmPkBgVnlg5kbi42y72z0Gkkh6xDorvwYohru6isD1uuGS8LwtHScGAFZ6dnXh
U7mC4H8Cvk4FOuQd8f7oS9NbMK/yx55TlIEy2o3Ng/xlBnIS4zxylYrxG7wpC31d
PTXWdWV4NPFmL+AgQzg2cKL68kIbYL6vFrEjfNfgOkaWRfSx+lZ6EddXaBIikTq+
5622PRXm0vr0zKkqou/E2xnJ28xFi0VF1A7GUBUprqkCV2M8V0EBUCVsydhlf51p
nc/EwnaSFPLEQKFoYoKk2QLOXqfQ4J9CC4mjKTgmRMZES0xcV1VDwD//vJI9wrxs
BRPDmxD7kAI2wUdisjcLpBAeoIlJwyI5N4NhNVKC0zaELM88LO5R3ErpRO6WKYZ1
dseg9dzM0aO84AF5qomGkIzdVdLbPFhEzjJLy2fbStDrj/6fn9+klhMexSM6W2bk
xEln0SVxMw/667mFmckmVGeuXAKL0sG29lUnPt7BbSXfnxd4araY0ZxYWAEZzlD/
CFrbiqsYRz8MXkkwDNja6dxzV8/wtUy8+IbNTMRr59VSvAtpZEs64F6YkeTGVXfG
PbkiFh53VwGSvMAEml8FXVolKdbDbRGy2WXnjCONi4ORIQHpUJYTl8mQN3XTPPxe
fnmYOkh0iy+XxfqcLsLrBU4trJ/uJLv5pRwxF2OjwSqo1MeWO7BbtrzdZYnaYVQk
Cva7s5a5HroGussOM2maI+kgzFb1GdisfDrT2kXxvsP/LH72VPCvXXnYrhwbO3AS
5+Q1RJvwYvwQddf+FhcRC/wKtU0q+LAkpCHNErrx07JUlCxo/FbfGI9WnfMJrzKd
Zg6U4ysq8U3CLT6KJi0hMvU9Hz4xAnYY3eIs7zKlU19ODrVfIZswlla3drv+Qp82
7iGDkhWVBr6Tyii3Al7sxRg5MeVGBwYpGbkMbV4VB0bmo6/imKPD7gXAmHz/qR23
aTA/KKsgjJ/ucNk5gLIOsSUy3+8VYfwFYRN0sIkEYuxFXxEzAhTlxl6jSsMfO8TK
yyLMh7Est6CaUFc76ZbeoJV6JrJh+6NNRDlncc8W3EyFbyRu0DODGrfgf0nR7IjA
m1F3aqVZFQAghmor4Gwl761KKN7X0OMaJjLPw6iOFt92ipgEZfdMviXo0OXhOFPK
ZW+tdFcqIy3tLXFA37opgu1Rdr/MQGCABVP951pH7zj7zeiCflIt9CdI74287f9J
PcKOIxu0N1t/Tf2MmNO66HQxqhqPdS5EEXAaK/UPw/gQF8rTn5R959ods9ng8fC2
YrzQBR+6vG+3yySPTwxZIhlf7XgzwbxBOHC9X3U4H1szE6YW/pMEeodVmiBjUSS8
2XGRsK0h3x1mo4WldboVUgz2RAJASBK8etuTW4c4GLCpQUMDkV+Nd4YhpfeyyCO0
232WyQc8TiniW6YWmBqgzotkstW3lT1MGR+QlmF0ostid0FrnSNJfb4cMCd7HupC
/vbpz6mMy3A4FprP3wzBEXZx23Vz8enVFchFYR7QTlfzu3jbqnYR22PSaPSOQF5w
VwNQyqNrjaN8v05Mo1IuLyiE4d7rnNU0Jyn9A+7GcM3cyMu6Ld3BUMe1iW6ETlxk
r6ay2bx+XUNzgncg5qB3l7Y2ML2VVsB2mmFEs3FHkhn/aRZoPLhFBvCh73HGeR6W
RkvT0wumTD5TNCo1RuA3h1Vk7UkwPhk7dL1L98PSqzVs8p7vbNNkY6XNK+HwWibL
2PCgsHpNpLrAsACmCM5Qt5/kOmStrqSWhzLod6Hqim/MDPqCyA1CVFvCEq2uUMYk
0WHITNeZm2+dteaa/37V4w/Vg27X1XkQjjutXkGCxgZsSfVKUE4QcpHYAnh+Dxfk
grLcE3eY+LArd4cANSkrXVc/Sp37tOoPYGQECImDnH+FSjXuGjUyYkXjvcRRkRsf
GcVitm1YgTZt/NMSmcpKITjIdWlATnjpenZNqi4yQG+042ko1NgVVvpplPCg7xup
DTXkpTT8bQ/4cHe9Y3G0feSszebna4H/8OWCeV/2i3pkjLHMQcMOmPBD/2ZDrPdu
6zBI15eQc1QmjhOviS3lQxxsoj+s6E30RzZo+5ijDb0qQPepGNyADVWnMlI5XRki
eHJUlqPKWKjLxd6kxTfIP1bE/fxVSUU39spI0pm6ASzzfJ0D0JBdKFDQOctMXjRL
j57Qlq4MnXiYYh5R6Icbya317A+WXiwVY+B6WlqrBmOV1RbTKtwVGd3EieRCoZkv
OFBHVQvC+G7qw1yDXXDkcVtmRwlZ38wcedWh0MKROkgczkcA8jakTfxoQ7kefPAf
hJSctdmQmKe7F7ivT9wDMq6fDO5tnN5FA/KFptdqxy4UK4seR7wBTD4r+YXrjnu0
i0GG/IITa/ZGSG2yl018lA==
`protect END_PROTECTED
