`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TNlK3Acc5EaIBIaVGIciC/IpnHXlU3ea6Yd1JhnjRxeMxRXFK5pAYtGv1SXB33em
l4jEFQ1DBMdZhm7k3NGCpbRiht0SpVc2S6R268Vdxxl95ky9RG6rYhKMsSKLXOJt
qhbuN3RqCkk0DojmlIOG0MvoZfNdso+3mdFV2hBs+su2FMI8IB4dVb7KsuE50HIK
l9/v7zVH9tMc+i4l+RV+R/NGb9q2FDZCk7AyJRwKUHQ/c4pV8ZvkouF5/QYCZBxt
+c3CTBfrMl7GddA655nGfzg3z/jaqIlPt8KK9ritV34aqgZkYH8H/odzCYtDfsv8
+U0hezd88PRuFZHJwSlIbEix2Twrrs5xc+cTDiWm8Hi2W7m6fctFwnca4YOTw4jo
h+RVYk+0AnnrFO8ZofWtvU87CpyJRuqus0jnyiwbp1uoODAXomUkxlhGDiCdFXL1
nBaO/XQ91uQjY8WxA5Hj9CqNI3JyOYNHK15XjaFLvRTXkVsaJkSFO6FV1ADpyox6
/CEnJ4SUd80do4IQqdP5SwS1siTBbhrzo3RuqUSlojvi6xqDo8jTYYQ9fQ/21cUV
x5g+lQfb2Ox5jrMtKhnsrY2ZOeUN5spm1Im71mxNtTkzcQJE81cb/EosN4cFPVg8
MrJtLSaGEGF6IljZGUASOFthRRXAb+wEKjl0gXnVsplpsBCgpvsfzIK1Eg/60mOD
uzVSZqWAO3rokYYmUFDNMxdczWzggiMxyWXn5jEFhz5CIF8Qet+OpkWqFKhbulBZ
8EL1qR+MvCE68DHygWjrSuZCSmSd0JRIxOcG3jcPskDhPdd/TjSvnIlxZwMHwkJh
nmqUiyKxklnLhfRjKth4zYbPawUQ7mBn2gWL0Ja5/oc1QyO6S3iy4d6QKEHkI9Mo
cK5Yam71FPJEKg+hmfEuLEEov7jaAhOQbRdUXPKcP+TXGhOOnWe66MJQQKdEbYbk
TvcN0CuT/T4E1jzGA+olUngG5zI2PTpR0xgXJA5KNvX9Vqd4LXx2VV5uUMRYmL9U
HePKlzQHKeMsdXupAnKEItEVkMQNrGSH+PgmjAJui8TFfNSFZZ6Zmxpx6OAFbYzj
j+y4S8A6bMJ5qh/e8f59OIvL76TUS4T9CoSCvkx6he7b8Gsoh2fFUuftmSh6BUa2
MbzhMHeHqNGdnvXnwRTxtFYZ6/cNQTba5aT7Vyk2wrdz2McLkGWl2PzslNShtWWK
O/1gX/X0/Y9Plx6EJEupHodURvogAFV6ZuqADmZuhApuYObJR2RhRxV/EM6SHspH
1jZj8cqtnhlMtmw8+K+w3iJTlSU8+T4M6uLCsyWJHWuVZK8gpDNG028gE8zUbsQR
TRMU7Yo9Fbupxzqjmmwo+75NSy3bY2I1cLuODl+LUbYUOE5jib2JTso/+x8Q2flR
0+H+I+E/5EnJBV2CUrKyFXEhvPaYhjhw4cp+Ws9czwchVHEeki08gvvbjVXvC85Y
wdIwhVhmuaD+c4IpNDdys9hCidS1RNKCmxixUbsYsAM/MjIgACCvpaRbNAnw7cFE
ut+vr1fDpDu/vKNQEwP23aXmLX17nKZj4hsQxhZ8LwcE32f5ftlc0NOCsOmASMsf
bptTZQxe9MdRbVvq55P4yl2uc16kdxqRKYF+VxnbcyTLCU7GGgpfjUypULS1Zru3
zsR2oALs/8n4paWhjthfzQ8goLlkxLycAOH6lkY4yIlLHaOp+i4NPKpdWYVn4OH/
NAQL7Fl6zAjMV1Q+4P5Rz0pKQdZtEfsMjbdxZqNYicaUu+YpXsDH+diX6g0IDZoD
/bwWjhsVa1VTTANoE1w+YwMlIBzfnmoAFCqwH4jxaJQbAXKjFsjBL9mj7GQjEpSV
G7EfLzemmfTyCfJbTF6Y0XMVEB+8Nr/H+mvy5I+2ZwlZvRzmHHC6qd8tAtQTC4UM
w2eHALiRdVH6sWdrCcrylTV5inmU3Swxe5WN3WuqeOUv9/USqWisZ9wVkQaWChIF
NT2hKeOUOI/Anbt+KvD8fIZWVWm3ZQyjwRa0Kd8NXKfNHG7X6aksVhHphd3idPJu
F32HFci5SZj5qLAqEoa1gyWSF1/UIIKnmUvei2xtK5g7xGLbSyun+du38iw5g41M
Oac3F2oQFcZ+ChS7/Gt3po2Z139vM0F1RHCv05Db7KxJ7Jm0sobCZNK3rgJKRmOe
6lHpdIaqAE4gmcd+uOLpJpraWqjvcGTSG+Qd0dFbaN5i823rb019NYxtbg8tgdXg
za1iB9XmvQwAUevoEsxm5dv1bGLedXDupkQuF6VcwYI=
`protect END_PROTECTED
