library verilog;
use verilog.vl_types.all;
entity STRATIXIV_PRIM_DFFEAS is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end STRATIXIV_PRIM_DFFEAS;
