`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EoRa9pbs5u9OgVJig1scdAxEJiLrERpbnGly8tc9bJa8k59YLPOrp2yie+yIc8zm
fhDwS6khnZRRL5T5feYKcq8Pp9UOOw5nHVP7wlLBHOvXzm32j0tICnk2tdGQtDev
6Bz+rdPiHe1sXTgkIIxdhflviI8497I3GQ9rOJmGuRpwwNhT8u11pBj+dlyF4UKV
VG19CmuCMhgeJoVhPWaTd5DvIA5IqD90ftYgHaVv/vC+SxuyqqrfpV43uC5aqxMA
Ti8CYUyZ4NSg+OR6YAu9EOElCGKiefvR2BCJyGjwY4TJMVDExV72EDffdTr2Rle+
w+tqr+iwmAnyXOGIuR0LblnpRQZVRvGRYFZ6WElBSwBSTos0+WDN6cuiFVVvq7tV
1XpKOPPbS0SL24pMOTWa9yx987gALFHN/Gj1vHykT1fxZjXgDcAeNn8uK4AV79Zm
6Hw8UQtaDaQaHnbFxmRirpOB7b3i4PlHbTf5AdHSLzpOY/rVcc+JuMA5cvaZ/FAz
Obh/AzRVJ2Gt2j1IYugL50VkY8zJ/w0KG/qT8KhZXuijxuI6WvgaRVR7ZUcz+frk
kFlh7XRm/5m4P+OfEuWb7kGGH8HUB/rsOFHzYU2mDXCEzirGjfTU1wxYsWTRiBct
OBAdSPgRwNTZC3wlOZLNjHWrSBAt2WGhEp0HZkqQNUo=
`protect END_PROTECTED
