`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DQ5vQ5HabIwaXlo9r2mN1m/t+ey7h7fRjMDfehKkZ7i9d3CxH2wX8XYvOllOiIfq
zUNXCp72MphFtytbOnmvf+qxclA8S9nzNBZWsRwOGeGM9C9NV/F9xwjTwSYm4IgO
aHQ44Ylvil2LwZm4RWu+h1JcsCPJOda9dMkP1sj8+cJYrs1NgKKzKkYcL2nMFt7b
u+SN1dkcCGVlrDmoy7l03/9LfSTslXTGMw1yAi/q1CJbNf5xlihBJa4aOTYiVozP
ZjnJUeDnwsmetZQ01QQ5M0X6tO7rf9gXxa8kK0diJrVQi2C0kasazm3shjveg/Bv
wPRyCpO04GPPLwGAc/PVsUPfxatcTX845XAfgQFjk5AHkFmMwy9QsFctQI/iKwbU
usXPikZTAqKziU40tsc8jjoXKdtFvh09gqWQ0TiPDr/HyUCozOBKlJwMnDpq9K7Z
tV5IgHkWutBIgUIMNSTpyh7TJ7idaycQ84FEMrkU1BJ4VdQEkuYoon3sRMsdFALM
E6s5X3EYehAKp/8sNvengOxGV/F/M0/qJrW0YnzCMy1jDi7diyB4ZwzeGxtSDBeS
sQCc4i0f6KJR3wefl1mFu5RvQsIXXkZ4N4H4rVngUUdvnrw9hhthL9Z17SMwkDA+
q8LTqi6Cda5DazTCriAxK7zYi7XWeOhMAE2wIGUm19qV+JltjBckkcgeJMDK+Bar
H0cOhmA9AHFiMv560PtyWtL2qOwfDcxYsaO23Nrl2Tk/wtQjkmHweDuIaswDAj//
SBwIsee5uGZJ3oZ1cNEYosLBA9nj/dVgFTl7t1IPV6V+Kc2LOnIqkwHRV/aQ0XWZ
cB0gU+6Q4Q021gH+X496PMigEPQKTLd46wWGBy46lXZ6qb5J9e4pkYxVkYDTastL
RZnvEiOuE1Slb4qUCogsBE397AHWqGTECSDKkzE72kFOBQ2c7lN8g4nU9yAnUg6P
PEHIkx7ZiXWAUc5KNdsh0KJPZtsVBW31fHA4d+54M7vt/0XiCoabrsK+1/WUQpVx
Hx/k2+8d0Qk4tl4Kqzgueg10A5mLjYpPOrj60LJK9Gx/3d95q6Wj2NMmWyDsiBTU
2GU1OAWmWJvUzAFMBPjM+42gsiMKbWMu+4IpDgerl+MNbX9LwEjUMYnjS4XPqqlW
vK9j4vsxBydx84xVFI2ZiFDkUDk6ldbynvkRXlR4OrBXzF4BsB7Gq+sLs/xtXtq7
r9znAe7xPPgPEgzPGsX4jdtBs2gBUvj8TEf3HAMnOLarj8PkplrCE6pmwlwUPVJ/
xqSNxUbMWSIPZ+oq1eLiXSeo0xifFyuiRizXx3/SS5KYYKRQ/TqpAyR1kr/E5rmA
vzTVwaUbrMSaYA0m6AYTK9riHaxvj+8vkf10CkICpqlLKVJ06kQE+VEzsR8sL9U7
XSW4rpb4738DMfAI0y9VFQHPYK9T2V3Y5xHHj8IT5GCRmo1W/BwgFT0frSnzzPc5
lZEieOSWGJrMrUjVydXEATGS4HKC6EawekQmLSyHsLuu/ZDIZ1nhgDaNNG+LXj8d
d421TzQjQqzaj83BDfOco26gy+s0XNIWLDH59LkyuxTA+ZTN5bUxg3qjc9+Smu7O
fdXtT62pTOt9Qmd9leknQab8KRomdFix8R9HbRV3RApbvoH5A2y0lQq6mLiTGu1Z
DNi3FBW4Ijrsm6RwlQobg4nrUi9gkDszE2ELGsiQx6PoAUqWcC7yuJukTFqnn6fp
A5GEPpuMv1iFm5gnWa5hvIzq5becWKqMT6xeIvROZkz1rImfyxsw80lo/WOFAeDj
ondtvi+LTvqmTCxLDT8U/aQpuR8VY3Ir5xkH+nXUtqWojaycwBW3CjrinbKvP+8d
YHo6WFFvaDGC8LUsPGT5c2D+FYfIr9yMEpqUYE+AW4RyGHFmklklnim0aFCVlf0d
OEur/Dli3I0VoPIrUZpookjwMDCHSEAbA6/37Hqp4yhNsbQyyTqeEyVVwghIdmp5
nc4pZwD5J9b5ZnEfXKgAjCRjTqgsOUQJkV3csk9n1KjvZMoJZj4X+iCjLmQQiZRO
7Vm/EDCG9TlvIwlVRHChDMjUzqqRvXtQkqR+KrUFTSC/VYIHpapJ1vpB5tpeWhkV
mwqzgf4XYJxmbscOAXPjKopycHZ6ljH7ZvWDBc3AZ/884KFIlKace0xNOzzJoDYL
ganBMB4w/WSkmCWmfkUvPdzFRxTE9aEl4fJ8jpYmLivadV20j3HiVlpILq0ZStcW
kL0ZerjsvIon1KjAXnval6oVWbOQqQ9QmeIA8S/qbovXH420ATrXewsP4dfVYTav
aYfNTl64Xl6+hB3ejOW3F1dH7DV9vrnPSCcSrkvX3MVXewYP3NaBxrtv9CBIS6X/
tQD/y1OvwLftroJPuMLE67BDDLTibGdjoaAGYMjeI9PkcsvkHjtKKG0dImZrRDrB
FIH0I6q//GnMZ7zTIbTGr5S8UPu9DMCKYdjd/M3QykM/3Laspjhcb7hxXX2iJvcF
/aPERzcr9TSeC1dEvSGhbpCMC+zD84RUQZvSI17sgEtu3KIwPkOLalJMYOkjZKGE
fHPTmcmHgbERv0AqFtRBOsHgpSYTP9P7znSN2Ql4Wpg5WRXPWR4ioWoU/iP6Gw0o
WgAmerBW+o/xJSdxQqnktVZdhidGsoQR1vy3UtTctVHIFrxxnbfXZy8tVnrXpslH
1f6yd+l4Jq+hkWn6BdY8v8BHE72N3yjcPQ/zmCMm5kCRrjQBfr2ydG+eysBy70O4
Bv/BWvfIcM6o36950mTYag==
`protect END_PROTECTED
