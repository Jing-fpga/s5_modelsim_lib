`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jqokzFoUndvYr4L5f1Lh9hPRtpeTT8zvjYwW4v5LlohL58xYQFcBlGAfxZPLRK3i
vww2r4lO4pASC1cAB5q28ALd+VTySZP3BD0kRnXQ9gQcqgzktI/SNGYq3bm546ZZ
goOWvsZGzMkohcHVNXPp/ujgSoVoQufIFGDKy95NgfKbeGP5eCuBfG7vH11/Bfff
auo2tQ0KXDe14IxNvVrRVmAjL+/2hHIIn3ffdx4Q9aSFjHCWHtVt6KpUHVhQf8dl
3s1qczJ+XckR3GOJA8oh8F+jhkl+XB8vGimIc2aeKpxbl5gqlRf/wj6DEX3Fi0s0
tbFWZKXfnFEDPdfWbAmy8Mot35CkLvjKpeEnQkXnayBmzC7bE8QS22jOtMyIkcZL
dwV8p6H2rKFhMjn/8gwvLNayiwX5++Sqb3GJIB63gNkDj7bjOODMkmXIkFfuCIvx
AfOWSvIZ8/BsMQje8wzOICKU5l60Ift2hbG5zRN8m35prFLFlTCV4PouOSP7NR6O
tvgaGiQvz5R0JgNxbU8eaakkqnjginChGk4bxjuRnm+F7mRo24rnCa2Qlh3pmtFk
YrdtK5zd4LIdT4YM8/YXvDQQN/aCBc4uc4mpkNIlA7+Y6ficMdIHFOBXVD0iLzHk
XCoiB3Y3cLkawD7zb97DeFr8PdpaZhPW8Ua7i88J8pVmqQFr1ipkVYfE1RCaVjpG
gRYvR++kUpJKL9dSYfDbxvArm6QDXLbLikFpBvwkMdPa+PcjeOkCt5fVw8HMaoxw
m/8q3u4Q4mt6HpZB3EHQsAMyrofo2yjeAYJkkjKp242YhxUG6AlsrmzmsynBcaWi
nxI+qNUEeVVKr84TMJz9vmtIMnhGAa5QCpY9lEiSieL7FbOwMRVPsNIQ+pOyn/Si
zP41pLsvCsvDEvjuZ5S635TmEH2E6pOrWqjShsU+TVfyyw8/KTSsExVY2BGRyWiV
nj4vQJJYzHOMWMDSIEuBoHuubHqOyI9Vh7yDZjC5iWXRK3ew2rHnqTSDYptllFov
+rQfiLbrrsjgzEANOkLjGNtJH75MgNEbJvSPEv4H9UT8M+AshIX3IdSwoIE+jqgx
ZyAX0CZrxTyN9IznxJdBklUt5RpVt8pSdtj90B0hM4f65wuCvE5ssf8McjFHHkmj
eLUM+xv3FRcX3tvAwYMAAY0Kyj6NBWwtPDLKy93yrigYfcy8wMFZpBaPSY8uffjG
GM7DpNhDjxqm26U+tJ/W348wr0SKBkFGwiR24et3Efs2vhG7f4NY4nyJdgODNvzV
pWIImBNqqofoxgLCCM9gtVcSN+ftO4BGQyCn4S3JPAJC/Yl1IaWxAF3/EwL7AJKQ
MTNh+/+koGBQBQQPNOox9QeRqw4sa6l/zuNUm3aZ3FOn3g6ifyuokRLd0aL/qU0R
l3nljmRUkfNEikVXp8CzaEDvIBHg5r7NZLLI1dBmk7Q=
`protect END_PROTECTED
