`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XVGUW2qi+REKe/8UaGZpZDKuKUc29HgEXitbPkvNawBkSsx5K7LeLiL6Wwx5N2rU
nuxrrG+6VIYWcFfJhVwFCpdneYG8zmRMk1OQh6luYSMDOW3e0RyuHMCh1j/IbBiU
Z8A7nccwT0joUvrwiKfSJRlRvLPKFLTH8iGEpSGqpjV0ZyFZPBPh9cPTpTPmFwP8
YJkCDV15lz7zXFLIiTupG+9IyWBbvU6BhdiKAa1lnFPMO5M/dwb4bovxKeGIbr6d
ez47gll0iK6AcRZCNd5zjc3dKNdyMIyfl79vtCPzkXp9AT6d9Tnfd/5zNzDiRWjs
ClL6tdFHXSMHKaRAU6ak1TWaerT6n2N7ac2/I85HWaq+22I+Lk/JA30w+0G6eVx0
esLmWeWljsveQk/1aBPsYpSyjDM9qmV4lN7pUZ8/Q8hq6lrqO6TZZBzQtJRZMQ+O
MQcg9pOln4WZkegA6ZAOxNxVWNzIf2pbdqHk/rVf5EloGCQpkuk2+MVPcaiFZDLQ
9gx53W/viYX4S5gTapgrdPH32BYjlUMZp4isaeB9qRuQCz2QDVpwua1vxS+gTRQS
J1KLppLjjBYWggfXTSeBtYUxWDlQsiMbPaXeCl5pfaC/poM5sd6w/t6ilRo9TFqF
oC4/XsnRHsI1zepEGFpjoDO8mSczdugCNR3aoPQ0DXGfpbSN6FzKCoCy4ItsI5Iu
pB9iqUoYaoeHN+ZP+HbmMserVI1BGaTWq8Xks24HOMiIaBK6io5ILiLjKdQdu6nT
Pm5g4XDIH3nlc8TSY9oM1g5cGfhOBKgZLJvV6Dnese2CB+MjP9Qh/QdkQJNFb5JC
OBWRJSqKVszyytVvGbY6dsx5vtJcW5AIYkgvE7d3oUASgRNZ67Cee3GtwwODoomN
VVklqaalc+7dQISr2JVb1L+cRSb4zOo5qX6HPxMBzYLySdIWygx+DzlRsiuBg7kQ
ikhZWdXRFa7hxrzkjIXuU5hSiU049CcADlbHusOZvAVZVOUB+EZWSCmdaxpJ7SxI
0F5Y8q+8cggv7cd3TzYqVlWOKQnHy/aLqLr8IQd8t0imlchu1S2B/4an24CKmKen
A0YL9gvMoOu3igd0Ky99ioUbMgK2DPGG1Nr6g3TzdOxThLbzlVp93xUCeeL7COOj
B6NwhMyZ2UEsbHE688w+XQg/KFdf+/TR9FeQXFNX2WdSIlNKrkz7xT32UH6bX050
ZndkHZrZIKvO7DgBGoT29W6iReKlwof/wajYcCM/PuVHqx9NA4sU0c2Ph0M5hOwn
OeSRqGQRtibE0tKcaM9RKsbfMPHCEmh4S1MVNLbrfll1tRu873aOXhIYVpSfZw4f
r9h3PaelhbF54FmUEt3qQTQZKYH05EXlA0biC7vf4DI8ufzm7kJhzVzH/hD4iugX
p1FLdgkvpwlHPEvF4ZCsym9KxEUH4nKKlBzjpfgOLGv9N5h8pEfzdaKPkwDGgjoM
cGOYNEoiTV2SLZlDXgn55RA4M36siLbwXUdcsCd9HNrjLSlPrGen50H8jTjphl8B
eeG2fv2OYmBTwqItorB8DVLldmwLOSLIVjOXTvJNvgJWASXXgnMl4v963t2rBAkH
VSYVDm9yVRdzjCTWB8YNnmGUIqgCERY4IH8PZ2KvkoB+KH8jPElK6hoDac8iS/bI
P0A3rKEFcI3wVeyYw+5YAtCKYCmZQ0NxE9DLE6RAELx9c+f1hd1GzANAIoYcGZiF
yIiaGjdxDCPR+np/lQCJ74KmVHvCmanve3J4P683LfF18DMzwAFpyZpWtwhxB4LB
5SVKH4sGD8O2Qllr+Cv2a0HUesC4m/Q3HOfkmlazV8IWYKeF2lqn2FbNlW/kREnP
+nWGKlWDahg0nFgrn0v0vg==
`protect END_PROTECTED
