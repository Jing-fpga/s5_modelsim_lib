`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ISUYNJIIcb/gNa8yGrNLBJdhM+LK+9C7sw0dNwzDiMLuntF7UXgMLJyYDJ1sBbvv
WENbO2qxrkswQrO98ioLoNxUx8qD8efkRi92W9mPBpYWgScjd0QhcEZeEcx64SwQ
LLGPgtxLzUV2LpQYqi4/ak9yS8OXPUukVzqgNwx42PuiiIl+Rqxc3PZtuA1pBcEn
hJahp4XVjcSJ2XeK8et5N4e6yhDjpHxF+jFdmb9sBo5WtHBcEfSL+hi0JuYYJJ+4
rIXwf6x81ZiFnl+THbKj+PY72r8EOeaQXeAmr15ChUUty16R41r4uJkL+WTbCvhV
0T6jxhRom+peTiA5nJMEmtktbGEtWG36n65CoFJ5SzBb6djLsw78xvDr9cL750RU
HZjR1pYcvJYWGtmYu0eggxhDn/2+wPWvYM/u2x93wrg/olT6nUxw/qktzgZE1y+w
LsizX7kOi8SlcRFlReqCXPER2/rjkKhLIJsGT5ATaFPanDojXYLMYtgJIVO9qtAW
F2FFU+aZ9lHSYQAxbERXypdj3lAD1jfQMVQyLPSWa+2UH4dJGKicLjlpLmB94prV
ccjpG0K4V1oEFwqqw44hacE2nPytaAHCVoJDiHAV9sNpRM0x/YOSfPIGg/iBl8cB
dyOF6N5w01E2IujEPaM2+UYDt8bsOYZKeCuvpGYaYI5eNjY69vRa/j9jfTtnoe2q
b4gGHwU/U5O1iLrc1GcSkURuC3MiQF/0jSiCHkcF9KAu7KFRwSLjzsrg+aBxKJkC
TkRbwEPpKyu4Susf2BXPiGlQABgoqdP+y+0F9Cv5XZHIYe3OLm0Z9oNQOpP0mnB1
2JlBhBFS119Avx03ZqUo/Jrqo2bVi/dw9TVIJwx3SSJKJ4gyaHZqSxJolz4xxz03
CS35kX4/k9X8u+TlvnYcVldRiNJFGAbhgDjRt3jjDminekXjp2n5OBT+TBZUVHTf
vG65KkFzBmlKowQwrAklwLtEcCA6El4PfldRmg2tceCZdY3bn6+y96h7jNECV3fU
Tj3QnX1mGLm4AFitbnJuSUXpQ8/kNTZi6wsgH0Stx3UcCmW7v8LGx4/pBevkDZa5
2bwgr4jTiqd1PjzAOa4tTmd8OOHTWKKRvMLxkfBJizUOlA5K7HWbpSS3B5yBtl2d
0bKCVF8WuBFfTFEBVhD37XDTb7S/z5vzIjTiaN3GW46nUFp2MnCFPCHmogOrlL/y
wZoQQoypEaWNmz2IOqB04ioSCxz4ncEINuHEGG0rc3kyOWXoOOuuu6VlMyL4VH+3
T32cUJDEwR6w/wcSiet/Dw0Vug6qKdfGDxhIlOvBfa8pkvGQmE1dMHnylnJJGeRi
+Dm8aQV2kIWOXJVS5BCqKlQynhyPcPChfhSO4/6rm/xyNiYV/Mw0vAS2TWgURQEr
2u623akYb86Qvj9V9b0Wz8yB3qf/HNZBix4aAfPP7q2CNmBls8kyinbdbxCop/JX
+0XsycP0MgtJN9fS/cj+kFjxZ5+YMzCxZQHuC7tV0s1rDS/aPSEyRtvYH/E0fh+P
5xSchrGKi9aUixwwqAJvL9aWYDLsElJGKBjp2JFgGSVI4q0cmsRiWdw0On0/LlA0
mfPN/xI3ZECLyg0BqdZGkiqIovVJN2R296Fc7/EbUiu3DHTRyYv1KkZ5mGSz1gkP
G9KIGo6xszxarvo1zOiv9HsuKXyJTvClQGWwqbbKwqaOmp7SpbBcDiy3gZkssjhQ
73l7R7QiW/iQcnVm1Byq3BYmmKgvf/L6FXFEVYYHyK5Vri4Vrsj9SpprhtLb4i6A
faFs96P8vvBzLUUj0BJuvS/XmZ2LYob5qz+crV1O4M/tmTcoTuUvwOVTBCqyxnog
3YAYCl/pHLYI/uIiwBkZnI1kX0AhfLiLVR6bzO0mtxsCRBTn1nm6p45uwQBw9QqW
toe+JqIaisQlPtvxYBoJMUYzDGd2ONicdvec1nzkjsBcSfBqII8tpXsU8sICLGif
BBF7Bn2NU+YrAR/FGUe5fvoz/QaJBNuQJH1cm9CSCLJ6x572hcD7A2b8IEhU4IYm
Wp7E4K6h0DrVup/YxY6kEveb42dmXU8IlWA4qhHEVwCJFO/es2FYF9YcM596bVqZ
nipe8h41FgIpr1osQFSrujlUraul9oxxbGwbgCW2EtBJCHN/CGbjVnHRQpgHrU+R
HlyFr9OyAk+xxxCTXg6kx6m9GQsM6ZrhDsQE5dgZs5QYkC1h2cb9VO1NNDUduXfG
O/ZgDoLt5D67vc2gITY3w9ZSNqx+Jj4WfvUVSsgtg/H9C6JuO+fT0vsvARAl7vhO
EQHGOziVmp16XbquTy01p/zeeX81DKw/N9DU0MteHqPCIokPGchJMHBMoA+GXkur
1QRphFkixy5+tE8A024K8N2zFhIBdkpzlx56DPvQrh9sAsUfzmSmsRVK4PfBAdCo
2tVszPC6YxtRo+JotXKx2mfWMKXms84oKG+whMPJaRpaC6mzpJKf9P6YGXHTtpdg
ZCupnnWQGHDSPNx+iObqgGUVxdd+6N4ni48zBsqAtXSv22wGJDLt+b2pRutYffgs
jNjMenPRIRNw8zEhDh9cTXBBR5McYxvWEManuzlsw65GJWkkxXkxqoPfDMGAqUeK
iIFc91c4QXsG1dAm/eCJg8sXJ2DX5/jP2MbVGdr2eA9Umz11Agx0WkLXeuqmR1aC
rUIM14/TepVxjf6/FfJLwhusbgJgezafDVY6ZJMsGa7aXf22HlBUA4Ym4E2uTLV4
PIFqRbVx8j74XEA4LXIfnzs22Dz13cxLC/euElPYPwHeau5YVqN+px9gYLPz2edQ
nHUl5S8dAhpR27linS9Z/tA7bZ0DXZ7rImvLqBsNLwY=
`protect END_PROTECTED
