`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ym7oc7a3YJuyPDbaEbzrKZALdP1zS6cl+U0rLgtDjLgEQYbp1qqic4zSiv/WKr0W
sp4+a0Idv0PsOWjlexKP35IVWUsNNuZcQcyp4U2HlIiUTlN7qCWGFal1g2Ja3JdW
pUczOv0gczj1Sslm1l7qCYHdn1azYgCXn0YwyJnHU486nOtIwllMdQ7yu2UIDVs0
lN+up5NJNMBfZatJ/rbs0LH5yk1fbXSlz4tGq1l+bEZ9ZrOR/uH1k7Oi7ABHylog
OLI/kf9nVn9gpUxLFZfzHfcEz/H0L2RGR5ux0YyrPgREeACUm/mSYdPO0340qoFF
qtZw1HlP+Bm7WR9KtP9bQnBn62Y4wZpGrTmkJHYLREJxQRLMhz+roQSV4Af6vfnJ
ETEX+stLhz2MSYVbnK+fGvWZUz+bBT/D6tWDGiTmYVW+QmblkpVUQgbapCG8iM8v
/2KwgUHbt3GmN4ekEWL4Fb+DYhZTCXATbM9rnGCyeEhocp0lFzxqzp91c+V0ddV7
vfXzV6C20NJoM+hvOwtVpEzhtB162C1cYJmigmOn5669l99l66NFwBR+X4ORG+m2
2GvpQqslXbKKZ8kJOV8NcdIvmT+pbcS0bTFQtikq1VK+ZqW2BIHUrsxqxlwIY7iB
QXoRodkFfcSA3IiRv3SX86QLjly00+X02WNwdqCEmDwK0VwI0HYgw5lkexq9l0c7
6gySCqpInEPKkvYFj2EHM8kKuBTKCUHzfnXz04Uv4zI=
`protect END_PROTECTED
