`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rr7p3AXCtAdXdh6uq99J9xu0tQVkzY7E5N7M/i+JUIgTauIXy5n9yuRon0FTD/Bw
CMJGt+mR1IxPGa9zZot9rcwShe1n0jHOiLH8dtuPfbn8oBSOCq2doQjc7s4Gzue+
37D1mWHvpciqkvqzZwLRze0hI4hZLNXKJKx/agwXU2jAI/R7EFqG4f8BvLwLYvh6
kzQaq0Y0eEkR7TJvBEdESFS0PKYH2ix0gQyimSjHv0FxVuK9GlqFlKk3ub0IjlFH
SDkvghuuvrW3rC+HZ+JQGtJVOfVe9X/AbRHeomKCUhMaggNSy3BeYoAInkUBxv/z
43rTp9s3k22MCKPr5a2zbBcM14b/MOuN2O8b5tu3RZDMWMhUrii9PAAKAepx5rNZ
uLL/2HaGBLTM6YWjvrMF5R2oohBDd1A7jIo5J33Fu3nWfwWON8rTG5LIKN+DMl1y
rl/qXgdVwEDdlljp0ya961z8DpzjeMWZm10JFlwQ3fe2ntCkzOEqF2reHrAKoSw0
eM/H8yA9Xd1hD8JQJHttuIQxZ6+GLbeFXWWoJc2lwY57L0y2w7ezswU9F7Vk7/zI
RFMqXQ8wUjRaPwTlPauht/gRy5aTbpz4XLjyraYgkNfhTEKSL7NH0e1s/TQHG8GZ
ehIbeEcDLwUBNolzBpqPI/K9s77v2ML10TcSrWT2d9VeCNQzy6yCkkQkVNe7zZ3h
NWNpNQmVzmcUVO/C4x0JKVW3ov7AEOv+RAjyDgkL+aFnQlYkuFGbE2/sifOk+Oc/
vBu4+eaz+R+Unz5IOdYpIbLyFe+syz+nVXwRtEsDFmcM1HW/y0nK8F2WuABw1E4B
w6Nf8N6sKGSjzTvJ7Wus1g==
`protect END_PROTECTED
