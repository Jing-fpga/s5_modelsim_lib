`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qsrSI8fk30wBWY4pCs9x/ruoi7t/XmWq06sGnKX9etV+PHVXgWKFpT1zrWNJziY7
vJkMCMeEkhQvBNgXd07VqqkUMAyxiTHJGiQt7kfpq5FRffbcV+s3PSW+NOXt16y7
c29+ozuKPW1I92VFihsFf+xClUGIlEcKf/mIhzvXE5NB0whA/24NxWqpQh/WDzpj
gVNQQocAfTBFC+6UwhEr7v4mP0TTdvkk/oy1qqSkImDJ33aMQtCaAzLv/4EEr82O
7A4xUNpGvPvcQQc+x2jt/cu9cbYkCAlHPQN1nGe1gz4KdLuRfndGtW49CBCxJS9J
Hp5iAhosUXl5GgLnmTMk6rWbeWfFyQQQXnm/7QYWM85cufriMaFw87U+X6GSjb1B
0ChcjUH1umVpBiv2WjaQzM9xA+dLylsYXTCt+LVBhbwuUHrEB1q2ZO4csalflvNe
h4Xo4QPAnzawrA7HNFcFNsp1lvqG4XFzYje9J14i0KehW4iJEGbJsbhZw1agPL7W
/B+zJJieiBBuopfRR5gdCpYAAu0N/ZJOpbUtkpozsnTa90tskbbyUYyo/Ixow+Vv
ds5asilb18DCqMGgq79iOjMrH/DUG4oGG4EmMZNUw2Lryj+mqm6YQwEA4A28wKGX
J4M0z+eLYMmMmfkU+9MesSDq1u+trokmc6GQ1sXXSU1gB1ss+fCT5+J+23BrnYw+
Ujofr86201l6ze7T1qjIux+BDts4KR7G0U5CoDd8SBcyFrQcgAlEjR2M1/9jUgQ6
V+0BEcB2ORBejGsvUQt3IrvGd87oQpn3mfqPhq+YYqFt2Tto/edhQvwBWoIHNnar
mqfPDF0TfKM5y3UU7mILlUdWjvPXh++RmGq0DEh5wWqjiuuNTvR2BI/6nSYLcMkU
atH8lc4kUfGmmdC/MSPYMzsQoEkXu+iK39eAJb08YC2/3TznX7k/rAQLSHCajruR
D6YQLB7TFQwDqjCsyXbJ8FikcVaZPneAnqj5A3nC5Sg6Q8DvwEgdIj20xJl36t9r
X1i458j15hw2NDH/xEimQjUB2TE/9fxGcWVvD/+09cUgu8jYwizE0cLmBnRVWjiJ
r74V6WKahPl7wB9Uavv5YM60IT0K2Lmd9IpAXAYXzQ/3oLnTba/7o3LXLTOBDuAl
j53YvRjXrD22Sg08KGjCOtNcA2E7d/uh4euGmDFjx4kEeenWtmRC8kW8R5h6Cal9
SVbw/Wy/XGLvafCEORqvC108hIlHr3Au72Qz5iQakJU2HYMBT/PCBIk3eEcoAcce
ovZxK/AlIkePbOtIS3VpzNTJQLAXPpQ2KZdrdHzaJM/oHQIoYteAlrkg81yZ4J1C
eu7B6kSddzqbviVPF3uhCHM2LLwvPVvS4KGC9/gcdWa/NcH5dG5qSi5fjXQfpiGO
g6GTgJITyu/w6cHZB4Fbys2RRdaWNgQ8BHZ/ywwtG5hDQYfgbcO62+nkniuxzeNl
mATzYjSVHFrGWc+G7mWqEL5SU7RuOE5g9wICTZgfdZjNPO7Q68M7gqoAYAaQz+0V
2/HeWPf0YgtZog80T/6BJyhbgl9FGWaTrJ3CUG/yliIeS33FDQeNz1xWmjbF+LP5
dVN6vA7Bd5yLYeKOFQrej9b3NJQr0NLFCD0LL1Aklt0get9uUQIBYibf8JNwOSpM
pOQgViqKYGS716TBt0RBXTAwr4OEiwdsDfPVw9zKIxw7FCbEvC6Iry2mJ+WYURm1
ETvmmFOJA/8hHsUyzRzDZPIZWh4QhMTHeMPIAiSyhwj3r7z4asSKaTWY8j5Era2R
+zn0iFm/AoyZZh6cQp1Wosd+ObwCoPd0825ejDSWUOBKqVX70ACV1U+pvIyXtojf
WEyFJFYd6X62iFGCzoF15ZwTWGjqX/5jfWupP6QsjHDceK49AEe6FvvfyjdWO+zk
ds9I0V2VNlktzl1sgBbJ1VuSdF6jC4I6hrqRIVessL1xci/37L2imobVfEkMt3n1
0OUGTASp/PKR5Wu+YTo8QEJuj50B3MnBNXyH3tDRyUuc1ziOA+OJTGeF9nDMYVBj
nDZ8fCbGbDBxv3TVmWll12O8Ro4qbRIvFuStOXj6zi5dtICnn7/Pxx2RtgtlQujQ
E8+EcemCWOI0mhkls9dFX6WM3SNYktdUg6UhzhXge2lonm6xXt8GWcti2r2Ni0+O
9VAEmeJye7kZcA9zMUA3rVCE1xAQNWUpj4LBR1KscNMS1AkgyrtLh7WOHz8tfzlc
vv644e1yLonFrLH+iFzaenkewLOcvfwb3jP9l2ly60ZtKsiyOk4kTUuFOwcc+Wf0
eONCBDsYq3lynnyZTZml6Se2W2rRsqc4yEvJ6rYOW24xhwX7KZHgxq8abys19cOy
ouA/Q3WTYO68ZlmFTmHmOvQDdhJzhlldeS6FUmzwJ7rrfAnY3qcjpovRit2H1GR8
dTkoUrtXmnz+EtWcmoGAyVbdYM28Kkc4xvvULLRB1+zE9IXDrWvFexPNW5ofNUej
3xwHghZDsb8zQ5iT5oP6jcReMlnMQikOggQ/63nsdDrYJoSGHcFy3DOvga45ki88
h5nHZ/sZveXzMBasYn139Nm5srfMDl9AayumJoe8L042DKhDbz+KOXil1N4gvOfU
sFgu18/FZcoRSyK1kDvTvluhYb4lEaAZ1OqvtiNc/qAGOrwz2f/7W9wxjzPWIrjS
X57K0IEof1+Ts1gXLHVUV42xB3xzdI8Anvhr2DFY12VCidk57/8Brs5J8wpDsO8F
FsODxH7hDyIrIo5QNje++j5ejwmOJ6Zhex+yrCn29rRfKutx1zV2uEjqG90LXwze
91e5vaLYBrYhQprWpnwqV3aYO20RovUh6SICNAOTnFM1TlrqpRQ1OBLOtvPPqG79
nJ8IKFlxgLdaIF4BtWlRz236G+vCpWsjWLK3IUU9/Wk8h+eYbGG57y9U2XP49wfp
4epwDFEz+hy7Y1/HgRgwQKY6pd/OF1hBrUdkWlIFcyKjxPPMVF5x5FaUriRsnHd/
wlddTyC9RV5tyYJSMxVdkbh2kJ/fAQp/Q918K0s/J98JBASZEGTgwg9RfPWz3p9i
grNaNVsApIDl4vL1DnxV+PijVwylSSuNSyeDxg/l2fWCA2hURC+zS7te2EyRwlXy
6uka3jQQ0VQE9S3HlpbNL6GCDjcSij/fJ/ePspbzXt+ip/eYBZbBVNdsN3eQAbPe
yn9BfIABSVgO096PRpWmYW19ucHytXOBaBCvuXqb2HGixtJRx1FWQB/ZCBLT9ROL
fxNYXXsP7pEZDTY/HmC3RWJIv0g/LIuoEOKYn/XX7VeFUKebgbciRKNsnjvUguBc
Y+0/THs15qL2najZY9dep5LLiVaCbM4nuhHRpYiAseS/a52piz3tBLERTeMRliuf
8Z0T2+XFtd0Qg9CBnpRcqRLzr4vTmd3xndkgE68iAGCFjtLMxIXE2aYkLLYOOBJJ
ERtLw2DLs/N7taIgbdse7sFEreFGBgOxmW1Scad7xle1Qt43UXi7Otkbpfw29zCk
OvlEHyC/O9vQ/IHmzSCgmFM1xqkjFOv+Zz3UB6bvPWJCDJz4TGA07h5JTefogwm0
vO8ZzKW8hQp5qGa/kYeC+VxENetdKi5EGuIgEd9/HBGh4vHtDzvxQ8k5fb8g49OF
/E5UiB+uO/jDGeTmY2jzidYhjgjvsQKWLJcvNXYfUUYwHJTkT2aWzy5qiAQzkmhj
GQSCXay07dhvDo43ufjUbXQslxw/Nrm5+jdTu7+YTXRN8w6WTkkeU0nSGQ0pBNZn
LuCcZNUF8wK24wAf7+iHzY6Nv+XgQ67WHC3et9AgS2kdnRB/ZwPBmXi5Djk8JEvd
xnDHgOvNGyLsi/lskHpoCx9O7EIOG1rDwUazPhE5x/ikbvmVJEFxY3xQrojPa8D5
9Y5r3DHO02hx6HCP/pN+7653/bmPOkb1nJ0gVUdUSSSuVjkLZurlMqPlPlvsFIld
5p3lLd0sXW2PiAWuMrILWYtWGvrMmcTPKBlC7w5twikbhg0bp6vybF/5murtBzCd
qmo5ZuuUPrBAv7hZ8M8/lawpJJ0mq+YhI8dR1Mb/rQXk10GJ7cr2VkIMMnkPpcU8
2OFMgq2y2VnU8IH0+WJlp2BhByoCbhPOriblPt9I4MsgX3EWK5FoRRbi56nwYhTM
iYDDM0HPRVjhnzXAu8wm7J3kjdQwG8iDpVUNBI5w0BowGFP+b+sR0ehjm10VSh0s
smRuMJ0KQzqwuOs6hWGubeORJ87kASpgvieqBU3kp3KL1skDGOA7xuyg7NYVpaF4
y0qPPhS7XcG+twm6pPPf08FRp26RjDp7B210LjAYn9LGa5y84Mj0rd1ch9xboB/+
Ij+jUl7tjTuT4eh4ozRHMJfG9QCDqy2l36oS740pibBjijzIbEMqyC2u5t0xDcE9
xl4Sot1Bi8wp7kIEw2dqGnoDMZ0VnO0qw3QW9qINFDIRW7V4MCmYx+DqGgO6UUC1
diZt0a70IJ+X1EBrfnOXzR8LfLV2gn9F0PoPqwfGsjFg00ZL4qI26WY5QN3Zvcr9
2JMKYVm5XbOCYc111W2LB4Tp6KWn6+FSUk6p6nsksy4fEn3W/SJBnO5bpi/KTojq
k/aUhIK7dLr6DvZl0x+YLxdXwYcvdhiEVklGj+2i3vm3lnt2yxwRgDmcsHC8Y7Mz
tBdi846vMPsnhy2tZ59/BmIx7/WWZi7dc/+OtzvdtxMtRV3J24E/s6hN2LQIB1we
A0vvow6W/h9/3IFK+itUFoG6fxVeW7WIkJmLE4SYpoUp6ov2OjywZnBzFXFhb6rK
OV9VUh0ynz0tOFiMVkuL9auIeC4PbxjOeN8TSUjcl6ncS7CR7SgH5HDOJ2cTApfT
pqf/greJbLI4cYeu126uRc2V2eLNqAPOev3LCLcSVV5DD16RGBJjkathA6nIkg+s
rsDeURXi4j8wPs/Vz/2cHubre7M6HsldamExNt0ZrHB2UR4x3V2+jQrsVKn1XD6G
dWA1h5/GfoHrXs8VH6pXGfFNUsYDi5DTG96Grthkm5RihpetaawwccqcbPFMpiEL
0aiyxyUfsG5Hju0/vJ1exAqaK5Mat2mb/isWOs4bdsM0EuDlPH+yVDa2hKiOpv8H
PT3/BZyvLHoDr6ZIcrgOSqYoESUJzNYokE0CSleZLg9wqyb8cijcWOlPXwOkdmVg
WxvEaTq9mPv4xsntHdeRXCfsfCKj1fdWjNec5i59CW6PAnfJcVAQoBVKCaim0ADp
RYyefJl/mWScb6aqXaeu65Oeqn4Fpxew0wZhhzFfnS2d2833D/e7UGFXULKN8z5U
4q0pFE0PvvsI+iAL5/cO8nM6ib+6gYfn0GtjRvdOuVGo6e0vv7hV9BQFXFkghASb
qLDV0iNgA8YmxIPkYL6sDbuuxZEpm6Y1LcVKk/36k9519gBMVxGYvzePU0sXJlKC
ploFarrewMy+lbIYPVedW6ZAIt9Lh/6jSM02poBv13sLZdIMGlAJOBaD5+eT3OAL
ayBIkrHyIPhho4hb5sqNqDNvwsf8QLQn3JMoRfxuezkOzZgwuJzVP1Zmwlksq+VJ
m6vqyr5lBvJiqqZoBPHmkdqGjlVhh8MNt08Puj3/tAA5WFzmpEYn+HfaPTY5fLs9
gHH88Z1g43Shh5ZfVaTuK9bKPIL/r3BexrUx/otOg3dbykMaqQdj9dG2Xs2XuzHH
T1zYdAqOy+sfapnjSclihI4f0BzBFF+vowfyr00E50LgX9IlbtTu62MYW362ay9C
hqJ0d+moT2F+RBM+f7UHb9WolUExIZAiENEG42jvpDWV60299JhlxgYh+VnhjcKP
vzqbi7GmkgDYJBPr461ALwLMa82HzLCDAduuxuruiBEjNd+/GJSnd2OJnUque3fe
G1I5gtXEMapD5htLYZLEBKrYjegVphrSKGZxybcf2Jwp6j/OTo6dqjnxNyjLg3Ua
b7SgQf9PVdw7HG3K4LH7UYo+g8dsn0wLlNhizQvccbNYNPb/GChAKr2AoHWBVV8K
O3ENLlb4LgUfvUs6FsSrc8zRxWczqEwVZ6RNqfypw79Ggu59YHBPzvpyRJnQ3yUS
ZGI8IwdUzd5dFvUKA1xnLg==
`protect END_PROTECTED
