`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mmZEJWoQJZh1GAViGCH6YTrFEapQdtlHoHzRcupe7cEXu8dZIw16YdXSnU0+7b1+
6aykpRO2M9+F/HtKQ65V2YbduRGyEOMB9onDzc4QH7Vwxrk7MUsLSU4NGE3mYFq+
m8g5vFOG2sCgoG3Wm0bgEk+RxDnw+tu0ReARLugr9K4eZQXY4HPygxR9tjpzxqvw
LfctUuxcAt5bqqnnBqfLYz4FhOvfqiSSYA1UUJhlkO3vQBFY2iNVvRwrqMCj9h1j
5kwUBTOgU2cydtkFrUZqiCto6+dmWIEsrDCV++sjdgNEp7h6SK6XXOIwBt3f/m5I
GoV5tKg7JAPnn+Iea3QhhPJARU7IdSb6k7J6qhnF2+/7Q4emq2Vu7MgKQMQgz7kM
+DIYYs3gPA9gxFJ6v7QA78qyaJVTkb6PloUEfHnvmIRU1pTTk70McfsixTDRFri1
aqa+ASq6bQpHXuwX0QunAd9Qq9/Ozy+KF5bsisbgCcDhftnrqJp9CBodHrp1N3tc
1CKo68CV1PRuZcfKxWZNh2ADyRW06g3MZXM2KXag2H86NRVvRjLOun+aB2I462vv
kax9I8lpOa94FDUbu/R/mhVr+nO7Pdh+j50RvwFZms26FuTm72YfPAOsGCD7ZaIi
9v7obEf/X8bb9brmuTio7z9EOLF00a93/3OO8sNPRuOcj4964V6Q10vywsPK2y0g
L/xUfWrGv+bzUivPHU9bRrXq60SeYwXHR7myluIgauh/9obBMZLVEMrGjzpTuZNY
x3xnDWmwv5A6ZEKGtXVwPQIsz3gpzmyZcWf3PuQz8bDyQ/nHLd3U/llOm0nv4Bae
nQcVltkpk/LWbjLPk9MlUtjhi6ru6IiQhTxD9hVdieYwro7/aOQupklrz41zALgY
KyhP2bnTxgujuaHwn20WKe4yPBKcDDjyuzc8nVtSkdSGeOLZRe9duxWll3D9Z3Oq
q9TtpqrH07gb0ho9pBSJWPYq5eG5SbZISIaUJ6TsSRIyZg+5Fd1I/RcifLEYxhf5
5qm8y8iH7qnLL/LP5e92kX+0TRk6fd4utienm5vX63dHyY4jR9P37/6Oj5+l8YOc
sDdSD17hBOhDwqrPBDSIzqtgp9SAjwTs77Yb9ITlV40P6y/KhnQWIiiKmMZEKLNT
QPrBBavtOwvYROVs4XYVH0sJETFwe5pNB6zWqpO5Fu8=
`protect END_PROTECTED
