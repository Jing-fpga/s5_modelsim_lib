`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9RjLXQwv+Iv7+w8ChdG4ZpMWGvNgOV8AG0nJtND/JMkgW6DRkDeZT8tbqGaK8Yu8
C4o/ilg8TlYsa8/TZ8uoZ8olrBrvCmi90/uqQqWp1ix83HVSU/3/C5Vf1oAxe3UL
2J6osxQs7t6JfTda2XF9ZyT/mq6uRW2ct1nPNe2JJP2s3bwHbH5QWeXFTwrG9Tqg
EkP3FBFaaYNBqR6ZaDdTQ/X9KtKPQ45k1jZejrKUaDentHcap8BItz+qQpjlpQzx
K+eZKL+YfbqEbm85hDarb6WkMHCFyS5BitRDSZCLxisE/L3ir3l+ToZcg0R11odY
XkelUE5SdwdcKPND0nLWVwKcIHwN4KquzUYdGYVzsPbpsbUZWjcDvBYheicJotcP
9FMvtPbfIFdlPdOmwJ+1XVeo1bD+5azBR6fdk5PmZXnVqWyZLWVTyG20Ce0BAYNe
EogDpGEv4jl7mT5dbl3v0ikX/7PgkgYOg6Ta9OIjsDgO2WNOADfNtAo587aSoSol
jAHI0ejP+pxSIzN/2lATTgpayV0GyIXnkMeo8o0bJo8olUrHvJiP1G62PEsoyGy4
O/ShFBTHtEvra31l5GIQEwBS9qpzAfP7g6kkwmnG/WmdIHztDfsm2zsu9M+Pnjsa
jF9sQtb/nCyvW6S0XdlnJDS5WQ4g/ZBB+uwtqgZqTguPGUTppFgSvMbUH0B2dxZR
VjbqFN9eBVCnzJGam03gyE2SE7LmN4QVmXPDnymS4AwoAJFdiJBiJJM85D3kGvoc
0YyBFIEbBUAg/s8l07qtbWyGrRXLdzvaFbZktXN2u0Dv6DC4N0k1iMTrF6uOIs0c
jrlU3qYECFYNuDbn51tGUZuNleKN4XNrTOjpI0r91ggEszjx0XO2HNLFTZdiANRD
dHtjZ2/l0MG0lHUPdefkFlCRrEs5X1q/l07elfXJhHff1sX8t4qqIzLTnK39V3JF
mlLJWM8dalJK40a0RU7L8k2i/K8CC+inVE9RGa1cM2OtBK6LdgXhEGceblIwiTQg
V3exKeao0vYbVczmHL0FaOI/B4sKc5hDB8m0xqymesAwPiKJnYCPf6m6dD6whkP2
tXE9jPspY0daINl6qJ5H0xkg8NPcFOfdqX8NSfNuxbk92qC4Ma7hi0uTVJ1PZeCI
uHCptqi8hMiKAQK+mzcQVOGIQsU/yLbwFxLYQCgvaNUpfJ1kKwvvfGauK1Fx0/lr
hgxPTKQKwsC56WpArepeC5AvyFaGEE5EFnStACVqkNTFpzo6/1kzop0HSX0PrLrn
ddrkn5yHzivrx0q0rRtN/GaDQvtevkUkdS3ngkM7GWbmAhDY2Wl4G46ijzEVSaQv
z6tw8mowPKj7tweHnortitchJNkkV9eg4RkCI9MXZkTtdmwnUbhDVyHOqspORxot
RXAuan9NS2MsYuD9GqmEVQUIy7JtlfG6KMD1/W0GGlWjPLJjsSVK1mFmtfOHr9md
PkEdxH/uYn2vLQCZedWcNUlgd8Oe3C85VXHXd/Dk6ksL4xrACXyzG67TJ6J1gq1a
UYb4JZR+N6C66cwfHYMMJs6Vs9AMIW0mW4ehSYH1j1qE/uyEt8rdxsUZzTcp/85y
3JmVMD9TyKjBr3omfyh1SdOyQS+u3lujRBgnKa33ds2YRBZEvLAlQc0mYOPG0pmo
`protect END_PROTECTED
