`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7qYB21LsZqBGuyJosCYN20Dc4a9VFkeBYzyTaxB8adFEUcXtt+g+uYf0ySIwMpl9
zmRiAl0M+haAKfATNCGMmfsGVxUDhdwpZvBG5NbimQpiEm4FmkrgJleOMjxnb2NO
TR6tr1RlyX7fv5TAOp9nXU+7wMswYly9rbIZd77HIpeMHcDh1YI7yN0rgJ3SFi9/
dWUHi3y9vaYvEpnnab1D7cnrMzBTAP5HWmqIt6HXdYlFBM4srkr7RuSPPKxQM4ww
37JEea4RaoxEYewKHSEbeyZ9boeUNmhbZtcbLLn7D84n8MleYSF5j/Oi4WPFDqOG
5W8hLajKiKhA5MGw6+swjB0ats06QWWH++DPxQKYQlfV4k38zjOFVrs5QBjeIXDh
YvMxc2/xcQ1zQ0udseXwb+5Z7P33l8jG1rnui/cE6aJKXbOz+TwQshK2TJ+3lFaB
P6PCsEBrWPYFII8PT9YwJd7t5tMPXelzK4YpRhqG86g=
`protect END_PROTECTED
