`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IgbOXR9VP5BIyU7ofymlV5coLfmsj9r+enWji3wpNKOBRyvfAF4dkYnYeKhXXohz
+aWfO5fxy3dPn3B/zdXDskEDpUFlGaU0vf9Y3tX89AzFliEiCnRxUP2kdVnwGd6d
qno3sJKCjwGTC9qL5t0BknsKXRpg1aHeDAt/UOoSa1vkefklFsyL5dAws4Chbe4S
5IWn0oOqf8jVgL9rtC6eyBDWaMI/uFKxmhXg/gQa34H+NxDuSkkdngzsPAd4R73c
QblUq49wbcH3bSVYDjgU4FhFkqh2ihAe50Yi3fYb8DjBDizYkM/zqShwlU6GdC/o
0ptc/WSaHu9zYuGspeUs+QCGPgg0RaJd4HANFVSPB7FKDOOIhEuCowOJEWy6WJ80
uftdHzATN4AOBo1Umu6eAUwFqd+cLsDUh6us+1oonxv1IKT8kXU8UzhwxxSiDlfp
qLaCImUoeSQwnrI3hktJgecVdYFfXaUuh1U9k3397xPUJ76Y2WtUZ0QmoyMAsNlT
czLvrWJa/CK9ScwRlmzyGKAg0YDWt+vdanuUEy1c/cPEdEMjiHNjBTILNXMq35dn
aJOH5KK0Z5RS7CyFmOAwInc2gEaLBUfGFbzYvcG0NUauEEwUPnHr1K0rSlWdT89T
T2f9SCVHuJeT7b8L1BuUCgBjc2hgDOczr2q3dISArDoGSPC9rwRwMYngPHfJpQnX
ZHRGDBKb/EFkah2h5iQoXKvtxrcD0Oda8Q2On6GhFli5Y77sh4FllOX7mbFbR+L2
/elU3/h3trPcK13Ab1GhV41H3IRsDd8d+Y8GKkErXxUmeHtyBofdxCx6lxtLr4x2
Eng536Y+TjAEYB7BiYCX67yXRfHX0GsRt9I6+9HfvLSCvjATl3BsktdPtdnI0vZo
DOfExGjRH3DbBSQAHCywPj7UTZ0N++u5QnzsE1gcMco8Dqbw8PPyfBrYyNkrB1II
j0NmlvZgVJ5eVOgOwlYMeHad9ZbD8GAmBuD2QNDYLimkiCp8CQWlcDFkfFpVe84Q
JAkSSZ1rFnydmbq+/TU/M0XaFFOYm5lbykWIOuHnvw7eas7DKO08tc97cjHy9knZ
olZSltkqmBmPVgK4uT2PyvvBg7iQer19V5plS1fYS3ukLR9LO+mv9EbxGXdWYnsV
cH6p0QzWiBvrVA4VVLDHkGE3+uMF3XSRkmLTJDBIbRp/mf4ejOOkoYD3PTG+ONUp
ggFHSBD5ZAkJ076Df0O0NsY5DYyLYFfMlXL1hDsLXJG0sMghQ1D0wAlN6U4xLh9L
viSk1Smz5Cmzk7h7x1LEEIbgYrfJFG/kJmiqQoezHdV2XCTq0pZeZOObiUa5sBVg
NKGVGzA04D/3WlxdyhaR+4P9CqHadks5zj/hyY2Qt/kDh97kmTx8f4Z3jtIIBjX2
y6oGTPwCyxftbftApGU0HOR7Bw4JeoegHmIzXQOHnzyjDujZ9tapTsqM40X3HXHk
qzqro7XI+WFdSctqMLUNqc1d6NNLCW+bZR0di8DykU9ucr5Jol1u2+rANNWdD4wh
vrJ8Y1sWqLuPXXBftfywgXb9FSrgr+k8bLHBDyr7qH6xGkFicz1ny8yzAU/8zhVN
jrVibzbncbEVU0yFXAug4R9U6eM9gvj8/dLVAf14gqAvxqjVoOgezUGbphsU0Hio
+ED0mb2HBXkOIOdqafiyhg9XU3HSuiKm2WimqXs4Vg3jhtSiuCo3xRdjFSoAy+re
x6UfmZCYsYdLXXDZxg5ZRlM4jvdG0BrAph05FbHP68ivy0GUvymVp5aFi9XtHu/I
3OZ21bpoizoY+CwOnwFOcwrJXxX9SPWpZGUfzxR262H0ym//8bQ/7V4K8J3CnnaZ
ts0BTtANUz3261Q0T2V07Iq45+nFhAUJwLtVdmAQSdOfSZ5GAitQUQmxoJp6eULP
E6xdtneil6hLb7+ZuaPu7I5sCO4FRz61I1JaHbeNoIXiovLsES4Kv/LXAST9sbtu
WYc5XLqCdNF/DjaftYzgN49j/SmVtDdtNXKo7O9TZiYRCAxn/avBiIZ+fiE8M4Cc
R+TV12LRwEtx8gTqeLZeMpP1DWB2L/i0zpGQ7MpE2hvseQl1elhalgt7SY45AWxU
881C68BGQ33WIDoHKs+a2+C33znY9T0ZQw4yjwmaWznBRdWIHc1pxASTZOU+fNma
76NzB7830IfUPDdLDyFKLZ7mZko41h3VHMHL6/aPQXMDt4eEERU2qxfgdvinGHSl
IE1oBX1etWqb3Nwgc0inhMwJGTKwKlw/NCsIWo9Vba13bvppA0vpTEDW6MeQF/z0
3WlFxw4pm52qStYiOTUsFJBrHaM14/pR2VTIcSKC6XbONi5OkZ300KtNjJIE7ee3
AQDHX3fX9WsMA3qgJqLvKyduXy6xIpfF+J8xEcdp5Y69AHYYcYKixkQw+a1alYND
+Ch4pH6IIwOfrOu/kUsc8tqcstZ4yImabUbOW252RF3rGDG0l1LWtDfKINsqCWtJ
X/mCt3N3MXTGuBjZ5tBNcgrbLQprPWib5qo82vcjIjJ8Tqjm7S1Zzl7h9ONNJyfk
qNNwVJrH75vMUoDu2NTG0b/AHOTE38yJTslcROq5t3JC0/p+t+/+Z4ze2RcZ4FmY
f3OmXY7wV9EpR2Ilnbgdk4VC1mTIwNuZvhtp42Zxtdk=
`protect END_PROTECTED
