`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rwk3KeX+P5szE0uK0y+QuLG291zypqul6KhzGjLGtN610Kc5kMCq2aduwVQtK7vA
2sbqO8ENFWQXlnC8xH1urdBs2XU+nJcHqzT1eaZsJbotl4gdPw5VCF8XU/IwgRLf
qA96F8BcMcc3HEYsFCL1I0o/hSCBsxLeW/ON9qvrSQ+noxuzURfi/WNoA8I9CHoU
jLPRZ/TAPyEJajXOev7EBqATOg+5VJ1o4mBtwFN+cDIkIuW0ITkoHl7o5kqnS8IF
HNu9Mr0s9AvV9fWJmkv3LA8wKvzHEMvVgwdHPGRY+4o/fWJKL5sYu2wQK8ZzDTb8
4xtG9n9k5wgZxSUo9RzfXeLdUkc7WN+cLXMemlUduffiKtfxJg8cwQGSbTperRxN
G9dxdPMK2Jge3cjeO/q8Z4H27t6THHXFHz+VfRU16B/GCdPyg/mtqfMBZ0hssspz
Pn0P+PwzW0AgRZs7HnfGaI44KJC/p1VohLzHPYpPge7UU6C3zbVQxeJg7a6hY0jJ
19VYD4AIvZRXTdRyXDdHWXpFLeyLCPDQUo9Kv68jmB5Op5DCKcP+8EZKHry5yVI1
6nY065vb7omH8gHE13dhZh+Q+lDIHpwV0m5o4jO6eACV6jdVFn6YmU+3nMtnaIlH
MnXditZISUtrMcWV7AqagzdmR2+ZK2lgvevzIFDACZtZb8lLIg84J3tfupH09RcZ
gait+ZYGMSUAQhvc/1QfWGwJgsQ/RA2xIpY75CESlP9tc3abueNKTYn1bIG6g23H
E/EeCTLmkyK4pGM8yZuXplUJTHqkX3fpVfdi3YZ3yqCbXGVa095gdf22dTCjo9Np
tyDtbcGpnNQTjecAw0JyMezk+WI2TmRY3Ndh3SgISiI+je91Jo677Mi/jhexH0uq
usheq/pBpT+kiyfRy65WR7pxXh41QjFBjZvhTCxG2vjPcJhaL1XZ3g7+LClopZt1
NTs8RGOY0dMpA/EZr7qmHlCUaqsfjKyhXH2Wlk1YSFDvVpztD/5kh5MiBNomNOnz
yQWU+8VzSv9MjuH3SJZt+DAcWX1XLhfQdIB5/gIoYhbNAnMvm00H+yWdhIr1Cx0e
q1oIaxJ1Q2W0Niqnq+6/WJ+Wt/sCZ7+GDi5esbpkt+GBysdHYQTsfu/yExipDZQ3
jR9zqn/3/AxBO2S56ftcTX1dWSSw7Q3l7Y++UYRP8aO4TynLVIqdcx8X61V7nHAZ
0Qcip+iFqZeSXpQR1zmjsMfZUB1MAnE3zq6galjCNcuoOXVixxr4T9MU+sGy9Orr
xGAcYKAwg+LQR6bipyZ9Dg4dlBz2EZfWe8aaj9mBJRG0B/axB7FryETq3xNAv37u
GQlGZmSedlSL7lbosaG7EwTzZORf0NX+hMLw8UiNjreoe3Qa4K+FmJH/8z7glG7x
rhGIWh2xdZVBGf2DHtr9AU9T7O5XAM8fHqKxhzaea2YKDYaYX1/0pmJiQC3VjvJS
Q51oZSl6dEObsCj5aLVffVLw3TAToYJiBrueZNJi6Zr+My4sD0DvkOUCFtRekFW+
O4HZZtg2LVZwjJ1K28FUEjQ+dNKgPd8s4XjYIg4ptTPt+zBONKrOuek+Kblpbga/
2CCyEn3dYvWL8mLPihTlKzONhxKZtjw27L0RsD5wyOzAKT31hQY5OOFIBSXIun3N
HJmzoRvlWyb5p4EpBcH8BIrhf4boYthVgd/k3V3LdsGA8ObKy+Sl15xv9KEUHod4
EqFf6yr2J2k83KgX65b2GMtiRg+ofPOX53Z5J4yNBFhNOAecrwyLkQ9cPmUOcF3J
KK3Ev4wdIn5TKE5A4y9C5O4zzzdj+9a5dj8BJzKliK1JWFTiHNeC9Qq85oDx4yId
0+T+5CfLJYpXslYWosEUV7GSKRtR5pVgFbLTsNXrSIJw+DeGMdviZfPmReZaEltg
R470G+K6lj8S7fUuFQSCtkMKaafCTwbmgK8IxM4iI2jF2YUTDh5uPuFqOZwtJA31
Dbs27zV9MTXnzAUYwx1qVpcEoCFOJRrFBbe07YyrsGeKsKVPcsT/VfEpwP0GhFut
Ja3W2ZI09tpgJYaTkQOgQHIeyw21D2Y7J8cMalmZkSJGVRXMg1eHp0kD1CB6zFqR
I9uuatH0/UmSTDqAlNU+T1A4uRxuejR3JrZrQcPMNAITPFQJukRij4s5abiNvnne
29cq0Xb6sV3yrivax/DthsZTdDw6Fjch49q6ehelAja0wwiJeQev+i4DM/gcv+YW
X0L9dj96MBqVBUF/h2pY51GrFkuN9oLR5NHsxPdYa6i2ZgPLWPjgwsEAGBSFKweO
lHHXOFHYVbNgGK27SRTuaDD72Jz2/XIkXwM3P20N5hIuUvkhVZNfJtMdPyjZRDf1
PuhjJdVaiMMxSeVKOnIVVl4XUkpgvVnCn8w6PLisbGYrbMJgNou94BiY32vmohiN
VjE9qy8eicxHBCv3hdd4PrFVWpAVqRNSQEO6sar4vFxgD6+Og+l/Fzkpxaof6EuV
/0gZMoDnc06SKkVVMvx5A6tp9BLW8cOu8oxEdDmp8Rc=
`protect END_PROTECTED
