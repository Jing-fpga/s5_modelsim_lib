`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3u2N9UGKFxs/I7wZM++yTQm3Mh0/mqBuvZSIbIWGQjBXffmDIshqYQQsEXd+E5F
eF3D0gKgDLx1Ud/RrBp24h1IZERj40M5A5MLne49XSqsZorYG73Iz61tPL61u87g
Vl7lU0DC7FvFU0lzC49js2p19ZFjsav19l/Ift/MJt06f3Kwd1aDF2B3IoHa1QMa
AnWlXDnrKZnnMnTvhUgC2eALFdT5cIz/I4feZoE6Pq91nDaeJ8I4BqOeYghrAnru
+4TkGB7I01YZyVPEwz/AGas55Dcomyeyk9lpg9kWYziTEb8ADkumt30EIDuCewkl
l+BJVTjt6a9u9yLlxoj/KCRvkYGCXHVhuzMaEMhUsDXmbgsue83b+KYia2IFVm3Y
uER1I6pu8DpeIzxcAk3Kw8+Nk+wl1FgKqteG2rzEJ0zQJ1rNqb5l4nPp4K7FQu6L
zND8NNg/CgwgW3aIfJpVl/JJWNuIbg6xadnOF9EQzLytu8p88+iLtocRjDrDLwtI
TPQcnrrFMNhmrra+nvLQ2kc7D6t4x1iWpBqR00S3u70ncx7nIRu0iGsISK9vejwL
uTJ04zM4IqKPKIhxgOWM5g8cNncmybHk07X7rZ7o3qQC4rcpBzqqIcvMpKF35bX3
8XnVxWS43AE9M8rYZttI6YP/qfJgrQj14PMcQu2lwmNrCPHSHC29ZocA0jFENCEd
7CGV1UwrVMo+oa0PVlqFjGbTHW94rpPHx+PPItYHBM8ge5UiPHzlg2f1yfZTmvbx
o7TwzRRBDoMP48/0y9ZFhZFwLZuwMmWqvMpA3oEgYZ7+lUHlepK8W9phJ4MhDRax
R/YklLu/5LJbOPe2+V3FVua3zScfLUSzmKwabGaZ0kVJvA2+ujOqP/mhy/aTGduc
JSmlIKAStgh/jl6+xHWOlulBmVnkX4yFHRhZg6KDBkgrNSiAgdyrMozWLKOyGU13
WTNkAvQbtwodnwEM5sZ93vd8+KkjZ8D/3nN7xtAHWbBqA7vFFAgWJHUdP1V+3y2c
yn57XjEhBaoQ0hBV2B2MmnP+YhDGUqv8mT6HGvr8h8kRZXC8rI2+j8QG/R3NdrGQ
HlmQWg08N6vz20akACxCGnuM7iUwtT92N15aIw7inXPBACt7fb6kp7WfbO1VBRBr
Bnk2aIcuV1hMD8dUdom9a1ewFuwTT+0Mz1ggNX5T9qu7dpPYbWw+/4LPaW8yAzKI
zrMclsD9rvpI86q6lMIbvhJ2K+T/QyhgWFr5XuEU+VzxiNgBAfZWq3SBg9gHhJva
NYgU6950Ig5aYqh+oCAWouMpc4sbkn7pX1Tpx9gv9obKp7gLMc3PzhpUv/9Zerno
B9dkQbdiynMWyq/7OuM101Qp7UA3TM2Huw4F3/wDV3OfaTwC4jasdnmdDKnwftnI
SO5tt4zEGGiTWyGYKdyBGlcizFM5R8AS7ro0I4jRR1VIG05r/UhZzyXZ1XJpCKEc
qLdrpQnCfaWRaI0b48CyfS4qDhJpJe7O33QPuCrlouhnuinc6krFHnyTDvZBvz2q
XKWdNF/u/oiKAJ0FZ4Do5QHL+rHkzbBhKAKE3/JoCYNX5e0b/nNbGhoF5Dc0hAPF
VU82ZJxcWIpfpNr4Jds19GPW7F3Al+mKxm5FzR9OYE/+1pQYMXP6xnRVePsbmFpv
TsJM6ys5wc97GOaTPvDMWuvsTZ4A7UO5ddDfk9/KDkrQBdw6PyofT4KcZokqQet6
CnBNKtv0RTjherDJCVXD5zA66vJFyIftujjFHq9KbKqqB9RiXwFMjtPhoZqijAN9
7Ur7Kq1AA71pdkW4/5lRLVPfHsrIOgquiA1XTAHVhgtErnWQavBy/WLMjqVjlAP9
TQmikuoYOXIno+HQM1q27yC+J6MQPhB6kf4x1g5kGV3ppbJVOSTuPyLCPB+ch/yR
GmidZxxbslino9L3GKUWKdOO+frXwwHuHRA7FqzMxcm30tZqMg2wbCtUxTfuB9mg
9D+J8chXIGZGKjhOXOiCe/mxK7hpHldQisxPRkkjgKtaNtpTnCuwtUU/qH0day+h
YGywAdh3lQ/WRetDez3rihp4U9gXIvTsvwjNfuOkg0zcXOn8F0vqa0ZW6N+dPMg9
5b0BpUBEtVbqtgZfhD8TaWqKzMW8VlEenF6oYzPhZuD1l/NDaDBbIUo9WbHwIm2e
yYFscoceJ7jr4vYVVl1tt0SPzGezA4umSUiIokYWD7rPtvvNZ1ZQw/V1LsCwfmHs
4/wSJZEnu7Uh37QoiE1fKwl/NsWccaNTo89IZ6b2tjSJ2BzxesyvhZ09Pi6fJSZ+
R5tSYCT1UQ05GfQDfqZFC9mbXAgFFZs66ksjms7N8+RU7T7ISuYT/qTGk+DVmM/C
PIXzVtBfQFRE8Ggw7B483W7pS7e7UyoqhwURCNg9XjL3afycX/mxkhxrMmgBJ7SF
91VGhbZ6qoCRdErKJW70eAqLUSkgH1ftiNVx9lbTAHrpO5EbLXTLd/QAmaU9ya8F
NrgkLjijd8ZSUY69NvW7odPfHk8IY2QMs9kTPThcpd2/R9WcEDWhdKDFvPv083Uf
cia+HI/4JfpqRGv1GTjQd+2lX+GfDnQtkOQ4QKtByYZ7j4T8lomH9ifImRDkai6A
zzTuVl4GUbDN3LXe7wiFGgTRk/6NyVjRfmSx2bOyc5Fiv5GBH+wuHjTiHcLNQC+6
deASs8bSIf69UQpmNLBEk+iM7oMCvHMiPLOT6fEui5DTkkDPJkoOJ6Tyxo5L/Sq9
2q19tP2gKLb3livSKa0mZIh9RM56cXqZ/2xjVFHali/dQXRhEN1YtfJNjxaFc+fY
hkJ/eBtDb9UvM3NhUybGhLZ4SIAvsj+MFevuo983iLAtEYhFqDM12m9wcAZLbzm7
Qih3u4OuSJfRU0hsNoz4FWqn/y3lLyvXd+q+jEASzwbreOcJIa0tG5Ia2y+4ckPm
pScztJBpW7F1UbZaOu+5h52a9fZC3Msrp/5wjNr09D7K5Esdxjpgq8Rwb6QjtDI1
lyP0RvAZ9+iIx+1crp6RukS1ohaw87KH4ILChpgXFr7/vQPp329eb+DCS5u0uFud
YwW8HLg1qZB2WRXlcQtFEbtFZg5gAvruDI5hcE61eNvNUJ1TVZZdPbRhhEGi0vaT
QLPhhJDUREl4FjXz3c6p/I4WfYSVZEzUUrgu9RId8jK+vRy42YFfEfJntwBONW9f
aedFIfp5G/e1w6sXDMqQMQAOPEIRFihzKLibDftc6JcM5rY0QJXJ33cm6nlUvgmq
9apWcwoVbdFWmFq25WjwbsY5ioqtwzemmqloS3u1vaxLnBzfPnOGUYPzTHQZdgVa
NJzoX7QKeVCC6NzRQhkuOZdtEpTsWd+MXHcXvQSK5xH5WFNJ9hpYrunxY9u+07cg
6gdVwxIndGxyc5iTYhpcxEdpg5+z3PNhqKnuuQkkenv2pWlFqiHCvpvUBKjs4grB
6q9D6DQNRrDZakgdbFMYPVBbtHiszGDWfYmuGONrKfsETK+LmsxRtS+2rs0MlLkT
sRIYI9EgsYhimP18A3nHZ+KkFz1PyXr2jHok6hBYt9H76TPcrhAMKVGTM3Du5rB9
ERyGK7vuTqUoEOdpbIpuT52t5EEaUL+LMpzptxnrkuJz+X2kMH5RosPAdy8r4eQK
qMv6MiJRjvtHFXD+de1ygnasz0n9AFsiH2bkOr1oYZ4w6fKFsFY0vhsYlb5efoKf
Hfw+y9X1U6C9hxF7LS5HUv4BQIIKVsGLwell7AKutcnJsd6CNghlFIzcA/lNJ3jH
lMpjG59+rO9KQEqv81ATaUZnJeoLOQKYKrANfr6NG/tKvTzNqGNY9tz0LygOgwOI
PtCGVNhWYZNofRfbu5cZ2DaC/2OrH5EPtd3a4Zzut+E9zZzaik954EwV69F2Ebz+
niynr0eVuwgVzSLpKZn8fulTjUk4YhKZqVUjHFmSxXOzUpH8qGddvQnjYSI56Rsf
Tt5yixsIkwFBmGMne0rD95EGSQ+V+/zQE+5R3oFbT8f3twOmBB/vNQvlS7dlxQHO
qO/skurpBDH+ikFE4Rf1E/qfvKN/3O+h+P+I5GQRDANqmDj4cYr5D+63t6a6sstc
4R7D5TcWvbSuwYUr7ykg6EfAVP7qrbucfG5+XvjGu2tGmZ/YkCWmrwLUGtvhogKr
A5hPdsF+EmBsbgjYWppQ7uM/umBcWQywwMoX9pNhL/Hnpmc7Al6wQDiTiMXkIOwn
bhI8CxMPZyBDI9yabXjKH1ijNq36S6m9C5gchih1SAVBbQKc2RfpXL5zA+Y4qoLR
vl1lE+elhGzSdfHOIPIl3nS+tKpOzO8vGQk8t5cScivvNpTMrmd8TXQx4Xjtu0Fm
HUCXl88JQbAAxzOWYCzoavTw4Xn0RGqbhlgIEFNXmfwDrpzAkc42okiMQVLquNOV
+x5Lw7jEkaXUoRQzbc3EEVY3mCLwG+jYmG5E8EXogsEj2m+RmjZgrtbpQsSR4lkR
8UMjdikpCsm2Qe3gVjdsbsYzLP/JrvleRLXYRVAT3AMPXnt9Ub/lTrGhznR06QoF
RTneJQIcGj6LksUes7LNY9Sla7miiRYKvTfXQEn8+yighUhuhbidW7kKW297KdJq
Qn5UpmwHLAQti5WGKy6jVgqRRTjflz+bxbQDbsvON+Pn5iC9ebGPjYDF+Vda17ev
FIK3BYTMSGXJBJA5S8zRjZmmBquHrXBJm1HWBD20boUHPCEuZ0T6ZpCbFc10xUHy
bl94hFK5qCaOGIazRpqt3ljSZae8tWXP+OI9p5aMceVVhaa4mVD7At5bOMsg6F7K
mvG7nb8JGYXRi9rodD/9dxTkRCTocG8VRSGx0Qs9mrGCIMUXeNp9J1NbRdfAyJOp
Fa6/xCca9cQwQE2ZqsosGWfq4LRF3SFzy7q6dGFFy+RaJr9gBCxxZ+CGD17J1nWE
TYLi0p/t01cBKvjUXZTxVcfwDtZM8XMt3bllgXschhobE/2EF9sDd+s4ta8NVEPu
waX6w4x7bbF9LFaFYNWKunf6F/lMmpRTZYK+VF4r3w9gqIobDh65y/0+r9mS/A4B
pIA4+crakzr5r+g4qSKDs/HekaX3QBMFIUSxZf3IjvE/JeSfKAEoh5tAtIzdhvdj
lOvvZcFjh0l8DQR5DrOoCHMf2TNrxMt1bnIcAzI4mdeLK0ynzNoNW7v6XlCXEqf3
OtYZDoYsIR11ipchrudbMGQJVcDGru1qWxwAjZDJV0b77be7XyQDaKX2aHnTM1C2
FFtmbOzWsG9ysVjQWcgbc3tM3A7ZdTWIrluzvtNBpYxJH8UIj/4mj89KnSYVS90t
3pqjFrwpoP/AdY5aGbVgIQCCuAcS1849rU4+EHEfOushZc+Z6jZBaSbfY0ojsq2y
5k5X0yGV8AAUUZmEGbijIwZieiDcfAuqN2zIkDJT4zCfdIVFDubWqziuqaLMAA+D
kigJqsrQxuLhCNiNNaZE85eRahCJVKNlpnuXM8jiIe2C2qe4/tEyYwt7xBVClkt4
2SnOBZDBhQYcHzUDitFdrqnGrjHkXtJm2NetWZP2sNMWIswalQnvSGTumY03iXR9
HALVZpGORdZ9J0tufoxoyud1GrhYZmZdXHlenRRNlH+/cFDwzpGOAGgHQudKhAdN
3IhBPWQ1VL7Fxi8dsJtZKdAmJSPxPObfQkc1OhXsU52t15iwuvypf4nHLcWUGzRr
6bmo8HUMXo58NIfFzlt/pFSWASmPPwD8SZn/16Ok32Y/bFgRT39PjrgqS1e85cj6
E7eXN6V6Tz37zqD4c9fNEKkoYl8K67xWmSIQFF2G24OzIegK1ZDA1zk1mfeq/iN5
5qvcs/Ed5FnXF8OB7NsD0mxloGuJQHZJWpBvQJCYTJVmJoAc9V4Gm2TMzIcprx2g
sPeXM/iXpQqzgFO+rB+kqMvc9LFVLXFHwoExBPWrPBHrZ1hEES4caLP28Kjt3T7N
afyTqZCUfyA1LdAe6GlriImWXt+a1vpsvbYusxTcJbt/Oqf/6BjwaHnVCuObosCZ
WlhUckzWpBFi0voDb6wEOhh8Val1uyxVyJIAvHIkhmnv8LKmIuKJc5SohQc2stKJ
kvaOWfmcXjIvv40LxBWOFa/F7ApVsqs6b5Gms5gFlDhi2mqDTqNrckX+lxoIPHSl
WK67u02jtc0kmRsSuAR5dBbdvX5wHIMZtzDhWxJJFIjP1Kv+ijZCcBNgLPk2nU78
B+IC6YBZ14BBx2dDVriAh4f6Q/PdZpn0G9wvlm9YLaEXL9fMItL4XA0YziJoNXWA
4YPewoNZZDXgk3QsBccuCC21k05cBvUTLKopFzgkgkjyAZqrvJGysanJ1U1oD9Io
Jqo97qavQQi0sMfFD19ZLZgSfDwmDpSDGV8KWtWZzhAeUqqWtADMZ6VubitXAET4
+AOzhJSxa7JLIK6Hh5QanQbxx5htK+uNqq7Z0NiC+unQvCdIvwFlVaAWcAySFfOh
swSDgDvM4b6M6YOV4+Nz8ho+aPKXjZKz8qgDVLeZXUtoIoMUM/kzzfMycSHj1HP4
XtKXZ/V9Hq5Y0caI+0CV8QBHlMbZbg8HSVdu8YYqFm08zPY2yeuUCxe+Lga9qm+f
lv91rH7ABFuA3ymCNc4XnNq+bm6INaBSoIRvA/WnlYN+4GilBTvM+BeH5hQ2SjUz
HVWIdOVT+54ouriPpmY6g3/BN+QPbZ8OMyhonUUZCr/vf1YG4pzEoaEaqFfS1hvV
boUzrMPb30CmLaQGUKlBN6cn60ToSrjNuEkdmkEn/AlR4VvMKkj5RrwmKBhA9IHE
ySdD6jRX9kZ3F86fEYjQ31GVOizYKYb9djdBivzEm4WMkIkevZM1LDt0i+JSeDdU
Os2AacVwXlm0W+46+DqTeNl0RoJDOLdWOZVEhsovn0IKDHgno97YLpMzhtZ8gVFE
4aahaOH6wiDjWN9yZ/kEvIo+/wWp/Yw/M2b3A+46CtZLMlSGUWhIH4IbZdgNl4nb
0SWj/BsOc5fY+cJkPDRmJr+2xKMwxuWON5l7p15RzIDPhtTivEr2e/Wm3/YQw/jB
2BKkjA89xcnQYMDS9jhq6s54/HJ12AYvhGBj2ugJjYXyHo1MJF2ct88tqVF84rgb
EUWvV1FKnGSf97a5HOzctOQ0m9pKNjwD4Yqp52WdztUljoz9ttxwNW2yTe+VGHMs
3Ia3RcG8qQdDlx6BP14MdH35hsEDa4NqTmeF6eJbA1QNs6zuYJ2/dYT2hSjAwNiq
R1h2K73tY0Wr/HwAZWUk002jgUbGMEIJa9/qsA2mAPISK1rABJbceMCHzdFbchZn
MEZPOdD1lAT8NaumAV44VKSSGx2kJKglr+WGJ8yxYt8e+YB37JUmceq5BmzaIV5S
WS+PF8kMOhEg+OKcqmyQg+USH+eetwF1tdikVZXf3B2urRpEBYwCBf4n/E1dweT5
8wDAdSy8qt+aYb2VO8D2ICW0cC/SURiPXrINOMouWOuV5WR1PBmtyVx4n16m9V89
9y+kDJqWvZmr2X6VfbjYIWfplOMc99oWtej3UzUyiZ0ziVtm7/Gix4JivAnzFf8c
Wo6uUDcHcq0CYDwVT5gMAYgD52sQ/wocFFx3Vq390yicTIIpe0HnX0Vy+v2XKsdf
IRiMKxnHmoc9xMJF6hvHx6mOQQNiSF/D11bjM4lbzHOZRndJSxrlM3rBmEI2BfvI
Yj0EDlkOn7NmLcFPGlMmHb+HxI50wR93kU6oixvUgDus7iYPvBH9tCW3GjPWP0m2
aFNAfJG4Grptz+zr/kKC5HVvm33ScDUR0Beo6Be6sE4=
`protect END_PROTECTED
