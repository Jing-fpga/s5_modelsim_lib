`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RKk8qf0D6Po9LdUbKQJnPraSMDo5quFi2wmDvQIhC08sZiV7HH8OVZovmoxKgBii
p7H37H6XhRSsjKbyh/uMJC3gqR4ADf1lsjeMEjY3cD/jJH03ysYIAHZQgpYJXJEl
s80eUcXqGVoHp0gx7+r7KmwJwAUE/LwSyTs9s8iaYvjBQb9opg0slqo7v6mA4DoV
yFVDNJF0oceJMKPziOmZhI7JdDbMXOqWOIaMSnFykCTTKxJCy1JldnMDZwudiKc3
osm7oj2mRoBOMOqZ+4O/in9L/ZwJBhqBZQ3CmXD2G/OzaawrOox9OtakCO0584wB
Y9ruAR27PejIrms6rHhE1TQWT4ozDntxaI9Kc131y/0ob9RXGu2VFHfKSy0irnnC
+eF7eMA7tavzYMI2YJQtB/weHI32oOP1jHuXMOyiMu1xBv90Y3FpX1vy67WV2cny
q9JWf+9LTwW/S4qXi4PvA3COzlzRRKYaGBMfP0R5PG6q+hd6WMhGR8KwI/RgR4fp
4I7Ogu8QMkgBgIhqI+WxZUxzh7RZEC7NfBBm+wIubtzNRBIi7NCCoRuGD5odgNd/
kMziW9addNWYD//H6U9/Cz0sciNKCHUV3qYkTVNZHqJQd8T8MfnFwWP39R0X7/bf
inXh65YarZplZBMx/C4gWa/sIeJw1TqoO9ZEcX9a4Sb30m2ACnMLwV8I1TECFE3b
BU0bFwSM0dqGBcOZkpIF1AahL6rbuE2JnDIWJxB7ZXg86pPb8y42zY7BQiQNMbKg
SSV5bxyNbAA06oFnIrrCmtxqN1Ww2N0CkpZX/SGIHddLqkHSBbw01SZHCZApHujs
wNbktULGNEHjkKCOvKRRu8ad8M0W04AO3lhwLRRRzNJz4cXj4IhiuoZWSTpdvgvI
mxS33jTqQe+ASJ7kOy2R+Vml3N9oZHuzHVlfFd1tQV71iLapEIm8QfSyrmiXIbmJ
wVmKKvgjuHs1fNCWAn+4gpaC9hiS7wHtWVDlLgjznmw9EozWabC/7iQvEXE2kDKn
HBzcjgj6ymAAKqHCm7/vvfZah6YrEdCrecC18eXq8w0lrDHoSNwkXk2pQWUmtSyU
RIRQM1U+L1RlM7xZmFAnrk8JiGl2fXQAsysQg2GHL8s=
`protect END_PROTECTED
