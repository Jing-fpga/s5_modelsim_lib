`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7QnX33cqufPKwWe6mtIzBFB0yQqWfYr4jZ89SvqQ4x31Fm7Pxll4uE8rIavRrSas
qgQ8c3JZL4eoGq+wUNGXOGccP/3ANYeid1/bEAQlCns7um067ks2dosn16MbA0fO
6jvw6+F61zNQmOx7fcu1t3/WyDRtx9YF8ZVQnxkD6JgDpNrwibL3JQyGjS0oLIvr
y9/MNuOFjGhT/VCcgn4jN0Um3pLxEHhHIjLna8T3VXwQbkN1k0jwVUp1w1qZAG2d
xWIm1JmOzRZ9KhhFROiloc9q3zOv8aGjKw2je7EHR4HEZwMIn73OyjvCzTxoJUSx
wRhsp/FZ/6Tm0FrCQq+lLxju+eoQHRWXr/q49WCSS2rKWQ3a98Pp5Gczl0ia81E9
IbOlHZLf/p0oE9Mdaj8eXOETcGMs4wId3yBtlCXApgQMgoH22QWaPbVt5Q99Z/fE
BbppS07oH+sN8LKAzNES3b1crnso9nw2CZOu8dBTqoaYdF2po8S7bIIbUfg8OCPp
9DL41MYf7ndQ4RfyGTKlkAOZ7VzbRKF7jJGZU8LX+AmqCUK/zHEPJeR000jzTRXI
EvX0AvUA34LikhmxEmFkhA==
`protect END_PROTECTED
