`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ACXT+V4OcimAY1GG0r1itWud0AjoUyFVREIxiU539zdTNs8Pfam2MD8fy1v0o/pW
yOeniokJAbTdfU+FcKg0w21ysSpx493Li3asOddaFJHTnDYk0JcgtFG/QceGHZ25
84QQF0NtxRtgZ2410P+/pHLZyBfJeVQxdfxWOYB42dJoPAeeZHrCE43cDsM7OZO2
gkpTGUQWYliYS4sJdzs9GynKJeNLaulX4Rgi6jFhCnhalDhYIdx7EuQXuFSR6yNP
3gyNjZRb7+y5/nslpLmziYW4PCMsYhkohqe0hXFEkm4gbn9hXagDeRApi1npESYS
Vlihk/TrkiqQFRPj16+iHOeObICiFUKk9zIvN9imjNcgNODfbpbqJy/UGP868FqW
vmQPqrwQF9QSZXQ7T0opOwN0W5ZUxGS7fUGOYIE7+Fro7wTev2ZzbqMmjcjaBteA
zITummdLBAI6YvyFaXJz5oNa0STr+akHu7XyBW5SmEZRChOJFdtds7JoOeGm4z+3
wleoJ2JNvbCCODga422O1GfwvRmoAFb1WtBK8TyIA4toQS7SLiZIrbF8IrO3l/at
oBFWllW/ar7ZqyIgIK2RIOuVi3KuRFAshTZkLJ04vCOAFVhz1qkkqaERUiGTQRlC
l2uxCzs50lmtdGnhF7LsFI0PTd/Zsek0fq1OW0X+rlX7Y37rL3FgUwSy01o0SCoC
6qsALlzTi+rtnXSCOlYufLsUM4V5iTn/Q3jc52AlRaxH42uBHHEm/IyhKJMqPtn1
Y4/KZSzY6Yp4ZSlcYVrEjSDpw5oJJo7p07BE08nbsScPZx4BdMcdTmS2E7rtAoxm
XHcwndi0ZqVoMOIjPzrGgWUWzkZ/XHt64TcWPD43ztg+3Sb/5rA2Tm/rgVRCkq3s
VcRjuDvxbNFPm2zNhTRiUo8ogziNZcB7BfFaN06WI0/9gIahaSsMdeYigX/NClyO
uX4j+TmGdGGJeITzpZwPUMbi5HYVHerQnzQl8SHQz7bad7tSkdvSIxD9AdIPgTX4
BjPLmy/cQnx5iZ0AAcjSbC5yy/NpEtWJXSP8aB3VvbZivQkhgL+9IIYnjmJ1bkge
a92taaQVx0cy2Erh6ZN88BseGlCUaqdTtMEgJKgAl6QAA0/914jnrMUljYjNH5zS
It0uX5HOvGv8vC23Zr4HWeNuOPZlNXrJf6c8ZkRr49TzjfwHWLVsmRBbfhHkjUb2
R2H83MugX/pkPIuQycIahNPcAHlx2GsRYrlZDH9i3Rh2KSWOSllhf/lGES3MVISi
EHAI/MY/q0VxyDGYcZoiTQPiWo2qDhqe0xxnc7v+o8oIgv5YYcuJ3wxnhbN/eiKa
pitRNHoNLdk8/YGth68YUEnhZ7noZeMrZDPLAY4Swu6ZkWXgKTk3whGXcCza6DuN
ZMnJ6I7NxUVD3UoInqAW1Hzk7WC15u31TSyr2jtpaCQEb3ui/f7GPpobka3AJ1TQ
fu+UuYiwtPxteKRgCmNrZ1JRfr7P299AbDChSOrBqiSdJNiE7kWI4lVaIydvyO66
KYOUjQTn1/QjlpThasKav64EFeXrRDWEJZXyUqOJvrFx6M8xy5dCcGb5yd4QgCRy
klE5hGAFArbTkiBcbH9X00gTMFGUJZgzB92PjyTMVVr3F8Ly+qr7hoyiRZfu7g/d
iM0KpqAMlv20xo7Srh/AhaybBlp1rMAeQVrch4xzvNwkL5emDp80hhATwTrrwmYV
BPlCKfHnrmGVWMXeEJlF+aWXAO60wBpJeXWCEX8mzpy16ITTki6q73mmn5Oyfrze
6pJAMdJXMSs4NWakCealnw==
`protect END_PROTECTED
