`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L0MK5PO3MkqSUk0g7lGHN2Xm4wVNmAfteoNpOwTntaBwsqO8ZvtjNv6KCidGNvrU
mdqQNi19hn5tVfchtu2I8xpLNZG4ksCHEk1UV4tqKjO4TOJlDAYlT1wTZk34q3DD
WiW4MekoiYePnpfgMxCf4I9he3CaVdWWwe5KLBxu3Non2Fd1L2qo+guYxnqj6lnL
9NZ0Jt5c44aiQwZDngRz7BhpN2fGywEpUs9dc6Dz0+fV8JMwpxWzUA7S4t/e7Qjm
XdXoVtF+3x66PsbnYZGVPdDEsD7rcPUc6pnOCi2snMLUrBCzJAj8yXdSpf7LKb6N
DBaaoeDpkast/vPIexKKA2sUX9sHIvoKSmfyPEPsjUJ8O3DXI94VR9s6K3XxcJNp
9OkysxZ63J/EKiluicf7wi/Ka+lDh+9kJ4GCI6pR0Y7dTVFAGS/rBW2SXmD8KJFx
I8Z9W7uU9nvRz+Jn3gEE4Q5elgtmQLNx7lwMFyHOm/96LLnQLiILJjTTbbrJqr5G
wSbvpGevqdhvgGbruV17xW+B4HquQuO9g3tr5mcjahK/VF+1BTkoGnORviZXNq7C
+k9tw8zDdgYNZ9yT7KWq9XpwZAFrXmP6ejueQ8tK2Vt8gtEMuPnmvdEw9BwFo1os
qu6KkN2yZzWA1peRFEUTs2RXZfuOefuPp+OlGOOwufnrlEjfytIg93OhZ4RkDykc
uBfrtOuR67jhUCRU/8sbhUBdJA+5351dySvGiirMSfavq2grApkY4O1QakmFP3DZ
Vn/5nhwXfNAoFa48AGkCttvHCzmn+BDDwyTnBNXRG2Nbx5o5qVEXgRZCeZDlb8oV
gxDahi/vcZtWPjnRS+Nd6aoBflfhoRe11DV+pD0aAJgL+E6d06ExYw0aCMB6CRyt
ZoO35SRXID1YXb9DJCZiWtGRoW6rLkQLQvWE4i3ZVMg=
`protect END_PROTECTED
