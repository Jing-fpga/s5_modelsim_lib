`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ivfAFfx0srLheCCNqdlD+lUi1xBst4T7LYdyVTlFA7Fc7cMNAN6WQQxe1xMpheJa
WJ/Wqcpozq9c/YUfslOvNMYLvtRuIwOpT2SrRzx3ffljKXX4tKpYA+GmkCsix/P4
NvVZk3McZlOsPvc0E19Ts1sBiBpzCBgGHfCAbkwg4E2oavbgCRhrbYYL4cDQt2Xj
GK7YKWCcm6YYQcoe4SNBUsp3cGPy/FcaHHiEmOPIid2tnyJsd+D8atw9wVZnI4yj
tUYCb+wty0yOkoizztmtYOfZlMnWZAi65KUAfXlPOMAt4acMISxKzwDa1H+bg+PC
pJbIhb/72KAVnKUOE9HxHLxmXruhvcRg3e2kFt/QHdZ6t4fc3xpsDgGZRZ8uLJTu
NYszJZITcdx7ST14PWrPtam5f+p20SdmN54DUXzJbv7F/FC9QFPuaSToFHNMuVCC
6iRyEx53PbZVwCcZzr4/wvBoSwEGfi1i1eyQlrVfosr035mTjbE9qcENRaFDxbTg
aqQwvAIOGhqg7mhnqokpUQWv41GO7TbJkNKfdpMTdHbgmv6ZeUKgMW9MnP8SVOJc
5HsuNpLadiSxYmDX54rjamkqpAE2ZYlOdNFL5ExuV9ucBaqQe0wx/wdS0lofAbsl
osB1rnwHLmPgtEWwfmz5vASafw4wjbRmUmPDnao593SFhB5dws03YsXDt2P3875z
b5nuFIh3j3gs0uMQ+R62C1VAGdqsIm+NdI1217KzC3ee5ThRsva1sWrpsrLx8hmn
aD3/bdfYqZiW6VslmGPQuRrWotQENpAE9HwQyiCnag7EsOybpqJZ9rjBjnH13QJS
B+V3uTaNBIsBRZYB3zP+v7CuCwejbgsrwmLWw1Zb983GLH1UPQ98OveB+7/GcgOY
46D69tXI0yqoK9YkCua+zTu4Jg0Dmp/op5M3vhZogZufpeJTQ7QSKwIzzZRh4j8U
3ZQGqBY8NxiMxxuNAxOYq3NPCZ6s1kTzJoWHufX7MQDlIpwuz8VbmZWqhNeaiFRP
1YN1Fnqd7r5AnElCoV/FqqiqkV4P/hzCNEmMtnIh2X3t7P2Z0OXeKzCj94Skev0K
kiM+372lW4n/59Jf03rN1/Y4NQJ2Myl0Jxz9HOgmMa+GfSfnzAEg2OoGbQLtq+HZ
zvNvIMXQtnwspDkFHtSkv2/8dON0TXDILjr2KcbdDM5V9KQHWNVuf1IuKhRZilFK
afm9+UkHmNeaW9m+pjQOmtH1mrWCu9wFkhIYukfsBDJLH1kyFuhfppo+vZmM9lwr
WlodIi17Y7E27oGqxnVBALIA2pJqeJslYZycbo+WbLCctAj3tYg4kqW4AC1ui44b
PVu2/gAEXbCPGxOYrv2snZb5IyK07rUNMARm92GHsYG1ZVcYHKGgXPeb4TxrJQZO
AbaHiZ+tfkrjZQ7V/v3I+NwJ9jxHlJBgntgxXcZVw+H+oFu0SzLbpvZeGuz3Fejc
/lm2vkp4l/t6kkwDOI2cPIb36cfa/8MQw/MXddZgVwj/hGFGOkJ1ylhSVedWYc94
5xwqO1k+k8y9yS5uuX/fd1o630sD7H9zRHqsHC+q9WpCFwyuOYzyUgmFuQv97oPd
YjAvqKb2296KP+mpR6ptTo7SW5Gt/AN3gJp95LRxdcz7Q173MIcvI4ND+llWx0jF
4hyLm93U62RU8IilEHU9ogtl2sNlD8OPb7Sc/rsQH1QAXub34Z3YVae/TWvJHTN3
N68ZZjzZwxgdpF/N4obyKzhifbDq6UJQW9xpiRN3HtxqVnqdvGcY1luOYiUucs9u
DKArbBV9Dk/gLDiB96ffOwu1RiHsa4knYQkmOEd0kkZ5RWoE0HWiZyGnjMRtGfFW
eRvqwsKE3qoppJ69t1vZKiVD1cYT4q06DNJYyyqonCzPY8uOkRkvdens79FCGvB4
EghHdkc54s9DDAv/SOWw7Lnt4Ng5adotfLjaX3OVZBqF55MW2gFWlMXJ2B2uUefj
BDx5h23l8X9evvmEhb8I8umwUQYVkrjFQ8tT0CSXgrpDR9oPRn3CGGH75cHg9nB0
yCK5o+92WHOTwA7DbgPHMrL1fS/LWNDu9lVZH+d9c5RbXsjS56hllZvMeHWGPpQO
zFefEchOxe8PwBBcpEdn3XMMqpQeS9g0LMLrbR3wH7OFYRC+zDsV7KwWMzT7eCqF
+n480p0vEL4XUvDy0bY1Mo0fLaooKIkKjNFObG/9pit/GTbUHze3JGNpf88YElcu
JL//a+aCy79UN3mLtr6Ovi+gZCVr8OLUzx8lpP/JoD/HjWCwmsbCGA5Jvio07Fpr
4Vo12W2S5OiXla9P1JA3Xr8sSjpHUg9EPqaEk0UGDV9uBdoduBidb+ylUkKu3Bq0
5qUSlGudMlqx4JcjnCZshlt5+VrXKRHiTZTEf8SWNGiGf4agOvE/qEglyLJZSAII
UfP33W0pGqUGmvX2TglYRHFU9MdHQRJGWLfD5Msphtsykjn1flAUqb8DSEso0iWb
eosPrhhWbpKDtOnPvQmCVRTmwc6vUTfa1cDsaYyrgjA57tqq8+kg8kZ3gy0TE/N1
5ApojPnKFrlRokXdXAnnG6k7yTInq7KTh9chwp+wibHIy/uzY0irofdVuRGTIPJH
/1eZWo/FTL0EkkjsP26eIIWJaxn7sRu4/mdgi9KXEoBvr/4kppkaMU721hyg+OIG
LleNSjoGlVa8zBby8kDLvNa0ftRuKm4nYeXj9PQ0EEkhc3xmEi8cx3bzyauoKw11
OvYoHisLepF6b3rbtD2qboFHjpV68pHY/9uWQOpIu8zySVgjWOHAgmf1JAHiWJA0
9GUoipEYBsU9ND/5UeINEygLvYTC2gHtHpFPzMMhzW7mYbFh8wAllk/BtHq63hvh
Ggcsnq/zcyAXkB6TkJHzrlfkL9+KKSrXOrMqIuf4ngUGE7PXWPbEtTgA9IrYAGWM
E4Awx99MmUzzBSwKjR3keGoRZJ1Medjz3hX9cJJuHTMBXGRZzitsjZ9eSYNUadRr
dHkNC+JIUxE5oTA4vCgW1Gr1DbpZLenPAFurr/NaNZ34MUTu3QG+OtbqE3LlGGNZ
m0cOZwdtvj0vsB3YBE/DhYxxRHq8aqWRG4jbeulq2jAqyL7ePFr70LdoCwHpxrky
j1bCQjLxPmkPdFxl94CfxWqxa9h5emC+Cjhw/QdOWxBsycUQcCutgmtWFcEHHvEf
2mp57C9NTNeJO1zu8QMatuWuoTxVmf/le4/rAIG+s2IsM3rzKgMLihwZFKGf6WfO
8/tHmDcGOd6YRPkZwnBf2Fa/KLBB97eeF57JNdMVAWQi+WhusFnVHi1vbZv29tao
cQGtJ7RiHOQFe8rqIk/ZZwYz7059f5WlHSqA61GQWou3cDORmiyfR96lWM6Bk0lV
LfCQavOQNfq5QZferguMQKSStnKR+AYvycKreddnCM1v1fAQ4qJBUFQrui/Q8x2w
xwpzZoGWEC1tCK87ZVmdgJUGqO/KbBp/yqgE32Sbxxs6PG5lEqy1/SiqLo3Xk0cU
Zlzm0H3TfsFIB+4DVpyG7xdzT3cuMlt1deepIrMrnqswggD2tINciQJnZqycO1BP
QpF8RorXy6piWPppOCShnhhVdW2+j8+BZIWK95k0zgczPz7EhMej+obEbUed6d7y
D46gfynwmFCAJ4lLfKGR3733SUNCXyqF2spBkzzujNGi34winEWGKToDPzF57mmE
10K10xvV2ngCAqUb2ZUyi87KprlnKWlW8MBB7/Dt/yGMc1KNcxPqipCLt3LX0/WV
sbWtnWILm4qmujnHzdtBHi4vgnwineufSiBi/euYm4jTTOBpq2HFRJW54/WV+CUK
i0CA3DfiKA6EMdNoVrpBymODRcJ1lu2Qdv9Jw4kuosEMeAEnLW/5QRkW2gF0wZuD
ruD4yDljuD/+NDuHh7a5INuvVwpQBu9W2cHUzMXcsBtGt7JLIRnHjEZrE0CPQuzU
OBlapuuVNWioZ9WoFF27gNqIRQ18cZRyKtnSuKc9Nt+9IHPY4+CAgpw3gfRtEf9d
uXgevNKtinO1oJp/v3vmobBPCtPqeKub5XdBc9dcteqIG4Iy9z0CujgkPuTOQBHH
griaSY/nd2xdPHSJxZOTdEN/YaRZRm1YXXqNXWq9kntXY9epPFePyzmk22exd51u
XHqlf+s5EFFyPhGr7vco39ZVadruiL4HWvGH7skutsVZTdaoQYpOcrmF7EZWFBF8
q7/LqRoETs3Ny1L6hDxOLGkITBUzLflv/oM/OmqT4dg3SL6A6a5VpHcXeJIJCusx
J/vhZG2fEHTPX1x2GyCgouHn9iLb4Pj9fBMV6jOvi7JMTnFjun7rqKV7mxk1FnTS
k+NH7bL9r/SYmEjJLZXRtVNvt8M8MkyFK8Qc4BfSvmHoVUyennGCrjwXYDKsgeok
Eh3jKZfUjrSaVbXv9cgQ8GkoO4yFsgg0evWAsRfLezE+/ohCoQTCVBzSe8nW/eUO
weJLFtPh4YBFbZYD2Hzj5R6q6dP+L45Ro8/FhB0a3Rq+0UyNB65EfP8Bs3w4bOEC
zkLtPNUlsUb2UPSjGgUznzOcLJr49BoosHREGGqjsN6Gi+X/iWhdx9eB54lUeaQW
mNT+dTcGt7JgUgY3XC8ZqOe+zjTqB1NWzxm4rbzG4nPvmtLeL618ykP8eo6fIg9+
IuSNTzKGH8AT3K6U0+lrcDxMxOSIoCU74CevR3hr7V+QVytfibgNSryMeqdGTV0y
qef/dXRtAnPo7D2/g81+6ne1TtyKxPN+lSVDzlV7AUYAL8nHDCFXgG869QrhxuXk
PGupqQC2+srmfPVJTVjYXjoSVaGvF5KMmddgZKUm5BXLZI+olvho2Uk6FoWB07nQ
qXMILiBPEUsPeRFZG3IzMIEpZI4iZWDBm8EbUFQ/Corn/QAKYh68w90wNa3TpOcU
DvFT4I8GC0CZDwoepLig5ZMUG/5V7awF6IslhjX0q/FE/ALmM1GcJPELESMAZiXe
cW2MRu0M55xsnblaBFinj5iKo2w7kvEdmcyDy36TxfTSRHyfNCsikTKVDYsKU6xB
fm/0eSxeAqiK07Iqh7n4Am/STO6IcDM4c4YIjEp6XrmT+Ft6cMkrYQukBaK4t/f1
FQS8UV2V8tPzFJO3LOiiiiwM4ZFC2Cg7HNJFuOvUtmV6u7AGOIZeyaH6DfV1JV8C
zN+tPNfJNLYG+2K4p+Ha1PKIu+xwJwPpGVeqj60GySfkFybHWT/9JxlhNoDnFG+7
Z9K5sPNUBI1SOAnuxrHKr6AuyxHvxHcOne+jXCS3YYdHQgA6eIKQUe501ymuSGnB
DsxF881d3PQQLFneIAZ89DDIVA2tH8TgDVglG0E5PJxzeoUFjxSZYWr4ZaQ77IFk
sSMDkS/NRfHi7jwfdzxq2EbTN4LFjzz8pTho0TIU/8YNVo2OoBI5tPaMz0TMUp/S
44AXQYCJq7yQYZ4EvD6ac7hKnMluSM96udkN7MkEMyQx7ZSqJ57oxSkKs0U9kMcb
W4Out4lUelLU+cXDS4L8VmTylLcgI0x6LbAACdSzcy81rjMja002Kwlzyms9D2U3
MUeKi67JipfyPh/0aJ0f5cdun2jbaZxg/REBz2gxPJc9e2W0f1hu9+xbz0uJLMeL
n2oZdOpRxq5uf0o7ujPmUffhHwKCGQN5yFu33O6/sR4unTYKkREXN0YdgUDeYaiq
ps/QghOQYb4+w7tMsrYAPIoMJ/vqjZQIsIFzff5YxUPbodaHpZdGlfuESW0q+JnA
kxLTrAC7djoi6DA9thZFlsDM7TQo2pO9aB1QJ2sYzFe3ryOjV1arG73pb57kchFb
qHiSA7i57SJbX00NMl5XyIdAn55+6KTZV46mNNA+dzHHhuRSISYvIFOPMdHAMue9
BU1+0Q2bvqZgUlFWBjNSLjTuGzBje+w1HXiHRac6qHBzWq6pAx3UVhHXyff2a3rU
lYU5VWWm/r4xR9B8asPMj1allbvYFPSJzajFhTDczodi41PCh+1mBF+rWVg1GdFD
lqUQuhmODuuIPU3a/Aefsjkl0sYN9d0o9LJkYjkQYgTtTo4BlZlWMl42DXy2XnsK
0BfmQZ7dTJMyp8FXPOm2w9GSu/8FjJZkeduSZBbUr2yzija67zjwkBVuoSceicJg
J9X142aGDVwZ/DsX2wvolquhkxLxmlWV+pw9jXWB0A0+JybLClzXJl5yoG+g/6qm
OuRSLQ4cikz0D79M9yn44w+cu7puJI85evXWR1puVF4mgZabbvPYH6GDM8EoirPc
kADdEdMk3e2/DV/arJxX54Nr8LxGmcvvDB23fSe4x0vJ3MC7TUei7WMmpufiHxwC
YIb69oHX1zqGbdBmzLazwye7DzpN+FzDO6SLZon6GNqBJtQECPnyZ7eMT+x7y3ih
JBK3OiKpBAN5345klsWqa4urnfejdkCreRttucKGH/OgC8LAAb/OAaRtQ9IA28xR
ipi1Q1r3RLRlS5Nz3lgZB1j+2MIpuw4vYClMw6FFYaSe3eMvxVMIbInqxoy5f8v2
0FgMkVidcGQNF1yXpHonWmGNlD2775o/RWHhmh/8sdKstTfiLhRatnwoJXEWIClx
9eCUZQvvsk8GjxroEkptQ6FdyP6qeVV3hJkFCSlU79UYv0oOoxleK8xDK+YUhgvr
yXxpPFdz363Gy9IhW25n1J8rCLTMdshscomuNstIZ28kK3pT49znSS5Zr+nfdLIh
+n1w6aJhXeW3oCle8447/F4cWOImphBvzq+AjVUT9yQfZr6ieRmq8m1vTk/nhKig
hzvVqDSrksFp5JsQlgDYiA==
`protect END_PROTECTED
