`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R4N76fOPM5XkUtiaHoy/dGKLiKqylKAMioueKRMnF1w7FGJ6NOx5IHQfvGdMdNWX
8pDg+qEUMSolbqWSjga/QY7GHU6oLHH2Y6VeVvENQK7BUfZr5OYa4x0NlBW0udGR
RMfBz/X5gO4SMeaBgOYuLPLKRILLsA69uyWaAr0RhE0reVr5a0EYu9pyA2JA3vMT
Hf5Lceg6OrRuHuDhVPwFEuVDnkrZ3YTJIF2RaBpf7bH1GQ/h+CfpDyAYYfefqCwj
4Yh6rL5Vw5ni3x1votj1gfYK83pf1OgUOSfdku8dvCe7J473v3B3l2mkfFQAKbzd
XqHP6yJCSCf8g5ubk2561MbASDGnY5EH81fSquEH1280yCPKOuxHFwIPcXHUoSjO
REjWHQizNcukbZSTGC1rRvXHOPTxO8rpSp/eZY56rOCfM/hxd8OzPdgwhlJNNxt1
+wrZY8btxsUavlC0nZLs3oXgeyjyOkLNCjChRbMvq6rO2yacLerEo4FugyuU+hmL
CpPVtehAtJcV9U3uBfK3A+KK1oJBlWby4QnOXrDAwfCe9fUWC14thexgp3KlsOTx
eZHYs/i0feftMuFAKHc5/8ZLGlHUQllyYLzQ0SR2jJEbW5JW7779GaeaGAO9avlR
UPZAU75vv5aP5B1qb6eezNRBIBy3RSED4AAxnNGiqaqdV1sz9wL6HkC1BHSBapoU
0dweZpgH/IWBQl3F1atPwwvdndcXIZD1fvq0RNmK9yk=
`protect END_PROTECTED
