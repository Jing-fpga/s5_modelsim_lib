`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XGk7MHhyqnWvzbkWFfohTzZ2UWqQOEM+bK0KAudi61c37F3kyoYHY3x8Iq2rCNX9
dX6G8kUxEsI46AV1zeSP1eYA7tsthQauG+JG3A2Uqln1N4Ufgz4ay65VH4c66MRD
VRsbo30VnLrp2CAY6YUQMGyYg+sszxC4Kp6+4+E0IPQM+b0K+SUGBWz1pkLCcDhK
KIrwzrJADrbdsere5Ba62Zq09G0bY2SsL8ZcWc0Az4NQVRv3OdKHh7aGAW2tfQu4
bj+rkdmHAZ0342ufqcDlEvqEMcUh9dNJa+6/q7ay4trnQE/bIxi3PiUTnVo3LnT1
56h54zq6ugUysd2KFa5iiwo1uInEi9QtVgcwvGNvrxtJVDjboKHQH6Tz7QJhr1sF
WF6Dio1Xzz2b0HWQ3Qn3Ok11ZHTNwOvRt+sVzkVwxeX2j+65uQ8uXsCWnOyx40re
HVGHSnR58JdGvtnrQlLWTV8rqciKR0hva79kZ7eb99NG3thGeIatRx2jGA5S0W1U
uPLYKjNFvTbQr9BU2HU4+wJqh0mnEO8FwXDgbbF8vADF7hh5eW/cQo7hfgUyhiOH
pLUXGGx4Lw+caOmoHwCSeEzAPGF4wfG+QcXjUqjYRLDEsho24NliM9Pg1nvcvQaw
OGcHMOegAzkG9t/RhGWItWJLVuii59QQovG+ET36eXzq4EeopkYljoWjRXjBkzbu
W7YBhGYoMjNDn3PHDzSjPzb+HuMo4TvKp/fmyJwlqjVjjvkL/X1HFWpNz+asEHdl
WAMSJ0P5v4pF19Clhec9nlIp+W4MIbFmRZPyhbIuqugxf3MEMbosSD8eQJyzekLZ
VM+g+HtRqfK9sHHip+l5WxRFJ4aM/5X481t5sNaTtW0rtgzhtgRVCQAl7kxNb6SD
quPgQDFqXCzwjKKzvSeYiYU9oajZMx+q/IaXomCLeYITyf2lakZW2iYNPofEvhnW
Oc9VHlb9fJ7fDxd43CNieSabgY8nOqcahqS1Pcom7bO40vUL8LyMsdnhUkI8pPUI
VIHOqdXKuc7re+NWTmO2acSwYE49UpbkIjiomX3XcocBeYm8wipD2UJThm7oYdOz
5awtArevjdB2OBM/wscPi6VwayES/ENgFo7HdGqedX4jO3LaaCeYC4art+algZWB
SsilmgnR6qI3/i2b1RZygCvC4GLn6sFVwCxzGGz5rCwj4kzhu0TNC9M/oV+bHrn+
in65FAYUQE+QrMSJcaWsdhY5bU0mRxtTqG4I8s/hccZ6JDXgU8CGu8kOx+T8fBxn
MK8Jfs+zmEu9BXqHg/bB/EbK3EqJSSAUaPoVJUp9r3a/tjq+w9ZvkZ9o5zxiqF2B
lifWxaR7zGpB0ML31GN/1y1mr8my/njDi6xcZaz8Gr/TFL8d0dGATcKzmP7cYIsh
j41IWgnx5DvyKnRMW2cI3z3AoPuQFosWj0R41HHn4Ywjd8VS/ajeTd2PEriarC9r
wQCHLwNAUc9QbsQsra9eUsby3ywK8Iu6Db8BszaWdiYMNjQgB2gBImuB1lmX77mv
Z0qe+uaNdWONR8gLog/7iactH65li0YHPR8VegueR9pzae7uxm4+0ypgPOSsJKZ5
9nn+zkOG9fw/JfcIMFIX1RLNXzzDgOcZFi/y4clatZqoLPl8DYe6P2516Qfocc8F
cw56cm0knE+jBWkLW1Cj5uUhBMm/cQufto7qPYk6/o248HYmYhVzF3SivnLRbXrN
mh4M1oSRmWMn0tMLaAb32C0LLiVjjh1sE/60wvv7Spi9AYPq8L5bcykEIhITzX+u
tEgC/RsVQbE8t1xivv5TQ1GLmiez2bY24kjOmdcJS6ESCwP2OvbqbfyYl9exdpQC
aMTDn/eURlAUUb3KnjsodF4jIQikdML8XYjfHZi7h+Ae0suLsy0VEvVddymFbX/N
9fUQNCmL4dxN7O5Vw20LuIohIhZPKIKSf5pnlvyKnCdt50W2BBP3GX9oPGXseP2I
`protect END_PROTECTED
