`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fTjzEznI60ShDbSYi5NjaO8yQHZXT1pnlgi2QvG14Qs8aWH+aKkp5KdqUKzWjHdt
BZPqMMaumh0mEFWFm63pYBrQzK4OXqx6FGRXtie48j0+CopKW0bDlaczbQpa6S8q
MmZGyxdgZJH6fvbnDsvmI7di6YqLxF/DNvA5EnM6WjLVsQxy7Knqlf8aGsvSqbvD
6WspzDSYKGHccfjcU0CcfI3MeKVhulPETz+y3JgD7y5wtzoJk+8fN7rOEp7D1swE
vSbYhCPnnbRz0dpj4H6aNj9mOWpwPr6qkMyqFoYhcrnhMOjJNFWul/9oUMNj8diu
GUTYzEwrJFJTUELj3XUHgI26XnqugJvTQ4hCTv874pHgk8gbuhUo7VaaA9CsD/IA
ERmKkc6j3V4QulBTf/X7uTRmmq+GFtw+gbFnanhjYfh7VmR0N5yr6uyuwo7xucMG
GS0PHrVbCI0b0JtvpRi2dlIetKBSoGWbj+IlF0bO+VI5xc7FhfdnXJoxeH4nwAyg
MtZx5vCuhatOAvcwv/ObJDzkbfHxk+NXunDQsCzXc0lpaxm+k2EpVAxDnyZF9SzB
ga2651oenHr5+IIG1TA2HrpPAXgjpbisPlsQnG64Te4BEBmkHbYfWkHIILXDYwhQ
Vl5G6x0mLmSOLhAOlKkJqSWAyGIK1V0d3iF7cFmlBv8RMtFe0S4fQFEG73MuArJP
ewxL2dOVw4lqSJhp5/5bcx5HMmozY0HTKyeAbkUjjJpFAC8h1HzPa4tTgxQM+9Z2
1X27ga6fuz1ZejSU6XYkGc8dNQ1rW0pKkyTxIpqi5zu98flxlmzWIK9w+oV5IwGm
`protect END_PROTECTED
