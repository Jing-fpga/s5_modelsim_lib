`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kU3RxrzQkDcNcGa+9ySgiWwnxx3Qn/DVZ3prQsoJckUWdbgbVX6g8JVWOY8q+t07
psjx/v7KxKGIG6AnzIJ9sBiuo007Y7zEpmM3HdmvSJIF3WMhhJWJkDUIFCfuMnkl
ieytLwulSa/mj9RYIFY7iFkIEh8OKfp9njvOEEdKOujvJymsTvu1XeBVOZ12EYTn
0EWxDhMPk6mcEpv6pm/hVhqBGburUJ6xHGohTRjLJYRGPgJRkmX2he2qJYc+vYZR
VePsD4pxlNCjghZWqvC9LL6USmbof+T0IjCjHaSxHBlVwObcPlfpTzDDyZHIo2X6
WQEtTGtrxMqSWiZSAqGYF0rZ+NON2coCR6o9PavX6ObsMcTWu31N47F5YQ/BRcyJ
z9A6RrJFOHVLkoWvoK/D2BabVWCv6VmDT3RSbvPlJQt1cqJi+S/SHe7b7IYQu66G
yUb2A3vu7Q0Fi/glDzQr0bWbZDViWp15Tx0Q5OPR1qtCvr8rualq0ZVyHJv9Er9Y
dFjyjv0TvhvHkSoZnznm5MjdF6BsA6XO5x5I/yq7eirzpE40Z6wtDFKGuIMzNZBd
vUB4VcFPm7aGstqPohuIwq0Y0YZJ5bAvf4IKV5htNVWUCTJQUnvHAVKkti6v7QYl
ih8+oVcUD7Bh427U9dvTBqXPJ0yLbJDK4G6UmgKba0Cub8JQ04wCzJ9kXfr6umAa
eKngRJN8/LZSqDlPpXCrxO71eJFyOTNmwF+NFFC4vHyvYQ5smOV5cXlJUf+cGwUp
IlG/SwpakBHfPGcqyq5dwklpMlwzShBG3sMKesVq4ldKFIOZvw0lQ5fIxJS/VbEW
zVsupzcACyBrycrSQmdN6PPOK5ZOwjYkQhdZrsnCyvWD9ZMBgIQ1T1qvC6dKJ2WV
N4nTPzbPe33KxshnxLCZkaLuyzq/8rJqPH1idf8nYpLpywAIN1GirciXiCJ7EvBr
BCT9d3bPCkfhAYq2o6C11BfzWBENgREjSfs9JPuktM7AbWjL6AEECbb5QltXePZT
j5E7x788x6yFIJYTMTFyEC3PT+BpLL5NmRUNTG0yLRK3f4e7TrxeCp80tLy68RPj
7Bkjd03eVJeh9d1BIM1lRnEq1E0+jtJ5S3Xdt1egvw7dw+ifwy/UmcaA28dtnsWH
DKjlopTFwuBh3LLkKyt/PmKd3yNToleK5V2w0Uqrqi6tv2ks1j5wGrnoPWV9mReZ
MbkYO+y6pafqFuhaD1w1ZSVqrQezrBDv5OTWMv7IclNzgBiMTWaMd+DHn7ExCx9l
IjILnZvKmbYEH3qboTRvorxYQyKewlI1SwtCUWtg98QFb7mfuyXcRwT0g8Pvfbn+
q9DZJ1BKm/98gd2wQOLDk93mMJ6i110EOiChv989IiBJTRm0HC7cWWqD5jcA7YX8
mltiPQHO6eVDnwHPi0FEZRJX03RBx9/Jelg7EUMzuthzX5WpKLBQhT+cRJRP4a23
oiH7c/Aa0TKfYAn9Afvu7FHjYenK8IQ0OLevrVWjHzLGkTfkNHQtBaLGEboDjnxk
IWykkcGsaVozpb766wJK2l4Y+4wd4mI3qO90T7UDhYT8ZUxnygbUMJacfBfP29wI
`protect END_PROTECTED
