`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QLteXZQLRMXDudLzlbLNKEK9kEPFh9HufKAcuCLPXb2EMvK1KJYLmA+aVc/Dse6f
gESSJkuEAESvh4HucpzHptgBdWrLSp7un7UuhwqEAiOk/zHVPQ12DHWge5M7bJJU
8TEVjVFoD/NPfKcQiGiBZhbPtrvwOWphGkSetUSqe0r4rwlr+26SBDWVkavaXSRU
o7LIC0H/2UxP4vJ6p+QqvXvdOqv/leM7TQFnhwrt3nGCLPD6UvmniYyAyphxbo6j
s6oZGl9OQhlf+oUQEwJ47hYVT59bmirQQqWpz1H+qGRRgqnapDJDYSI+HP2esY3V
pNCmwCAJSH/u0WHLltkkoDUtq6i0nTmBUsFIDY8cn49b9FmEAzAqEQXI38ivb2fx
oPT0yNS7HkpZjfvYVa9nlP7Lq30X/Ev+bYQYQXSAr3gxt4NDYMQbML8WZO3qEh97
8CGnL5nuEgLBAe1LFn8AJRKZOVIH6JBigJZ8qUXY4G0P0R24w+/vQkRPXlWXW0el
JlRJWTDgvnUBOtw3elo0GT2D7bHyEa9DQvPvJUnkvBqcdPRjxSJUOYJtgUWdcjS4
eiElZYzB2ngLCH7VYa3OHvPiwSd9mYEsu7TwHKZep9P4IB4SLqOc1RvhYkQ7jTQS
sQW3h5muLoutrO8A2W5zEcEKFG5s5x4o9Ukm+vJRfGqlqBsodW6vND3/XtUmc6oP
f0nh49xYYr7NbNXjkauqpPoZUTcrTK6jh2cqEotyYcaJuBugCTV+v/a9rTDltfMN
pH3fm/3GeJEIK8Ki59ubuFFhXYrAhlwFfxCzbp1pPAx8IcFn0+iVENI1fjCYxIRi
gMK+9Luq418DscTsIzeMVQiWllOiBqEppBlCKFaNg1iw6Jmt49RJ5yl0ocSur6GE
OG1KJ3bh573dKqD/v6SWr5D8KK5FsdjTV5JMeQdOm7D81egPti9CsGxrRmXPp48b
f3hx2Xl/i6r38vgUQ/byUYhflnAUcBI1FDF2DIS1Cnnwry4or7qcy2iqeYVIasbC
QuTTYBChuUTBYEFw7u+rgyjK/1y7LCYbZqIjLZB7W7Hc565qUE51JIpxjdSdjpja
3QArPjoMBgUYjq8JlfMhlSHoXX8v3Wuy8DdbAmJzKoDDvPo8n45DfBNC5lGuwYCS
iPByhv/hL2rSVt8yKU+QyzjIBBBw39egQBFPyef2Jrcc/CAU95Th7l3lDhzpqywm
jBlNgGaR3IKpQG+0R9SMAg==
`protect END_PROTECTED
