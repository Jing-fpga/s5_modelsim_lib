`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HLh4YiS5JChz2EWmuOxKfClcOUf8QZGQ0hY7p3x/svXuD4PgNZhTuBS4QzXFEcUD
qME0V0kcTErkJ8HmZR2ePX1DDd6zDn4AY4sc//by3MJdTlfsXD+trLqU2SrA4qxs
qJfrQm+f2ab1oBb4uaprl1MFodzkDBW1IdcLccw5dl6xE8rOMEamxXVceSw5U4Y+
nXjGP/cBeF/6axGgKojh0PGtwr3rEeHZWVge8OiKecO5L1aPyGsFFixzjAusLmQm
clyJjKcx4BWvLFWgOtGrxPy7AB7pBsYArEX1e9Z2q1HKpxFEbZPIOU6J6u4hmgit
8dsFRFuE1883hqTFLq44nl2mSUV0eZHNut9rD4DV13luERf0mcXI57Vv3XzjEJBh
5r9LH/4PzFHl+wJ1tV1C2y2W7/dKxS8c/erMCfHIjWBfXf6UDHZu5+UqGkbH7Cs1
S7IyuBLRdhayd/S7mTLlr1CUJcSWe6wL0KDJJ1vHDAnaEiZWqlwzp6zVCdGkvq8F
uTULjSBc00C8kdSzSEfzG6G21W/pdyf904Vo+Qgso3RelgDfBLYcl6J5SYGwkCNq
ByQxzOywBzCVpILvRz0vgIigKCP3skIChDcrHku930BcsfJk33JablmfrlcmiDN1
bm1hv0oAbRpIfS998tlJaJw4ay+2ii4TgwofOB9AiYBBtRCp42VvU32aD3FlMFvf
2CbzpA/XiPsP7+0bHomq+4naRfZ8XDWU1xaSAFk17nieGijKtp27bSj8NvSlH5Ug
yPeEQxwS1W+9TJoyt9niMjH79d8qzsKWBAob/EVO1rlJTg3YcZ9qDYSIrrmwkUv2
/dxZJeILf6KPm53E4305Sw==
`protect END_PROTECTED
