`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dFn3CBIkINDFOVGSdR8IWGNPus4ouV7DLD6gR8/2rYuib2Cx7luum5yD1MxpYuB/
wDd0WKI4r4yunJ1QJpxe2V1fkARNVr6mBnqyad9JdxH0NRHdGw3/kcn/K5skttmi
3PQe4jkVVTnzRxvvMI9IU8GKwgZO7aSibAIucd32bSPhqWBs+d48WV+h0tAapYzx
di0BFSolr3qzeUnMIUcUANIVDACIHk+MNxosroBJDxrJJpz5m2E2bBPxPclo0aj0
prD27295g+TI4v+RVIqOElYKBmEDABd6K3c/VvIsdN+6YjyBwFimmlbHqbJ1B2fa
dd3v0FyrMHZ0dOVG+/jFTzqYXX52Svvmo0rhRrX63Z3rpGdCqXKFBNHJCaw0Nm8r
/o+tHgNQ3BW239q7TlUFWkbphASygIPlkg+28EdWZrf7Xz4vafm1A+dXZU99f7LE
kpRX7Pb0BTuuxH00miDZoE9cLyWxTnSNFGOB0EZjE7LinoCm3SOW1BAW0z1qZLKV
yRrsq7FM80J0NVs6o5lcHm4zfdP0PohDircSTB+ud64lyQPmRNOHg09a14mx8bvn
i9uQ2qRmsz5b4SFdUup8bLsc01wcIOuIkrMSK0JX/zFNQJ+iMW9LIvgWEYRJWZzp
KejGqMtH4ntcE85yWacLnDI/oLl761Ox3F62MkSO5Gm6xgSrgmcqqEUnZ5bOt276
J/eGDj+QIqLtRm1pafw4GlDsOoMxsuSr2NRZJJBfx+d0Zb2QlZWqcMarN/t53OJa
KZYh+23TgAM1gexj4YjsWJmaNIwzJNyCDuvrt1zrxQLRODP5W5BuStFsqLgVRFVN
1P3ChaYjsLzsrcjEUIUOL91s8d741jhc5G8eCR/1F5cHg8/8LRpJ/iSKusS1i60l
IKz0KEOtjkCk2Kyex/mKKNUxUPvcHYHs8zPdQQKrnZOTrDYzcMN4u8HTCupRuc07
Ia3YwCM4QkgKmN4aPz3yUEEL9U5zb6jA5u1lh04gFSwRb9AeOwh2OavyOMVKkGEz
MQkMUdyAj3pQriVQYGt5tTpcyVct5umRKLBC6JWG5RFJ8ff5HhKtqYqozhDog2md
ZL+jAYZk+Ad6FZiDkBSv9gvZSsN+Y3gNFKVk0iSKhZUlMaF3CzkrexEWI6PHoLT6
hQ2EfMSM+buV7Gw+WJ9Joxv/g+J5WWpLqVQYZPYQjFHQvFQCaTPyRUbbkx3dfKUH
/FFX0ZzLyHbhsAo25EHlnFz7J8bcsLcwCFeqTdb3vasGH0LAK7jq+h7JzeIO0EcF
3zPI/HsV33nQeNbxGXrId9A8I05Jci6V3atvW7GLrS/dV1LxxiB3OGFUMrJGRpMz
38EKmRd2eZo7HrHr4g8TG7nbp9eSa6/EFDRG7VourSwTBvep2AmRsYqwmQmCcgr2
0KFBroz2hQMhDe7F/1i9d2qVdPdaxVbqyDcbBlTmLf7LvyJUJxIeYo1+fm011wbc
z4JaVr63uEnC6x35iqJIMdlDCpql2PVe06nEnwreNzR3Dnkdeyc6quJXdI5F22MF
lweo503HoQdCJrw1VDf3ME+ErBuqnAtRJG8lDFLF40FSOcTaJ6c8TtC9vn2tMwpB
vzwlOOqa+HduXSzxqrwMZ4iiBr/9gX+07uG3q2hv4vHv9A/wPrjqEdHqRytYm/BX
LoCFEz/QqWcLniDC3i5mTv69HHotLQrWff7U6j8rSbMiI3R1R5bg1D1LrwJlo5lA
U0cLFsY1WDiTITEXV4TSj+iDfkpnurrV0cjPW7f9NeURm/etcnRDDcMRcvULDguj
j6s/XodQoAuDGjJnw2mBAjmnvZtLgBRjdvlQB6QjM0egH4+X3d/09QB2sDVkK+F4
Y82FFfuqU1Mz0xxVLxIVuS3/GjoUKaY8kKT3yfW9hvQsKqwE0t56sh1OAG28aOQy
WBUrhozFVETmJgEkjGRRBnwZiKmVacaGlqRk6H+nTrGWDErHIc9bnH4lK3JJoKZ/
Ewiko9r0pkjeBT26qr8sj4aNl7IVXlwGChVcO0bVkZS1hw004jQKh95PUtZO1a6A
U8Lxw6ROxXSoGYQ7iJT0wtknfCMKuymjmjbtKPqonR9g7EIWe4SQxd0sINGOQRo3
dgu23Lowqqy54YBAtM2Z6SqBe9yPEgZ6BNdLVKOgu7VWOGu64fj/Ah72NuoI78z7
GpWkIztzGQtl9uOhfpFsFYnNFq+zzCP23zVNLHBzEmTyqPt4w+GrpTyf8XXNvHj6
yYHqrr3tte368P4Z1/NPp66Z/G69Q9iBHxjGQuh9DuR8g9BqzFvCL1QPu5dw1ATh
UtSK6PSFyszYHSf1Ch83nwUHQ+iQmt3VPE07x0BTu/xANGF40230mkOVUMc5g2uz
SClI1grLs/tlMi41xBe3r82almvug54VihsdInV5kyXnxMkxVTImiKWauPxiZPVX
DE4QF74Aa4LZCw60WadcmKxBDsPQv3HwJffmk/wD2ltpjwMrHzxlfncQUkSqZ4Mr
mNQmNmaVNZcUiL9gmYfbBVw2bQ6Qn2qrEeXm7i++Sb0Jk8rQDSO4PMWNxzbOZ4q4
DgYUYv5f+GEueoK4ZXVBBQlUB3tTxAEae4Ktp1eY62q1k5v8eYP40H+DGoRHQydI
P3ZgUg1eu+Z8b+GJA6hyjfbHVjBy3CgDUcaU0Q5yQenpEqOcztIGCR7N43Yct2eb
uBCs/Jf0AYyvHIKoreXsJEPI4IyNHmRINqCjGLup8t0Xkfk7MyQgCbvIZpkwDXtd
FKfDpYiOdNmIvaVdrQc7iWZ4Z/UrvjWBNTONTfchwP+OxEB3ejQXCig+9bdoC7RV
dJtE+q+ZoJeNLDkCWTqFUt0nTQGMsbrsjkgrlfaVHfmXhArsPfccVdq21s0BmfnM
t+E3UmnMeVWvYm18VBXJxZFL0WsnPWGt9FBmGHRBwS9TKiO3wnQhobAlB06z4QZI
NGSlc4eiFg8RIcySN/uz1D8d0iGpWRTkl3YOHAZtfQUUqvU6sVVoROcjd7iJmJuC
72RCzg75zhJmvx7797j8CAV30JpPikvy/Y7cptLy7apTxt3RZDRfeMjurFIqntqa
KxpHpEiLOOflqXQw9SxldKcZQ/ZJPJUUFfPKBTKaDI4ByAAwbDY7MXIwqz/2wjlU
PafpKFkvNWeSYXYwImtLXuPUQ0xg8B90x/gM65c/moSiEY6gddTWx9vHHLei+2qH
hbafDrK0ILeC5KBxDrhAA0cpkti1eI67lQG4w0pOJdsvvuYHz8as7RjDHqsNNkfL
Yi9ZJ2WvIi0DR7NSBwG6/ZS8N0Dqnxu+hdTdJflCu4Zak0otiG9SvoHE5KUZPyqa
XwmIPuVNy0lGnOz2pejpQf/KuCJZezkoriQfS172RE/YzGFa5RLf9PRhLz3VjdZr
LI43tYJQpDLmBHCXpuE+2/KgqEEm+Dqu8TGISCLTcAgGfTu88+PCl3Nv1EPMlKZH
GSK+owDXhLffJXG8M1nLxO3VlHZDsbHq0U8BUHFutowf50mg9aZ3OseEN4TFg2ja
eGeGIgnEuok5FtndrCmHp97j7lJhN8gQhnA9AwJW/LE8QMYiHA4odY8X60GYpS3P
9IplUTJl60KhoqNQKwug/A4Fmrv/2u/zwD9Ps90cpvocYtL8t2uq66vjOb8tERQO
LroaTiSP493OnpCCkf9TmpNObRKQ3VMHnavcZCF7QLF797f27Q1BczyYLhSMOLFn
baQQ3VySiFw+D7UP8F376Kyy428ImlT1/dSHhuIhp0LzBAotkXM73EJPhE5VEZLi
8WjlZjBYi5qWzxaJUS1MMeu2L1mxYogOV2BWWXT7oesU+MV03PTgLEd7KZOsCME9
IKFPJDTy4z43OqJgHlHmTZrrlHmspNo8wr/P2tbffuoBNHKcpfAuGbHz8y7vY2bB
5KCal7NZ/tiw/hY5A2Fv3d6Cr42S5y96xeHTJikdzQX7aizJFYOf81AQWpONrSid
I7/kH3lkZr5Kj94AmEbgyXmCn/bxnOhmMoyOfnb5ygkXNYJG1/t2bLMyWXXGTsbv
xijBbsmi2/+y2Ajv4UF+9+5kSyoS1oZvkhdWapUkfpS98rILpblbEvZBBabmgRUc
y72ZG9PJGFcndw57MGiiuHDh2CrpQvQ4x88lCPg8GsRKFFJxtc27QRl/BSGo+auf
HjMO6HkfXTvih9EEYGhUNw==
`protect END_PROTECTED
