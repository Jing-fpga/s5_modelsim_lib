`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZBcmmFQZAxH3PTOi0DwOGpA0HFYlQ7W7DYImVF6er8gOHagCjO6Hk4WwdajOwusV
qSjLYAxC7itfOJUKMk7q+yz2js+pW9Z8eQgpYNEFQl35Pue3YrYLGkzbgGYoMIVz
u74xgXQjK91zwLPs0bQnKpkCIxVjyvGC72SR/rZu9VOleMbkNPFaAwig2wLz5WvI
Z/AE3gHQdXwhjQ72fe8K+GZq8Hk8/ppIE/R8VK8+ffJSqstbkDPvsCu8+b7Sb6xu
UDpn3RsducvWCr5Lt4hkrQtQ/cgyIZ6nTodM1WP9jHSeHevvp01TxxnHHgeYCLdd
pbcw6iq9hfz9Nud/N1EL/wXdH1DgsjhWdQXtZT954cSukfD0hNfPbyHdwzlzVipf
2d4dG6pszyPzjDfuurHiqQW5XxzjV0UMrH+WzLF7t8wWsi6Sj98HOnPwQtVBSZOT
rSG3ykGzj7qNs0nXuuIbTBJkvxfEqIEi3ufcsSwYI/XcXi5KNuWVAbdUiFMBMOr4
s3GrTTfGQh2uH0j0DYZPxaXpk1dUDAnQmfSVzA4vBAveY2srmDreXkSVIwHrtXgV
Wx1niCg0vkhChPfYhuTDliO9DDEfGtMK4blTsZUSh2iHOAoxaUytMoNJ/mT/gpqy
/KiofwbLlPWiCvhhIWgH+K98Y7gEvk2J1+Xlm7e+rPkaruviO6l5dwCLSjet3XqY
OlOL64OVbgfvPonF3fXkEQmbALV0k+wM1oeNPP1/co5DKFBQcLtBG62+zRUJ4Qyq
hIEeTQGOtHqZmbdb01RVrTfwQegsnIEBe1VeyS+14QE9r9o9zQg7DT0GGrrcf0vf
caj+MRoZWx3ZXr1hLziboQBH6dl1df5n7xic33yDij8yZq/19DeyFdRHF1lilZM6
r3W0sNputuhMbiWaoaAuwkzwBLOC+AjpEzCzVmg7ZfM2YoaKXprOpNumMR8mKrXV
OBzGGirvk40kLW0VklynXDxeLUwmI3tyP/akexOW5aHx/xA+x94vkiEW/+nwkWAy
G4S1qD+fd4nePpOK19yr1VCPXfVORM/Go+NDvmptH0ynlvqx93nWgee0xUVr+G3E
r3G0yQv4DkVLg6y9keKX0PsxwJDGAy4Jhm4xfecu9gdnNnoLvpXxUDL1yPIK94tA
fomRzB2M6OjZ5vRfWSpBAN20ogClrMnwFTeM4MR6k0cMoBiT9LyNqlnzSXCzNlh0
f943XdmgnQa9Cjjx/TLs/cbut8GhufKx/SgUIoakRPPLjIQArppuOa3BZE9JTKK/
WqYA94AgM6j2F4zLrGYyeDBirWcmfBPVcIWFUyRVTV0rHVcYuhWS664qcO0eWPrM
kgnqfX0AfBlexPtYELSt+LYjbpeQxG+0JTO+1jnYtYyBF54v/4ttNfqcLFzQQmNk
A55PeREgaf2k99ptEKZkeRCw3lAwi60jwpPNPLRoBHbxPT8J+eyKc06J39PeLSj8
pNZhQ3KNdKpbiS+XBGUXUXHihki67A7p9/mswrupdL+ytEytTL1QdPU46jtjUybf
Sd00biYSVF4YL5SGEvaxyROrlZ5HxZA/k1iey4/FrWuShalMkGVkmI6vdyfLIafl
/95P+E6hzkT4vMqtS8zjq1h0YWvnVjkJ3Pte+rKKGoZYeSZqGl4noctZumyLe6Wx
YfvS0EVqzg91nln9CV5CZf6BcnBe8Ta2l1cJ/kC8atSYWdcYrPQWRcGOULFr8QEH
XJ29OPlpNf5t2jS0pLQA+ojOTPdHNQG1y+5/fRpI6IP8ZWzdIAfBkGRzYe0hDJaI
B9UB0B+EmMIpOlVIrrSzbUY+kvoe6x0YWmVBYIVaeFjjBr8CypjRy2tGycC+lwkh
Ifgk09lgd8RMR3RCtwMbyj/TGDCfWOKP0RUmyTnn+oG+fon3+TFTLwny9KrQTv/n
TqPz4+At3bqOkogQkh8ZsTd5pqY+Uf0jyADVhethSZHFiy9ljPqSDuGJJMVSNvfK
TGA07pzj06El5y/pdnVnP7n2VffSlDhwUnl8FPTI6B/IB8WbdxH6wZbqZCydIuZg
V51UGcfIGW48htfKs6/5v0ykGrASuF4LbgYbXjm3ULYT07k6D+JSxkIMSwhP6U9J
LqkJElcHxHirb61TT4hy6T/Hg8skDgE1e1vYufFQVC5ATjfkfzjpL8Lpdnj0RlEl
nvNE9FIPoiZqAlmME+lHdJypDxOU6UCgUcod2ykv3Rp747bgZ0SuHGpFz9hgYrK3
dutZjy3unBbt1KxI4SG6Ch2iGF2kpdLx9WxfudSOZdnOY7/G6nne+O3sTufDkqWQ
1G+uji1xyFVcgBB25z/5mzVd4YhypkNyhtaiWQUe+n7u1UefzvyDySpZyWiWUB2V
xOPk5SZVSkDWwYMvHMk9v8KuRY4QDmSwPGjAYFI48QQ24Qau/AGkJZJ76EUiaPgp
ws8gF0Kb9iqcKHgPvygKbSYkAuK9tZSXfEo1b/iLP1uBjVtE68VjNy7Xs45nm/Pu
gM4kFKU/4yLtAGaabgNlfU4zGyaCoh/Q+C0C5J1dpfSLUEESZUKytcx78e0+vY3B
/gaEJlNoCVtuMow2ycYdNI4J1qkMB3l4Lddr250ZXGp/LqcI7mXVdCBBn9aVUILd
cLmVyutU7GfMyqBZRpuFQs1lwLzP5aGhwje11Ewvn6oGKdMu0H8i5HZUgBwk0bgQ
YyitbGMU3qq7HZ8WmPD2sUEJ8+8dOJLZ2mCyzt82xl5rBfzooUcscoDg0gSZ3wJ4
m9VdzOsv2HY9IfWXLTv42rfx0Cva8ni+IoKMAZVHzqGel6HR+AdxHvMkeanHE2Fa
h3IcQtAwR4VyB6V53AyIRavKSJZLeymr4HYkh4R7aoqEvxfoTBtAeX87XJzo/ju1
VfBfSDneHCjaWDUkaRtjxMZ15M8jcDktG8AciZJ0uQBcIrWacgDNMr6uDIYycyS9
LM/oTrAslp1AlkjdfTktumlMBA7CB26wQRCEIFKThCXrrs+eLUcHbpTeyyGJ0PjM
fvd1WBodqADQ6MP15siqYY1wy5kdUtc5aB2umd/I/GuIZ5Tn7AWjT2bG56qyy6h4
/ZlSvko6hlZQ3mQeS1p/nRC85MYVEOXbVvgqp+dmMkdNaLQFb/FTsF9YsE56Ith0
WPHrgdEzW7+Q0BRfzZcOpDIlC4H4kN96F9B4rBTGT6Avzd7BXJJ3+Em0imHxM3/B
T4btNTeEP0LYs0GIFDyM5c+wvGN1fJZJciIF6AEon3ezYfgWAe3Y05NWgg8bPIOG
SxA07VCAiCx9yydZCPDjsSsO6zL75dok3k7A7BRGoxmnZI9JDw7mul821kqCdFgX
7GaGfosLN0iQxg6EwLIsoty7rrXwF9k2N1GTdcUh72uT+ddqTOhIojjjko0dVRG+
RXGpAOaFuVQMPqLoSg7OrH+iA64zs8OfhVSdzTXcx9VoD/i9NaQIgXta0MtZwq5d
CYuY5qncA4qNsdLVQS5IjQ==
`protect END_PROTECTED
