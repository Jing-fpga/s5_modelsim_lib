`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gieiqOxi5EI2+/Svbbp3bt0Ey7AdI91NwwN+kRmHJVc1lvDPFjEOuedtk91mBvX9
ahhxYYCI6BsR50cRn1ihN+CteEuqOlnxugpezQq417WG5XmEkmPYMqhUTtjYjTFh
YiZr3SsQsRyeibWIjj3LWGVkbuyub6lqoZ9xkXM9BmpD3WagMTpXeS9eNBYxUaGX
fIVkB/EcERkqdHS1fikK8C64VLpK5IHksMD9np8qUEFKPLF2lfSWxv075f55jUBc
YjmAjtqKWGuuUboA6hQ+bqlpzftTEX7yW3eIWCe4dHmEem4ji3nGLHZW3OyFZ2GE
HNiwCr9OQTTVLv8APISbjq1nB7ZZUzm28K8m70DBkP1oSye4uJ4xVzsYQKp4YHO6
PTR4XYXJZYzRsEEEkPep0O0EDih3UTOGxSus33hHGPhEoKecaflDyB6YFVv2PcQq
ZorFfScH6VHuaoRmu4k7FK65bYecuHY4kMdlU7XSvF38DI76lvz5xrGakNxOStpN
3HCpmGeIi72jlaCxgb2qLu5d44AosSEAW5fcPH2eFQlUPCtDIk0OgECgVm/4Enze
eBG4GRVC+xZark1d8semZJJRcYInhqLNvFdJFvRhBB4L+iHupcZ6vlYWFRwLTPir
7e6Ke2nZYThd+PwEV2xgY3LS+MsAjnhd2ZmjiV7dUr4H12OtH4W6edcaj7nVKhiL
+EdudwSJjN5yihCORRO0o1yNZ/diGE/GV+5WRIYZpDKOexj6m4cqDouZEO7K/D8j
VCyEIoJbWA5oloOdpejrTqM5TTQe1FR5HIyJcAdMISDUYTCR5i1BP/UTHWfzK202
rhrks/L4zh0hcM30SSWtYMwG4x5hjxkqNyueIHro7SdpijYCBvz/jsus3cJIVzmU
pCf/tEFvItY2KyZQn49/L/TFFBWoPsHIbvxC2QfP9nd8G5jpzI2Q4wU/YUq+Psrf
NNLZFVgofhSvJJCAlgom0onWCCK9npn6fKH3L0rrb+YV3nuXj4GJF3e7yArTlBhH
cutyNFlGYeTvXHXyTa6fBUzZrvIQkkEGdzD/kgyuLosoIRnFQONMfx/92Fli+w++
FavIRDt1Gh71gwkoU8FiavjIBI194cJxIhkr3xHaO86OIhNRCe+uba18Gv7UMRDq
6Bk55OpJLxsddvBxorjCc/SrWQCYlAw4vCvcbgnJ1KJ2YAaXfzp9ShNgKBdjSs1C
ZPKaJEBfIm+lF0+H4qhiVEJ5YaKE+OzHHrm3cK5jDD4Hl9N7VSwNcUmtwAtj7bNs
mX/tTc7puoni6HzbPcrWhbeXpUdvB0p/wSwDNUtz+GCLCNGfPpTn8iUw87lyJ/60
7MDteCDG4SgdWY5yEHKjp9juY7ydIO5Sp7xcwGmDpe1zkpKZehBaEQnorx3/4ivd
muJduP6SIOs1lbY1/+ybPJNxQOrehKN+z0b/KnChyYBHwVzAJzqaJ8LOJk7TpOGK
KZZ0PNAya/HjUpJk2elSldN+v6e6U/0XnKu+jNazz2xORbZjrDaJ9G7akcg754LZ
hEjuc7kyfTrhlJtj5gw5QKMVJehWfydwZOyvNZfYdcFE1ZPAclVARCHG2tXOKvoj
ntheZINsy8rBQo5P0HVY0BnUNsOOxg9N0TArqrBLSmWATsvFSIpVYcJGBSgcgFWP
0kU7REYrwY2Ktzgz0a+oTg==
`protect END_PROTECTED
