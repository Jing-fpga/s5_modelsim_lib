`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tc2xSUAYm3X9OqTI8QHqlXu1BWJTFfccAeMHCjxvy1FEF7qBxi9Vmlhw2ePoiTqj
Wdf8omuegHRwXpusQ/15wV03ygCLFNJqksOZgYCml4mlsHH3QZ+4/xbSP7ZrpXU+
6Ub1XilshIbN4q4E8C8SoYVr7/QBnBJ9sDyu/iVCIVJmKvZXIOsxdewn06a3CZyq
tppgoI9Qe96grOx9X0FQr148tzKBfXO5OZ9wdkRH+Ohzr6dlPfX7r7dhrmrTWgZ7
K/UyG9k20VQXIDkJQbgupEFqNieaL2dew4TYz8PObnOhevtYNXW/iUvP2h1NUFVL
Kz0WmksX2fS7+7AXdGzCatlMxzMIiz5Nzjq2LOmKssO2/WmU4a9hIJqTznmDpvDQ
rCo7G24w5m2Xn9wpYELz71nHR0esolq3Rruk6cBRSTAld1+deUH0wGvluBJCGz/A
VTn713XR2qFoeiGu8B2tg9ngM9ip2lvP2aOltTcIdYJOmiswnwDtXLC83ST9IZri
UUqxQxrkR2HOySwqixmVkhmHLGMcnvca1ArvSrepIIIkbyqrmcS6jNAF8PC6g4bD
c903JqPL4Pel0O5ARmLsyGf41jpeh+Cgu0pQNW75eaz778Zbyl42nJiGWtbVw+oD
4Ln5cbvXApf3qP7Kvsojg6mXPlpdg+2AJE6E+MqCFv7PJBXmR10EIH/CPB7nnDSo
abx8Qx7QryB3GsNXGE8ONDTNrgUbtCYJI9SMjbfzbhayrwrykLUf+olD68JGZCD+
RxhL80p4YIyqqWzZP7pmK0kzM8gRhjn6cTHk4GMaIJFvXrdTRiNTfkx2sJnelSlJ
w4PwTdwA5iVhYHwJBednI7IxWyMmXnXvZVSzn2noQ2DETowl1mr71Dv86h3f3PWz
fbrhqUDSukBXhcBQPf41DkagqLQ5jPpHSWVWE2xiOsOgTXD4OTosdiodIClPcJFA
yBcVD6/VVXJHjsA9QNv88ahQtkeyJkp+yFHWxV2+mDKredHeo9InhwE1T2n6G3uH
vZ6e42Xk206ZxZd/eCkqldEiYqJuTv5pMKqa+WXr338+CQuxBe6z/Uwcs13ttM6I
A+2QcUXHvgDT1geql+uSXkK38Lb+Pm7uo/b9RAzW7PPIBlXnUkq5W+EInASNO3sT
BuBisWXq0UTdg/vkIngPIYgXPm+yCjdD4Hhld0kkb7K6cu6xCgzsXHB6y7DedEwf
d5FKTEoqLAB0Ec475RRZA4pxUBZw0LquyJoAUwApPTjN/t7it5zG8fmLBkNKV1iY
GRzMFLo/aQJTC8SoqSwT6oaF89tBwpUg1IAHdI8qMwx5Nuja9PlCY+JLnBb4MDxK
sZ7NNvU2AYBmevaPdxNaEJVwXhm9WjSSfdw6Bs2MBaTqfHXGpOFpZgBK6Isjdtlt
rJD8ot0THVTs9w7TDaxrGApuVigqCcxpiSH/oyTpqQ+U+Su/ZGPNSzavc5WCs/vb
cl98VgWcRamxLVspUvYQudN8g0SiN6Kn/99587zoLghhsLjpsJJ0dLE99gXj/mjl
jq/hHC/DbzH1DtYBouabpedwUXqFYDmraKMN9cpaNGbr2NkmOAXmstI8Nes1MR4u
423bkMFZLq2jf2uqagwbQV08TND1wj75OrxXUTB7FYO80Uj37zDwRzJOFZAmG4A8
myF75Pj+chBflXktsdbM57AOCamh0Vvnb1JhEy2oCxF4hjTiOJnTuoeUWxKSU4a6
jXFvsG242TIdC/EgUvAgl0XkwnjlnVIVZt0HHhQXb1zdjLy8rk7tu0h5fuJZjbOK
oujWXl9vAjJGwkW4u9V4fccrt1+uMDrfgaVHmkjVH/2QVbGn9v0VnedhTkxhLLws
Yth/GmvpMQtaZbwSEEgpyKm1cSvFmBim+8JeIR7GAB4gYTOUFnRAfC4VkW/ZtFwT
sCGa4/u8EEjhxmMZWp1KwBl2edx0n+EadioDu6MfRvcAQmbQk5oewvruyC6yAPyp
UTBRQ4IWKR9L4Gt71PvOzbrbahEaSXrlJkrgoJMqQ3D2bNABCZrMUubv3umuer7a
XeMDEZNjVx2bMOOL2POI020fTi2hbAsAmzywgA088VEy5O3Zd9/owl8xOwVAPiMN
d9Dol24uFJItQBANI+DpC04ZuQZrolGzsUg1m0ZxullllLnMWBpKqeL0ZoRL8ZnB
rQLeps8i4wM9XpTbIk78Lhnk4AMt5rlqWFGoFtYji0S7rbpsLZYOBUmN8MyPBgCq
fm6B3wFm3JBWN91Ssdff3qo0TugGU41PdygobeHWvNP0wARYeoJywe5lvau/xjjP
Oe/ufe/vlSYkryhwMqucOaoiPyHARO/qbw+LdSWDL0nAcH132F6sztGZ2UTElCqu
2riSkdhtfez5Pd3CInD3eAiZo5BzH2t8nvZFbiEfVUT6e3zKkcd+QBVQfxvaLECc
vxjida4Cz+PNyZKANASLY+B95kwly8aiOJ1bsIVmuhxwRIwiiK+qCovc3KFXYzqi
ZeGuScH2ZYzIc95iediTQBj+DK0bVlOUefaCj8VOy4sNdh/MeGqftTQ16JJStgVQ
7WgGXkUtDy1DfXpVki/AFqasIoDOIshKC8ZVEFRmK1psTfnpENuVcYKtW1FKTP7U
dVdQdVdqxsrW/XHtjr1XKVE84CDFElficQUU6Y90bQqmCyd2yc8mLrJLQ6I0vUJ1
lcrYXsBaoso6LxI2ozDRcNRSU5JD+2kfe5XOPSavHPaFLONmsKfnUec4M0hN4bqm
f+fK9wd4bVrWcoDA1cgSEOPbVTm+Kl0Fu9uBvnBgm4OPruuTjvIguEB5Vh4DSVvF
lNpClt+niIyzpKRxXb3uMsYqxMXi1b3rFHfJald5o7VYsaudlIRjrX2t2HY+8z4j
wZPukquI8WfADD/NrUnUorzZ2YwTzop6Roeygh9VlAFJPMJ1G78/8QZHG/2F8ws6
sxe48UmzQrgJelDI+o73adz4Q52u4dUIYKId4EBf5jiC5vQPeu8RP5+TCzKBG8lO
kScHBKCvwpXSjGNynVtjsqUMukZpyhAov2ddK96yZ+vypyMGw/p1kDsY/0rrJcXg
pt33yxpN77/oe/wEW13SXQu+E8g4E6XIGhVj+NWMtxf+oDuO1OwLAMdVCrLkzSKB
FZSaxQEx7NN44X+0cCF7MG2iVob/63ZvSupKbYUHM986/y/7C60c+ye7AU9C5ytF
3rfWl9G9AVMtMlXcIj3LEWtriaCTrpQuOC0k2Pr8+eQ9StUxGH6+H61w2Tu9bnqz
wUZbyKTqIRnBCfOMr1Pndxos2b5U7fJ/7qKobwxYuH4bMyL7b2SBzdAxN5FI0QBi
vSLsBn7LLkk/0ESYZSR2/yDLrP0RGWXg1Me7H9DL9Imt1UeJTRDjBa/YDqG+0Nxl
fLaWmyzjWiVsnt7DSDSDYyI0EL/uO/Q+FhJE31d3A0tJ3B9l/6EOHNu1u2fV5Yb6
XmSAsFbBnM7a/iSHiahl6dN7fmfVoFgAkB0Gj2aThrhKtxRTiYaP1OnHxmObC289
+njINmQnawlMIN4UV1jpJY/nsU7crzVzyeENJ64P2DXfu7Bcurc5FQedzTeONF4/
kbupIr6kTVU5RJL4hEu8QGCiLW1U9V7NCozzSX3+8oXX3NT4Ol596OHgqzBQZ5Rx
hkj6FIF9lYyeAnSGL3KLNv6ueMFXnCkBmVBfzO1X2itLSRi+Qp2i88qdF8voUQAB
9BfIqwPwV4OTtfyBaoTzpUVDwhRNZO1rGtTLWW/7Vx7omtIhlRfQwO0CkSJeHFFP
5EFgH65WOXOqHcPJCscwhU++kcEBmy7znKr1wmxjMTDDzf0KPTDAtua4zmDqWdwe
Q3P1OV116Tio3aF3yd3X1DDiLz+1Uf33a+dwzY77749Osx8KSHoiNbV06oDWvojt
QyDDXLQnPNSBJ1Y662lXj25z7EZn8eY+my6GD90Pi5Lx+ItBS+bWMKLmaL77EFMG
PEc+xBDWnOeZnIDYculZjhn6xMqqekVGcg1ZFdOUbUxJB/IRyBi8TX6U1vVPe/We
iT+Urs36/3hCgfMrC6xxmBFhSb1E2AqIgxX337r1KfOE9oEXZVOScxpklu95xcJa
egYa1EZypu1dwgCE21YD8GY3DtUn5Qj797wpHRRoLlXXNKA2NLVWK5byCi1gj/Wg
VWyf1Y8+BorWW8YaTW2Rc5Bh/x3c31acvwrnms7kqTow7LXYOhfEbORB4l3YHdnJ
+PfWzMkMfoNyFEjDgg57+HEZZ+1tb9cKCWUEbu6x+zr/N2rCqsOyYjW07rTRgNNz
DaUT0VB7VqFn2nUYleyiMuM9m8DmxTGkGG0I6kpzxKdK8BS7fT7zDAA+GXCPXi69
NZ1YNRl/+ugLrAaBfkZoZpD9PGl7fokElXyfy8FMPFvTvjemVnS8wQCBox8i6EXu
eV7u2VcpBDTlOxUP61zkoUu5Ob+Kz8bIIjLy7KYb0R4heO3LcFPACoYH+Gsfmqse
tZ4KkQueX4CBfOqgbZpslFqJOEh8Y7G2pgsT4BuO4bxGRvB3uggDaBl4P+0VzZ+n
BjwN9jLIW5aq6AY7yrQEXJOlpwO5BZO2EHjqorMGL48SQlQupQLnKjr423f2oidV
2JSFm56MPnzz6qv19p5ijfiNFSaFmA4+9ZNn4ggBTV9ohl1Jlzfs7T2l4HhAQmCm
YDaacjuGui0hEsRCzSW1PZwgw1BxmT63HJoXAH/ikSFFu31766NXpvhj6Juf5oC3
i+2NYqSfdtKyfj2xMp8Kn3xFlaAlDU9twjXgBNvNnWlzzCMRVolYdE0a4AaxzMue
LrxTpzJ/avn2NnFPqz3QacGERpFvsaubbofrePNN1EuPDg6APhpCMr2u26i/CLfn
J+wE83/Bg7iBySbvqv7o1n2i7rxAzSb9CFmx25cGtbEniVY2zLdX0TUtFIRHTiJr
/28t/3ZEcXKHhb/eHkDE/9qB4sKKteZuEZAyWkcRfyekVMEegTfmI4cMcKeuYwjo
t7cErcSjMHQyeB/PX5m2XpKD2fDSF+N4Cy7hrZIYy6hJVNL1nedTf+JPXGTZSYbR
sS3+8T0hrQjhX+dCBdlQbaN9gtmMx9siqpy4qZ7I3HoP2OrWFWU2jeVUCCQ8S6O2
t/oypng2Afxk8bnOm7X+5S/ehvRFGDQrC2S+u9vmD7Xxfg9SNXzoSgu8Cr0i8XRO
8IgatAlfRg+Z2NHMelvPGUF5YU6bas+QzR7+YWYtORuvvc7ZALdNZ/WwwZ4s1Xh1
YwP3fWq12q43BzlXEWXaPjOegds+qu2RpNULiXgIndRumqVJpFnWKsljZGXr4Zrr
gO7uD4Kkcj7dVKXa46FLrCct6MhzlU+j0+Y1TrwZEmZVXPEpi4/BeRvoqUrz95Kr
8jLoch3x2eeIkNqQKjLqFM1+nqvgtCcN8ayKoMUUpMfaUF5slfx5dcixvOY79iju
1NPpSEujBWCzEQ9lzHFArAddbevZh9rUijTnybkKjD7JrvxKbTNwUxFAHLOqdGhz
vse3XD65mGjrv1/uLILYA1jgleA79EP0iU1LYw6pRr+sXDHL0/kA7PuKTS6dboDS
TCQNDtpWx2C4tJVo5xYHCKhWzvBkwH0x6/TNq32aFnnrsbwBIy7P9DqzuvL9AAoo
2AdM0La5uVZ7CLxs6m3Z1Emrx0ItIqKClgddNoQ9TADVvtXbMHl1hrBAO687M9aN
RNQ988Nf5JJiUGi+rXCrZTfdC+02X3DMJOMF439N8uB9ZmJ9t8kKmUwBv4BQAUwR
cr7MHncgDjafAI9taa5HxDiIZshqbHFWg9wu1Qe5IEbmARi4KlTpLYgsNBN4jUd5
htgyk7Qno9KacZmeTItixCA0BiwQsQGr1gij6u52VH8jJj7YtJC8CpRjAWoc/WRY
lJYnUhKRN/xENnUs4jyxOxZnMO4nstadC7lMBHxTnVlPZepqEI0a4CsoBOYkzvWJ
H/VKLCyf4k2OsHKLJ9L8ZI7StcjldYPJC/V0uA9vJ6MW1lp7nDT5v9sK61tE1qny
dYqMXEY2F5FGM85bgHOcaNjcquTqy+bJXnucFSxnEd+QrqlSg/x57F118MHUovDD
ecUzO0fHo3QlL0+d+WMZ4RZx67jTe+kY0+avlepy1wvZ60JeK/E2H4HtyBIV4C1k
Amht9OSVlKattyR1Geh9uMoeKaNTop1ioM3APoPHVLgLh7GLNkq/z/dHfV5ETjRU
UnX8RQjhGcb8K37x+pxVP/0Vu8EmPCeDwfGXFxYv/uO+r7xpqliBtVH1Z5OgDtHH
9epRdHAVLZY3d3bQZ8c5HGCNn5RfbX0qVYB402grpXQFMYB0MTDcL/CbnOdklpfs
E/ZciPqZKdSaq0vy6YuC/fnQxZbxM/meezwoD/kD/bfk4oiVmuNipEPHZsz1N5Xq
iu4ojoV4lU6rfB4Y0L9UGxrJ8uXM2Hah8daoFoqiXNjDHpTMRRtGUlcTV4ivKqNX
KdIjUUlksaNujZOxZ/CoZTQCuuXDMX8kl8BYejSyNDQAZ9fmkVdRw9ar8j4dIqQu
+VrT0I37PzlonWT+Z3dCCVhGSulUi0qP2XZYERSJkQSgPLmuB9HRZEU/vi+lGByB
+AhOJPlZUJBKuDvkEzdYSNQ/9srh3wIp+iyIDyLIMOGH87+sNXOBha89y6Ktappg
/WKgF0/nHMzXVMq5LgxCe6UatgUrnoRGUQyRYgLEggb0GcXk0ZXkrSp6tcDw7979
8AF0XjIL8inVS5Libw1v4qp8CzjZLWs+M0Gq2iCB0WyFjJt+Dpbi5e7uxm+EFiGO
7nvKTRaDh1AwG7A7TrocZuTJq5IJnoRbUYqQd0BQXsV0552aaJMJswemmgoDA2CL
chS5h2T1gTTRwV2NemphhlKBIpILsx4aXZxnEYa7Z7/lC7ba05itNwimblcM4YRZ
koHj6I+m3YnW9kSvpa0iKP0MwxA37E0QeKV5FBuCzCoqN00ExQqwFpsahhN7eDjY
/MpzzxMTh+WrnwWzTDpBx6TKOFgcKy/sIGCH/WPTPKWaUOhkJtR+DK8RfJF+ZvrO
LN3E2E7QDGyQZi50hmH3KmWYujttVBRsvNqRdFlBmdLB8WhGhsedTF+/T21s65BL
qq7RcyEjv7zyLFRz9cC9DI8RybjjvwdeEFYlKEszvpQ8d6SgqMXo0oaaN0WOCtUf
tBvbxy+IA8wBvmRYFFK0gIqznsZ0cvYg5CsxPQTs/jkM1O8shbIV7cPYtWMXrYG6
N527aY1SD6TgJjXFdpMVWfrXhhnPOMFM5wx8tuYG9qUM5Hr/eY8rD1w1HNLtlmwt
VfTQ9tligIjAe7RiHl77p+aH5sXIlUW5C9uxs8Lj+UFN8C8d0LfOPofdPMj2SKBL
FbCIJKcArKDh95+KLwhg0ByH3RBlUj/9dhZOATbcMpoIAVqQgOled5j8SHFiv2eK
fNjQTWTUmsRbodwYH5Rn+wwaFnmOG8X0ujgitiCUNBiD8Pj3q9d0WnJOhvNlr5KO
IEsAeM1RFIGQeEaAhjeNJnEixcQkh0x1XIm1IGPt/CHS7Z5cxakZM0mAAfDSD+bm
zx9u7+z6gkcWubrrBgBAQXlnC4tg9B0rWWdp7e9PIfXCW5Vtp4OvV2RiWnLZNc5X
Usiz5CGrRcb6yY7Aue0d5XNpQlurR4EneUfh+ktOXiJoH+RbND7fE61ydEDlQaJA
JOh7VXxcTtY8ocO+dsMNhwjepdvOaLBZIIGDP9hcatpdIo/SjmCStldBzN2OXg94
ZrKGJvmrvRevyr11cc8N0+qX7xOPDe6irmW6pPrkf3+udxiQI8vGT2id+bj/aghj
JKyQgnj89SM5tkaZH9r8XYZaogNmGWAI5k8XaxUflKNJOyAC+cHu08obcZAUOgr/
7TSn85vO7ALd1kkZswxuEdx6AQPxDaibt6u7WpuDe9qV/ALZ02LXCVR3gPb01ona
WLa42IdddG0PV8u+zM9wHIGVn5/1qYoux8jG+OaUP5cbXvyt2Rb22mFBoDxVEIwV
jhJf4cmS+y1JBDaMiEZ4eMo1pNdFL76Yc2JMJBlBXu0+s77bD/JKLNpoEoABAKMu
yVi64VeXkJU+cqDDtc/cw0nhVWcC27dT51ry97hzjGB4+lsQBhrrFU2W48XQ3igh
YopZnVWPtmQ9O6+VvYDTu9k2rcjLYslfVwcZZjCSH3u5YdP2eSncavZdyvS2t/Oq
R88gF+vU6rc+egyVlPWH1yHdh32eZg60vmhxYO8aD9h7U/55BUwByovmk7LfuQGJ
vmYgmCm4sYNMnTXs2NBAc7Oqag5Ft+HBwVROAJZnkf0w0sDaDeIFjjZzWXf37s67
Du2yt+ScbBilHYbneRBq1WBMy8xACgMz8lCyRRtcz0IlMh6iBOT8wfUuJAXQTvpD
mSvJIhiR3BF6YlQA098PMdmYPTHQpehyCJ1igaMa2jL+ncJ9mqsalUr3fN+aTd/4
MspXLqMPNDdBS0H/Qw2QZmH0tEnLFtAshAFgT/VSoHhkTIYqY7/J2g+qJFo0wf5g
A4/C+TfBzJwxE/IBmrFnXKmbPjBpDtSZt7H85dCGkfDSNBBngqs5WhxKDRrcUZnI
v6/NFAwudHNiI81apTaO+PiiQjaKL9xuhXawuquGsMqKMTYDHLIk24wf2UOTpugc
GEmb8nyZBQsfmpNI+znxL3kVa1hf8CfIzvAqqKDGrH+SQdzm6yfloW41wzaPGILu
cfrDRzDS8H1yszf0GYjpwHXPWXrEwVcHcf3cfkDkdUrfu6V/4ooyj6X3ezumtyPi
rX0EhlxujAvkwdoe6fiLgbNkqCq1zQ5lgbxEJ9qNZZdw6/de5Qso8kWacL30UCFl
VMehY9ficrZPyhCyTup9sCdtK69s5hjH+mDnUILFUJHusGe4FkhVi2LRV2Tt4gbk
ieZYZR0herF53WOfDCbTWIdRtg42gf6RRcPr7t8nOIfan4gYXwpf0TwvjqZxI5wD
eEMY2NZxt+uUoaDXZRzRHUcxl8CCPXuVizFI9QHgPoXIAlv7x50dS6co/sUbD3PM
bkRY19tkuqwfAO+FUnbQLlGF00f3QCsLvlw9GoqAqik5Scy32cq14FIFKtYlNOET
TpU7jkKfM/xz0TEXGf17+F1yHxGaiOCLlGNtwwxK+aMI3Lwf5ffWqZkLgSHna1oq
ssl6p2n+OElHfNICspQ5w/fECsxe2Jd1BuhXdBP+4Nzq6iR2q6YOEkfKKPa9CAJM
iO3pnQXxtu3VTz+7fhMVGHhgn3EnF68sBeYq92tycJow8cVIfNXWiqpxk3Dt59CO
nD4fOi3ijIsROryaU/5ZxKPCcgLeZRAAlNP5ufLPHB5Wa1QYd5Ki9o7wc6MKg1pp
tdfBi1NS3G5lCzME56tVlbui95/BR1/ma+/P6mT3gK8ROPX3JSymSxbQ9vhB1qwK
JufFwPuSRlOfYsRMISl+bGwI4kiDmEOWkCSxWQfX0+r7yCB6ovV630MrIqttRSi+
rw4sLSs+TYPKf8OrrNfm7yICokhyNFbHfj6BAxsP573n5hM+vKDu3KsXrryud9gJ
pD3hPtCEMdKtcTAqAOtFvnv9v1aiCWrmVftyMb56Qyi/+GQi13O+VeMCObERQYul
qK8Cqjei0/9il45A5885SKpJ0RpqKwDCby04l6Ze7umFtkjWoMol2/f9ZbacdPL8
1JIKdjePZwqHs7bMvoUrR3kTyj9dsw+0W9pMZxJ1wz9xRe500IJttO2/l8LtRmdE
x/B0NoRaEhTb6QFEAJlfzlORzh/8XUMvXrCk3jjJ3oJA3zb1GX4/rm19wZboM0Lf
u4u0Mt6XwAmuo9+w8DNpCze+VnqZ/7ccQL+xAslCvcpFYYUjOcrWbGcIMS2/yc5w
0HeNiuJZWuHi9jZnNiwR+1GV6XOopywwEGJ4tGNzraWSnEG4hY/unz6AZYD3e2oj
ADKqal/Olymt6zFXHYNtD/Br6QmZiq29DYczkAR0/Dr2VsdOw8AZVUxKWRIGojFB
U33Gk+7iX+YV88x3TO09g/IchTQTAneRhwQ5M5NjO2QoufPkE55rrjFo91sCcPqh
clXD87QRyvF8RnGE/0//qTCYLi7l14ZBemH/MLyZGShL3DvtcSZKV1kCF0YBcVS7
AF1BpcQngM0XDnrb5GwEowZtQCiu/KqqY/5AO4/DdQPFmPtE1xl2mbW7azCKDPqb
c5kVpaixi4AUoE60PNSkhX4NJ015I87OpOT19eFgrIekA4/iMMB4B4MFUyy7MUL4
RCcnPx4K0/O91s3jSxjaDEo0AIbJPAOD5H/zGnilbMLlpD/m748Nht3yqPIXEva0
06mfVvSxWPquo+1CcBe3468R1Awa5bC7YkoDOQ2iBKYzzKy6KWsV3oo0+4N7B3Lb
9+eJTEA+53Pr2+gxYLj8Unc1sxL8+BVSttRCgbcEOrF8sAXYKscKux3KYUSAuW38
ctuYXanZ0GiUOoA6tKi0CNdGmfUqWZ9sPr1HyAdCyH6lg49VfQkvdyE+O+LpGDXo
nh7SGCxvnVsQxZ2H10I6wz3ni6EhhV1rBG1pByljKXHidNwiH5jp5oDCna+l9F0M
oAgq0Coy3cFJEcGcBsbPdHFu+CmGY8DGB/NcDYVVuCUS8liiNQYR01jd9EIwdSuf
ki153p4gMOK93fMc2tMqROHGk5GM0+Kp/s89FkLf+unKBapwCNsEl9ixN5sqlbnE
UUJQQEgakM+HGeqXUGAKDm6XuIHskuZcZvEts8MWqqlTsCWNEcg+x6mUIbNJ0okw
xliUwdb95EWAHPQjy4CJUVGFRRpxH9sdjFyrnFZlGWt0fhodp2WXBRRIf82b4t62
sCdQ/hrYzp1w+h93GkWLR8y+Tj5+4yxVIUEPZaLgKluKtZ+FL0fyuXjuakma6lFn
k1FRhtf2Ug7QKQyES23o85ZC4pEhH9h1VPZIFl1qyrV2ms2vgOMmZzskp0Y/Ry6A
05HVi3Cku9qTF4yFid6lOf1LNGy/RXbkWI4hE55fZBdPItfR3jTGDLEKhs1i47k8
LX7ejoT94LdCaRKdHQAqYi+j5lXnSHdqEol9uiAUqfZzwN7GxvrK8v3tqj5Fe+aG
ppLlAUQVu7H52sVfIyKYl2K9zZJ92E5A9/b9p4qmHXcvb7rD13rN8XpNz9KO19jB
NtKketGxO4rH6sNhmaGH0us8phgixFT95unJqJfKjkvmwq47fOxe1aR54ULgLLvs
ZMb1mR0FhnxiYLDmr7eoMEIvV0LGJr29uAfbDkHseSiw4NXIWpgBLsCcishFQc/e
rjpwfkn/Cqzv3sRHrZEVtosu+uvD8meJdewyvfov8TKGDbl567b2dxLddIi7rMPs
WCYZihvXJVnUAbA7faroTNzRIL2C9j7NMLRi2Mz7HbaM9aNiGd1UBat0HnsTG2Yk
ghh0lgn6MGk5Os+Ei1Fe/71GnPqbhDYooYYn6lAo1DE4rVrI2e1gaLwqRfir0CR/
wzoGxZwcu8T+fXW6IO1nr52CDX7VinU/kwBryTSJt1emVeT7UMyyrIeRV6h8UfCL
MmgUsWGtSvCQr4UqAYJBzC8BbleVY7GRXDCfSkSCdHTAFcmcpJ0HXPv1Az4gL84o
njdA4ePdykUJ5wcLv3NReUVxVsCuCWDqPzQkN4t2nZDlO5T/sJxf2IE6O9tNrk+C
B/QbgztndiL9rNAR/y1yUzUzMSHLO3T6ZW8WpXCmP23mnswrij3ZE68YmQaiw1Z3
WAlsaDg2K/TOiifiwMO9lD2sGjyeNyQc7qdf8Wo8WpUB2bqNZhbwYrBzc1Az6L1m
hh0cVdNTD1M6Xa/VjleI7eXeqMFEyYfx1g1aIHGret5lIAqGFnCnumsNWqbr14IX
/g0xZyUpsnP1G8vPDfRwmGyT6FvSqVdLGM9Zi+nzo2eGfsli3xvKGSO9vsEHjYhs
BfJYv++eGbpWXIHRbeyPaIF0MpY835AwdQklMvRkcyAn2JkCa36q3tYmUUgGVd6c
u5+48kXerz/p/LVcuklB6w2x/w4K2IhpSg8nr8g/v0ExcvI6JUNtK3dvNWx2NmJ4
H4gr1jx10c8vv7hsno39nIjdFBnZv20IUgQ9l9AMhs5/GQRHjarQUEms7no1a/c2
99oeIopcSx5oPGVul2WJhc924a5HNqeKBsHFomPvSA7qkxy3JguutboSsspOcewk
KoKYAln6d5spy4zdRlHj0wpD1DSxB6drWRYU+hysIYcBH4B+Pv5VlG5bOVgvZOl7
X8mINaSLltv9H5RG2+sOpWj+JKyZ/IOwaWmZlfIrKSXy2BCloOQtOk8rDBhmTpAM
MAXXKVSTQUuk3cguNkCBzUebiOGlVGExKCPNzijhgRd1grCw279l0M5UYBiZBc+i
ZQ31Gnwj9nTkhkOAGcPabEUdH6G+xWQunv4ysF+2th0k7HO0v5YkesOYHCoFVDoY
nBOPM3Lmkk5rclQ4MGox0K28pgAes2PVwfKFINp4Z/i0AVaSC1w7mX924r0GcOmE
lJbBVXoJ/1n0vp7uD+Dyq1tADnVBSGGBMzHhCcIXAfpRtQfaeuz9IeF5FrPg9j2P
glYeBBVZ8XnwHopDut8J+iWtXDkmAtuWfX+PQMrlpRU2hjKfqwRHdkQa1NmnAcyk
TZF/dfO1wL+UlUiH77IjSMkeexVn7ApvgzjOxi09qFQEqVck1yQe4bhYrOpcOEXC
lJyJDdkUzXA1fVRFuNtQSn+B79nMg4Hv2HLCqfaJIp21ctXMa5gD3P85zqCtfKck
ASs//e12NTkRB+XBcmmXJrp4htLxu338LS8Kl/NzNnm3bOTfCBGMmQnDXMQRNvn6
EqkJg53xd/llpET5m4ULRA7JWnWEWscSZyT6C/ZEX7vo4rg7WAVPdOVj3/cwmoZY
AA+wAKxr97GTV5MJfXIlhgErVsPczuCkSMbsn8Pb2cW297Usw8n6bPjP9LHdiIQ9
W93mtDzwn1AMDP7ryG9onH0yP3X4I7+DS8LjcXDx6i3W8QyOgxFNDbjws71yheqK
hySKtumcXQw56uXJLjGYx5ec4Zyqlbuu9S4Aq0tCG9pXWhWSaXpOor+MCVYq0EME
pvsp/6rlAbxa4KPl173NOtX4o80cZE3pmn/ueK4K3fecsZiz+xWqt1YDH3Z++LW3
/uHm4akt+WzSt+YhuEBQC0gMsTdLUs4BN7UKX2VpPFHSM4QlIUuFMLtpLnjVHLwc
R0IOk+Ny/CqxTItOZSO6B7/APvbwnzO5OQjOZkH2QmYkeBFOteV+F7x88vRjvS1W
ueD8aOFwlzFAYNAf6HpztBe7fLskxxK/C3uth99CoGJefSLbS/PUpb7CIcNqduOk
Pn3X+uYX1+hMsjVn6dSN16kofXUimcwHCbShdboGPzUd3GQktzv8fcBsSU+HTv9n
1u1mvjXbgn1JD1dclRTx6MDHS0nsEiryX+yfvWsr5x2FoRD2zKblSNOmI1CK6rJK
ZVg2jjyFLIeZJm7jiEfPcY6k2XWsZDxHvz3JVcpiOe4tuneBkWjYo/6eXzG3J7RJ
bS7iF1auiQv7rY+a57QtYQrdDO2pdkSn8CKksUzFns0C+wxp/63cGtQntTxG59AC
ySQzjfwBfQ0QDRPo8aIOyWxEKj8/5+lldjdtOo2w1STAnaCaTOwxQkUxalsMlQS4
9LeV8HHtZ6irgCJtQFjxrSa9nV5NHI3AiwASXkaDpcV4Znu7VlelA5jUUuuHN1dM
cGFLh+Rb0pdAw1AT8H0jNLl3btSwdGvlt2BoHvwJauUI7I1BEEwW2RdXXCdf8BI0
GjMXsCnLj5/QJNDGTkUl9HjRNXOxP1+U3TFT/2SOlb7ePVOya6SVuO0so6mBOuUN
a4MOoX2eJjo/WxRSr8DPGWCuYjqNWwvDfGjk4c3tpPOUYQCNRQiBvDKJH1Ujxr8r
ybUeahYeiGbjItpZP6lv901j9br24X2qAFz/T/ZomAZ4ziiw4arg76eCw240107I
1J1gRpQdD6oSO+Xjds5dvai+bYIs9Z+CAo7oLEvEI6gyEnn9ImzTcpjwKlDRPlEH
4yEGJx+pDlWdfHhzNnvCZVVRQhHKqEDyCLGIY0dLOWnk4ZnR/XdcIbJQEWgU3QxF
O+xt++OsLEkAaUfswTWaCEYCzjGKcKK1zMc7n1LbtZi+YEHB2Hm0RudnVl9wVj8a
xBKSaussBVCYKhhigdgbffDwXIi05Cip+WmP9We4MP29crTie82iYi2g0VFhmyed
tMVQh7T7djf6JZSYv5s6K+y30VOuUQncfzpJ5VUnPmkva7SB6MsTzVcN4zPdOUmN
81s8e2jS27u2gM3jLNhSLLHhruLbb3jYcm2Dy94QvWxChejzilVLUygmyFI2WS1E
t355Bol5n1TDf6cMb7BJy5Bct0AGZaA597eq62KOr0N1ZtjM9wGkaI8gIhlV1OYU
RiZchKUqHmQyTwEJXwTVorer1Jn+bbTaQDyWLNTG00aP9pLtkrRiaTYMUQGMkNXU
foiqs3R5ehQbtASwNLT652uHgJyLMGpR7dr9q1B+xG76q55A3evaqyqR/VVDiqV8
FTAJEJdRVRfjDdD6OMKWtqjLAeCo0rvt5xMZxb2MZS66MX3HL08T+isWYqUNIakB
vTfG+gS4EPuzHXwRnj13CYaD0jMPXycHqAG3tvFppCEJDIfKxZYDUepZYUyt3OzY
e8e5v/A7tcXoFByK47xGY2e8ATjY8iEqU8qEitwnKZ9V+XFXrVad61xK4O2tObjX
d8rVDTTMpTRxVxkBZtHGoRZZU9ljdInZ7KkcRvOA/gf1VLAczD+7nuzJMXtHuE/3
PQxoqPCHh456ayxjWBbtQpSFr54b0dtviKGXfWHSF6FgkddJvR55kPOMSEhfc6We
uSl62QsdoST4kMt9+UeZuMZWwinmzbLhDd0oXEVC1f0CJ5jicDAz/RhlUXKJC0wm
9wCBL/cuWD04xem+Nm8quGIjBWuNCJrl8El51qbEk2/2C3xpYhAFXvrC94Qpu2Sh
6gPayieYRM89SaewBAtXCmGrPcSx1SGLk7Ut5CMBadvueCYaGBUbLewzliUQR/w0
2u9OURfJYIsgDnNEsDoYpONvjKWUAxe7peGjztoErMK+ObtAqdYqAs7Cj2FISKR5
bs9q7UY1i2dPA8LZ/VCecvWSR4qVMtWbaRIn+ttgy0TRW75+U4objueIm9urhLQh
yXN0SNCXhY1kVg4YKW2uYwU1+/8KDjVePind5iKmyZwQnxJ7xsyFjwlT7JXQr6yy
2roNWXjNFRKcZx5pbW4LxyyqgkMiRnDG/Z+ErSLntIB3M/cgIARiTd4n79OejlO8
6DXN9bGMevNUfxg8VFj/HtWua8gAuDDskpH3g5M8zNHftC+0Y2MaUj5YVMWD9Cgw
gPGj8f46/RB1UKjU4/Fo6MizNvpTTCGIOPEOoawt1u0NLMEPTLsLAqekd4Si1oLi
e52eyWNrRym9jQPXhcDlmJPUQk7Kq21FlbI9xBUw1u+9dumg6qAe8fGbRKOusSY4
zP0tddMy3IXafVPqmrSDwrz4crg+Ljk+FN8CpZqr6ws7HTmG9Vnox5/zaNTITfKz
aPHBlOlh+hM6NcsVULo0DZVuvq/vMOmp3aNfZTaWxMyAvTTcJFrB0NB21rXsqc1j
VLGrFfIJBrfvRslL9cfzyMTaRHwleOugY4FC+7yKYKqFvABQWEDYhPkbkhyCZOto
BQj7PcmAg9Ai9d2pd7YG7P/npVgLrLqXPTsNBFLAVD+PdZxUApaY75sMc1EhCDIx
Yq7FAV3hmyK2ZVmonICx/JtgtUh8aQRNgTJzVWy2APsGJxt9ivJV+aCvDw8b1IIu
DDK3KKuDiKj5S7X8hYKgkWd+m0dTWoHhDQdaUfzv8ddny+//WctBPku8eaSSZQRX
sMroaJpeqpVvzBYu8hMggJmmt+Y4VbhEq7O5EFiwbRQ25/7Yw/glRUQsCtxNRLJD
Vy+UnMon78TDytdAUu+BdbIHtEbTBPixV68Zp+GWkEJNx5BXbp8Qr5+PWSscrwhy
uQdcVTfrpi9+DWy9p2wo7R2b2tjrbmIt3uNod6fth0ueTJ84w4404u6lHfmLK9Vc
TIjlcw5f1hIuGXj+yNNdmmylSrHArvAKC+Qz5tuR3SfhdDwbriQMWSJSxWA6p8oA
cOS0VX9VCHQLc6bHWmBgtsSUnEzJ87vKpeNi2+4LUrwHpvc3DudnyCv4eH1kRw1q
Lj17JnlLCwK/Bg8m9chd4E9vnYuC7trnKazGa83Ck4wZ0ypBq8RuwiyTExfqC514
JgAnskUPp40VxFML0SvQsj0ciTGSJJTg7RIM99v5KvW8PFdvxg8wofHWjriIn6hL
PG0pXs4Me28twexXyG2P3MjdjSVG7D91kHZyer2xYkXBoc+Dsq6bfuf/UQz3zdbW
Qc3pdT/5/CBIWpe3sy5OE3a9co+E5f1sZqiXJfrKPWi4B6iTWE2PAsa2y/jGV/9k
SBYezu8igkVOg9Q5yKqGJ1+JoTMhdiNpJoFugvhnkx1yaXH+cu4wM9aD7u9z8bJk
OaXHI1mdfut/HzW0Dm43k92hG4WZnphTEKoja/vNrX9qpdEMhzgvNpIPCVOIXinT
gI5AByIbmbRzsB8xFpta0N3/kw0yZyN7nIXb2IJLo3PCR6lQptnJbKQumLO9RMb5
tfZbWBV2pk/qVhq6vBU3ne9Adw9RaaJm1NIPaEp9Uz4nq6ITrqkCs4onM+nqUKEm
XXWBuz9N20IWqguUhEqtRUearQfXro1+NkgAShih0C2Ff9rNA+OyhV/SmlM0AyD7
rNeNn9tD3GPJzolnuaBSJELo2Gd+lyCprmJfVBY74mi6VGVIZr5nctK5ytmCxj0D
SjQt6qt/86xZGseiernWgdMcl3vEIT+zB4aLkt3BhRjs3QmwONs7dqiI8CYB7MZj
ORmf4apm63gGBllOJfppEq2BAREW1tS1AlPpM180BRiw3zF4/gWJcOqVXaosdnsB
D0I/XqG6oZ/iiz2D3rehhR9mRBbmUClFTyTDRGUKcxqHnfH5BwwTI0B87w6l9o5b
Kfd47d4+N4Pzquk3Zfa02xHSCehWDnn5MQAcleiY0bNYjyeIYobi+dk3Kanncw0N
`protect END_PROTECTED
