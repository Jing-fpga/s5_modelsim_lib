library verilog;
use verilog.vl_types.all;
entity stratixv_hssi_gen3_tx_pcs is
    generic(
        user_base_address: integer := 0;
        tx_lane_num     : string  := "lane_0";
        reverse_lpbk    : string  := "rev_lpbk_en";
        mode            : string  := "gen3_func";
        use_default_base_address: string  := "true";
        tx_pol_compl    : string  := "tx_pol_compl_dis";
        tx_clk_sel      : string  := "tx_pma_clk";
        tx_bitslip      : string  := "tx_bitslip_val";
        encoder         : string  := "enable_encoder";
        prbs_generator  : string  := "prbs_gen_dis";
        tx_g3_dcbal     : string  := "tx_g3_dcbal_en";
        avmm_group_channel_index: integer := 0;
        sup_mode        : string  := "user_mode";
        scrambler       : string  := "enable_scrambler";
        tx_gbox_byp     : string  := "bypass_gbox";
        tx_bitslip_data : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        silicon_rev     : string  := "reve"
    );
    port(
        avmmaddress     : in     vl_logic_vector(10 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        blkstartin      : in     vl_logic_vector(0 downto 0);
        blockselect     : out    vl_logic_vector(0 downto 0);
        datain          : in     vl_logic_vector(31 downto 0);
        dataout         : out    vl_logic_vector(31 downto 0);
        datavalid       : in     vl_logic_vector(0 downto 0);
        errencode       : out    vl_logic_vector(0 downto 0);
        gen3clksel      : in     vl_logic_vector(0 downto 0);
        hardresetn      : in     vl_logic_vector(0 downto 0);
        lpbkblkstart    : in     vl_logic_vector(0 downto 0);
        lpbkdatain      : in     vl_logic_vector(33 downto 0);
        lpbkdatavalid   : in     vl_logic_vector(0 downto 0);
        lpbken          : in     vl_logic_vector(0 downto 0);
        parlpbkb4gbout  : out    vl_logic_vector(35 downto 0);
        parlpbkout      : out    vl_logic_vector(31 downto 0);
        pcsrst          : in     vl_logic_vector(0 downto 0);
        scanmoden       : in     vl_logic_vector(0 downto 0);
        shutdownclk     : in     vl_logic_vector(0 downto 0);
        syncin          : in     vl_logic_vector(1 downto 0);
        txelecidle      : in     vl_logic_vector(0 downto 0);
        txpmaclk        : in     vl_logic_vector(0 downto 0);
        txpth           : in     vl_logic_vector(0 downto 0);
        txrstn          : in     vl_logic_vector(0 downto 0);
        txtestout       : out    vl_logic_vector(19 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of user_base_address : constant is 1;
    attribute mti_svvh_generic_type of tx_lane_num : constant is 1;
    attribute mti_svvh_generic_type of reverse_lpbk : constant is 1;
    attribute mti_svvh_generic_type of mode : constant is 1;
    attribute mti_svvh_generic_type of use_default_base_address : constant is 1;
    attribute mti_svvh_generic_type of tx_pol_compl : constant is 1;
    attribute mti_svvh_generic_type of tx_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of tx_bitslip : constant is 1;
    attribute mti_svvh_generic_type of encoder : constant is 1;
    attribute mti_svvh_generic_type of prbs_generator : constant is 1;
    attribute mti_svvh_generic_type of tx_g3_dcbal : constant is 1;
    attribute mti_svvh_generic_type of avmm_group_channel_index : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of scrambler : constant is 1;
    attribute mti_svvh_generic_type of tx_gbox_byp : constant is 1;
    attribute mti_svvh_generic_type of tx_bitslip_data : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
end stratixv_hssi_gen3_tx_pcs;
