`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bWPSmDxSZo8MsV+RZ51E2p3dvQsqfohcuOUL82iZB5OdynEaa+EM+aeXf5JO3Zu/
HpKG/Z0s4yc4u59JXSfctnkucllTryVjKbo5aeGC8/7AU3g8++VjyaCzzsR8O/Nj
EwRj96zeMgQQKWkmaKM/lOOEwo5Loy8L7BUDOaEA5FSfYQT3dOojUmlxKZVPEnZW
y/gz90OGi76sR7nIDJWecBsQlpoQNTs8xudeUCgL8JeMXg+uA2NcJoXiYNw06OMG
quND5n/oyfAaKWfnXjsPM23zCI7DQV/kNTxcaIW7KqKXfaIBv8wyHKltdfOrD4nd
2gS64xoj3BTcnSbIL70X0s7Kkg0vACAyGAnjrcGkaVGzUXK/h4xa3D+SWiVmBEd7
CDoAWofkV28gfurnPt0TQq+AfGm7LJiJ//psGJ8maATJCAIiDfLcVoVS8N3VFcBN
VvyZujHtX1hkr5oqCE4sVCtL9FZTGlG0r6QVLeTPR4uc5R4MayP8EupFXWhPKckr
SblFcXOsKHurRqX5HpL/xzgv4pIqOAjtoN5QXuEa9b8Z6WFuqGt4Yu24nQu1M0a3
H3WH573inU+w5P0I0jWhInZL83/XqiJeLRYKz7fRK1mJi4wqSQLbP4S3Tr5iiAk3
djJzeLlDo7YZxUi63eb0Bwgo+nVQiCFNBrTDjxj8ziJK8wDGdC9qAYylnZmxMSvM
5K839yXCG4phw08/yyKYPn0Ci3fsIfOy/gv+WJNM+mCpKtERib6qGcLxt4WDBRGk
mNB3/ErY66bWbr2ZpaUy3MU1J2bD0tNsVRal/eaKZ0qlFlJDPUb36R66/NyTou4R
Xs33kL2Nmcc4ic0l089FjyIOaCVUGLYvOFS/sn6q3ElzXJhLdziQxqIuFm2Me3Zc
xx03KTfb97vs0EXSalDNCfB9NmKZn9weX0EJVlRJflENJoQW4ik99Zv1LW2cwlcM
H8KTm3YGby4Pt4Vsdg/N8OXMlYyfVb6ky7GDJ2YdKEjDlLszrWK6xGAMTpJ/W9vp
gaGnPa+PD4D9qEcIUkqN7HBerok6ntyTr6YenPwE41qjRePccKikvUNtlWfTpcfV
fxi2xNmdQ3TCeJ3WcJyB6CM/8BQcq3Py2F1qZwQv2Dk2Bmv7Pfuwvr0By77nFrHA
Pa2pi80TSkNEcMbh1JkW4Spo4ya2X8iqS6ItdwuvuA1qZWxO7f8hN7qdX6NHPm/C
gFWfRsheEpQTYFNjhIcPaZy2UblYd4aaa+YJ35Wh2BaKvwNzhTk01WHERAUfrY1d
o0XlFKo7TxDbo/trR1fuRXycCiRRa1qXsypbhoBMCPT2c9VWKbJGmBog5qiozx4O
rzsKkmhoClOfIC+4dS8bIqmg0Lvh3C+HBGbM9MChr2LGEBoEYC4hAJtYYkW72Wss
/7vq1QokQ29yyL6mdkBgrU9VqIo64XvVKQfOPktrLyIViBA/4YY/8LKNevZhhfU2
/H2vYD5En5PxZamxm7JiUCb9BNecJOD2SztsrigMgjYEG80nz2rlP3lxwNscr8Vo
FHCnOYRI9r6G4T2vfnGpnOjtKf9yV4p5C/V2+jcvhEIcHY1LmFEX2LlljdhgPFKY
jKpPX2F1n7VaWnEzqmypIiP18WCN99B5MgMkG6sBEPKVbWOEuq+a4O27VDDq5kGg
nLtaK7mPnsCEILCXWZW36a34clhHbWYCHw475Y/Y4Wym7w1J05IlKaz4UVOmWQ1d
ZgVkXkBaOW8oj70ZNDcCT1lCGRdba1WRPnwuLY/QLD305FYvlYmaB+4XuYKRz/CW
aAPJzoFl3Tn0kiZYSFfOdvz5HHyGd6omal6LwbuEAqeDSBhO3M5QfRBf63dU/fKe
4Ff8X+kr5Bfd183difLLb+mTP1zvmMhUHeXWpcDFm0lZ9+609W3IIz4EiLa0+tZ4
H4cwHOmnfrGXlWjKGLbGdtCIXQdxiRJw0C4b5HXmzHRMGzGXmzjjV9YQWAiz3JfE
Udz84rT9PqPGR5jwZuNmndyShFTv/7eY1xKNnC80SLXnzCrgKnnJfrZcZxgEb6eq
sl1/M8AXKWE6SRyrNsgR1eejAUokL0JrGwOvBojtpVgGrTz7KP8SYslXD/hveMQD
P3QPNaLL/32dhI0QQZsbfSLST3dq8b1A/nx830m0t8Q7wPWlbbKSxjZxhcjxIqDw
zTJ+LxbKg5UuhaxDFouDCSd8x/f0r0OTqBVSJYtuhZtbgdIX7FSo9ODQpSnGhIgm
E8gPpKZQgQlm/WfnSXa8vJumgXhhiD7oQYbHsLIaRV6o9ttJwLAZz1ag1a+ro3W0
e51t/H7xsL5AxsCIGif0L80YOQrodU3kTkXJF0SQzkt8EB+lz2p9E3+hU+URCCc4
7uavHaqsMOHdsQlrMNrMB4XwHD9H1BMEkIzfXeqBVR9Fw60u7HVmPRrd65yJy+PL
1iXM+wnSZyIQqYHo+AGBhqADS5qUfa0PqT3UG4vJzSeE1qXT0jhRTlpjHm2iwBEx
Lb+KtqR1xjQbtPoJPWPgCEkn6YoaF+D2vb4a/rV9aweZrrY2HoqlToXeTPVpSDNO
hxz2uUwczm4bVBnXQN/0lyFUdpOqk26EWClUSp8t8GUOXDVoR2v88MooliHmR5ev
cSWtAqI8PvZnIxOObglYUn2+7Cg4poJsZPd5uGatKZwlFD8LNSDHIJVs+4fRPQ65
61D5UIF+ntlB4lcvu5w49cKP/7QlzBvqxnhzYZ0q36+tazupb4p73EvkgpztBKXJ
S8T7Ov5ecLqLR4u/Qh1H8np2k3DWlZCQ5uV9XVGLtSEk8ewvObxNOPhAPTvV2B/e
5rDyWwi0a87cH9qewQIq2jcpwaHu+Ytysq24WtBDR/SnDUKB0/aN6olVVTuAi5oO
uxbuO+QrRZOfl3KNl7Su8GHO/xK7fbTdFWEUCMtUsDIKq6J+X811hTabn0uJ0PaB
CCQsrHQiXTT1HN+prt1HA/LKFMo4/qAmERqLTXioJ8Y8dgctAHLSpTvhFzQq9lW7
JgXtMzijD9p2TEkrT+YjQ8/6aEky1MODsekRrdk8aQqNJGtSh4zVFIVchWSY6dLZ
teDArOaT0GXkdA0vjbJ2Nan3Jj1bR5wazPyUFZfufBAQ6PW/iAFoqGniuz6OCTNt
xYtrUkX2wWGIEk18StaLAzR1Zhi05x4NQ7q4rQCRVfblfn/nrgTAGdX7EqRS/A+e
7cS1S74avyLKlOXZ9NdZALIss7aCQAZa/ppuw45YY+TTFwvzMhlkwwLrL8j0dzYs
5OXlQXDeQ31VcOAHQBdQZpbyR1AdhtpVcvtN62/U7BhE0p3e8XDkT/IfSxMGq4pm
lqS9ZdALqBg4RfwppcVrhxKsaXz13UaMvYlcdQWLwsRG7QDpwfraU+zCEGCCAnzy
qbVI86wKGI9FZFapVmv9jcHA0oDltWlEfswdhM0eyWet9qfFcaRzE+CDOTXIrOeO
Nkd4yYrLUYM90MJePP/H7/5GUgeNVSVxeUV1bscNYH8jfIl/nbIWDrDvQyDe39Vn
dAurQYJmA+NbKfCoLuek4G1K67JAt1nmFs8LAzTLL5EQtKkAAsftkM3CGmm+Aiqs
/jm3eadEAwjjgPz/E6w1eOhef6IRWJrmRRHz3k3ktyDJBG3MCMxNaMtJIuCAnINt
7/zQVDEuCaILBij/bBz2TKYztsXNla6nw0htaoyE4YzmNpmA+p36knHEU4vRN3GE
X2PjQvcByhOCHOL63BGG48w7PFoHz8cbhOORHNHCqqVigfkD7XA21rUsWS0cdam2
B6cKxKwD5Y/GqD/N0NnIiay91uIKc1/Ijw6iex/tgHNabjgywajj6nJ3EJK5H/SX
EKkojWlmT28wYDBLITAX4rqLVCjDSIfm0Me2V1ZgrTHNoxV6BUgBlgXa/WDp46w/
0p2MZ47LoRTWlnlaqDrtHG7//ILaANbtiokui5V3ieeL+Bg+rpgQRwfEgRKpjn6H
wkMaNSEzJaHxm9t7MvFBdogH3Qvc00pApzLl/S/JNEtLNQVBgbgwsM/+sNZKnJGi
BgeLYgyWsjWdJqYiokHThI0kpezYCT6en1ddojxl6oSJVXPAXGg7Jyq9ilBzISoC
syJbjE9xTixPysjCI/z9rt3hpCDCE6jLu0xVblz5uKI+lP4JTfQLV1Dl6b0EENCN
Rxv5k++eVnKBMr7KkdqAtKpnXvwyRjHu7+hGCrRGUB46X4Ei3SiQOLqVRgInZ3e0
6Sj23emsqEJi2aDOwZQj+XIZ6CCJoXgCDYm2w8dN5of2Cls8u9TpJtpJNzomZGyY
5hAtqK9O9iMhAILvAJ9T1ta2XfcQ7tq8UFIv0cXBYGgmUIApifp5mVrA6ISPPMqX
S4zH94cmWLMjywsZ59mzXwIlMBIGW5wNYy4cZmZAtGQD7fn43J7bPa5BU8L00raY
hL3L9YGInra+jdHW/xkOMNNhhpEGta7VMJWRmiZVzFrYrSQFmcrIJQGEkZLL5gVi
leHKUl1FVTBFDZoUfGwezFMUxFOLZJB3O+66jfgqc+7865BoI3taJD+CRxNA5pL4
/jr7Zwn6VjK1MMa+wlRcpWNTCUxhHVD+SQoHm4Q4eowoR7SVB8IK7fWU/bDaHsZ/
+vyBzCgQux0EqywQ64ATe0qC6r3dFlsKHRTwC9D7L6gVpcoXOjo7g9TxbDkzFDoo
cf/biQlA97DRPzajvwawu8cLWlouS39hNIec8N2H8j+TY4SYE3Ph1g7cEI8BhN8z
iAs+topAy3aA5i8bbqiBWIyQY1XhswR4fwPhs2rn+Pk3dzkIN2kiOTSNQAeV2h5J
On+lrDB2xLSpUUsOZcJ3bw1f5RkrDfDeXjt6MwwAaeiN6E7LC7NrICyBixox7Ef4
GIJx681qFqrbytnNf25HzHW3RcUnPY+hM3NNsIuktdAWdf+OIBR75HmPprt9Ccm0
M/kT6mxPqznpRSRZjOCITpVjM5ZnTlk5O3GQLSKC+PcVoCSKC9UblWUEUqkmumHa
3+mCbxWX4Yz38RwQUSyJf7nVsCvMrvh5ttjjLCBNK8CNtm+E91fkQBI4LwGKHhRB
RFE04GSYV4vZtHoyTYU5dY1TJ4DE5nZd29enq7tS+zK/p5RQTfH1TkOcd+IitYFa
AHPwgfXLxNGb3YDe7NGHxH+MjkupM2EHKGRB2UzgoKVwcKMzkp3JcH9Tby8kj/G2
f0uhAXosYBKwukB9FVGLl96LuGCxcGWIRCRxSx4pKR4wIej+qKAhb1DAsgteg9PY
SWbvEM/3G+bbsXMLpme5wJsWTyhj//9QJXfnkpZJgeP+lY3o07kovzoyeT2DdPj9
uLS90mj3N09re8ZpkNJjbUWCKyENBUtEJbr4TjXNQyDDROyBHjGBvfw/jHDEV76w
BhMoVTqpHTJJ4wI1hCz3s6XDkBBx4ZVs/5VjIbKDAABoBl2AkDH1wxZD4O8f+D4v
HyrsYsDhtym6L4/paKQ2tyI6NZ4oklGhY8F4yAozHWYc/p8uUElCb9AR2sFbXix/
FAu8Mz7xGp5/gjdHzIAapwnqq9SKpWjWioQcoMBFlkSEGH4md8KRuTDDJhlPAfpl
y/b+3gaKD9YA8SWDI7Kln3xH0bPvo/KU+GMI9vw778YsSX5bU2q1gpFUiIGR02W0
VaAphPaOT+crZyrs+XGYQ5CeTf+ZyFu2bh+C2dhQ0uHMXDJGmWlM8S6Y65IUpd2n
xiDNxYz7CcNSDb+9c3O7yCRx16SxnJOgHM/BqVUz0nqYVgkzzogWxdLMl3eNZBRl
VINjooKcQ9L3o2m7+nVs9oNBKR7I1TV562ZC5dAQPjsRC0YTN1HAWPMpdWA6sYN8
zsEXt77eHPlKixHyJ0tLp5o+J+GlH3FBZPWgbtbe+3UegpWXsxiNJTCjJVfIXydn
k/WHrPR+WsafB/ykzftiUftABUHqGrAHMEJDtnEAAHs24CLCeosIBtCGNVCuyvAs
vG9dZJgD8ELhduZFBkduhG3shwF8fyYxxY0PqMkz5X/IjKAQcud+FwGnbIMtwj1E
1eArz3B0uJbYR+6dDvRqqvDOOaGYt8DGG2T4Zw/Nx0yFE01Gs3nbDk+tuJaaHy98
mPRrWN9+vKRHHXNc1ZLWU3ogLQhG7m0t0ebkHmJ8A5GLm3jMhUUYnI9cnt3BuQ9u
wRgNeIKlzysGdEgEEFpowc0iq9V17XVF9zTqwAlG1Tm9i414VmQGgifmZTJbyBCv
bhUdAcnYf4EOdFKb8xe/cgW2gbcow3FXkkEzOWqJjYVsnZ8/69N93bFgXrUHQvpn
DxRiFvveuDHDDnC6oo4kstvC0bwMjb8ZrSNGz/WQK5Aeq0OM0xjDL1W/I7XpqFd+
LNsDR0nv6nnqw/CMYOKBWWefu0lbbG5G7g7XK4EXE+5hQFNo0ygTRMXTbD6v41HD
yB1li9UB87boACYDep0CHzJKpO1/S10JBUXwJJpGgY1uYpbLJeQlQxy1/ORXBThe
IQrrIuR/TC3r6vm3nJ4VaYRRs2FD+ULsEtWPuhoOimvwHHevMKH3NHzN00TLoLma
hiUKVpBUsu9usuOC+FUHgab9DmR4uRC/8vTGBVIfCW4jG4fRsBlDlN8JEHsWG530
AoqiCYI8aiTa2VO8gbYJkR5ydM+yRwyM7oQy9jTYYDlxdAyfmtNnG45po4URPqbb
hEFGFhJV/hQHhRGsXRgwI3sQ2XqeryEGBm11AdvMhPuy6S6dM1YYFjf2v5zSQSse
uA0WDUBOos1JPlDJifGwpKuNpY3AX9ZRHjGQE78dk/fADs+6hOZ9ngBSzHmO9i5S
RB+GzevD1UOxsQ42thWEJEtFq1J5MJHLjII/MJswnWohorl0ncT2XgVPFT4nukbs
brfLh3XV3YX1MIRm3wgHVlp4JJW/ZYGXI1Dl+eprpqAndCta/kiv64oF2uGDCEDV
qpclnfDrfbE/vCI6htJzJz6bx52379raGSZT+9O8rehuFhv8LdgY6ziVl/TcMYIO
dAfciW6KjGRniTVc13Nm84fdpu0T87TmomxchTJY1xZS3G0WHE9WGmYWMa9x/f31
7V/hfl0/9aGFWOke9EsySFYWowK01gW2UvgooHUMDLtqpRk+E1wjaGxv3DdobMbm
Sdwu8nQ90braa73DhAUxG5UMI4V3khwrKcRwTJgEira9WN4Mc6XdKaOP7w10OR0E
VmtIv/YZY33vKjmKoxXqU3QCIGTwc8HqBOxmU8JcdlrhJajHSf4KF7xs3bkf2QyW
dhxnhgbnfsng7D3d/YkvRol6i7PKZ95huLsqgDS5WHA11WOAwq5b56+xQq6vRKSl
CIvSS77xCt4k1TlPhGFVq8KsSY4O1M+e+a85PqXEgNLMBq/ZpSvDDwwLM/hbeygL
GNoAow0Yx3Y7pVBJBv6QQ9Gc33wJ/WS4lA/ktdgHjvYuq6GRkLBHRl4DYRYW5t4D
Nu52oFZS2S+TIw3rUBD58Ie/Y35Nf9MD52wRYvpKTp/wIJ0FH6pEq/0CbLzMziAM
Z1MWl1zC8Q8hLg1Ay+935+DhQNvGFWQTOF8Cy1aYiiBorBuIY8R4nUjQ8ZUoi8EX
E9oAf3R435gOkBmOTw8z+YyXIlnlRv3Anl1uXWh7J+WMOtwxmxARhc+DN8IeTZl/
WO+ZWuL6WVmzDgPjFHd9HRMSwNuIvRCvJtH+G608EFwh38FWqUXmFZUH/pCJNuZ6
4U5Hikz7+9sc6xu6Gs+VVqkGrSHmAfCUAU5pEmuLU4UOdWkT0jI+zAmXL1UDWdgg
0MnhUQOSB+Luq6VmG/QDMU9UbqzAvmr4t5Y8TjoCP9d3uERaBTeyG/7nWKRtDxFv
co/nMfTgVbVBmY0QZJhoATjCK4hi0D+Mz210fnnZPGntkykHM3VSHnVm7CsaVmA7
0Jl1a+j8gKSlXh6WaeF1X7sdUN64GSTykawLUOrDOGsiYBZmPbPlno5RPYoDgSNB
p1WnjuhnihAe8WWAyF2yomjmRZjehrnszF8wQHBhx7Pmbg4OCjz6OkF46ry3eN+n
L0U/JHRdDc7/vbgdp7JcD0u2mVVhGcL4UgXgPMJgil9OC6jFe2yMoF6tRKfG0Aop
qQFrNS1cOlmaI5lR3OyqBzqxOhXNzs3XTtCoyeSz+xJI2sxta//AiylCblZmrQQ/
5arRDycSj5Utf+qRvoUq8pGf8Qy8Sp6wBClVmg93xm4FXOgj84zhxY7Zv+yZKMkX
lnKQxR6pFdc/DpKRB9TD2A3QxsuTVLoVS+aVdGEVyycr8yi3Z05aNkkMW0r+VoBH
yvt74lu5rS3nIwiEkkA16ngRX+gNS/O4DlbpxHhMb4HCmgl2WsmVcqxmdAqEVSiT
Hjp/zhOwAgrwCupzH7R7M9edGzliA0UN5h9WDLfLrSmMmIfOe0IOq6Z3FuQ8vLki
S95MsZLGfge2cjzBILgEWMVLeU/2r5HURtk03vRrFSObzjwiAPSCt4LwxHemORnC
4oLGO56whB0rsLFLWWRopCAH/1EfMQ6ChcLMVfUYpkaQCAwbGwUaC/vT5Z8jmtOp
gJwLZWxFE9NEJxmdHCVKyysMxt+I+uVDcuMkdaEOcD98+XGU7Bs5vVNg00xhFAjn
AthD3WnOKvXUR24avCjomQt1y4eGrm3+DfUW3tSaqsA9+ZHBsFJqCUDAmmEV02h1
+Uva6+YHfAeuBagUhGzCumOQ67EgLdiEiT9mI6Lh52JaMP0xEMAh4FlCyG6N5u2Q
OF6LuQq3QM4e+Yl1UFJJVpSGM9aYQcWE+E0D6pIT361fDNoFDrMsthO0QE+JaFhP
VWhAqAXH3XZ85NbtP4G9C53I8pipCv6nRwV3wsKT7s4FOH/D0b3hwQXx00PvcgVy
m8qMDMN+zekaFfQ+WziUcMAavq7jVc7ThAp2dKflt4IwiWh6/dSSevqKDIuos0X1
xFdhjIacwuQP8sOKnlBZFPeZ9JujLSAOA7KVg4/z81a5+6MEk4SiCKQvkFAEeOiW
QJfkdZLGIWvu7H3mUQHy7IpMnVQOydFhhJZ3NUJ8+nqKSoYseTTpkr4JnH7PVg7W
NsJ9i6xCvGnEDkqb+zgiIPp/B/vfeWNFAmRE/xuJ0FyfpPR8dE2qvVvK+tRjRNlO
QfUGBl0W/snjGwgIJt5NidwDREgwqdh24i8V0zGOq4UqynUzamq8lsqSqxNzhKrd
OEUVF2/r27KrXxZzvPA2z2TYL+EWznm02uMfk8HytOoV9wHAcx3Xrc+wu0SoHJPw
A1UYRDko9eqGpp3ayHxTCxoDNrrKsM3ugRwU1GEK4CzANCqjLoAHibqg8GL8xaEh
KS1hATilcUJUDFDPFu7HvsNBqYzbjZOxA2LLMS7Z3ARWTtEGX1/hLonFugTARK/F
ghcDVyhNSD3ql2U2OGqJEQFSgARP4E8SWDQjcSnmZq+2XEmBMLD+y07pceiW45wk
380WYN/u0AnQ93xQyGjldO8qYP5Id6UR3usQaEX55e3CylnZWflOfPDb5dm15uLz
1rm71sW4fq9djlueI6wVKJ4A8IbstpzVrPQB5Pszvd597IddBX6gb8A54+IOpMe3
gWcnMGwASdQQHWKBcrS6seQBCd+H65alAoBiijhVYYU8+1aAsKEtDkD4qqG0NFB6
/PsEEmjoe4ceUK/hyKUH+ysKIRArPYbPb4J3HL21pfgSNW09Kg/OdKgnDpNLwVVu
tYYO5zNByuiDHMc3u8pxADgrRStZZLMsuhSFs+WyuXj/KXupSsd9Fr86QO3HaSF2
9Au3+rzzvuUpqyqNXIgQaV/qiMEF7FmhgaoxLPvaQShO0b1WccvWhgRJ14JjoVUU
lVudU/TZufao9WOm2GXB+kU1q5xPzDC4Up447x9rf51TvxCLC6KD+6o4oU16noy1
jXAEOocMroNHrYCHOJEAIJylteYwlyQ5DdkjUi0VNixl2qyz+IhxZOg3iWJOCYov
XyAn9dh6xh3cU6bgqxkGZcKQxtu9M30NOQHMYRp9ZBZ/2WWEG5zDFxSwZXMaW1O2
QedHdlIXvQWM3+Yh+UMTJKKlBTTYN//Q2dplx1ATQmd+zs77Z3S0YQKRx4Ei0ZvQ
/VSH0a2RMF7yguAM6Vt4jBIpiQRrPX3CJtOQ2ozJJfRsifyfFLusIZIAB6L+G3Zc
1lxuUBA5IaT3SGtsvhi4AIyvoRtIZxxnq6kwB8OnFbSoXkV6xPShuad+0OhwhYnp
GZQTBdyvibWnGUQbce/izGT88YWRD9QQtmc+/AjQknsq3qZEfh74aVBh+ObqaQtR
oIolPOx+x9XnfrrwbIJPjT5pp8Vq41/RhMQ1fjyU9bNxn2c8SOUPtnL1IIcIF3EX
nEdPXcl00BZLH072MgAGLdEI8CTFRSU0/FetYg9snsg+zv5N/X2E8wAtVgGE7URK
zshRQ3vCO+u8abDl8xMCyAZBEBMsCQLU82yekWQHWSRz3G3gweIu5IpyulUyuh5W
vSaaQQsZz1wqaBiCG29MKyRSZ41YrjeN+syFUs3qCvrFUcVUS6+JIvio9vAykY+p
zA3E/HIGSR0mbwh56vmKhGBiGdhb9+ZaW7hv4q3mm2ueuHt8EcCwaC/2UTX5z7te
fLcz3xqHI8YBmvFGgkqPDEqn6CdQaT7Jzud0GiDcnttLYhHM3Wv5G+HSduCZWWr5
Pg6MDqI4ixOa+FwyZ+9r7Utp5vs6em8JdDHL+DDrA+9scq3DuA5RYQHTPI5L0t3c
WSg3t6jt5joDsjxo+dvWA+RVxQ2ajHqckCyWQl8jeiMsjxDTqqj9U0s5zJawFx89
fKzellMChZQWXoyrLjgd2EfsmGJb6woy0FKGIcL7OR2cRJpdxzMvkEnTjDaoD5pv
KKqcWeQpFeI2APLNoZAUGjniK/FX8EYvT+zcvUfUPRoi1D6Xq2ynxYGaQAIni8Bi
+ZvxDIexUU+PNM4XR8HZ2+5Qi4UFwihSGyGmSATWhF3Xtby4NK66a97bw3xWZw5z
pFtL9nAYbzkZHfzwvdwKTIHLyCCuJgdplKs8stequ++ai+8DHkYU+PdezcHYCMWn
bRiRAzEh6BFANH+JzFvifFbspoyy6mkkAU83XRNPs4NPS5AlWy10zp2PujwD4Khy
LGU1JuEBN7bL+JLdC3BZBPBbI3m2CxuBPUvoBGajAC3EKTmhTTdEnPte8cSyB6Nw
BDZRpVeqaSJMrME/baRMxiLSnPxrEeKHcm8O+5uLSU3pzngrWyidfKTylBjPv0nV
inv9qI58+nYUza/BIBO/tPos6J/p4e4ZLRr+am/ZKSVKUC9D34tetekG03lFWyic
42OJhns4312rKrxY6usmu4QSTxLbR5GVJBN9aC+f+4Cz/uYeA7E2JAMrih5p+wXf
Dhm5HbMro6BEwP0P5DEVYQdSiVL+EuJuzZjK16K3E45y3KwYoWSqTth/6lTZcrP2
bgA5V5/z8VMQngJhxW1IyPci3S70IQt6xm+JF7PAg76SzpyE053HmcN0bmngE5vy
Trk61OqIZwAGRxeJj8ThF4WuUVClcu4bpuvdwKRNp2ypu5AzjL+IuVKt4+3aNkme
azvaOgQxo/8oqauG0phhV65B5/BijAR87VUoN1mqpk2jRg0RnQErxfeXZX0eQBNr
/MwWUEuBHQkMus0QinYNMx29dT5u9ud1kvr9nJyRW49m8A33qNQxYtpsog3HHna+
aGySIY7iDptUmwmbhIJl2IHibHDKd+N8EM28R5PdNbGXwj4rofN/ktOyJxNwXlR0
dJ9LXzDjeYFZRUJx8K44XoawGzYQVGfcniOXr8FzjEyS67VLmV7S4RK9Cmwu0bOO
s7aWItlKUkUtFLIO/IlOKlvMmLqf026As4wTPaqP3aThVnS+op/B8INT/Bs9rhyw
UsJxzKvbJyGNNOEfrM5Y7Hog/EoeFcxRtmkE5TV+9GUVsssrBUC/Z/ztHdi6WX+x
uVhCmYUafiwq8+0VxXshQBy5NdkBt+CH0qZhNQ0qa75eMLiOCSzsNgzO54R8df1m
R5TD+AXtazxlc3WDlFmjcd9eSu3QamYkPKQ5ba0hV3p1ERg8sHNA2iC1hmnEldP2
GV8IlFrZ7Hxzb2FgYwzGUIFsPrnAhesoyaCUsSDh2O0xtq0zVYEw+tZ2atqTphZd
vaArdGCY70QJidQIjTn4vNw/pcsgYmOoN/xEZxgMiz0ZT2HLcxQNnUOO+phST7pH
iyEBn5bE6XqZ7lUg0aFpMMX+EAYUO4bdrVUMDeCG7aXilvDqYlkzfbZD7jhD0qB2
GfNpVJtj8cx2YDNzpRH+sns0O7BsqOJoB2SeEiWI3R7AmPF1awVkiNIavBiHtYvk
7n/tkiSTW7vystWh5HZWULgpNERkTCxM4uXdf+KqOZVjbC4JaYQiRglHhbG5hOxj
v+dz5GW74JdtrVXCXNRbTCZUNQQUD621HWrxj1ykLpnJMmQYBBCWbbzUpXAcdTmL
yAM5QBxDIttfKRzpzLieaZjQCuJAeZjaPjK9dcyZPliGL4xp2YdDgT9oyRIkKGfj
D3jZxq/qnE8r1/OAWiisqt5iGerJSHgfiG2LJQJAeXqeQaj2GEYmBvWD8OAuaWl1
Uh6sKF1QOpqPgUvOzWtl9yPYIh9uDX4vBNju51sSqJREHKZCGDp8VIb5vanql+U9
A8nu0ag5i/nbkMHl/ZhJ66ZGzA4XODI8fWN4PwA8M0aPreEVG4h+anPEnjnEK8As
ybTPODUotS80kleZf3r0K0OgGMryKl6wqUpcqOYy7BR7jlaDy/VMLbiyOjRzVzlH
UCszAwVu7RnoIqUDT3P9Eo2j7K2e7b+8FGAIHZa9Z4wQu8RDsoNEVSvjP9Ny0zET
L7ljSa/BMr2cRS1l0ZgsqOrLpjhRAkDavv1vepbHtb4kp+Np5DFeZFQ0u9HNQIFv
OaPgspy0DIcCELmCIoLq1nxZe5jiluHS0etUHApiOCL9gSZQV9E9bnb0nmWxodR6
OosED/1TPmQH0aDy8cHSaAGULHP43SHDdHKYKWy2TZ62UnztiIPAdpST+Lno+AIH
nJ0Pfpuv85DEL3G3ejKMHzTk6xeijYjg6b8LxDapvR5skNUtrPmPbeebUyntfPp5
jNjJvH3GEFhQijT+2ku1dy+UEOMnauaQExW8a+GMuAckdwOkOCWol5UUCu+OlPaQ
jWmRjSPhSjhK0CXI08O9Jpw1NCEY9AgqowA90UFL/Z5arab6ts4CIiPrPYnsFiEd
t/kUFPX6h8MBuhuCTLcCb3OwYX70WbCD7oH6zJuh/Ivul/3dqCy+gcAQjK55j1mt
DV0ctigEzUM0YzGlYoVjjaC18E2T94y7JYF2+v2d1NtGy1ttfc1/NOI0JquJ4ULy
DDqAUTQ2cJU4iIagzAIxMPKitY0FK8tBTPDrZ+wnBg7Uyg/fXxQjIxK7fUg/32Ym
BxABteLP6Cvn3QEFWYW0cd7iqQje1KQh1Pp7hO7Jaxm5xXJRblCHGUmDn7QMI1yt
hH/tqEyoF5rGlwADetc1Qo06uSQaJpYEF+Mvq73lVK4KwIk0gowh5pdy9UYlosHl
iJ5XNyKPozqFxwqKpoXVIGb6qR8J3jtQCYjkXzGD3tILoxn/U7MAyA6FA+nK6ZIF
qqmSCpb1pukgsKpcsX6WKxzD9NJxIk1TWpLTZTWnabksJcO35BYy+Q2ed5QUWL1E
mYAo9qpB5WfhGfylPAgNid84KAHiUeGSESmSwyy6FpexhYKMiT4Pw2tDAHsC8iFV
flmzRKPk7ny6LUhSd5L4tWuaam2m0tLTUH7GziwFo0qZmeiNyrCTLWAXqX5eGjkG
WJFtfSVwOxGtyODLDdhhvMSilc5mwz6zIGyCDU+8phY8+Sf1Ov7y9yaJJ1zR60+D
l5tUpAjdVAqA3+5Tl/CZwm8NwanlDQawJfPyIltSaFoeNGIufDNbUQzjXz9UDfCV
J4G4WsxA9S0b341YdxTUyuvsJhcHVZyFc7ZQHar9jT0CRGCDgj/94FLt/CRN3tvV
vpQemxgOmzcJoK8Yw/WATEzgKbk27JL+tJaktVmU5aYtlh3zQLq3BXGTVC4e8UFw
xupdkcYdDztVJDeu7681gfhQTLmU98AqwCkjK+NbV7R7U/z7U3eBNwiRM+/gUcON
2LoRoRa0EDXSyIdJ47+4xOQrvf4QheJ+3jjVc178pdNhy6RccYlRCAgCeVsdSYYF
vT4M34XdqPo9GaVjvE7UHGtlmejxON8usm9ZfXgl4X79yMPoz8DOC8MVo9wj18K0
ooSo1sW5Qru6SsCuOrCGgeLEvAAFebUe1/MvsmfNXFwEV2gqnSQB6xmStLPL/dW5
ZKzFOxQpkMK4c7ApQ83SDHXZv0uogBoRWHRkEgLP2TJOA78osVNqQBGsLpcE3Aau
YmKYwMI48o+mTtQOPItKMQDL25U0SOygi7xVlZE1ClURlX+edcOCxM3H2HfpOQhg
6qHOYuN2Z4lqZnUEa5z8AdKYRhGeaO9bf+OyMHUU4TJB3wyPDkrrqYCrVcy+6VRP
S9YDZAsDWrFqD3hpl346oo309mjHenCUZ5ba3COIzZl9jQBqraA0WNHWe2Tg3Z4a
gnNEMBjdQOPrBSWKzzWo6yA+hoESlP6v0WFpWxf4y/HxnM/QLT9cxihTyuDLlgYo
Oiw3+xaIGBgr3+TmcO4vferi1WvnHqwiW5ekl1GTYAoLtseGZM05HqZKhOppUelN
jYXrGQhYVJaZv5dr32t1cTDLsZBxvnx47vk7LtFerE24UFk3BUA7qWy8PzqsgKyC
g6IGzFYsBhcPjRO82EaqmvLrFQ4YHXzD+mikCJBSUksHvd4QXmUfEvXtKJkohBFB
J+bend2tGcd05oiI6Gfz94a3RCOaTzdy+xOaOkH23G0vLGFnpfdSsIUETQdg0RJ0
STpy+E0Goi7P2FiuGb0HZa3/tuIYhYb6n5gWaaaiYVKS2ahBBsTdoAHis+toMaEP
4JAMcK4apCjAZu0lXljrolsDeFW1UyUolrGaHIw8cLwu5pZI17MWOyaLeu1/4f7L
gVo6xnlvmpzxPF2W7wKt5io2su+JyqAb1SE62mGlh1LkWZlLAX8NsOWo3hZkLGzj
Fvddyn0k5+QBTvu2lhi7r6KdEtcAceT6Lwf8RXkmvAoyv0l4oOcewqdO/IPabqRS
cQyDs0KLAuqsMAjz02mGvGo37EJKjYMxSmjEieTxzLz+yJ1K5QIlDLynYv9vRvHc
9jHgUqwkxRGKxbu9u+I7wjLP/8RGJVBTygAIyP4oRlYu1OlImtEYSLbFSUF/+5Ty
SeauJctQerDMMXJgdmT4q1FLIJdGSqOZzE/dIm+mjeDr+iSpKJRV+YjdzZA3M+0g
BRUFCw1cm+jm0QnEj9A5fqeayID3KWVfclLpckiEZkaET+wXxF0u0RmVqxHAGrub
1Ap16gRPuWWy0lKavw3ahN15uverV3yYvJ248AEwUjSssW+v+n8hWszFgXWgb5Ga
qatViJQtTkooHsOVs2c8R4nmNKUJ5ZRXIeEwJ35/IPfrsRus5ss4QoZNwCszWBYO
YDdPoxbTSa1iNIt5Ls5oBW+9TB7oki3YdsAQPJe0uOMEXFuZAVEAHo3XA8c7ONFo
NTaXnWxfMCQtaCkQMogDk/T5ndX02SvjhX5kpq56SHBAEk1WmBitgzI7CzD7yni0
9Kx7IpPr02HvQ7PMCPwn7CpOabjoVZJXaKq+H3oFw2AjK9Q6hjuc6s81rLu0hXv3
yJlzfhT5VP5DgG/1I9GoG5TtUMWXIwqm0YaIYRPDc6FHBN8qUfVGEl/ohigLClN5
re+DzTEbdP6gsf1fL58kTwKd6QcNoj3ZhwNU/1T02Rhf7KIAAkfOUByoHr8tTEk9
RUP85CKRR3FDrs4yJAi2fdTsD3x2FOyGhyKfUik3unTRLiMMDtZLVXBFPpnKto0S
JDjLduYMv3Q6/OAjn6eAghPHbqpMKJiIW+RZIJNXuGdgFlUSwqGRjjo/t6uY6lRn
xyhIYvOCNzzh54rOlYKyuvxqFXsA+E6dBEejyP0TtJ7woS99XcrzGj6DY+hl/zyp
r/gOC1LvWCWzVjVjJAmK/OkA1FB6EmeWUgHmRtYDBJXLje2zzhF0L85UJ9DGtJ34
486GQWDmf4ScVwM6/DUdMQzfezaDNKE8fM272Ql490p+PmBlwlVy/4qMD1ZeGLPw
E4x56Rh8cFPEYuktkaLtYYiBs+OKubiCrwpeY/dKWcR2KHFws7gyxmRk9iv4Xexx
6Ph2oqCeoRTPPzPxCQMbZdLXW0yUEgAC+5dad0V3L3KaKZ0V0w3ZiB7kyvF5hV50
8dz0t9mrZFEnWoi/1+KqJjii2zAcDlUx+hkCznkQ6JQEcMWWAOhWtYWnZqap9Xy9
DJa3n2koHP3xnHpysTnRoiwop2ribkRKSlIRPrI94f/Nriei5DRpyJygVDWR4Ebp
cVmAzmQuOQm7irL9d8s9qF+WmIVWz1emr9kmQdsvFEkF6ITXjNpodYMAKweryfQn
gEA5XS9cEd8nzswMCAyD+t6QWIlc5wm28gnoXYj637sXhyBENfNKGGb9rNpR8qrV
TF+kVR28ZNh0Qc8y30zerHDXYYCFqhKQEyqqwmCCcf6k+qlsHjkIwTSmgklJDKXK
xTzqHxuqQ6M63u154gwYpRIgL681HR8tdu3q3z1z7erXXz5hyzEDcE8qeOSwoep0
2XstVROLIlbFtYoQuofoasGiqqmUSVPnNvq+ydIUb+DyIVKrBRP8zVCsHEsxIHys
veNK83THNgs3NU3rYUV0S+p1NJsONNHf/CLy1kqna9HUqw4x+Qky8m8NuVL47liC
ej7dGfuAEn7ikkohfuSUL7NAWVlAEgsCUu92VkqypevaV7BrT+dT0J0lRr7DrF/g
2HLlZ0Rd1Wq0ilDTDDN+u/A+n1/1f1ORqxiLC1J0JcyLssuW84PYahV9xBqQiuJa
EndfeYz7UKL3EzCTJ/cwkV0VjH79IQVWFBetn8XzfnWXMfqO4nFcVzvpPJbD0a9G
MKFmiU8bEhAHQtOSFy9GM7YgQbruD9xeh9CFyMow6D4CovL0UpKWXSBDWBm93p2A
7vbV/oZndL7GJdAMPahxLfa+hGvPeF1WtJ+LGtAfdbVWdH5huIeA+oelcSHkXiJY
KORPJpamBfOCfM9NvbVZEk1tJ1cqSmPDeAWfBwu5DtQ7i7Mxdog/nQ4mAn3kw2XV
s0R92Zf3y2P1f6fGr333Tzz5jJ5gXPwgYtc4nUaZ5M70ti59V4i72ChlZSaMOd7y
SWOB5ww5b87Tr5442cR5SXytOxtOXIIVGG+8KbFAaE307XINpWMMWjfMqX9x41HD
UoNMrh3ud5mNlQJhpUmx8UsknJkDRg14wbrUKavJ4sx1JHeA1qhL1om0JQ4uOrTp
cO3dRxT5gw8lw3ugj0tpkLxHRoHSN4lrHZkU84A0P+Uaumj8eVRFH47CdxrqcvN7
n1TxthyeKaoGR/SVMVXePP0eGJPMJIyfdoIoYoPisp3VukABqoEGRV2NglmFl/h4
88uj6Udem2m7qf8kY7Vl5QGDVXRkR0nDVVQ8oK3gS5mFBts2ifxvE7sJ/3SA04Hu
AZ0FZuXT39JdxKMnP3KWkR5q2EoZ4h+XRZaIKkVDhme124oXMtKgX3Dd7cdXTWYX
E6JnmVnGHst2fqhQSwG21sf9WR07pGvMh8NsQIYPOEZ97Lzn6FgK9aqth3mSkgGh
kNxl262emtK4z8rG7cCj8M1ap58lSh5Gn3G2vlAlyMjVstiSdNLbSUHZeBhhm34L
DEq4lcosHnDT4iQIeLPgums4FOTYdO7pEdAQgdhotUcA1lEOSQXhOBQEIJVSmaqK
Ene68SkvbYnIXcaKwhyJf6PywIwDcQJ171hO0oUVMPZzdIc/qFp5Osj53Baw1Z/M
ZftXHEjV54dj8zU/+KiyPUfD2XmWRGNDNA737L3GyA5UjntUAn9QJF0WWj+6WGwM
g8XfpvYLa2Ts961JZke3vhPQIrFDJAgWGYGQWeYRx09tA7xZbedG9PL43wXn7J91
nrtXln5XpHkyL+P+O9tielJAqFVIPWkV+J86XS8aeg0eJg2wuLxBHGxvbbT005Tp
HbGdP2531fGf2y7C8N6gAPP/OhlscaMK1Em5hFL2opv92M09vnhDKi2IR1Ivwv3p
ssSzWYIKXnxRGKYkUGshADSXbfuDhNj8qAa3gQVgOksQMRAcADv3G8ajU+uKSTkX
iHpBjEoshquUEbfblPaXCvaSFR0ffDN5j12qP6QR/OYq8rpgwhMisouH0Rz8mwlu
8Flb4FT8wDS4gYjuP7pTnclxa7npjQaXjjp5BMhdX8+b/nkbxHDnRvxdQfWNK1zO
0OTOVBxbg+6KtwniFSFxT2e+O3SApj3cFygI4e37oDj9UAPjMAdBtXkB1T09mzpb
eRpzXe3MsLtd7+4rdEYV1T3+7uXBHfRKyudan+7R/pHZOno8rqY2jIhuPjqYZ1em
mV91Dl9c55dvXX1t0rityoqnguu6czwW8aIn6ggaDyzTjuiAKLCL5kuEV9BI498P
LrnjJ84vvlij0iVwzRj20oAIcMHXTYpjkpUCUu5ekwxYTA9e80HtH7vAMCXvki3d
jZwjuHT/OhkmEbtsVcS260XSmNsmX2o4255NIdHH6n3cK2qT46ViJiedlLe09IC7
XN7CWBRrVa8fpLhhnd23LO+3M14If+xSE36HD4uC88mSfsxrAkldFg3th/eWGERF
tO+yXdg+uh7ym4IXQ4mcOc1iiv+8pzZ0PHPCKPcxJNjo5/T5I+4jMmFHGCB14Hgw
6/Sw0SoMcwvxADfGwXWmSpinqKSQ1j4O24OJE0KZL5rIhiErM+4T3KNVYc4Bz43J
A80P3klL4SIBHQetWndOvMfeyrLKhMC+YzN9NX/0XAOzku+jQdyVnLkkxNYqNJCH
MzMRCrPK0G7TKCVEdQr6f5GhQ09tvwVwmVryl5xJZbsuwM+3q3b0Bx1WNoImlVPn
0p1BWhaEiKJay6hyfjYjtTugpEQATNbYIjQZVGllVA2WBVPpgsvsImEQHD+zW1rc
3kcVxpfIcxf0RpYScgWHoausN1WRxJgj476FwEEn1Sq0FA/UnjmHeyVaUcdDzi4Y
i9w6YFOTottvVoAy2OrlGxulhyWeWtMvh9n0psN4Y2GhPMI0q/lJ3yWGHgUP1Fo7
eOHA3/vrVEc5LgzVEdgIGAcHYRjp/aq1NFG7DpTfRpCluAlDV+EEhxeF/7Q599h6
M0C4VFgHChKrvACgrmohzpff1Z1eq4bBYWy3KooqZu60n9n+2CDqWwaqJzb0fSvu
Y6B9RLl4yhFQrD+wET6KkgV+rItOljBXB6IvdObarudfIVnLfoIWmqMBNe1NWGaq
Obt2KGFskEtpueOyFHS+lpu1NzQhbk8ceNX9QCZnPqRdwfkB/vqX/yKzqHLZ4hnv
V6ncHpUTEyjk7j9QJWySZd2s3O32m4hVD+Iwph8tvjzby4qbJ2lavQW2zxSQJwep
GbxrkKbowqtBIJXvDaOq7SPW1Xlh/NH64aIfP1jWwhqoPoLVpvo58YuRMKeaYS8h
2HOy1aXHIm30FxKDhQGAPvfjfb/L6bRdyU4iLlgnw6vXaiHD86r/yPXvzI2SpzEg
pqmxeP41KMyxvw2BtePKEpTOLcxedLAbr0JNUHVvgJo6NNXqDuzQKDQ4saoJ8kCQ
1I4OsK9oI3bnZz0U9/jG1tvlJVd/Be/X1fpL1xJaFhpbFMe8JrxTopWABychYisZ
mg87u3tgWE7M5K9PyI1mCV0ujPGf4/uF+8ci4pAfbZ60gfuqrLtQRLWsInoYdY8M
SkM7P2zvPkok/dUIT17SkHmvdeaEqRorZT1n1vJHhP8kY+7xCibygsLAKtOnwtaf
1cLK8wJE+hJWlE/TD6u/2RaNAmypXmj7dU3G4+UgumfTvh/SCwc3HJMdqb7eILZT
IUsucXgAB3JVeBVF6hXyydkQJlaze/wyqkPiSxBbUsK7Sqe9BAEI+5WlGVgsDf+0
GiEg6hmXvrBcXzl5n1HSfn2jM4bL2lQTe2qMfEPuxRc12D8u3LeUAo8CChFCwzY7
1/aTuEmk7mvS9ClhGEJTm/kWpVTrHMpQOpMlJNvZoGcIsug3it8fFDm7AFiRFxmP
Izti1IlrGPUqBqyDR7sX5dNcqrr9AX8ON3wrwLJk+Mhivy85+HLckThgp65Ax/jw
K7nklcmO5VC5u2/8dZ46DhbCQaP/stUmAd5AABQWoIJrBMIcX/7mN9pCDWMluvCK
ENAsfZrD6j1X0iJSHCgUHH9SXYkawej18REFex3HTi1hsU9xspNv5Tt1AhzmaC06
Epw2Q+d2q0RGAVIS38DLggmmY2UUxZtYE1h+O8yYu1EdK+qeSBLQoclVoz+GLS2N
uGxT+3WoiO4tmy6ho2M3s6D24KVL4nEV0rsodZGd8RO+s1iK69jAYvljcUj4R0yu
gJCVQE7sZzjnMU4CTSMIDyGhcL/z86xf1SF7ToZsoG3mjzo5dyZsDxTWCCSv6GV9
69y9gvw6WOfthJ+KsFIPhDNIyPrqYFepxRId+dngD4CdJbEP04suALEzdpGizwCG
TaeGgLxaIHol7tTc38AHO6XKh9EvGgZKyIHrvvaIr4ICYUpe7061W7LAwN2AVGmK
6nKO5aZ3WRaIbzyLlyPkRUwUpyBrAUIkhs+WJAWH14Ynx5SAhVWbEPrzNRF8NQ1W
4hf1rBkxIM7ByiLpalObEf9vKyMbA5aOrnpmwAd7V7nyDodCW8pMC6akdqAxsuAm
AcunJpWp7GhtwpQFi0N/QKzN+HkLtoqX28CSCotAJjqFVMkfTLD/UilfVJnNfmfj
+r4Qq19TISg/zHStqeQDbo5U86lbnGp11b42o/eKHdhpizWaT8P0UmlXI6X2UxvG
Xi+315kbNKCAPw5W2ySoQiIL9SLRnjGgnExWY2WQv+gf5cDSsqnKg0y76pB9uEiy
WS88zoJRp0LslSWftilt8JrkVFUh9MGcN78KvL5LCJRbJx3N37dOfJz3HgNdBc2k
M767KOx7oTCwsLRumVCdcFiLWeeuDJl9TMlvrOaB/qSqoKORwAzj5qB9NPMJb/8B
h+A91wYdSh1BWMhAItWvV7X3KD/qkW2mMkBsXQvpnuDpmpbefQBwI50xVYVvg0z5
YlhcLiDFMke1k4k/U2uS+ctfyTHeA+JM1AmyW7mXn667SSMoDuecyYwqRVpW+TaS
VUT6ZZh5A1459vf5eJ/PjwAxZpcpty1VW2m5MEeT5y+ndMbkHtrmL1c95AvWKzJk
Dm0s0lY0cB+KoVWJul0qiJu+18DWbXrQrMUDpCPJ4DtDj2J46VTb3NckVHJoOA2D
Yqf4uWS9maJViXcptf9AnrVfDQsh+qivzXrueiqOxX0EIzJzSOdd54fpz3lBCGa1
pC6OpfSDtDiZr35bjwdR17v1t+L5xilfVS393DzVzQgZnefjDEXdBl3H6QCRqtXK
cteYPErV0rFwjE0+Izdwjl0RTAxCFjb+tL5rWEOBITMiQv7QsT/nbnXYGujQLlCv
0ZujdtyNCBZvhV6Bs3rCQpAZcUWsUAPMmmtkpPzm6DjgUaaWk5UZdjbqu3pFDPlC
9ptWmlrs73MTXxPkN0EhpjWWhsB0akswDjgZiXa5YfveNSfSk112U1cATAodTUnA
x9vhrq3ZOqbkPh0ewdTuCF36RrYQsmUooaC9xDl6w31IGsrAh/rXbL9EfZr94TZ0
JSf7Zs3YN7scGnF0EzHf71fSm7TyLR2SN5LTFPEY8qhqKYGRijy9NjshHSaelPKH
Bb5sSK0vsbtAcN50UdvEig==
`protect END_PROTECTED
