`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x9/RO/DVnMNYNfDSwMDK6y+QgbdjCKSDrksHlRORYmlTFLf0AcMBnnsjLYna4yhW
vlR79/w+xOYnYfc/RIbPcGD13K34BdTmx7Gff0h/P5c9MuQzDqE/XN8dt1oJ4xV0
QDqkf6UJqU2jyHsQfR4n0nKfKERr5Hrsi8W8sPhcUKE5Tl7XMVjjJQsdfd65Mdxz
2XhLwG9yUfQiVyNAkCia2XewwohJORUlwQkKUXiN6XiPr94i6K6ohuuhJfM/f1Og
Pm6+rdI1APQ9L1YhTHjap9tciT48ZsLivz0keST/geyyMX649sW6kCGe9c+Yrizl
ew8xd1XRuB8O7p/9HFFuO4oFuty8UMUpXoAKhSueLOdz3sxKBfcgtgsf/qxF1754
3xk29s3e7KhxbcqbieeOU3B51qO0raI6Fb+2oIAyDB19VShe5LKJuz455HJvMc6A
cX/jOobglS+beXwG+pqA+7eMIH8i+td6zdPyFaAimwOgAeYyxaltaRdrmX+j0qZS
m1jA2J6AF0FKNo/UjaFI6w7BEfU/1mK6ria6WAx4qfJK+XIABgZNX9tIzHqZcFwV
+lCwox7jUi76GcOFNsRNU4zHZjUOhoiU6iAS/DJuHaiDrmPDeJO4N7PUWoK5RGvy
xLV6TWv3ecZcvCWdYkkaMvSWYt98MYBfXpDyKSTD7E4JEnY4FC8Wm8oLoLwn6DNe
wn2LaST1xa9owQRm57Rbg7HblxDKES95K6owr/ldzi7BCD+cGsCIJHXi8G3raP7h
5IsnnWg5bMVE3i3tH5/RdqxVaOF4+3aAagt+t9cN3MMZJhmGOJGUZCce5C5hlNnx
6YQVsgrw0n3nGTSvH5mjsGE6Fa2tbUiPbwNPyshVpJ9FWVRVmCSWSLFXuS1o90vo
kZGTeeKmTScv5Isjxahdi3hOA3cbyC8ms02RUPx5iqc2R0AA5Y8AFKO6Zs0qNwEk
110lQ/vmrhSNUKji1R7Vb241eusNqJZDySJ4+ct71u1WhdBRa2rONneQe7Y6a62Q
ahY9xUz1TrCkPJZ2od5OKSXNKn7eSBySzvNMJyATkDzB6p69pNbkZmC/B/ZQqpDK
sQB30Lfj1b66eGCRtOlSF+nfYF7vfN5Z3IArVjvM3RL/6ssh84SKlV5bo6mJ1X2g
X4YIEfJ3rV4ZNaSjNdmMQVVdP6SojHA4dOXrIM8JiXKBbz7nxEMVs86VJqEe1e6/
3Oh4Z7XZYW2Pc0MFePwKD7Upw8IVn+mqv4jeYgLjJ2LypmDapbB/b7wzyzwQ6TDe
Z9vgRtr0CMKRGTbjTppEGInCEKb+GcbWch/lHn0FQNtCphAGmC6nolO9WHDvQJ/8
x6V4f6F6j7BmeVhQGWsxumqC/0x6i56lcl9QficLUcP79/GOFKa+HVPuLpSa6btd
EMFAF5kolHPX7f3erQhwZeeKL6iAmZuq/ZrQgocEGYun6STaSD/mOy8MoxC8SUKF
XLtbORBtxPdE7gHa/hQkvh0mc1kRLHbMC15/6X4ewhtbhYxLvzvuZcY0uDnGJ8a+
cPjV60Uv8rv1LYmdtNdcXAO4CJ/YxnmZ7knNRCY7jKbeCnd1YWmRFMvEkpshV+eR
1PG8xfeq8deaScuUddW33HPAwiAyJxrWMmYU8+cVFK39PeQ4QlAPTddRXLpzHr8l
WVksQzkd/OxdIsehNYPzMbPCAMlTlPVpFmAJAACWFj0NWB+RfvE5y63eO9D3CSI+
8a4q18QeQBTMhUarNV1N2SQChl8ku7JH//jbwEwBrSQyTFUKUBGf8LUm0+c4dxSm
ZABYWpNXQAPisU3HJUtzsHNn6jut8xQ6PN2MBhR683UOFLa+evHjo9LSrQ7UdCEi
9oTq/a6pyXcH45aj8VNLLcbs9DH/QkQDcoes73rS+aRzmwEMotV8R6qh4iizkT3T
iN4DFqsgst5UJ91c47FMbI4aDnatANe3IhBZF59jG9V7m5hCwvKsyxP3niZEBsnr
2wVqILY109SM6eSslDXDegHpNIJUKpaUuAOkvmpnJkyGzWzvxgcdfd0T2CszKH+8
0lrF+HOXzF/pp+PV3EQB5YohzMwtqsKtF8AG3i8GFPuomH7jF902e3eW21C69ba5
qZg5jIXQ+5e0UU81x2TPcWIFzZ++0mucBlNklJqHsAsLHqZYl2KUgAP4UUlVJ5uP
hPs31ZwuINp7rrVprVnO7gnkKd7hhScxRs4w+T46vdGGp4indoAp+G4WMf+h7h8N
eH5zb1GYLVtL3+Izz51H71Kc1KzVpz4qt+ptTTmWfzvvRoF9VTc/xddZnJ1cZHhn
6U0MLwhZ8NlMnXYpaS8y2Px9yPhV+vgFlEeNDLIXq4GfJBd4XEEDi6Lmie9O5KDA
jn2ntzD8dwgytfkDWXTcMjCqd+xwRABH1qGajRmKP3/pu9jkrhWR76HfokloQVKx
eMq2ctc1mus+FTQTuGtmFYJM1YKGIg1DLs83ZWgjDjXhH7Javo1U/hbZ3FPKqVq2
8biTY6QQQea8ZHjPQou1wVm8jJ3WwT0AQCDOS7VDEDIEoijvqGHVLnuTYXq9WNCj
XS/q893p446Z9aDNigIlXS0uADhvfU2Ryov6RdRfJhkK6Ou7ru9ynx1hqoE2Ewnw
HlzrQFmYhIhpHiROsUOdPvC5CiAteJkVMK3ukxWcIFyNeakgvzOaL2y4+BKn3BmH
YsNDGry8Ise9LIB7A62pfMAIqOZ6de7C4JeIqrLqwNpM1hWf+9Kg4Vd1+dZ1uXsF
Kb4K3bUWWXWHCR1dzrqtmjBNiNHaLHF9mv3RGRcW+2IBLpfo4078HWSEJoMiSPVa
OaiYQkTFMs2plzodJCFmBXEAqS6BEqEHJeradDrjehWnQgh7xO78A9AL9RyDiJ48
6+8xs/vw9gMSt6VrnQlxDy10o/GuzoeCDf2RXN08f23RgRgZMf5oMyticmGECIch
a7jemGBAo+DtZ9i90Tcl9mm93d2CivOHuZppCBKwwj/AO8p0jNgBvBzKKFmZQdvc
c2ypVONkFr9dAEggfXIYXPsLaIlUdEqAn8vnZw5HaccOOFWwQql1+/J2yS59MYC1
DI5WSl5fQrfthSnL+SqDzn+8xu1pI4TiemVBB5c++TjlDE/KdEiZdJcs7uYv5dji
sdvQ+7M7gMR0fpKfPjUsL60lLPTN2LVa6CKfFBujEKdGo5+aurcKJcZNkrFMDnY+
DdnoEZK/wwL2qHupqaFOpcGMkHmZbcVoHaR/H3U+3psjKciaAIubh9vqrl+yzGNF
IFAwJtEmV8dgaQZEfM5C4yS7/gj8sM2HBreUNighv3Q/XVuZUCmqzTpoWvYJNZbe
BSPFVflSlDjtFf8PimSHO4vHjIZJFK/a+EE0UymPO5oowZll8S8U/G+HbcprYnWT
KqTcVF4LwRueQQyDrM5sQqIq7AJnpqQwLIBFJs1/+XdSPmhlV0nxwCycd9mpedKp
qQVk+RtAdcr3cXlxxCQdhkKGyZxFioYKRV4kfvOEzxew69TtKMZU3ZyUGK6JPUCf
NOhDvsNrk/XoRwuBnjyKo+7wcyumaNj9ifKNts1XYl/EvV7BxTtI/2VzBGBebcI0
IAygsZSTDS0dhWTZJ9zXdTfI4MKwM2ZCdDUS3NHlgqjS7Ejj8WWrHuoEP2JYyFYN
v2+3ehmJXmvVhcWphmXZxQhFcLPVpt4LEgaR/avtXf9it+YpYw6wUoIhNxUOQEjm
A2r5geHXSiFrllXd6AgnwXTJOBlRlccSg/KFH4zyZTNzdJAj7aPpN+siH95h/PSf
z33mhVa6N0fnC8R2e3CPlrpw7TdepX219IPbYZLLXAPvGdgLZWcrVk+9eC86VMML
++RIEcbIOvakBLiYdZ5LgZgaMEkP7oqHr06snD6oZO524+32UKlHrzxVSDnry3Xe
aYeBdHGb5JL3/XIcZ/Y9g2MqRnDw0oo/SQR3nAV4X72XabrueQKoXrdbIpsvmQM9
wYfUJdfzKZH/ln1OCUiK8EENIt7t1Y3ixcRDxVjiP0CH1zEEzngnzbR8AoiGTHvC
j+Bc3Mu/0GSMFJ3rEJA7wsp6phScARzYjWeBpJuTPkTugbzsXwxCnPqtfEAHID38
AT418CAaGO2YEzmtmP2FA4FvY4LLOMyiyyB0sSIZ/xGOIVxQ60ke1k3Z/9kauYNC
y02Bhk6NGIfb5W1fI1K4yvwVn+hchQ6SlqFHmbQzkc0aoGA1UadAe7retnZnfGrD
N8uXmHtWFTUiTfVXnz+UObfk10xPrCAWoSuoAGu//GIBLdZf+65a81fvVN3Aj9YD
Kcw773fvayR01QBJPFxAgS0lIEGk8vhK08+OpvhQ8C6fJFn97wNehIFLw7w6x/d8
K+NF/BhhYePLPu+MgaQEG3S4VuER+IVEsFOUu68OKAcW3FG2hFgfB4zhL+t5JbYf
4axWNdFv1S6vkIhGHoZgPqUpEIPmP+H7SZPZhdjAyGMkMlnU5WnDeqvHzYagv9dA
NlCuGM3JYx5KXd055feEyK+M5pMt0XT5KY3TPseoJHOSW+aUMIv4/XBdLPGTL5L+
jOPHdvr8ViyU8U3OpLOiyb6ZGAY57LdJg+pmZDQlomzblZ1Id3kvHmQEff4sD0P4
xRmrIqULglfXZavpNt7jeuPmwsqz3lPDNBKJq6EgyKOhK+kLtR29Se6xAgqjDJ4N
ozAVRbxFp1qRYRhL1ibGBts1D4+QN4zGKDgOi38yLsk=
`protect END_PROTECTED
