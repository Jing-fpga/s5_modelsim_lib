`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XM3H7ZuzayXlovAbtkP8Io+aDPBn9htEhrVT5POOxYJfG0ItJbrnkc00y4TjGsZc
3vDpJ/ru5sOucVJEHH/FHO2rClgfjgfuyoIXT1lpA6FJ4HuFat/FRSyNtXjQYvZI
mCx5BWwFdAc4fAtbdZt9GLv8TtCuFi1BHn35OXuIA92Xy6Cdw8UwDpyPHRqGH1AQ
pKC3tWDCezSMjfqsoou0MdxWffXyPUhoZZzPbwuH7Tq5EYdt9XtAgtbX6REgdG6Y
q95RYE+oKONUg9fafJWVd3Ju4tiuFdRX6xcrHdOVrhOOQt8ng8QurKm9bLaSbJic
jvlpiYZVyNpTsTPblM7kKo/Uejaznyqh/ldtMXFSPyFUNy4F5aVohCExGL3a1h19
HOpad7oleuYgUCRNlSGKS0Bc6KrDge3FXCr6IbI4e2ph6vGMozaiU78wv7Pim1u2
y5F+NY/MCRcbnSmHCFnmpgwt6ztQtsRwgtcORr2vI6/TmcTPgTQSLAa1ibmfU9RF
L1v55e/MX1qZl1ZllxKUueHlrhC6n+q0NSYe7FyFBbXmMJnyo1nt37mBeHBd4+cw
AHGyNioSaNH0LCJ+jVLyLh0DIyLRtO57C+cUkg/MhfYKdrXlCEkQDuafed35tu9k
ErSkSdfr/LNfxv8JdljEirQt4z9Saf0mHmQjXWK5jOyCF0l+EbnVQ3MaAzO5qKfX
rN4t0P+dLJrq09UlmtVnvtwLYmUGl1X1PWGqR3bw0d+Cl1AG83SuwtPJDNIAy0TU
beGuhJwXNDo70JOa9Mw1ytrYOhURE5zNkO7OYGUS4Y+hGtFKB3JN0g0hmBtJqS1V
aXNUyDoaV4w4s2OTriDA/jD77DVsgqMvmIdW7MpRUSuNZ9q7Ip6PNdz/a/SLXyMR
Gpafk5CszyV/eSt4QGCxZJrK7LP66fQARj8OIvDQcIJaj/H38f/X77nkF/5cIcfH
7Ws1jKE5KaGwvzE2dP4tJBk6kR3Qmp9g867sz9uIkfPeTABeSejxIVyr5P2pFHfm
NqyjW424Ej2bvVoj0HAPv8HGknNECRTy+oSrMu73yyxy2+5OxcZSyivY5jhzD5ld
cqzA9srwyxaALW4xpvGyiJjwVFPp/hDQNNsUPhQdHuw4ObLquFMCnl5bX0CH1srT
d+h/sjArHQrlRByoCIrJLz9YsxNw09ri+0/5hBzwK0r8Sr9glNWUFwV0YLzzDE7S
g3PMPptoC4lq2jbTrb79KAedbqxTbWBrm+mYl1Cnz+SHF4kkXtlETgYZihT+xKp4
OjmJv4QRN9/zHJw3vADY8osvixK0G6uPjRogepknv77jH/nrdx58W4/EX+RwXfNY
T+nSxv30Y4aDXHVs5qaAZ5z+0ReNr3ytCATbwgf7XWQSuAV7e518Js1GNUsUVJkz
R7f2dpaaNWdwwGFH/xBgc++8u3g8qwLk/8EWNfJYYgWrRukfdYlaBS91ZBMBbs9+
4XGLSavC0JrUDS0fszK6zhItGcqIQkoXRxUXL6H5+nxovKwpmGYaFTMVu+ulG4Lr
ZmxE3nMIB/nzvuFobNWuCfdBdAEmm2PbGENth1YzBJ442kUT45itDtnwrwmJrxvE
ASLFlvK3k+CUUQc93W+OActkbpnHoGtkko47U9o7tQcUlyl84WCL+t8KtIMOvi9G
CzUwGVJfvBaHhK+zylxNt0ImgB6WpdHqHT9uCY77aVDlBgmq5gGxyre3veoIMKg1
iPQrem1zZnmXXBbciCtqXex/lQTY6ESbR0mpON1HcZhr0+tEtFNE6jVZ4zsggmCi
`protect END_PROTECTED
