`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CIb1D8kk9mmSwdvaK5iHHkkXPSUWAlNFC6HhJFuCcgmM/hEvFtOiVyz07C2QYGpG
D8uBRMYXUQZNn3DOTKuZYL/eYkxgr/ss+DdaJhVYehQ7pX4J+J0MuCq9bpZwASdz
VeyJE0wzL4x/eaGv46a+kBHMqxTnBbiI9oUsXe3rTex1LwtszUnguT1nCpRfFrrZ
HMAP/+PSmAapBMSNiyvlog2rNEo6wt4JbcdvkMe58U6fIPFon+gAQJUFXVdANCye
YUOwmMNgxCanWJuINC/HA/qAes3QXTDC0yb42z2RsN5Ozye0AwrdDS1Iz4wWdfOf
q2oAX+j/aDQkxKCk2bU0zlahT9Z+QH0FXu5WM5M553hZf4G/TV4duuSFUUBhlliz
cudEpfPvBOA4t4dD9KtuFR+H2zeqVtZKDMr/AMqDb0GkgsKJTKqpX37f+QFgG9kd
YtP/FQxIFnSsSapf1g+Q0sPmVYkEYy70/s7ThrswRN8bt7StH6ED3wnA4TjhK6aJ
eeLcOMyPUS4Gpr5ney7Xkragn37jb7v7AqT00/hpKTAw6kHtVnumqgtFYk1Rtm/c
HPrKq6ok1VB2Vg0B9aL0xJ2MZI/X/W5NUM3q2dSTCGtGd4i+bcpQ9xK1D3qt5UK5
CxhBfHpQ3RTu913Nc9DuYNUqtiM/Gl5JiHmeeiI6mhvSQj6v8naEpNpToI6VSRBX
JF6t1ifTNXE0LIwqcvXeXyvDgcd9sGW8rt+4rCitKDtJOM85yPdENMutCJ50eJd1
7ov3xFlgEorlepTgqh9acrNITVCeiQBh9HlFCoICxGAj8HMxjjCU/oIzA7uHdFlr
f0wR7oe2Hzk44z382tUCk0hJDw5LiQd/mdFWaAlmC8kyzf1YLJ5pMCi4UWz97Ejm
GtMPnrBB7TTkOMuByqbkv5+uDVx+YDDDuuC9JsjjzXo0EwOaTrBREzAoS6suWWSx
G1d+t9MepfW9rQ2C9ns0oM5aH6RW+ZevxBdZYKy2sX88L20Leg4dahr4b10rY29x
BzyakjQ3La1WjzukF3kyN6Rl7p/CRvtIgfIMPXVGOLRiUWpipzm8GpLJUZeFha3V
tJzYW9mCT1lqfXZKfs46rNRI45SZgtV8HYO7dudAWmpuKjDoGcWtImgOPpZW8CUc
rnJvYmxAdDzTHnW38mqs0rKj4nzer6nejq4izTih/o1MKoV+oYOkcZSsZxLDHAVS
0iZm9BUqk3CAYMSFY/4vSl1K30uWu62TIh7CatiQ+cABFGkQSwHGrwNRVG78+Ob7
z6zXHD/oUKkhW61+QwO9eopg8HTKRLbmaCOD1ylMMn4YCYZRnwFC9e1pO3sfgjCe
ZuU6DD3Q0I6Xp/n+FQdiZSyFUDjHQeSPubMvaty3kTCHetiudW5nCr6BDZ8KSrU0
tIpeAJeias53wljpLJwSAihAYjrQ6UaPNv08+UXsDdj9lLZwrE02f0Ga6GlJQ1GY
TnpEb2SyI6GI93NiCOgCzT76XPyuDzQcwWUYOoUD4+k8tAHOYTS72kxmNluTjTBi
bO/KnSkXZUH+3TWETs2WJOdKjNybDPCuuAa9tehOQRSLCzvQcP8ER3PA/b5kAHer
sxOjNusSipsqc76eRjVtMvyeH5ZvsR33V1EsYkvFq1C1UnBxowCfn9X7ZRC7jvjh
zHYHjwf9PgC3m6nlVzpLr+yMN0ZkUBH2/yZQ0H0fFQouShq/3TDN1q8YskfYL0/j
5vjr30sQe/n48yR9kHprkYeMyN/ItTAfxHy/l3KSc96rcu1MlDweGAoZieINg/km
eWvO+1nmgJKR+LBQKbmWSDlfBXx1oPY0C17xs+1wljFgWevY3R1KJUOu6jZT7N0p
POpBDLH6pZlmr0D057ZboWk5TVlxD5GCwTz5xV4iev4B2ye5yM1UrAFaD+9RwgGX
BmYnnnLRvMG8964lgtC8jfGO94QaHMDSFwpRvbZEV5/l3aGbPUfln2VX7C9RlKBz
wt0vVvTg8tmNnt5FeZojh/J47bexGE09/5+c1bkxOn+DufgTpEyK1vETDWgv1DoR
kvjepBzlRsK1Yl4WKqzFaeN9VlhPprKG8C9v+cCjlxkbKlTWeRZlXu3Zg2vA+xbm
YaITYul0scuI3EldlaVxqtWcJ3tiNyGSuOdMKHBv8mIlZ5219Skr41cgECGYSlsm
aer7xoUZ35msN4xdSh+R2r99Obrf0wqnnH1n7d0eJlFNkSc54i2HfKnLYxhnK1bI
i6axJwTtADczzPCN47Q7RefSV10UaJE4BIFxKrPwjDoxCznm7fFqzzJxdefot4OW
oghMt7YKjhZ3Bes1rgB4w2ZWXDHzXBjNtta4vcBHS7vNzwSkL2+3aljPvXl6hlVj
D21lMTZ9nNqu5dB7T0wZeS6d2QBoLb/QF3ZVh9wQylREgRiFZaGENd9Bfw+5VXtT
3m8a5rtkFGFAg7opoDT6sJS6ArPxGOC9m7MSIyiHfoUCv2DAyv/EroyuiO1g/ZnB
u+rFN3D1vmMy/0z/x+OrD3youBZeg/XEU7x6fIqshD2WLy2UCOh4FUFRbmWyeC5l
n+95poYv6C6+ilurOIrI4sxo50WUkDQ7GQ9z4gffkR/yQcdjS/5+6bbcEHthU/l4
X0qs62aDdzlYsbzNz3Zxqr9WEdZz7kumqZcpNTaiIbCod6FGvJHva89NEgGjxtgw
Swkif9LvW/TaH0xLgMevPRqQvk/dn7q+kUX7Xjff9ryy+WqoK6ZTy0q4ogbAKVm2
RX62f2iBtbzbtUJUOn+bElHozsKl39ll/RGpKWilFXZd6boqwiPz/1TZtbs6ox0v
A+LSRgxCFP1JCcJYkjeyzMS3xFGK8REm6ideZzJrYfx5EOVxXAlhzAbXVkj8Qc8i
bUrQkU7iCA/oPicOkSs3WxnAZXmh04cudfln+6nBFC4xOnkE1uisST4ZCUkREeNr
ZVwF0ZWO02UYgoMHwhjcFxv8tvRBABdjY1/ClQVHFbWVCWCjAAfkFp+5EghPTR20
j2gMDjvT//Z+EgwrMeuLv1AMdw7hMgVpLSkD5fbxkBDQ2IWX2dUmEi2y7OLQum4k
MerkdcLceF4greL3n4nHA5Fp214fGfqwghrGDwLVMRaklxtW3R3OM7w11PeFrPAR
pujAGc1gHKlzAnK49bPbEeMH29se9SsA9qCvFVpWAz2UGVBgrssR4NZzRk3QuYP/
igeCdG/HbemM63Hkxq0lyxhyjzZ0kh7sBFJIa6k7fjRRnynikAX4K3oGPmhH2QXp
BgbtrS7sFCZqYYhgEQg5bMN2JZzAg7wpgt0Vz/pUi4zxEPwSA/TEGXLXvMAEpxzf
JpawEh7GyaVrzBYSyC0QbjxEa0Lfz+2vQ8Gwk4SOYMcziVrLLMnfhbg4ET3J8KLH
Rm9PJ0UB8fvgwS1JcqBQ012D4U9G00rfi6L78IDoxFOtYITIXgyLJ/Xrzo74I7wz
JP2tvCmlg8pvwDy5aMnHS/PmDdJZPjdbD8f9KBOZcbemdFA/Hm9ZAZmsunC27Zy2
z91yXJm02lqU/w7jljE/zuBjjfQiLQKH/aFPTCM7agVweEmi843N3Ca4A6Dp9jci
+RiNvaAOv4I5BgdOkmJ8XOwFRHrbAZqZYmQRfLhVR+y4BZq/v12REErL1TsgJ9lu
8PP954O4OfyixhPg95tu3IRUznPY17JiK3iczSePfWmK/z3sryTF/OIH4yIG1fHN
N66It0xrqMvBcH97Lpr8Qsx980LRKO0I2QsRpfl9uT44yX4L3siHXtIO4natPyu9
glTk1QsyHwfoHE9SqZMggtMLSepcc9hSx5Qfypr8ZK4kPDW0YEqNrbz9jQY/uVHL
4FDY7pnK3OUeSZps1zKOAgrq3nTwBBZUcDAaIS32FObwCD7IQ5i3ieGUs2RDBKXU
3016ecPo3klEchgHW2yhEtD6Stl0eOn1c4hNrkEFNAP9MnmyHwZ1ARiRXG83tPIx
rO4/9yvJKRCPtBUmvIDAtTsO3oSm07h/RwscRnIexEMzUdL3TQSf+66LjJvzrYZi
sLRveFigncUCjrFM6RlPDh2ZWThaqqUjqv5QiQOTUISxFf6SXo9lSjX9us2qp7/G
II7qM1bd0mDsmKVnxVgpoNi8JhgS7k1K5r63yWmw5C4nlC0v5l+JXtL9ycKR/9PQ
h0BQzB7Dk+N54bTd4CXqD57OH2dcs3q5Yit221qGLWG5sy+l6EQQf+dmhOrfAUB9
DDBrP0bvtPp28aXNpqfWuhFE6OgK7vaCK2XbP0nmM0HAWalIHXIvFCXYLPg1LxNx
4QdeS3KyzNDuZTwXKHl/kZXkJ6XuVbnqIunffjao29pPVzUb7Wm61kPmRt2vptQ6
OtlrQJLcJtTnJG2iCB1tLC0vydNrd1VJ5D0YOpkG6o6zetAqwrIwmo5hd4v+Mike
i29i6BYiCRX/texLpxbe5yDQt0BEFUju0n6T4s0ESEzF0QpA1+oXD4JBu3J229F2
hMvru8byBZY0sttcN7ESpxbS7tQsOHJLIT+lcaGZ7RgqEOT1ExTa81lOOWOaWdt6
YqPtusMcjU5P0S1PI6l6RDFHXPD4k7oQjU4j0h4j12ljhlBfWmyZNVtC5bYhdV4T
b2LpKpryijaezpV0o/Rj40i90qBtWCsigOP/iD3htGaOzCp/91cPvlxgAqPuaf96
pKbGYEBX4RecSO+zSg+CvRWX0/n+5oMgkgwymkl17vrY29p512B6MVoV3xhWZFkE
3cQfLyyJA26775c7lABw9gONHB+5xZhbPHe7+f/53w9RiIFX6EmwGv0hcpK03N0x
g1eJS1OHgMge98nJNXeWKZ3rOLfwiPUYrOmsrfe8CFC9yyaUxOG7uKZGZaoJC2Zy
ckBI2uIAs60tLzsiGBb4bXemlA2J5RaGpIzVbzkC7l9xzTu9M8IwLaC2M7J1oNTX
MYJDCRgxngjue5JMTqUUVnKZ21K6SuPYRNzxMiYnbOyvnRQavA46csYIMjrwlZi7
b727zxu2TW4qWYeR30LWYstqs7ApbWRZ03fByxRABeojymf0yIklv9AYNLm12aOl
0EgV3CMZukkwFZtzPHX7823QEoLJyYoKkD99KlnMj0O+eCEeGUEglWDvSypMKfGA
HU0VWlH33zwohl45vb3sqzw89Fn+KXLF8/PArP0bsWQRFK3MJfRdHYkrAyZoMV0u
kttH0VHfd7ulOBq5GdTHe+jEd5R+leQatav+rVVJtQahSOK9dQ/ud+Drdw2AUJXm
BbVlg5ij3UAzT8xme18eNWERItrE9e3m43EaNZTWFsk2MTd4nujtYe2OxoI62ZmI
tkpShgpA36LgwJWX+00gt4kxIW/2YF2vXCZ+afXUp3AajCoiKjkHCSMIlAQ74Lqc
lY36m++qwqCEQ9onAsmYgQX6ojUHG3SxZZUcQN0Wc6qlPuz9Lfv2VyAixaS0vFYu
i9pIazgkr6TcehpHO4Y3v6LH9DzqS7lJnMIVJKzjPFz3mxtyxi/V3Z84DPr3A2wr
CbtqZdowUh9lf9YbUWj9sEdZKEtvsKDZwWSdJjzttkzLVuWFiEVKbRkURGMT0KZT
213MSF2SCIVZnA/Zl+nsQ0xeBsW7/i+ON9BDfCG2gGDy0FydnFAeBIuf8LWNTeIa
9Z4Ih8LEmiw0VU8zwfHMAZvuA2R8728L6hXyAY5Im5PVSaIZV9qBtrvKfwsRLdId
tB3tLDvAryNC6K8Tzpx56MakKT+3KbtZZRIkPPRSWU1GY//P9KD5WtV8/ltEiXDR
P5mdR8AL6q212Cft9XAQKgae8vZGTz7RkGvF+0PYKnRuiEL2XOS0p6KJcGj+e6zm
orvvAKXsnHQl22AjNUBCfOnQQSznbqVwSoRqWdaXX0QKocVy3tWU+XeM/g717lQ4
/WukGU958dZWw+3xEpHryluJw9Xu2zw3cgTrbSJIt8xoGuJqfjbq6vvx48MbxXXr
Qxd99j9sITsKVODJ5s0sRZrLP2khSXUWycY0oy42c9vkLvI+mOEF3yaJqE4tKwwg
Vmf5rs1ci4pdbNht9cEnT+gcdFtI+2fCmX0P83Ea9CmlSh5kOupqd4Oktm80eRlz
hSekAXo3ZishLJeBb4rYQ97YDDIu/vvF7VQ+NEbc4aeCZaZfKjgPJWzbZOHTaPpf
0paHgVGm/bd+VGz1EzA3qfl3eHx1RVO0yIP5ClPpRqjnUvzOtDdTPR8tTb0VVZrD
r01NUtu2Da1B3MqDoz7Xs6CkPfFTehm6elm0C1SMVwve7lPC9z8+WAOe+CTpTJDV
HoR2225//40scWkpeubFQdFbPosFvsqM+IEHcc6TJQigJ9tlUXsEbD9TS9CTqhYI
nwRYDPhk1jZGvWYuKerL10Q0CIptF3N/BqI8a8blfoN7gFnbKhSigQz0S/jNPpyo
ZR5kV2Og/qyTWikYaZJQ+B7kW97qleSoiyTEh6LHU4l7fHRq+cj70DHrtiwxwHRP
N7Al57ARhvungNJYNiR1oBIvNNl2n/8PPC0nSNIfafjjRjYqXKDQwt7KTm58Y4jX
QvLpZgRnAbY1fag15NLXzkloCo+jBCR99Q0UTJRNt7KRdA2QxXTPL3EtxhlGPsMn
jNr457qongRpSeoBdkXqEOvVqqFkwJ9TbNtdSzqK87Q6Z1VLR3e4Edyhb7Bh+8q8
di8FUPS9l3S9HO1rpnrQbjLSZLayqZN2jMzBSecfUrDPxpDoEJy9txQC3KFArLOq
7z5ds/FPN7Ap6OraUvngIiXVL0ff4h5+nAmBk1K/JmTIvxXxQ/wgjah6nW85V1R8
RekFW5WkR85NgAyUY3rHQ2f7RMHPwVfAFD+HBS8H9Pd7/rHH4x2TL19FuwqCSL91
zV9+5DfF51LBHnUm6uXBcqc9nlJNR2ICZuITvXHEh2JYveZJEsaAUc833s8TMQGe
leyR7DVR32YJsnS35+DiLPPfab8vlqOFQbu18NqepPszhT/akIv+uTLKs2Hw7QdE
xhv769dP5Acd4lBYpNx7F+OS+/NiksrV2z9etCYp0YIMXltLjM4xcKsPLsr5Mo7Y
RLlz39eaUAjHVwAtcYBID0YnJpMcXAcl+EZdiylFJJz15UsmCYndMQbAMdjktVnL
TS4WDqNKKWwy/y1+lsrHnrK7mW+fMkOT2HUOIFa3sho+fco22aheFYV9v8n2uAKJ
3bPHGaDNzKALkf2rV7T2X9YP82qWZcDaqYO3/FEjGhQktczHAJ2sxvdHxOD/Rzda
yBaDtFfty97V7+LV45UIiRwGi/2apgOwhuMUbp2RIideSx7r8I2/Ch7oDuz0tgA5
i0sBDUQbxL0KgIju2H7o8cdGXC+PkAe8SEyDFjoG9i17W4/C/kLVBuu+lX+kbmP/
FfskdcTXyLTRA5LjTQPlSkTTVoUAzOALJ+AjPnEIMAW9Dpgbf0nYhJdKYGWLTFpi
xDJdyJIh1booXFSx40SeR+NnEgBMqe2Ov1WgWh1QJwxacWzSBD3zjS1VWrj7WaOx
P99emDQUk2pn5wQ+pTOeyxhRDRDSHtzNhXO9QCGMhiNKFpQPyYGgDTbFEfZvsc7q
PO0PGq1US/TCxoWAufDO3BjswwheXSZ71T8A3L8JsGZKwZlnlk0WgwCiDGikFauD
IIgznrmpK+Rg4/eft1GyCJYlpQID6k2pTC/nm86tTkkqKGrnVxaTY2ITshAXcgGa
GbS3jaJIsuiI9Z0VZDBqP3HIfBJh49T/SHkYrNBz/zjUmygPUbEc1mUPXRjO8OeK
sya32ufsQMiyrQbIHF9YVtSh0JNriVKjuwT3k3HhJydJ6tm/nfqPCOhnuhiW32Wu
YKYC84axTOIQScOHql87PFu2Iuww5aBY9Rcg7Bodq2W88GENW0nBE93scWoS/tOY
J/Tmuuhoi2fDL+bv3Ebf13NESdJkX3MWjnc7APMLEyHL4XcMdJ+h/mcABMgJkMYU
2Xxr7g5o0uOYGf93kop/8JB3+wSoXZFD/lI7aXjBe8lE1YMTB+qm8ZmLPYK14CCz
D0VZEHzYDyjSFD5o0mrF3ocnAgtX5yrPpwtQknwRRp6mDumIhne99897PeE/NZyj
OVIQDkm7iBnkAj9cwPBCf/DLXmJOmJHEkOOG5ziBBC8wqxk3EGHakOXPndX5rdHy
1IOEtkz+xvJ+lL13U4ohlKPJeVHlfOKwKXtluunEnlZsjXdieeZKp6xYxGAJ3QHw
Zw4GW66a4URifEhAiR1h+bQ5QCW2E9a8LMOvEFrLHJrct2laL5ZWYo2ytEJCPKf+
RV2c9VpLSXokDNlSOvr5ofe1GhROHSFhjnUwJ1Oz0q6sA/YkU2pCMEDprqqJLlFl
KVRKA9Bu3dIwlu7xDLJD4sCJ5PC++SJLbyUQWQcSmQzcUlHrWciBGK1BSuif5CUx
qAvg7PjSpYwggegFcu8dmLMbuxyMHoJHMWOovPVms78=
`protect END_PROTECTED
