`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5nXbDRV7m/6sqnpZajuzJBhpB02iSBaloeirjGbXHSjEUzylqFwGIN5xSoXn5I7F
xPeDI4JMPHoAcIRboJum2W/NtXc4vDNEFQ5fDNPOjZ1tp+upp+jwxwxNYg69NwQf
IpNFbP5akwSKgbDJPnpWKbEiNPL+XX1tFatA8MrIWHC73fXTd1LwM58hETvaaLQv
jI0ZreUx8v8omyMkMe3ZzK5w9uFQcK4xmAlKkFCLPfw5f1QCEf+Is3N0IoKUv2bI
vo5uXaS2CcE8TA98PURihsrFkZU4XwGtdSrQGoR6DOgxa/YWyEH9L8U/ksdYl/Iy
sfRWIB36NxhQhsWfI/Rnwg4gMySt+geWv+Q+23FWRk6uumwH0As0AIPmhnWA1gNx
o1SCe/IfrjNTwaxMqtKhVK6vXWIe13YylNlnunNSJHifI8eGmu2r1jX/mU6rgqTB
qw1bANf9+iJEZSPywxLGcNZuF/VMk6ewWhnyzs6TM1KxJutUfhzuga/zvkNsWgBl
9A58go5aCETlZ9HtwRdm7hLQqJAL/PVCEiVaE71EreA0NVNJO/bLldBGmVbYsSs/
NVKnKIuiaYG/ElAVVzjB29a2ot96mvgZ2HX+4hSBhibvi8LGs3FfwA3oO/o7Sj3c
yxTpUMDbTxuIWQF9iID4HjfRXRQInirt/8wTgOrd/L0Px6Jkz7H4ZnRXetypXKuV
+iq+FiYYwOFTgau8p0oPWOIjilRt4XF3K7wBZGxwduLkLyxfp9685iVqRnIQV1s4
KuR5GA2nzq4ZF/kDTcWds8l4szssUSxv/lowtKLTg3PJBkFeQQV2Q7wQiUm8BmkE
lwMGoaDXmgRUuOl7xYXUkjaygcWEkshaBlNZCPrnR/BJRkOkDnMRorfMpG60f9qk
0eph7vJMpTMF7hupiWnu/2jPA/FEWoVTG21/kwXE9IdL+aoeEXp+LS4XF2tcdPhx
BNcYubM02jkvd2fyFoo+30EVzKT+GzS8/KRjQdghtEB0DnYMpP8w7QSINIoE4hTi
o/Au8o0YyotMZvp2BBeuQC9BVRCO0GhB5VC3pXZqo7n6ncp2i6yPo2x+qQVYlxpM
y9j/0dsn3xeOONv9+bhgG34OzHwwKQuVnGxaB0akvg+VLe0wiJ58mqKbD3v5ec64
dqrYC5sdjmI/5HMO8DDazJp2oiAy1c0t14x+PFtc/jQljLg1hfptKSRWKnhttxPI
an4GrnFV5HAq3woyLxIWZFwQ6zT8711ZUfmoSS7jAPuRPSK1pOv0IP3sOaH66hJk
k6iH15XhTRgV9ItqdOhIqwJrm7+L8sn3SylW/YX6zUrwdAO/tN3kms84U5hm6wKZ
UJi2SiyMYCUo5InRykuqbZHWAuvrQbhC/sO71E1DMcD6hPXD4neXl8eD0T3hiHuD
GGi3hEukTCxX39ROFkL8UEPLFI4W+daHhr/7lxQebggYoanDvx6iaqElg1AdQehY
QUqNnUGY8O66sRXrGSIkOOKehGLBc2uu6FLBtupuVBDVy+aebbPnDHSZxoHfqYFB
TNhJHCG9bV3EyMPej9sfRAU90S+jCWYW6/2CJthu0xrUhUW00trrPhBAIaA8g0vG
4G2PEVD0ireTZzcMjGW79/TJXWyXrQoaKu2XAb5tAjbhPkkRaGYjNPKexam+QU1s
Pyfd5uZuxD8SKaGhFLoWbHhHYyblPhawZ2fonJkKxo/bdTPL1FePvHT6EKuF8nLQ
Fc4HOWj+B4ihC2txCZUlo2Q25XAXCZxO/RnazmymTtjSfw7MocEWeteH3ZnXDemn
0/t3d1vFGv2DWgSzZpMGkjz7621L9DBVSXZRqSMZEDudiPHxSg8rLEb4xBndGEbH
FtAu9i1WDBnBrT2Y+4kIVP7T38RSOYfZD5Vr4NTPaXHS7AG5FpQSdWonBjbkSdVf
wNmlBMGZ/CgUMguKL6hPmbnryhTC5e30HqDClJ1QpLB9j43tipCYy3gnarUAKAGv
V+nK24yrhHqaYPN0gCIqHCAz/MKXBOAIcN8SXxFut0V7nkDea02QpuLUCFy4EPmI
8lNwZMv2khNFsWA2uT+tEgOzAmy13jmwSGHNDhUqn10JgOrmFbJsVi5plwMzL5RB
GIvDtaXkeT4+HFKeTu+BThiw16Ik4LDK8eoz3iccQZKD0lXW4jwVpT5R6t/g5Oa2
8okXGjKxsD5esk1fb7GPidRJjiaHUpl586/zdUdYmodTdqBp57h1TwDNA4v+ywfC
LJXDUAfOkmxuveIwcJzDCGauCvcdJRMrUwPkYJtmunWgv2Zmo07a5Xwr6Q4Zp29d
DvLiBvvS7pwAGxTr9eAMjWb0SA1TZwkKtwIQhMMXwdaLtBkjomoXkyIEUaz+rDsg
2KzM72lCpurQ8yq3hnDRzxedHEKpuqrAujGFxBq5SCadbeAnb+yvhec8ewtmjxqH
uMTIhFJWDRFbEBzBp5kS0J6QB5XWHfF2aKj49azgiZQxoQ/o3MQQRKbgQSLHtkoe
dSFnzmNGo74d8Df3/XK7ez5y/GlSN/2RL3erJh2okmeGCMSapP/p7m9/+Re9cI0b
W0JqYdU58GLh45FMswjCuYQWTcywHiJGKPeV/7vKYD7HVky7ilEJmnMhF1YN/B0i
M3PSuQ5EsP/93xR2Fgi7+uQwkhQiL0snOi3DnHZPELe/ASANIYQ+8KRVIrm23PnI
ciArqLCW1JMFSH/oFGFF7EMc5LB9tE1BJE88uA1dHLOVipreJw1lZnQhV8IUIg94
fP++7cXwEf7T09+re5KUra5jqOOktksWkRuE5Jss3wgxIaltGBL3xE/SLKb6yHfb
bXpgR/RX2oV4LtiUCTBCr//UVIuhuit1CKM06M3IX+CJ6xRXK7km5miS+qBAhT+y
eHR4MTStDsGP8xerHJJlvTv0DGYgM0Jm06lIHNrP4BxhxDl3tShi5ZfHpu7mm/4Q
xcy+TLjUnOkAeoY/NTXg4Dh8P3Rn1QnSEJr3FyYiWM5MaoWgwdO2nePurRnlYkHE
eaaLlszDPpgRjcx9P1LMbgemQT6GavbcUyPjbIpxTudsVToxF+7AzfuUJ/xHNzLE
c4xN8gwawtNFeV6YH3XSslapZvPnM0dFtjkrE78/4DwqH+a0XvHeEz0FGwCwoQTY
H8aDCD8SiFSYw0I7HTbMEb5xOXughAi9opJ0dNtnZBzTBffGTFowpE3BbSzO+uMP
V7FrXZBG1+N9BaJAkA4vHUuMjY4v1gDUCBqUYCToka1PwZIiMh0Ce97dF6/EyEAK
Dk5hJv1wBhHoM/wVlqDEIMxS/Y1FTseTHUx5gYy2PCVpr1K24DHeuzAwAW9a6lwj
OdBwQDAivPy17ltNj6iCICoGt9Q/kIG349Xsm4GZJF9hwHLn7Pme5f9PWJPdMQNf
1sPRve/rjCbU/AfbBixSLonOO7CIpjxJzLU6kG8e65LN9tEm85THc9LN4G3iN4dO
0UegbU3DX+WQN2IpIJH1nS51qjAykdfzyDgGAKdoKlwm/eAMfIHSBCjujReXsfPT
54SxDy+NVTmH8gP5u2/sqLoVBRsH+NaP+WhNs2HtjskgVDoIbd3dElyiVCXstiTz
t9G5MGAQpiEtLU6VElb3dzvJU3YP0snUiNpZZvbAz6NE/Isr6PBRssU7+DF1HpAD
Elv+A6U2LRwVdJ9FhlVQU7T81I321y6A1i0BTey2mQ2BExHr23Y9lxjQcw+Z15F5
EBRNETTYOUJrGGv4yAwDmoAVq7sMxG6ZTZyN+H4+fGAl02grZeT2NW1Sx9KG3i21
P9oqhTZw85CC206Gs41n5H7X9Svd3eAm3mCR/SPjWvC6QqGnriX6Bjsuhhcaetht
1VpqgyPj9g8wywozTR8IZDbTxP3qoYRnP8DZAVcTda9u5F7hoc9tT/5Hdvv5Ymm7
mtwpP+eILPU8tH/5bobJj1y/Rml7Sq77XhOWx12INSQw6WVV6RGF84TqZcfpplSb
oq6x1pywRZObCAmUqSWuigO+VndEOTccC9leupC+Y+Nng3ZuFRKjk+1pdaAonU4F
nAKmFYnodgSJbCi3n9WLvConkjIi3XNi0T+9zCZiJ6fCa8iI28jKW7AUnEKywCST
+ZVde/rD4f3NMb4raK7++lW3gYYd3nwLR5XO269Jv96ttOYLQistQYmiT4UL11mv
RTw2TsGj7ueKBF8MXIPwmyWfAexOJyhTjSbmbE78OALRdbNxFzGP9vAmwCtSWV9+
`protect END_PROTECTED
