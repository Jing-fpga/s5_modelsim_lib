`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u4deG5axXQvgxgA6PPuMvGUIIfSSdlsDN2y46qTBmIH/+kccJfigFSc9Q3n2mzks
eyhPDe9QE2tW6+Yk0f2CwzaYyegPILjONjvyPbvBco0m0Q7Bi/423Ap203cn+ALJ
QZrQ2eBxpzHyLoVLVj68IdbulAJuj0YWJDaPpF3Mjuov1FHOeB4xTYgOgFWsyD8Z
H9yTEvy4XQ/EAasZrMtSbP0zxKZlTFukFCcNqhmpoFxLdAdewXYQZnWjrhqjaZPf
wWFl+21ZlBKe73ZdiU7VoRX0sSpoSLQEmGjbXv01NnUebmglELt2hpggpO1Ezt2Y
BcX0nUGANACblqg8lBo5+/cmUzsAxN2m0mcDthIwgRc2PF2nOaA+ytQjx0un/Jz5
JXXj39i0U3Famix+SFtAX3QUghfoXpVLDj28XDMoRlxgcwnkr9WFIu8uft/TYXF7
rwxyZirQ0lOlQGvOZPwXT8C1YiT8MLF0iUxVRsnWZq1/+qdslNF0KuLYIkuQoFdV
ZIvXH4UL8A6NehG0xfEdDiVIRldSqC/QEcIwvH1XBQzIV8B2x/X5mDQR+p8ZH/KD
C8jeki3OoBwmBoO9vQDcdgosq4NjWW2Vfq3ZCLUGm1yL0SgfE5P4D0guC6qjSJ9N
xAs8wiu5OJ1QwGHKwQDF/SGTVpriCsuTyyCjKUyuwJ2Aiq7wEfKa1wq61FQ1ziZB
jnCfhW97eH26+ppwSbSL5uW6F4BgX5Z3yetlkKmsFOt00Meog5wiIS7XjYGJNb1B
trnO9NA5x48oqJ6qoSsxPmDlw6owuNTWuHRE8pb304yarYb/czP530pdJVqoBJ2P
ctcDfQwdRYF/3V+jT19R1bm4JFLHIeNebilSxoTiHqex0QkNtbqrm53M1V/kJAVN
Oz0Z414G6j414pvxD8knEE1U5VkMQNgHFz8phXXOhMoEsWhEZhqDIydXx+1cAfbu
8Y8hqSr0AMwKsoT3VmXYiOQOk64kvf0Qu/L8Gpe+Ascet0okvTD1jJhXEv9Jeh3W
aAvXelkStzj18cmyvHUrVn8GhxPCp10tXQlyeukKs3+Mr9ww+I5HgI38zPav5gxb
xM7+BsDCupkbtIr24FpIcvpWxOR5IJQKxxq7IK74PS55yN34dDPApVTYokcZAZxT
0R+WYzY/Ao4ILPsbM9JNOIHR9P6J/GfdJyXKJBlXC6IxBZPSXN59ycLtgELguCXl
FWda+N6yLuf7IZ/Vq510V1gId3oJAAWHr8X5Ty761MbvQQvytjQzyRtFp6D1p8jg
JTAf3yCeS5udmKXUEkkHGydzZu0V8/kd/mhOAmmkSaZHOuJnIYo/bXp4p1wC3yPs
GKrN717bE6XXk8D32rWLHDA0uQPD9+5xCVCpP6Q0b2SJ2mygS8nq9NtLwkmjX5Nk
z3L/6HlxHqi69ZUuht00i2+O0IkQR0tUGd/j5xbkl9bzTrx/cGXFBmIRj4XFcCv3
2gjACHGIi9XrXG42k9FkfBgI5sLk1euHSS8pI29BJDUZwKV7KSXM07WO7B+5JNzQ
IGbW+2zMmp4F8PrrPkKvu+j53N4ker5E7Q8SjHKj4NquYKpWa44cAKukteTxjMSB
8+3nOSMhPsvmpJW231XmBEN6KZdrpdcs2WIUIFHnY4BLSOs9cMl83OxSnhw157EA
aVlRi8NF9em7sbAU/aiYqSp7prCSgocG7BSeYj/urLHOr9/Kz+T74vo5E0+s18ih
86bFcQdCcwwcI0XXHYe6H18LmiBQwQsj8PSVReVsH1N0gUjtUdK7YrRy1FX5AW4w
98gJmZiMKOxwSAnfjz8SR+fs4+rNtOoeHSZFy48LVsHuzyNy+3n+6EOGjw6+SFNk
uWwCX24X6QLTOVRjJR4Uv/Lg4sSzhEnwT6EVzye2HsovNTcsx75MBkzhXnl+TjBg
unzr24aZUlFcJE96ARpi8C7kRrt1DGu8MY/CuqA/6FDe/13fQ4JfL3K9WYo94W+3
Fk1YRHO7b+15cuyZvfaUACEz5pxssADXR0taQvDM97ygSWno/GIcSEGmNkf0Is+e
mEQekHz0Vmok2c34lN2DqkrPGIl0U9lsssemwqn98L2XbX7avfLXT/r5/I+zIV6L
JMPSzzqB26D8cH2KlxprLsz8HOaIWBJg8ILbp6THnnqOdwLTc7AQrWPj3yNUdeIf
jfkl66nFWvarn7xOfUyhYfWxV7z7Af0JwbiGqVP7RJ0jqidirvv/bhWf/t0bwQqk
PqHH/ev5Ixkxulc/+EJ5Uagg6mrQlikKoL5jkz5lFoLzibCSweRFF4BFlKZFon5+
c25Lf+l3DOSrRSbLeaimaPD6VDHz/15qnICW4UXj4fCccObSZm1KNaL6ngSdqblf
ZGYIsaHFX/+dnBaij/OWheq+HOQWuFj+d4znvG/nLbN6+GYkdEz7W6RPnA0+YR/9
1kCCGou40htFS+xhFZgMCV59qRAijEWRuMj7WDcF70eLJv8VwN4/4QR45JCA6FM0
w7KN8OPM71HVD6zKxsqxQA==
`protect END_PROTECTED
