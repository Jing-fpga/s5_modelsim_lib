`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EaRUYL62IHJxDqZdqFfhWO+GKyWRXkXwtMmMM9MQ22eAvMt0w4/nI07STbcCKLTb
wNARWvDi3hKSMMk5gH5ybB/zU99Mlm2ZSzHbNjDFLvd39ZQ4XBfhIAXgu1L2XAIB
YNuFlF7NyHP+nekfks8n57xVO+kGEjX/UnvZKJIia5E94tyx2HTHeATikdNhS/dU
9jVux7aD+vjtH0doOiODeSEfvsVtM6PtzHY9YzoaQ/4xkfg6YpjL75tnmW64/d9x
2QWCO71cNclulcIHbLg5Nn4VocJ1Nq8zjoTth/I7S726EIMH2aRdO3X1+ylle7AI
Hs3V/aZO8IiwPLMmCY7DLwM05z7rQZbQiZqAPzgBp/9V712AohV4IBooZpXEIIjS
YhFDJ/KO/n0hYVbvEdi+t5QvQ2TrEChncMvNzGEGksIenxs6M9VSmPPIYbSQigE3
fPgq9UnKnvsfysSiHnlfzTnEcT15FELsGzeiz7/R6k7cJnYewaUUdw89x5gQGL9T
V+TKLUXBUy/MxwqhBtUxyBXUoZExvuWVkkudK+YLwPupHa2v+popxxQp3rBR27a7
rh2jRUwEG6ns843ZWVYAArhX/WxqmUxrTI/TA/Fzsh6nrrfHAY+OpnDRPm45yfjS
DT5wj0GQjbBtME8+INyZ+gbO5gWI+GJjBJF42gnpOfacfeKs+PhzT8a/yjtUUBBF
h7mN57qfZ/7CKdksfOEtQnb+ogAKb3DXRxK833fRFRi9FbomaI63QVhlNELDk2KW
4Q213YBxAEAUYDmbQNnraizjQI04ufsgH9qvtFDQX3OsE5QeeV61Bb+90CzNxYct
PuP+bQsh9RGuF0qoFkHuKy+CntDP27sUZAR/xEegMWo3akQ5kAGNNSPzYCRfH7NG
XGPueUHJKHWKrhgh6FqYqndWhsV1OfkKDq1Ss6bJMA5zhpGz59AXXZV55RVPcEUi
CoK5V6ttz2jWE9ICNb/77oTGWVMXW1+fkVbEkTCXtqHQrS+GpC03fFEpsFsWPXWN
B7prNOVdLQEN0fNZdwmG98lkebFQlDiPJHTs//aM9LZ2aLYKwwpJ60zvJSIUKHbg
BfTqRYFy5X2hnepmD/UIg3N6Gu+wrMxA7BZZHNhZfy/7JCqjurjzEXXP58oYGLrW
Ua3EEkeYWC1qCxFmQ5/3CxLJsoG6U20/tiX0aznWWsvmLIZvB2Up3QnrbhmYcdbQ
uZo1OKPISOdQJS+lgi7ONPRomotOHOuB9MMfgDgVi1s3S73L8yYicuqLVJFGoM3b
LZGHC/UUmcI17foleY5c9Rg96uF5C/Q0GMFXq9EM3DGUKOqRasehyeMnoUxZ7zXd
UwGDJ0T9dpOd/w9RrxrOAX7mkGAJOd4nfv4+O+opDBmhiMYovHv529CWy2pH36fI
4R+69NlzYZ3G9VekPZfgr+dDUlSfvkIf2Kiu3PN+MHKHFG9JRHuQhy15vhYA7HRc
DSnKzr4YvBSxroRAj+GoyfInLvoTRwEzogMJsjPxQSIUx5yWbaA3ksM2AhAI1eiF
wf5WNCemY4/DY72HjvN7faqN568pRxnSvH6E5SsKc6u1PA6a1vMwaWj7WpMuHlLU
W7F/MMZDXtTePQ/XkJEFkFAOQWAtD9sv6LJSuIjEGlVCpDhy+UPfw7T1lnG5IWyU
zv6tINSgXV5mYgUN4jIGdQm3hw+4EsQBPu5TQnPVVQP363Fc+RNJRwWbSVdsr6QO
aPPzJO9eFHFny8cZ8C26ndkaT3OvR4ZkaEd27/bYFT2yqJ67xlI5fML+Y4NVi/V2
1ymUo5Sk+lT8aJV5UaiL/LnIASnjtQHlZqcyAZKvLUkIIyN6I0Ooe9kwt5gXj5TH
mSfxogINFV8YiTAImzLccmgu0/eK6u5gGa2hsD5UbmCPlHHEGR8/sTZ5gjGMJ+HG
3F4aBEkJt8w84Fzin3jlKoiit7RnGz427nALarbX09r3t/TPjUOji1GA+Mrk7Jws
L6pu9UbYuDgIcS6qKIyEkA26joOHjxxN8vatOVgObXKRNWxVbx0yikuLoCNLvjZ6
jgGmu9qCi7tsePiy1TLcM6JtTPV1ely39y3WIqtG6gFyvz1OmNitSESmyRQszonQ
WdmjnbEe0e6+MEzOPAqodyYbtVh3qHCk1nagQw5WaS9OTltkjLWwPChsnK+ns/6s
fcLjdVZygjdaVoEmn/+WtEGrF+aajs4EJGWyi+UTcgemvjr3Sx9hfKL6UoZfO1GU
QMN1zM8HjpTIIm0poCC7s4Ph5IHw5BQCMgBYkWkjd9feq0LRRcpOsc3KLC5G0Tj9
8Y3hFJtW4tSb+Eym0MsxQT30OUzI1Hobn+BFzlKS1Gk=
`protect END_PROTECTED
