`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QdYPEY0QeD30hdnZI2P+SEeV4jQ2ZRmlukvKoiORJsGXibUBo6hdnd/O3l+jfNHM
y8D0OhQVmU12ZrDqxC82w2YR8FpJGUHKuGL6A2wyTRhvoAwnvoNdqBktvlEZeuBh
WkWGACs43OwX8LCHZtjyop4gntcOc0Tc1+qHRduHDyo8//inbyzEdzamwY4UaZm4
MAtgUeyyvFVPlk0F9t4caNnISoHr9xlWCB8dDSfmLgMncHqzEL7dtqNV+GaJPIpF
u1gme3DG0s6qfd5C0KDvGj+mdv7PernuYk08sxJkLIwTuyB7NOU6tBGQBBBeG3da
TVbixqp7EBhoCi+oUB683MOwqrK8mfadgKjddd/I1Oc4vYLz96QxXw6wogwGizMF
/kGsPHGuvCN5vtIsh3lOn3BKjeWbHKLbMsPCOjvMuNfBNcoHNd1e8uaabcBIfrU5
+gXzUPKWsjPS0zOC+sxWTN+1RwNpZhO1CttCrJksapBIo0lgoXSAEHe6zQVPrOHi
sjXCwnc0ndr8s9KATFwesEpgyRdHuu60UjvgJTbezDyFUtEpKTNTAt3fEhjNsGfn
IsJSLnQcvvtve/pc5sHzLzdgXIOLnE7n4taG4c+ggy/K+W0BEU6J+H0jX3sgSatE
hlFFcpP0535+bAFVzRATsLHK6phTCp+4Sh53i6Da1fNOOpPhgSBFvG9xmsOp/HTq
PU+xkGc8JWZR+idufLZ9IMMmEXLhJ8ubZyG5MLekhY7PnG5hdPR2eGaKnMRJSj+o
09CN3vcjt/bBoJS/1Etd1/0ELYiwGAJQKVbLy0qZDhoCKcrhRGVgetV3di4ILDOT
GHgvErStKzDxx7GBOykHAXz+1/AROoId0BNYG1f8GZ6IlszMnVEswNUebs0cAPHs
aRQFG/kGd02YKRtEmgeDMcShMEOjqX/6Gjrr2dXTGhOO0Kg4FyTS/xnQ0y8gSKTh
PIX8PdMLuM1eVigalo9NdeF/2LoI/vTJFhjRfP1kWmQyjpaBXq3nX33GWNSG/VxC
1xuxTu+CnxEtJ/8tuuWrJZkf9fTsS8mA/e0cJWygh9bQpoHkMfOosp6VxIEJ7KP1
0OmtaOSOR9ExWDWSoqm8ImfxQklqYYcsOU/8BbDZQuc5+HFeH+Tsk2dG9x90sRks
02mX7PUtK1s7wtp227I/pNcU6rwu9VFXfMrA8/gazunu2k6Ftxp7VrotREPwT8e+
r8owwOwZfk+sgV5sxbAdeXdgmL4D961/Gf7y9/oB0io=
`protect END_PROTECTED
