`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i0P1Zb1RIN4Om1Q4lLMinnQaLRrFeizjzkO95iKUD4+WOwb2HaODbUj9NiQaYenQ
EqHmMgE+YwzUKMs+JzdWpnCJQuBwO02RkgSgiCnnvyTVz/Q7TPkN4URuV+cjQXwP
LCNvTL1qt2NkaNiHA5sU/rWqgYRREky+zrDxQEPQvgEM8mNK6vqLapG/m8Hl+0JG
UaNZb3vEB3v2CsDjxEnZNi5M76fmBNrVpHqtJLznR7MvfgFym0pd+Rqwwl8vNJIP
ydtL8TVnLoUn0Yl86hoxeT1okiCIrJaWjeyc+rHa81KWNhCbmXzUX50orIbmCVBT
v4PTRfdQl9RvAITlt34Xws99S8qhVyMTdmShDF0rW1mZoU8czlBejehedUE6kvWi
mFhmADhghQfZ1mvVF+uIurNGAeE7L23hZp9zkawy2T74dY2yrvF3330EDmC8aY23
nZJ7V0fFebHMts7tkivdnHnD1LjfIoFH5Pj4dDwDaAMk/BLJDqTQs2GapCoAios6
ubWvwv3vtiVpguw5a2EFohU02W0mHg+ooX6h1D+vW0bJsA1RxgmON4PZVUv4eEO0
vG3w4xZF2wvRtPD1PHj2F8ImoEw+te74IVHxqPMGlTfAutRPRrjSSgpYh0kAvaYo
fReXWvJKKQrZYFCckugKBYJl2mGWGnqhV7OA6wkMOFpr7asjCXVqDHA6ilwN8Lew
goI4OnSflwX0Li8AKwfm3EE2BAdP4Tsl8qXZjRB8fkAmHXKOx674k2nVQEEGLL9C
91PD4uZPV4hKCNILe962kFAswVoFyRxc8Gxa+X4AdXzWPy/7x+KV1JPxF/6Hc5pV
rlvEKy/gLrLa/cGPP0hNKt4PqzMwmad+CppaCHE446XnW04Lo2JnUgyQoiA9wl6X
lnugs9m9OO/7xxgBn5XxEqxm1YLPyf/nvPS0Mk4FIciJ6CvuF5Y6UmRhgRXAjvUu
a4q1jrqIX4fGvsHyRcqG/JsldIvCVJws3aYOJBXavmk22XLfVG9D8XudsASfhAtJ
qw2/vKOTAuhIejYiA0pxJFya9WGiBdhgi9e/bZr7gKby5DUhCxi36coOoYAarrod
5UmlBdLD80YqYGB7V6IJb8bv21C+wk6pD/HmFlY89AbD3uOIY81E4A8W3nsOPn2o
7r6IUJvNxCIRoiHErUZpQPup6ljRqEFbpe7hd4IldxpE2m5GKwYbjgIYPwwUMO5k
HpnKx9Qjfpcv0T3zEnhGTRx0AqjFs/CWWVE2WOlbc1cJ1zYNwJrQwquoIH3QJD40
/LZJYBEDA29zMRSdEOTWIQZBticQPQkiQRPWqFoQVR67FYfbd8+N7yTjpe4g+Thh
j2XxPQlR8Sn93iPYB3FDJ9zR36KPc6cg2k3gUT3dKaFh7bq0RrGucndkP4WCwNZ7
RPTir/Lq6mLgKOTkYHI98luEuM0GPk+uOQ6XWdQ1EX/WydiBIgjOYrKpwYrAmS8L
1Yhk9xdOP3mwXcgij2pSFKOeIEHXfu7w2VVihtPyUbPuB9pXsA4pV14N9Spzr0IO
QBx/zpwahG7HXDB5aqNHVxg4QOA1R3NB57z4CiRZPuGzQjyDAulA5iGPID4fpSLt
BXyvGfgg+PeETAHDDzHvDEWMKglF7mA4UeHJe1nRD0hiGpUFJVEM9r+aYz0Eyu8W
1c+/R/smeuauVVi0aDoLUW3r7J9keG8zjQViF8JoCymYmB1EYicVRRfFEb4K63qr
dXpUBWlqYyET1b63r/M1qoLVrY+ezZ6n53yhg4lvKsA1KVtZTS6vv1zO5XAFGZ/A
PoHnKzn4VGXOtL3Se4f4aiHc2wySTvlvd8AENx+yPANs4DcDaKmcwOC7legOY7sQ
GJWhxLkmPsoFwIUYgrTuRePo1M3PoqUrWrwl1/RMeDqSfevweXd4R8jinYOFeBMH
5IXsB3kcDki/eQzUqtDR+priON6pBVJ/ji+v3iJPzO32+OEzAYlxtK+9GU8YnNsf
wHhi7KCUlJdJfInEjRCCB/JjDp3P6hyw/GFRY79ESe0m0rW5J60HEuJkF2+Ytu+2
FjZg+t4Ctf4IQh3gcetFOXX4lQCGr6HERjPtX/OiAkSmOspmp3GVWIwZkn3UlmQb
XRNseuwxSs5mPGHaHMz/sKHc+l0A2CZ3YDZ6Me1Juh/KUhFj9Sz0QIIeceWpKt8P
9avlWUQqkT08xS/yvnIqtlufKThvhmOp+COlmjCYwD0mgTySYcBW4q5a+0G620ln
uk1JId/MhZQAPrGqewMdIbvCw8OxxptxQnxMRbMHP8H5n+8XnBWF1hiVgbhg33Sv
D410RcQhFUZNtltAm6ntxaHVpC3CGuxOxc+8kGOiP3Q3DWuTZpqt/2fftjPuagQm
2WeRgY570mpuMw0BcLHCQhDA/uucu11166Zhq8ZtNvDqTO7z/hDI6zh7S3xnERS7
e2srrurLKt+cbIDSosvoySpcuIR8l50BtQDllXO0GrvhuHYodfJ1lIrY4/dU87c/
n0CC1PWGZbWZnWjEA4vF0yLfXlouOW10SsE4Ldncvcljqhdd+a2IL9oPhc/fWqe+
kscGfu9IRQu0yagBUdMBB6qvEWEUldAaAEryp1C+HcRl9MGonrX3oIIRLgISxZvM
pVH7pxpppS9k6T4+2tWQYaPy1b3ACY2vW9OJh/LzRkeIX6wRXKX7fTVHtLWSqOJB
adXobq/Lpf6w2zAq+fbRyl6Yt1rT4V7RxI0SNjqH/gG51IeeUjLdNJjSvRqiq+v6
tWTEaNJD18syMI7riKoU4jwj4nNuRQ/u/adKlbBBx7oUonIOyfTaWOVnLzP/UD8R
QSx/4+qQtuLlUjFZlS5HSM+o/pDXjv2BTAs8QWgt9gf3B3cOaFtNyihR7aMynq1x
sMMenffVhz9LToPE4aZdqb1EBHgpteyNfmP6+UpdGnCst7GFpeZniFZDryzLr/2H
o25wYoOUyNiT/2RHbZ56NpGsVXVtQj82v2foFWbtJr0V9toKBlExh1q0S/pAlhxA
LLsfomD6V74+Qtqfrn7MWqGAA2xk6Wbu9qncz1hfwWuVzzp28dAETsjZNRQoo7L0
9BiVhmFJ4NtbQKd2yISfgkVd1HHj6cDn//Es/V6qVeTniZWCpgxCL9TiiSHCZ+jk
XJfUXuxLqZ0tNqcYohiebiFv9xX7GFkQGSAHbs744TXhWVKC9vmQsSPCVfrCZR1k
S8gSgkZcwxpHEBDPMaHI7XtF7GlaoKuN/LErChw/srpu5UCUlq2Wi1aJJhqUi2Jg
274/fGXb2D42u4eTJdoqidhjl+EYD9J2YqF/2mhqoREzYgl6VG9IcgCy7f2VTKzM
Qjv52zLDpy3rwdA2MI7spyV0OECp1+xiHK1p9aYTfF0e/R6qa3gjECVNYmUF3o2g
r8Hy2OjAtUJaN5BNwXddlLI5R+VuEpWL33ufz4veqZfAK+mmV7TutLHRce+k9sKJ
tCC+rza2GTgantmMONAe1BCfhHXwyz65a34GNfMvNW9YjTcho1dIEfNo6lzJ3OMx
O8Uye34MVCIzU+OF8Vnt28ueLrgq6GGqHhaXwEqJXJXvA2+c3GMef19t6HytiSsg
iREur4ry3LTLhWpOs0IszcbwpqsbqVNtKj61sHVYRkZFcLD7bZR/WxwXACKXQerv
7iNY5cx5Cf4WeOMBQ0ORw94DiqJXVFAwmuys06qJE2u7jek/lHKEyH5bqK0tR6ug
V7pvjzFG+F4dUwDL/pUJ2TMPWM+BjjLcq2jbpKfvamrJCcOmb8lYEmosylj/jPAZ
4Fo0a0IKZ9MtyaZfi/bOhg6F7teQwTrhOp6fm8zRUh8G2qhzeBD0BQPFpX59vkYA
S6culK/nRwV0RG/5mjBxdJ6xhF+COEO7asT3NUEbTX82E8uBv7gr4AXru7hXOwO1
VFyUGLEleFmFp+xGUHdKMRBuk4dHsMB4t2UySUcJQ4XExQjwv7FyIKu1hbCd7q2s
tNm4iHfyI+19R2NCW8i7vmVgv6OKQHTtyu+Ul08HxFGPF0xQcENoczhoCAhAsQpO
UmkX0hyQDeRRcc/1tjTRXq4X3lAHqfAIS3YP1InVvZEuOm+Cca/qLFwXvyrZtDUs
6jX7auSsUrngR4nALNtRlF8WcQuJSWGZUphnLHuaC7qPvXQshDG0yGJXl9qCo9kF
2rZJIkHTBSntczimglO00vhS9f6jBu+KMFYXXMV40vdvCUCXlajAoZe/dlcem34q
l60C2304Pu0XFsKXm0ImmB7uXqfuYuldvv01LS+9UeyCg7QEU8XwnoPpGVyPpmvT
j+QRp3Nslt2lNIl40ZJDCMddTO5OxKdOYM0msMoyewo/9MZET2xSIJ1+VYXoIHp6
CteGAQqDZWJ96VmiliTnKk6SC3R6EceAdU3p2F8tf+cwS3+GkeKDDWz82nSPF8bl
EJNfhRP02AuwoiSHbeLzFW4+s4e38UvtYlyolArHiaZ0XytKgpfuyx/SkXJU/LMm
QND6WksrZgBmcPzitcE+/3f/WNKJyWiEHxcz65m+sjDtz1M7m+EU7dQhKwhg9BCH
E1QVMdm0gkpinMY6yrzhEJntbiDOw4EU9urwhctenDgdBR+2keebDwJaERnylxpb
nLoQBo0Fg3kusJ53AC1oW0jk53yOZkGZ83sPH/RctK8LSUMQNuRJlbnNRDDGQbZS
9kQlFS/hpAIdy4pVxjwxRDbMcazUbYKq/NjohhCqRIVd0cfMEi2x5nofxIMix0zD
vSzCDgnBpt81BuxkGAdVDNqunp1eTwjyDJJCqCeIY3rtL9iZh2Tj280cTO2X/xKG
/aFqAogg8FNiuvduRHpPQhTJcHBMGE0Sk1niMnXS6hXGBpYSntLuAaFJ68iX1si9
DyJBW4bZEAT+8m2wmFKIKp4/bIvE0eEX3ZD1+pXoeOWMNgQBZT11Re7OGiH69Jmm
GCPRo/tQSGMp1Z/Ixl/ou08CkUSpwH4IveFt4kM5cQ9MqiEeVMcn3BZ2+0ak5PKd
rM1Lu2IPP/g18Me29lbL00u7W/PaEdqyIsJV160yDPfg60beZogjox7BDMGNqaJa
jaVgRbjPKnHiyoHA8yg1laWGC5gd4H7+Xd8JQMooqfQ979bvM6EMVBCGChp5JSTZ
xnC2OqybCHhk8JL0cRSVsKciTcEUrpafPczOxhZi6ErArRd9lHYwrCDXek3pwfEZ
uIwyXlo64aQC7L6ylzEiWqSRetKCz+ghA6rPlUei76aDl2SxSSYEDJFUuLXGdHuY
H4HV/1Jrd6ax+yPSLQUpTKjrGFZ8OqovmJiGfv98FPwO/qoMVUYZYALI0xD8fYKb
bB0OpIg8dF6Lm6V+fLDAB2PMXqU81iVtCeh9aywdg1i2hV+rnS7lhZX128meEtFX
5rv26M/YwhbHJNbPAKFDMQGKR0eeCJxefxxceZQiUOlaZUJ7gQqpGdyTsI9R3D4V
U0YTH+MNv2hppF5lDt9fEZ3fPxuqU6xYmF4UpsFb5zEykOZM+QigoySmS2rbFvRm
csTvl4CCNl9noHkk0tmWTvZD3deY0kgJVNdcHcDvdxK34tRI6l2R53A+kigArHMb
m2D76Egcq1hNU3wrhS/JGgr+dUm3bVDhs4pmqizZWhRJfy0u3DCgwY3on8Iiy0yf
S6GEhmZFDd0bSW28gYdHQahDN+NoZV0VPzdzv4nK4RgXWdRVP8PAbwWJR7S+vKnF
vl7R3vamad2gUXxr8Ll+VV6t8OYM4Xn5Y1hDa3hXPzTTsRJp1Mxg2T6T3YHos5MV
7pGXXLiBlAdGNeTI8YHKEzPlmikwmuPHhKpdsLVXG1oZrrbWDICjUmk4TrE9HlNf
wHwe3sjzzxu8gP/5KC4WK9v0rbp6Lfghaus5diLQ4/XE19Co1mLzZKrK6+Leghv7
VfRSgDlgB2NoFKHClo2RJArn1S7flgRwhP5u7MH1Zsc8ZMMTD7LwnUb0kT2iYglP
`protect END_PROTECTED
