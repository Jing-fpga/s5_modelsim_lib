`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qRA/FyuCzXKjqn70vFGwO9krTv7M49kI/PQo2ohJ1xJ+xYsbvZJsrWL6GqqlxMrN
33VsH9irzNaEcoY2tV8HFa18JoDjdlElpIkAP7OsuIkTDHSNyJG3Ss5AugeyfbhJ
dNFz0cYXJO8dyLDAcd+oxpXOTGXWEXcFrc33OUxlCTamNecBKFtcFVKdGopipz3i
vNG4eHxHeV5jsJPg3pm+0a5xf1uN/8rKUVzDSpPaRk/GvzCFFoaK++yCPhWIbT7c
nhaBSGwT9VnNbAmgM87E+qwS09ol2v1zE4AaEvNgLHenwOLNuOcef1NxgGr+8XTm
kUjY4m0zw4THNw8s57JXvLh74Ml9J7Jdl8RGf1NhQruVnFmr6a2LGSrSHLrQ0tOD
RTCUHN1Sgoss6227qy6XjJ6UteBfJrlUcxMWVhg1EFHJwjR56fU2KWWboGmgNBBN
3lBlX1Us16tTcO7NL/Lww9Ki+YUbODebHRI2yMH/id/zJtfsgNxnaK3k4q/4dpAz
zFzuHkbVsUQ0FFBbYD6eec/yBJ4ggaNrzSyWGPLfdYTOxALsScL83viH6K0QfGCW
0ZbctlJ++tWoTZoHAUQrsq37ExA2BgcW9Lhlq5TJN3FH2aPzosMYbcCtgJfHR98P
PakVVrtZTKm+Hp6U60Nnx8tFLE83vZpQgNx4Vr+rsjRkzW2UrXe3ZG29aiuIuYVM
UbZ9fek6dqtINMhZZsmgINuS0t5P0yo0jxA5DIrqtwm8T0FmCdYpXv5upmsSeEmY
mvAMeALqxIiov3NituqRGLI83campxcW+ZtgGAsJpKNVc2ixDLQVRozGOm9PCgyQ
zmTEvXGEqk2QDabJeg4JzX5kwmU32h1uhIoBacsZkEc=
`protect END_PROTECTED
