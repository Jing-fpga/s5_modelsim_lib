`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r8KoAq4qnVcqPrF2zt8e7BPxVZxb9mzOizG2/PH4+jru9Crgg0lwNTY9VdEfvxuJ
Rs8vuAGcV6cABY+sqvUAgc4XmCfPY8dhJ5nNrNQ3YDwlwtQQ4XbwqmR0VL4XqMHa
W7aPHC2PH8XN4Ve/LivZ2NNnZn/wl5KBecPWsMfEUyQ9olKzbPGHgyRj+RPhmbyN
hAg5jXhqrNuniEj4MIRSw7qOL/sbYV2FOhgxZk6rMuDIYykvcHQ7v4AgOd7grtgS
xIUvCS4oBn1lSy6M4DZgI2xYEKU20YDPpMKdPVUmZ29haAY21jLNDhc5zpwKkXQL
BKnV1GpWA6mKkVuRKczhBkUqz6bZfFiktLwjH10YrQmiKmrpAd+brj1QheEP9wCa
UKaWllhkvhKx4iOSWJZoRgbu/yxFdFbd3lWi4s8zW2yXr212FoK54S8hqJPIuFG4
Ae3Qv3lrlBbU3WdKJTWiEce6E2RYSaY1KhIFv2UFFdsN9vX8OW6aME+aLkgiLhoi
RpICyoILGmMUIMBalJrYkfx5vKqNQGHnoDgMv9pyFrQluiRsdKbI5piZsx5hyeOg
g/Es6KVGyk+lp6SqRSm5AiemXwkmdZRVSNoetlL6SuLJbOypJEA4WZ5Y3+51nQNH
S613Jt0xfs64ZJ4jPmb/wk6BQ2V8/T7VTlc/1Bio19w=
`protect END_PROTECTED
