`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oMpIMIQ86qtm/Eok8wRdwnZSozrdGQ7IiTSjZZ2y16Os1Kr+feoVU5BgBGSxqtHT
ULSTEyi7R9aGSbRWhZC+5whkfvZm32WNgogf/7oUT0QwHHobFahMlRZLZsMpUXE3
0xx1if7TT65a2K0HqGb01MYgmiEJJorBz3yXhN7+SwEnYhBbLUZqgsk6WPIAGQe2
ukMvT9vhHP653zhyDi4F58CsRqGJ8sJRD9aqN3Rhnk7tq3dYtrqXoPNuYxjiKbpf
QGeyDWGaoUd+yaxGjK6/fyypTtBkf1fuheuTU2ODHSgcVT6MCm4ReKIRM4I/Oaql
rZTf58SpKWGfh8sW7BF5jseSYoYB/4FlC/lS4tsYLA+UAqILKR8dFs8QA3DZkLup
d8O19EURg8mR0YAx6Eb0Y+49KQZGFS6512gGiMasGJbdeawfNf5TlOHTHzZN2hcw
SYpdbVn6vkWiDp3C18yLFtJ5SW4HvhowhIIJpKJXg7HjAS03VYZ9zaO/4NRZe/DK
Ne6Ea1oZ8jZTIyIA6VrDNw==
`protect END_PROTECTED
