`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8j2vk40/ghydnF3qoqaaeEcgFib/5x0/O6oUyqYr86m5MsZCMp6fNRMhhmBNTrBj
7UAAEUgjZhA4bVBWnFFeyYPEse5XBRZgouDzaMTnWHtJ00z+0PrOYv5/cbnv6Gon
XUIBNUjcGHixQOi1zP9gu5daKbXpuMNNJqF6h1O3R+kMMUUJv8t+/k2eg0HPmAyg
SUJjpwybNLWp+YS8zXOJ2LiC5jcd0x5sMSaIDvbXAyZl3sJx6wZv9b6ewOv2MGqt
6i+WWSoY3nwjwm7CM53CQJyba0kKDsbafydeE1dRsCIVR4NFKhNebsMTRz++4t+g
GGSa0szoH4yCIPamRL5DUkn5IESf2cd5nvqUaHxjF+GnnQP6c66GuK9brHXBNmoB
rdniQvLofuhItmapYRm2+lgZAkOB3RznlRrUR9O1t0T8zPDKgxb8lt2dqW38lkIp
Tz74WuKNVM5HpRRJsdrf+6GTE26pCGvT2GRUBiY8czphEcbXIzTpZFlFIs/NGnPx
/K8ANE9jkgYdaBReG2JgxsNGfrhZ+bEbq78a/ZWTwruCe84KvK0a6THORcRnUXwO
Epl6PrwyMWoDSbR3IsotiMxl9EmThycUA8E4evORSqnGL1+6PeqkT9JZz5hk0xXs
wzBo67yJdea6l8q3fqEjT/ElKQsM7sD6n+LAHY4WsRMHorHWHMGSlChCRRcMXaSX
jizsA8KQCZe0Us7Rk7Pq5VpLdo2D+zmb8EAwxbpk2A8IiVwoZAyKrwRu8iQ2L5j1
BUpg29zeqUzTzTerchkX0k7N0kuoTx1+EU9s1d7ChlkSOyBHBbqtLuRGe8lxDlgB
7NJZDMXWqyBnXMPzaCx145m9aMyu181ljOzoodQkbviwuq9RHRxm6CaqjF/SaOTm
KREYvFYTwfhWvIDOimY8yy61zzEV4OW8VVTn/Cu0o4oFRQtYZlwTnjIZF17FWKsV
7tulI7kujeYHGuseSGvIATDBKXUoacZ+vsK2guqVZnW1oi7F3p4oexOxCu0oElpd
uvXXfBlHBCSExzEmU3V8wo1vIiNzLYYvBMQxLXYBA0SrD+5fqw2Zox/ikimLBrbW
bKQoV3Q1m41PN23MtjmAZ5dzuJCK14Mcv4PKJYHseRowalAptzuyyg2A8oTXz5YI
lgQrQjQiyE8g3LycALVm6CkAO/uHEr7Snfoj1R9v2pCho1C22Vwo5XF0vduxTrAm
Pf2WznwV1gq2PD79qdKb5uIbolh4ARjuuvGi6FEUP/iPaMb3+zDxs8UKzccHiSaa
fRZJCfDp/GJw3/wvaY4y5jy+e4RoPaQhYl2p+ngboriSZ49VV6VDV5l04s2CkTPh
h1DQ9tlAd7oRaJNn9FpCDLy6lFRU5PP3fZhU5H1L2MoEjJS1gPs1x3He9wJWEh+6
WEA0fh5qAdRVqScc8hE+daBf81WLThIDj3PrNmGivNQmu3aZo92ZM2oewHwR+XkK
WZdA1uEgBmJpVDLea+TqSpcdfyImYPVdU+VZyDbXjnOpiCp7pGTYcxzE8Jn2VGb5
/lPgKgOFcNVdpX6p/uKNyS2Ena5Kw7LHj3fuJb7P/WvxUhUj44wMcToywCiOLpbY
sBnNwcPBotqh6/QQTFoPMfEXS+LfSaOIzu/6voHQqpCLPadQPqFBgyTzZBdpkMBo
id+dXC5ApBig/UaeB9XRerMIyrC2jZnI8wwznbU09dqa87H5e/AHDcUZ94C/3sb6
5maoHD+pOcdJjIZBcyafwVdM8cuvuZ1K7js+H6EUQ5CTf5eYcqG5SYU0ib4qs3Uv
+xnaW71aO1M0ruMVSWm5v94sl0aOXRqSeKXFWPeMezv8rPTGM8mjNhyoMfoZ7lP1
xEOOuv0Pne7nPxu1bQ20bidap6RV9786ekmfEGkAZGkGw3gb6r7i8ficMqsXwAk/
Q5+Vc1QyOuO5kDa6qc0ysJKE0dpnIUjVIu/kdACgGEGngpASZG4wEMkc/DDoKQkZ
ZKB/qHT7L5waV8qsGRXyQrEtD8CDwhv2cZOeB1okAWiNKPwJkH8QTwryfSKiZTQH
zzoj3iJIM8ot6sM+zrEBZH4ify60HOaU0LzZCx4FG2rznsJXPCDyBw3NPmdvNq9C
R6wiGfneb2paIbb2IwBnzMe+wGb3jTZNrFqqBvfejkr/RLOE0Fce9CL9ys3XJ67Z
QEck3SpuOY2+glJ1B4LLZSoyciK8EcE5nhkt5ytHP1+OZNdUtMH98Y7O3xbCJIvq
62Ws46fyuvjwvjHFzug1/+3J1bvJ9o+m3jVYJnAMywqIBx0PQiZOLZPqdku3slYX
eNsqSvv0TmqGXGxox8oM6TTexUDtwCTEPv6edx1Mt5QqP5932ptJs8BAkFQA58Nm
n3FHMmf4oDqxR2bBgGAgAUVxRk+cdpD3LY3VRjmIzMHBLnpOJy1VsAi8MS8HTGAu
NKzx7hcwPEqC2lnP7Q5YjkGbslUFyyGJqW6MX2lC80LleH+X0EMuMLngcVsvbEJ8
gy1OCf1ijAEvYv6iKrSgRW4f4mqRJoKytKjt4VMZ7e9mz1Rs+7sLwcLoLpbINnqC
3bHc8XB64eD4N6G1nU6hcH7iqgbD2vGYkVcCUddIsl7KhRuNWlTq/drpEnVhz4kt
8+ION3AzezRDM0gIM0ZrzIHegpy7lSvWJ8idfFIEjEeNLTODOZq+KCI1adsMQfFn
+ZiZZ6LOXVqYqZ7IH/I4yoa/GMB/8Dpy7KZ+jGqZo1P4BVtuU9CBSdB2TtUHmV6a
hDeQHb+90eBOLh2ku/NU0E1xqtP5+FQ7Q5pus9L+D9HL3ZCyCKtmi10Gv2AP2XEp
4Ew++mmgummNTmOGMKSWT/Y+OV1O3Urq7wosEJEjKahtDSelEKIdfngVtG/z+gfU
OKB/nRn6GIYxVquU18KCGI3UblnH2ShYaXiXhjpePyTRVGx5KnpSLggV+jkzKIlt
KOUaT6qvkpeyga8k3FwQQ8E9dPZV1csnXCMcerxeDJIOphM1uethLCRJhc6JU+tV
u0EbSB9SnAj1EiKYiyHzTNsQO545lnmJ3dNSPEPs0iU/GF12eoYR5qBHkWvhVBvl
zncRo0Rdwo686SKtgSGIMfXYVlYEYRYoZ+jQob51ok8nxpGNfaJ9oYGmg8VMTO3J
x2y/J32JtlLyWjFic5pWlpHBAofKTIRwTcPKm1n2G59ZBqAnUcFX0vF128CeQ3zH
jPp9+V0r8QAP8iCRF+zU8Fo2N72g1hL/jr0XXw5Mu9y9yTKgOAbzwMIMJoq8jyF8
NDF2R38i7q5tIv01qRsFtBMGcd9j+GS7GzyvSeRAHs+ezf0dC1IEhHfYOjavKvb1
Lh7FRB2EpvPjRvl0/23huCMwZHd5quNpTS7eHoNkJLzc8zPd9ofqqt7H2QnXeZtZ
wwSSSgRWzNEEcwLYnU915ct053x0y4VHnoaeCCWK9Yt92SKELaHI8aVyQLwaNS52
j936kJjh7f6iG7L2kQyqdmTbKe7InbnzcQJfTkQRv9wmFe4LQKwcaoqMDihMQgxu
4vU6GsgewxbJoL1FjKl10RDUnKes3xZRh7cV5WzxQabbbCqEwOi2gql0Uz6rVMny
LuGNd5cOhcp3Mxq0BvTJ6Eqa+CWU2Jh6i2nJgxoSwkehAUe1w0RXRz/YxvAgMtKc
1SNIjND47yZVzKQGRdCth+IUBbRNvFalhnuWTDJ7fsncS9VuMFb5+bzwvfn3Nk8E
eQpOBAr/cLSq+6pWMbrGBOZqKMpYCleBg4dkuldlBJbeSDroXL7dzqCgnojw8o2L
onStAh4STOs8jhRfnazgUH2tKMyaHVmwW4UKysJEdFOU4UYlgjIvIN9iqTA0qcNi
avUKsUpzeTd4tqPTF937dqLSgoqxg3mpkUtmcTpna3Vm5QnNcI152zTVLNu2IEmM
LUf+6WgOPkv0waXbt2IVt4eMPh8sv1gpf+rt7uTGkSUIcQuiOhYvt6UMs3kS0CO2
iZKKlMK1lNfHJKPpCVs2PJzS9+mE6CW/1wHbp5B8YpapckoPqX2x4XlhK2T5LqWn
tI8zFt5gFig8JYQ/nOXaISP4S3YPQuLmB90xxnkaPB+T8j3mgEkCp4QtlYSrnMdZ
x9rowEPIYw3FvPQYn74uY2IzIIAe+xLGpbrio6K+/jDXK5Zl+E5HyPjzTXzxZzEP
vBhwZ7qJxdPeoolT5LDsTtAx8Oh3g/akUaMI8aIdveWn/IJsAjOUWa+HErDecFyS
ERkXhHf0KTx1s4Z7/YTGsBQlmGpcsoefXA3hPgK5QbsKKruYczkZYylIYOW7VFC3
V3X3dHXAYjBrMp4FlWxkqjdRV2vmRsPwms6fKp6FiK+6cnlWb52WzuQ3YW8c7ad+
iL2HZT259NFT8JAL7FhGUeMnhzpJmQPPl+SEkVJYEzj+QaMyxmyOsrYMTB+SLyTW
KBpnb8kTNdXizHn6SZLoQXG91Fdk+Rox+eyQadkVgIPjwg/3hGdYPXbaObaqu1kk
ZOauH+4tkjb8cpZVA90CwCsF3avqm8FY5dKCcgSiPWI3dtxUzQnbN+DFpeCR9XGz
rWiknMWk1gM78hEqrKn3Qv/QaWE85oKJEC9M5lFkRipXOJCRX3r5t0Uds96gqk9l
yt2dSbhqEpTcapPupy3QfpXYsBj0HFA/iO/wrxfObfeCLD6JjsMu9qcf3XtYlt65
Z9FV8mdAF6p4R3Sws7sX5nFpAqWrZwFKAR9Y/p7/OOgF7wecsmvL5XnQip9dtI8E
uSyJn2xx993yY3jDCfOsMIheOnE+ZmRnED4/UKpHBmoq//qkgR+lMgq6SluR2UN6
yjAYVGjkpmf5tNFO1OD7RJmiGRnqVyoVC0HTlLTsptI8yN9WtX+OZj8vYACrkVrV
RsefFaVziN0zL1fSaOWTbh97pm6OOUlKMDAwp95FiXePIHMHzH3ckVdstU2Ihhgd
0FlU5utYoi0VWK/9XMMhlUIpaDzu+PRFtjUj2yr5uMwPSliLzLgL3rJIB0mDJQbP
9mrdxdaw6YavQPtOQ3OLJqUyrLTmLP1VzHip5z8l7+/dpug4b5yQM2WDCVbFTY3W
kU77gPkNeJv7mkCWh+fF0elRNjHr72tdYY+mmN//4zGHjh90RZzLglTyLzQQy9ae
XkHI7/Oy7IXrD2TCNZ6ijOhtXWY333mHaJNb+CZXeASxkA6azRTf5ENQzwSNAZNh
Rk8TANzdByatbyClcSlrjyKmdr4KgZzMZHIkXptBE0BoFLRwAzZcn5teFZT/4js0
+J6RynUsFThgCivapopoIHPJuvOuZNcMEiscUn/idp5TJ/Y3oJ8OYbxtOSh2GeTH
/L+Db3upgKU8GU3PCwdE85M50Xg33OKBbHVR8r6cxZJQ28bAb9m+Twc838Nbdd0C
ulfWNUlMIF16wt8xp9oI2jPZ/u91ELM/J0gPx6PXsFqs94JPWWtulEOjeiHT/+65
GmEvovFRMREtiR036uoI+dCyRD/XgtH+6n0/1qQ0iC0sYGFVI3DkUObwWNkrTwAB
kYNPlqzc9jEucDHnLJDrGGlkciwvgUcBUdkN18MkODXYuq61k4xadXmq8pR0EZ2n
xxqYgbg7zCJqG5HTIM8XXEq9aUKz1kjctBzF75FlZnr+xoXLvxO++E8YXn35ZZ1j
TMdZG5iQs86goRi1MLie1MbuWaTJdP0ullSXN4fjraXYArnPEnAm7QtfsVaIleRR
SeuKPyLGfSexk1Sp9sgYzWAic/lF8fwfD/dzGOqgX49JWGEECSSm3/xK9fEWqNoc
QOklyn5aaY9btcc/WO9TVy27QtrsMNZ4AEuHo/EeakFSm//8C8nimzT6lFw8DTbb
82Eq4ZXt7qeo7JIDlcp2lLVeRQAYg5G8Py6IuZKFeXxAzoWV4PZOznfcH0Y8QFe0
JdRxXwTZ1ROLRGEm7CVEmxznPd7Ze64/04EeB0VRUN52EipialO7bwI6WfUW3G9l
o+HufYZ7p4YjDcbao2TjoHozX/CvVKO9y8ZzzwEkjfCkNZ7I430hz9LwEp5Se8ZN
/yysw3hAj/+SlIR1eafb6y6kOBKxEA+JrYnF9WGCwYjiun/CevoQXfNYNFmgKKrU
4S+ON2soYrPtcwANRhUsVcvpnnwDRZMIo85NPISvM7CIKNdNMOWMwDKsB0bLsybW
Fy9qGY6VQYN5JEFBC5tX0Zpf2UUzsDTfjgkvMljz1Gsq/87kqJr5xnUiUZmacc1c
opp0Rb0Jjf50CSe0cITDIsAP/cXVDoW7cJK9yk0loBy4Lts8o8yQ8JE+K4KNG8q4
QzYTClTyE3jy/cdrQP5+zkxX0xC/FFvu+TJpwamgikFafbrf4jKwYSJ7ABCKOw3R
rgHi/cVfdUrmREyuLBWFh5H0lKooJ0lt3hS063WmsKJGIBYFM0ukpSm7CZnNy8mo
SbdPRaf1sYmFfkRg3Yc3+w/pFYj7uKI0LUCLrDvY+2Fs0VvMe7bDadahxsYkAMaL
l1Z+OS9jyeJZ9p0DkKoEjgrGSSR6AJKwWRdORrRmzWwiE1WwSV4dJrVcbRTNZflq
XrVIM7lnAjfw3uCFc3DMHtNlC4Ejf0H1FRg5CWS/bIe7H4XVwBWWtvfEVjQKcrhP
PpWo1ivxCNOAX3doSk8L65lvxgnC+2qCd2wcNZR/vt3eRLC/JNkJzxKEZSe9fc/A
t/fuT6Srf1YTL3Aslp0Duy/Y19XoiAMW5mQz7Bd1rrQbxV75NKIX+vpunL7gFXbr
PljKvztyrOZZXAIAzTuF/itLwhAPE67t7hRR3j5OFJ11M/0RxfDu2EQIQiGS5tTS
Br5RGxe8hNziSBntY3jRW5u5QBO70q0l4VefoQAnnXczbLFkrkIa358xhWEHG3Hz
451m8zvvfcnkb1TQUEoH+tCaPumSHIOm77AUdwBeOK5JADAQmdG/TGkO5XSnuk7f
UR9dY3LY0FLaiwC5Spz31t5CViJ5zRoN90wTCRFQ6rNXEHy9PvH4TrB6nQciOFAW
DrNXhiem4IAW1emZW6AKQs8G/Plp+R1WQwdm+vWH1xIFuUBSkya/x1cve3QKCp/0
QRe2UsL/8TI9z4WfoFVAsxrF4jLapaLGT1lQ9UVnJUW+mVDzDsANhwVstL7qah1j
QtdGrIc5byLVzituXj8Wao1ciWj4g9JKHn61YY7SmF3YDBPRd5xTclAITmjyF4a/
Pgk9AvkTf1rV7rEOAgT0I+pjhRvBNt3YjRUYO+ro8kuiBSFxfJJxi4F0EZDDbHlZ
vHpkPQTqyAlI8KgnHr5tQpluYqW2SemRiFVJcqqpEBAUQsJfO+8u/a/V+kGCr+5s
+z5ZQqDe02VKa8Aj2lRLNGgos/dK+ozPEUt8IBOMU9kJzwT4rxeFYF6kG7b1ruif
XvT4cT2QUAugHY8ZEqM9V7iPpTOvIg5Uyia5ALqphQAfEh1jS/VbYEaeLnZxDNgZ
vwC4dE1q3HNIGyRlYxn4Y2sNWO15WPO+a1nnuMgoe3HxVRvT4rB2QUcGiPx7BTtl
pacJluUWpKsPaVvIplqaBHyyLNjBlUX6mOM1X7xAV85AoIE8a1UNyx1RN3ea67u1
gDaznXGCsQRPirRrbDp5L+RVvLYLgOICoIppETd8IL8BFuqXsv6QNAQwH7RWtR9r
TnnZ1ubwrAFzPdagBgHrJNbhBdqpL63Nd0CKbfHnuDEk7YOKVqFAcKQuo0v7GpjF
fP/aHFFfe8SWMKnxfUwVXnlyNFymeAYrH5+KaWy4Ve1x9PHFA2uTckOQ8HpooLo4
JNmwzBfQwXlfDC2teQdqJmKjtColv3J5/5Rj0e+drurhIL550/loEfXHoTTAYFSW
RUTsy/VWV7NTXXr5Dv/dd4yACVq6UCHMK5ez+kwSFydrD2Bf198dveoyMafTNh7X
70zu/IYSAn7+s1ZMkAZSIpj5YslxBpXTrvJLtvJcf6MwZEZiAwWUyp0+mOVIQ2J/
irOSAVPBHgJiEolt8PlQ2h7ACmQW580FiwmCh66mNAKYb5X9K/+vOXV0tlkpEZ6t
73LvMOyaFymLmrlVX+XcsKRAqry3pLNDNdiQOlvyqxcSbJBdc9WxngYiLwzKHT9x
+RWpf34Bj9frDIFpAc6H5kVmptidY0ub7NOXy9NKpRDW+QcX7F4UrB69IzCxuvCc
KBSNFjwbi7SCOG+6ipYnQG+VAF15vSz+AzFVzJhDS6zYFqS3IrxOdV3x9v8ddbx7
CYV5Ew4Wj5zqoBgDUGIFZ3agBBeSR0aN4c9b6P78UNxugcgUxabk2azRCSJX5JDW
HrXqT6BawlO4R3FQALLxYP6KGDZEdg/RAHNVb9P3haGtRCiX8OKSyCX/iE20DWDR
uc3dKHcNuj8yJLjn3WR7VRNbz+ZzqgEuhaQ6z16iCeAZ0d1n7NSKKZw2tSCvs9pb
F9QdAwvxe4ALkEZkiZtN3fK7HQz5AB5KD2UZKg535Bf099aIcUDRV6p4eg0ZgSQ2
o8mvnhNYfNcjiWD39TVmcpurHzWn0ORQAMGQOH1H3azHb4TQT8sqJp0y7ydqweJK
d9ev04LDD99KTVgFHV9xQ0/2tYYkjsQ8irQ3zoucp4gVdmPLqtBW2E8fpLWH2BeK
WxfnSs7eHhf9p1B6KEVyPJu5a8lFX213jv4FpykuZlOPaYqMhAbaNlnB8Fq6u9ET
b0xg7IJwFPtncz7laHBOvq19xEXeybyeZQHWxOrs3QfWnSGO/mz2/WkmCZASRzFP
fp+vaRH9JoQ2YW8rZn9A2hVTJPOxSoqKBJ0OEKBqCUBETXR3jD5NKgrvdjlUF1gl
Wbe64PwuK3oFgPGC7kTGleMq/E6n4fifl6Mn2t3DDfWxUb9B4CHKrUlNld1w4e7W
zGopyGHOU/zEKFnRigwXj7pceNWod5UsAWc50IQ0sKAmv7HHsuF8Qi3FElQpinhB
Tj93pIdNNRUqP9wBzvjsFIxrULJwV55RVHiLYX87FYTxJF2OpjE9jDPnTF55Z8AN
Bu2TjjFCB7cadKCg2yR7+DQOubwCblSU8GeyFlbEbxsIiDFR7q0oFOEIx0dPPGTO
pV1ff1HgxMLLGhKMvbz8xo2dlRvYYIEX2jUS5TDKeGn2Wdq8ZNtQSDGdKCOp5iht
bZSg1czkNAF5yEiq4k2C5oLweqNT1AQOfv0Z6wwqflKSCSaMAV8E6mJaaKAT07pe
uuLa7ovnouh9fO/9lDTlhVwGC8j036GYnzIdeLvSXpMFbUmePhrZS19Ytfd4Bzfo
xPqXJKme3Z3ZUAjKAbN+TgkODCTujXiDrdW4NJAwLSwCYKBZaaf3X62ZNT2MVEq5
4yh9ny6rqWkVQ5h0It4Hch97fUfOwwTMYMDbep7wY/SpDc1fhhzODDiEi8qemosq
aXm11/m05o85r6OIw8ukJwdDq/DG5Y1A7KZARwuYLRr/wK4zloXb51riFHyT3CTz
8ibejrbaxEz6c6FUvdFmjRUdF7oxZomxQWfsWWOdPWcv2QiqmSF2heIuZYoPFKKq
dSQjLrkAFVa+mzeqmvF6xYSRYb/Xcbg+EH8+/s6bSFmojJB0xOI67LsS1K1ZdSTk
eV/tpLQirXYJmusjzo4KmhtACf9RkyFfWsZEAPfYME9+zP6xlyKQrEteEH0Wte4T
tFJVbNmUvwM1f42m0FzwBuhXcMVgfkMCjFEOImDYTL7MuAqyk7JleB2npCV9aT0E
4d75vPDfyLvftWNMJxq/fS1bqYBZHBIoxg2/vPXxW9CUcQFTZD4cIVC+5L6ikgCJ
/IVRET7QRM/tEk8NCr3Jxn490G4Eam/irfiNBbhZpGUcmGYwAucZB6DRaz7WrgwJ
ClmNtbCeJN1KtshHUTBgzFbayax2jKXBVd/qH8RtBS48+Gm7bSk1gwSjMj0rJYob
nD6xULslMJcQ58wAZuUsz1wiKV578szqXgjhfgErDJkwz1eBgtGTui9mbRaTK498
ImX7O2GdLTV+c5yE4atzBJKQY03av/rlvyoYyXIQ5t69GhYfW2vw54yT4Yedoxyk
UqKqVVvK6rKtfUMLZRmZwIhCAPq730su0mBPz4sigdGggQxir/DJfUpnFrvxSOjQ
Wz21SvRunQirv1qOiBzZRG07M1Xl15XPeKBFJ7IHizejVO3IaXpqdknHOGl+URmm
dyP29v7ld1vkBDX1Q2jbqBVd2CErK2gLbme99cxtzwLKIhRzctouqCefVc6LWUzI
l4F7a6BVutXNF10KGduTneqTFZ1fL1KTJ70qP7Fz1xTvVqc3j4qcYHt7m7ASGCPG
orGbvyJLJlmPmmue+Qox67E4lyYGOb9KvSa7C1Tky4b8nZJlE6ZiuAEXq4n64X1s
aM8e/2bTRCzzsEcdhCOV7kaL/Hb8PiFYAUYMnU/gac2w8QxpPdw5u+19OHxtQFXr
Sfqvs5b7z7c8Adw9q8qecpBhuc+z1StsrxyspwDomP/ml1UdU41A0ixwwuNeuzoe
fC95u7fEOEIi6t767qjWqQCEbkPJr4BXVmW3YpZaPlVEmSdFv/t3r2LCBF9vR0p0
xh822OmsYq+xb27V48XjDpTwP1j8ns3onD+BuI65jRyszCkKj0MUeb7AthidGMwV
pVJRbnFZtwKWF/mQlbz6GU6JwEs8fm/zsaCN2bFEy0Qc0wjg5eiDyoNLwIlsOAfW
xpEyJ3EnSskbFmllp7s0Z9k78jNGPJCQUk5OFHWvnD60HCcoh1x92bKTCVUNg9vk
xT+0j13fbv79zN/kwwyOViG0a21Mj/lSzkCHw0xHvTMoUdgD5Hwsylkh1+psHxhb
uIJz/Kjjjk3rszyOpC5TVbjrZKzihuZTON7aesHcB9knWX3eXD4QbjX0JoA60jCe
WNd2w7Spdbr2ZoYO5DrAs9DrfST+2aGmfz6ph7ZJeKvAOhrVD303KA83y7SnRrZx
JL1pbDAl9Q6mAxZdzejT7QWIhxd2gtJFK4zp9jGXkK7alp3t1azy54UVvlf5s4PN
AuFqsPoGbvQSjbY8iwgPGwXBYbtq4Mv9WCxgR0PuWo5x8Q4GUKcF8kyNtNJzWs8i
KK0fx9atskUI4yPZ9OrPiRA7PNW9Obs2hRzG7i6U4FcLVeYVbF5dJzwC2X1q1Sy2
47Gb4pTSj1zEuEE6erCEQYmUpOPXrMicptxViveBfbZ7NLqw5sy9CjLx4JiavU9r
QVpR5VTRi4fSifvkipw21lTsQ3X3I3KaNUhqJBvYUGve1m1xpz6nG7mqoOEr2d3P
PsBIwslvlKf/vRf7Gy3AE1Anqes0w2TjVmM402RtfeHy0EX0xZImOqBDe6v8/U9w
OANaHJ3Lnj3lJHl9vlQmGVbOQDoWFffjz48NFRBkKSgZ2IhKslgpO+T11MN0Ev+0
KHis3Ijf4i1Gjr5+nvLmPCrJQvhRf+KG+zrH7THV7iu/6f8u69dy0AVKR5POf5Im
KIVT250mkxwdyRLrLsMrbWp+CawUdNgH7sxGqt+OGy41Wz29hMn3+8e/yTycrxCh
u/MKcjEQBsJleSR9jOWC0nv8wUusDvt17CjlvKZRU3pJiTnCTAaE59KpboEIL/St
GCds24NNezBRNFDSksQfIQkA6bQCmfL8vdT07dWoUZassqU1kxbBa+TGVdrzXnub
w+NxhfY/Klq17pH+hrwQQpeIRP/2KStADdhh5WSPYE6+yyAAOIz/hwES/amaeE2j
SQ7d1SD2AWw7qquyoEGhK0rkFV8sqADnLi3Za92vss9o0Kr23IqEbRCIcqGGQZmP
h0DVa4kHw3pwZneTM9IQjMpN+PBdMLFQXmtKK9wHI24vkLtcnTRvvfsg7U08GjtB
xA3hAL0zyvMIYOEwnlJTTvD1o+g7xyd3GPKZwobSUMAPZmHMLrnULGsJMKXvVniO
O4biiZ5xp2sCVqtWXxFXF4FUbIlOyUgWCyqV50mYYu83jglScFqOilMjyHZb6nLn
P/BldVXkYQynBgokKVe+z3DzLnkH5/cj7XFdooZyNhFWToRQqmwDgwD6Eb/9qOFe
pocDdISXEj4GhTPvOu/pG2cKDgHMv3zWq2OLG8NSfMdz9ifUL1Xb/or6saSLA/cY
ZGMAlYaVOYPMTVYumzxBw507BOwee/uXaP2sbgYxOVvDMJvnh6czUv6dsIFkpgH/
ov7/UyUQ9eQuD6fKwr+Qo2XTUYXv4vLxNbCPm5znAk0/QlbGXjMpbm7pNOXCvxyw
2eCwlY3srScyuPbuNgLnURmtqU1QXtGMEFH1fOLUtQ/wh8PNgAIjtvONFHvgKsjK
LUsA19fy3/Wth1Zj6GOXF7ZyQOv1IbHNfksazsiTG4+U0xN/nBoFDULjnUnMaMfr
2LIygLFgarlDEmC0QOQpdWQCkh8zqbxlL3M4ObqBxsn6kpl+uurfffaz0eGs7F+d
oJGrFo2Ci20tcjOLOgXFQIU0jC0U9ZnZeh1tTBBm/43j1fs8ZD7g1i5omZ/chQ5u
lAtOFNbBPS/PpdTnFGFlsEsBW4UmIoR57T4wYF2yFsdP1o5HMznURhSO3FvjucpO
oEwm95QrfBH7U6TYf2vglLXRkVnMUdTamQiOrUnf2eexU2v9F0sBw22BUKHs2N4t
QPzxuIRBec237XvJBANI/4mrdRi7cqQS4+y7jRhHXCabVAdI6vg6fHuKnah4LEb7
3jSSGPQ6IChhbhO+tj/9O0K6MjDRIUN9C04QAqUu6RInJcerFIm/E9Dt+2hqHP9x
kdLgpjRitp2cFpbhf35kYDjFIGMkDkF5Yf33a7b1zJ90EZc2fJRZ6B+S82si3GNa
voyBaDAaIzgf7Re8zLpw5M7wi9zsWu7gLwaJRL3Wr7g91xyyOD7uHxqDiOiI3thw
tXxxQAN60iW7Qd5DM8QfCC6eqlbmXFT6NmmMp7BufZLatDvzTqMkmBjDBG/fZXEz
942DMIlCUwLQfVON2Z0DuMjIlmMplqA6vZmfrPwgz4srej2Fo6A/Wh5zulm+n4gL
GOXNQ9UE/A8BYjO0sivawwIsB/Q3bfK1CqlAH8yVM8zu0AT2TcRiuqdzG/4Psmp3
PiUvHy4JXj+gAJFQ3FcpxtqSVOo81wC2+YUb+b38Cfa+OTxgxQNvN0Vo0Xu7HSIw
GZMUi+cwCSeEMQNW7U49P6vaSDU2AXDEdp5TVC+wXx06NcF9n9+1CuOr3b24kNeX
ELUjAMokmyZzo1zBbNQdPLOP2z1qWQSUS/KHI361wQEpTz+kIovQbBKYIBWzxqFe
CiprTvYESra7D6RMAUd/kv9FyFFyws5x2vJLJz74bMEY+d6I4xTqCiY4v+aVIhNM
3O0IAvC1PISuxScnXWOxpxoC5pGzyePqP5/h4jIQt2Qj/BIshZSwdo/KMigDZ5WT
jwrQGkpTxaBG20h6tk/iViFp9XRJ3r2qxrA6vhB9ZreMFZGoj6ciEaUwEcXq7++w
byZvShIfwYwdhV49HIGztMumCf7+dyDFiMj10GRKC7Z7RG6ATOsqKtmj4wdfK7AS
HZQXs4Ec8/pYufJNxGKed2rgaBRx3FMA31fUwAhJAc4NNI7wF3BfkSWI47CS9nBC
SAxML7tjtukFEIyDARKvYCDGqTt2o4S7oJp27pv71bcqvamKDj0NfnWpozLfhZUF
B69blwVMQqgS8R8bWHIGRK7gvKxuDySpqcqy2bdsWzL3H5z4xrxjXnFBwTJ6pmxm
F6ws+YZgBtBQ4sxW8fano+lLdzYp8wFO4HimTzT8A/yrjQgcv5oVZIKlu3ZDn7QT
NxCwUqc7Y+fdaS4WsOmm6xrsaoCRyih9tbAZ3IlLiPn8lLpV+IVPK2L27cLpyRdX
6STkDTMaVfTH0SR+lWiihIhhfkDNZv6PK8Dyt0+EldZb5/N6ur3XbiC/2SKRJ3KX
ENFA0Mca/amhzfOX86f+1KHE8MQbf7Bw+jbQx0rkFPsp2XGvtyLVBh2f+CcV8+44
6WZQPcb4X5o1CO+DnVC5/aUHSWUUqo+dB8jEXAXeefe37GHbKoujNojLomSvJr+W
XUZc+3CwTKw0Ajrx+nrI6Tus55bRNbWbJthYFCH+6uoPoLhyDkZh5blEHExF4nXO
l8pFGrZ7LEOyP+S6sLlLmvhV9fxKfNMZnQtGo14+oZoTjaki81VFSFG1lTAMtATD
5SYVI2+MHu23qj15qNwWjy7/Fq+9CqcYKLXCDW1n7R3yZLalxR7enA1jiZEO6L6a
CpohGjf5J8qO0rGld4AggF/YyfvY8LR2M7HZMM2V5BMAJNwVy7MOpupvKQhsg1/8
n/Bz1D+Axr10VpCA1edQ+Nlq/RVi3EKQO797eX5+6d/ChVTtzWps0uLN9aBH3EEK
ZmAZWbsLIBCaNBp7dRbgkSIEmHYTcVTPTT0qUINx7LK586iliHt4sWHgg7Ct8fCL
hf11OvZNnXjRX4vxtcnq7TGcq9yBZIoYYN+cUPNljwu808ToiUb4smDiHWmp50ZM
Ba8tyoiEVTe+euCZ5HwX/nMUj7urFmJ7/tfP4QMJREcVcdCYsGuyJzL7forYCKve
ii512O0j68Gun1IOQJ/tBNg1Tv9gTz+JMCZF4/PJuEZOcz8xp1yak7K8SPvjGnqs
6W5feV33/e0Y3TWrcUeXiPFN++FyouSfS4hEqEqPQzkA5AaFSE0FeBuxKed+Yjmp
4QovkeY7sqdGzg0X4m01HjuQUH3sbxW6wvqBI/ifYWFEwNGI+OEPcI0yEN7oY70k
qtl/CVkisrm8Br5kOOVugMsnolfGLXh4+Pe7Grcg0xUxZGQ5nkPfVzApidADFnO8
Us5nnJIR4/2UcoiDuDhWTeJQ8K7RwX6oMvg06C2QPCMby3MItp3xE6QjEitE/s7D
MSYH1KPzll9tBrlvvyd/uPafTz65ePMENFZq+eidLX/z6AosPBaCoFskuAm9WTvp
5hmMmrltGVkeqXjPRK2dTJMWbSWnSQUKrtTdleWDiC3oQ+EjTJf4Y1Tp4zESPE1b
w9iTRsVtXcs7qnPj+ZlVIKlmn8kMsr2bk/riTx/JcukanmeaPJWQDn5tW+AKfkzx
YcwYlgW+iNs+gs4hkPirLxd3y9pTu2/rHT5ZcDcqktYPkv+x8MVnVOt+8s+NkJu2
jhBYI56YaFU4sO+5BjxJ15IRMuKHleEX6OnLqla7oXOS4r+FxSxwpUOeUlOM5OFK
wf7LG/ynaXTSkprZ/6ai9aPrQikEdEuQxxd7owpPzttObUCzwKj3CCxnyKJY0Crq
cIgGUvBndTzH/LKTZFswGrqF/3C1ngxrU1cUGeCSNk9Ib8gYwLRpmYqXl4wyr2uB
8YL3K7fcXZkwUE3TnTZEHHogzSALb6maHZAk+r3c5bBMX40ixzNF7OX/IbWCq7AY
/KLBIdYN1bmTVJDHBnRTTVb7W4IKmjZM4JhW4XtBU0BNSzxzDA8/EPMGYqsMo/2T
Mzf+RaLsaGsMAGWf4Dzs49cdJVHQcpMwMkFt9DRBt0YBleacfapGU+3yMXgg180l
dMWzGY14HSc+O857aEYXJdPfpcahiPLyGJf5Wiw2M7avyp8/Ih/DuOTyknp6JpV5
/smO+Q2INFTJciRoo3/zACPmIh/dgkjPd/H2lA0ml1VkXMvx1bAtqO1qmq3xzGE6
fcHSsaC0tRsDpunaUtYH6ZdTYChjWs8Jc1H/YgDZyepTUCFEPVjyHsiAlWHCpRaR
KutJhvxVm/x9JTMoLa0oYQY60VOzO2kux3bMtSCk+9rOgxuEwKmoH1JJLa1M7pi5
YHWNUCHOZDihI5MGb//KVnZ7XF2XXtDZVOMQz//bgkqBsXkw3TGgloqt8zuLYm++
C8DcPVBydIbnuBzTkLPvZTEZa1sEj2s23EwYKBOX4Rm26tBFyrSoO245SjQ4gCyg
HWWHTzZDrBvX5JvyH0qnflmPKX1nhT8oR6gVU9o5heia+TTXBzlard5mJ1RPJ/BH
6qdg6yYJ7lMLj6C/qSIdoCf5rnoYcEQ2efvVSO/GWeJvFuNHZeg+f20ubPOLfoS7
BRCO9P85kjmBIg9hfLycgm73pMIgPtSLzoGujA0s/6OhFtou1YgLu0put5Nke+Wo
Lm2HDXJXJLelGg85pDPLY8VJ9BgujeEz4X4RNXOXFSmUBwZXhSgpB/z7ZjfuP+Bh
roG9qGUO+f3E5JWktI05KQ==
`protect END_PROTECTED
