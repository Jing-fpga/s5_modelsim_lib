`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AOdlO0X39YaqteOAhh7NgoOwCWxjAaEQKThFAzhwO8vBd40b6f8LKIjMOB15lg+A
kNY9IDYIsVl/mJtjrVjJY4dMPyE54bG7OQe2UHhcRYPbybFcePq/D9FSsiRgbdvo
WxNyrf8SYQhGYVi1a2JuijYs1+R4H1LlzSjShp7lhnMaH78o1ZjQuxEtteDgnwwM
KoStcm8XVYMlefRz7WZwuxDwrJNqROPiwqvMdiEvboqPD1eOONHKM6dnXQO5e8p6
h5voofskqtgZ+R9OqMgfFeEZI1XIm/nYzz5KdjiJZh55LGlqbN+PxK3CV/YB4wVG
UH+y9CMX55nXi3YhpIG1Ie26mBvu9TvAQ5SDGhee1GTz3Kn52vng9EIAkQB4AHZq
Q4AhMyY1OV8QnhmTpmUBn7B/JSd8kecV11QsrlSuBm48DI8Se6lH+EbZcifZv6Oo
zIrzE8faBzTBOcRN//1anyND6ShEduYcT5+HjHFfPUhm6E9s6spKsB6tfDTQwx/F
u/izHYh0HUoZgLFApRCu5JrkdMO02yUz143J6IS6FMpuZv+z3R+WfhrDogeL4tjX
wxoyzK1EwiRpkwknaALw289zXHYWT7fl507lgBIKzH1/VYMxLeM7SanGt0wdRn7C
tGvgHlSRMGJbw6OhrnYkV2FQ/IOwDgBkAlryFM2tFL2JPsxqIFJhKj606yB5u1vl
059Q5AErNuJjiJdIKMmlhhk8AgKhEJkPHedr8LXOEv9YCWtZKhBdw30iiKMCfv0Q
gDB+Q4twFYkY7GDQNe0OYj9iRyIhJheu271XWhg2Gh/4/gUync/0oxlMZpr0k9Ng
C9ZkvFgVVM3E3h2IYJBNoOj8iCTF50OguIQz8V0F6HQRR6n1aXQXvnKIWf5AbLZo
4SImFqqDTXAeOb7u8x/YWdplNmV0o7jr6ZVvSafxbaSMSkxRSBd+MGTuf7xEnXNQ
Kw2uKMozaAZdlGBBBye6JRUfs365+dDvNN3hqguxfm0B+bshNfSqro0bKfSU4phX
5yeu6pIk7w9gjhQ6znxhwrPcLK718PwWDGciV+CoQChD3epYZUnceoeG18bp5zAS
xLWLOCJ1vnrK/dkvre6Bsl8TBJV6kcwPxxo0wwJRNpz6gf27hP8RM2Mv8yTvIO38
X4Z+7upLqGFsJfDd7ZRG0rEWdDU2s5hhqdT9FQ9sPt0y8g/HkJzwkElL9zJIb+gf
asX8VozNCEJKrHIVAIdpb/AUaS2VYB9cU/Y7/yfKM05A1ESDEWbCgw4ZH5+boE5G
obUFzItwBraUiECkooSXSz9J/+yPRhSbVz45sux5NAviNuMgop+xvB8s0UHa9HXP
9LXW8SpkwRi74YGXW92wg4OJi4ZqLSTMocslR5cYK6ZdS7Lr6VsSwGJZAoWwpGYU
FdwLqybQV4UVzkVJuqpb+TCj9LLN61skN/0VlpojILz5i2GKvs9ZJHU35uMeU0n5
UGQzLkz/US0g5c/xirYsD/J4Sb2UIHQ1pt4/mZJP2Jc2xnHINgylSpUNoIVh6jWe
KX7T9BlQS1KK5GLcHzZDT0mMa+CIVYPTXsX2bG7KQwT+gctf+C5i/sbPcSWKy+BZ
iNt9sfUxYvOkQEdFirZc+Gly5XPUW41Ns5AL8ap0rHAyhR0/0q7X5uj7mJnHP6R5
uZV/gmV9PT5C8ucr4W07Fw==
`protect END_PROTECTED
