`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0fFDfsCVLat3phK6Y5FYBZ9actgzbyTvsSgn10Mcshk36J+TKGwSOxKHemvzL1S3
P7z2qqnIMroNt9BHccEvTjzpXinj3KGjYZmWJNN6hHrj3l41fNL4XOuYSKDAeJ44
BAyH5OjjfFV3muHAfpY5t6I0p8vw7praSJ1AXY4QHf1J6RLUeTh+RghAkXb7Wk8z
OXQUNo7G+eFjp84RJWL/bLof7q/ZPMKhaQhkRJBAwfVBc6uPACgx87xmyP/Vk4Oq
xYbXcA6l8KIFT9MadjTMEL72O860UiEYHbF5mna+Caa8JzNdZwI0MPClKm3mYGOB
b1d5vF5XJyTCfMdwPrg6HBx0ILN7vqLpQBxdfuK+Y11NHjTxXDsHiJRNa4Rkj/mS
fZikLvk+Q4BQN0nnw6MCEOQFayEDB3Y+8xen4Mi7/XWcp38E5r3gQDDRPWBM7QKe
4j5vgkmqP7FEc02ge5ijpcz/26wJabcgwiFGLYONFBvt30t+M2/DhpmFTS/hICvQ
tq2SWhxeVk7JWwVupvhfP/WRjLRWuPu/l3YrDgHRlyfsYD+WtzX9YfN4mvjsM+nO
07LHLNbA4koVVgV45BPYOp999XRQHKmPzw7bT+2S87Mb/rp+pVMzcMp6oy5vpCAb
E01wKrCFSHYto4ZZeLYbt+5YewNaoA+gNbDQwdFz2hp6LjVVvY7rs/eaZWVOVqT9
7giT4HvuxRerqDKAdl97I/tcrxm7G/9EajIigBCWyoXHuu1/UD31VBHdfqbOEzL5
fS3isJEVRKA23CBjbmcWPz1+Ll5fvmKoUFQgmJBS8fEYt6KRmf+Gz5ggciZHp2/O
YSI+fs8TWSiEWrD4Ym30vOtFUV0pSjax2tVqamenztnDWIqh70VmF0PhPHh48ODR
lkEEb4mYlKTJ1twPwnUIZeEG/bD0ALMopXWYvKQ9osfyuYzdWDKpeKt8POeiBjUh
dCaId1cN8pQunTikoqL7XDed75IbvF8QbQF8uguYaHYbgJrjS0URZG67hvngmlP/
Ghx1TgzortmxR12EIahO0YWuE0v3kNBqngOIezvz0SO9kWF8DogLtSLFWzTOxr11
eBrjQS6OT/R14QQ/lauzT2viMD8AIeHa4+NxULZQgySCIeHHvfVKUvuvzrO2+Xul
W6lSqMPF1Aokj9Vi+ASy0U+QKnoAUZsLi07KiIulMu8BPe9qFPqxNUYJy0hEeVXg
BZrec9hUEt/wV71QTTj+Oc7wJZp4zJRpjP3ro0TQ95F1IFpEl7vAnGjKcvUjXUqF
f/yXA5rc759StKJuW/3noHjTPX7qH3BRRXu7AlNSeaKZSfQ2IZ3IescKqtJgssuI
d8QcfgzqjnfIb+0Ji2U/1pbz+wugEyt/XdrFXG7p13GWB+w6QqCP1LoPMu0ua3Sc
gk6gL9dUSDFm+Hgdo/TsIa3XtbtTbehG1P5CGdB4T8INFlaNI0I1lkSCRXQtv2Hs
hXK8J3VfLnLHBCHFzqnsuN6GAZumDZ1axnbCxjfyJ7pmT109LI2Tt85q8KCH0+nY
BJKnGQYkTzU8NXcD60zImSsRvOI3MF3244QQl7S6hnojz2Yxjkvv0UG1HtV8bwRk
xtCe5igMZwOboEpZ+7+xpp5ZfTkAqJujwyzJQg+e/3zTt2BFJzFa+lU2Jq7sWSVR
Y8dHVF6sMglRrQMDW2wdQvnrTKSB2DNl/D3D423ciJCD62efpFwsGXGT6H9uIRsA
+5jqQG1Fah3nfPNNMI+dy3uNIDpTbJuB41clbSMQFn1gjbtZbXt7KQfZgEk9G8RN
1gq0JrFc0v2n6USDNIy67zrxYuOeNbOnad1Hs+OE+x+JKmPBPQz6xRfT8ZmO9cd7
F3ifNyA0Hhsr/0nMCW/PhED+uQ0x4iNHOEEirXqHYOSlHHD7LohUTELojM6Mmrev
bWltPcvBXT4JmQb+I96MXKpSKolgILVwFScXeL/7/vpMFW7kfWR3p8PwkOx6sbnA
RMw9luIXaWaYuvM0drd0Z+U33nD3xgu64t877n6rWllplMjOUfZi0Su58eAt7tjT
Z9CRSC+fywAmAQPa9t6Ldzi8LmNWOCCDMt7fv8NtqZWLl4DJP30Gv8XP4DbWteQW
MuHShQbcPei+OhcTJZHR/RhMsiIH6+Qn9dhTQ9lpFiwwMFQgaGdU56xalt+7K6P+
912Q5df+5+RxfCET50r7encpVfspNa7cR9VuZYFyqg3j3zJ4neVjsBQtTLpQkkMa
Rk6V3NEKRcsc0q34iEXPUtU/fsZa2OuDHoxQ3w0+zW6bVjyQMem4kDCg32itBK+g
KH4+fQBv3KR8D8LHFghYaUEzEhZG0v4CWmyzwXer8G2deBpn349rzqXjdaFd9lIn
3vHaafhuZ4fngJ8WMBskBV9CG62OdIaCVdvInjJ483SQgUtrxcUfRicPuAwrSouJ
p7L7z281a4pwaMWqPEeQ3w==
`protect END_PROTECTED
