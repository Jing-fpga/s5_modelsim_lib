`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x4wXXP90+7O5IDl2k0I4e+9xt9q7h/fy7+uIg7wAQTZncW/byvWeqY7PO+k1Fp0l
QY90hkcVsvWUZojknI7jMm40uLVgwWqPgjL72LRm1TM69JSva9cBh066Ttw0fXaJ
+0UG0bHgvFgAZIv2BAPYiVRv2mDUYzAxn0Sliz1YN1YiuKVDPlv2Ehgg3Y77jOru
TX+ZRO8Y5dlxU13+U9mTOCTtSRXHRMdIWTsoNQXJKsogBA6nHwJJhGuVQy0LbE5r
JVK+zXw7b0MSXPt4+ZaAXp3hChNsGi+XOx5szTKeomRP2A6LLg/FV8aYSihCbxX/
kj9XfpkiihrFcmA+w/Gj/9GIuC4wuYpcrHk2M4VfJmGXbb8smbqs6rnBSF3puBCa
8OH3fOOLNznl0XzPXCFV0zRT1/kbejC2sI8/9IKTi6fWgzQiBoavu5SOIDnQs/2/
qGIsJFWGP4uEJvBiELceeA3Jfh2CsX2WQoHmjUzk4JNAGB1irdVyiPUOBr0CnqOH
javtPjpG4EF6EXLN0EUhncy78XplbZc9TKf6xjpcY03Q64eeMFYpb660nSeQbIRc
hLhO/K59Z1nRM8UmylVd6se7jjhE5ilWYSvr8MSW7mMZ1HO/mgY/fg8BbeYLBDnU
kMyGvasg1cEd7fH7h+0nMqAaKysWX8BIO3AePqLOxczbpJCXdnZ4K1umNRpNsHqF
ZzrPL3dya2U9nlv0lGFnMQG6uV3sWm7V7f9C0qZUpAUrDmsFudsqYexwDXacyXox
lybFScBDmP5M1Fo0oZ9tajFOCT8pFsP9QUOzXAZnpdHLGSImCWxP+LNpLKaeH0Po
FftW3Fphd271lcTb2qPQRJN3zk08ug5d94APiFAQosrLApBo+4yW/EOcsqkTdqQG
Z2t4uoa0B1aIaVSQ3Pbq025SZSda6y/U5j1E074HzlyeLgUZY0C52pO5s/ux/QCK
E+mZcFoNHWKYRG58sNeOZmzGzeF+QPY2t8/gTKCsgXUgQAuGdqEgqv31w5I1C8E5
LP4Qd6saVj454lqwsdIA+eRTrWlme1DZ0sgQgN96zVVU3ZCWld4+6MhLewPEqL3r
2oixQV6BFSAOn3wzQoMrx3nph/0TPMZyUzPsvhkbIeo39xGnfWUz+gf4VXFHRzVe
5yh0yZilbRb0URT+2535R3oMo90560k1g8WNVgQgCwASFNSJgP7GApEQbmRFZAA/
KLO9SwKJ9R+QUPJE03MbW3CE4K4hX4trN25BTHSa1icoEF+W+A1blmCC8ikv1BD/
B1FCt+KDDfEm2+4wFmLSPkGzZdB5vn7TppGajDh4Bd40r8RTlqJeSWNCbPaKR7oO
KYSTEuhF1pKnH061ghrWU/PL6fb1G3kqz0TAwouD15SMRx2wShtfEDqvrp/DmTH8
ifQ7oi+wUznu8W0/RwwU1jnt/Ry2D6NsMOBpmXVT5Gmyd/OMBoE2RmbPSHHS4uoo
BLYSq56UjO24a+re8lznh4xjGl/LtNzGioe2s4w73PPZTxzlZHKC0BNnYeBi9P5U
GA48eLGMeW2CC3rtuoQchAPzohAQK6vuwOrXJokOqKrGSUhpm2HW9DUuktNbHnEl
P9HEJbI2KopW25aTpV5QWZxxxeqLpf9W1rR/89U9YhM6mq2Y55Yd8ebFZbyC5vUl
8NK8nbl/w8A3gcH/OoXbB5OpKOHhjMib3zcR1HU5rJKbMtfFKYmhypRq/AA+Eyir
eCC+JesP3HctnZBUj+N4IkmxqOeaI7EQ91XECczESTG9Ryjd8maQwLn04nSV36B4
iKv3e6+b4j054E4PSp+HV1OBuPcKwbXNlxTB0ar3Fk0UmxLZy0TpJsmZzA3erqQk
zkCsqJ7JPWCy9ucRSZVUoiZw9fauUsCEJUq+/qS+94BUO+7x8oQrh8dVoQnKYcEX
Lcs+YbRN6lTgbyB2JCyomIh/nt/lk7OwsT0SxzXQrBoapVWg6aglq9Yg1S+6la05
yYNboSgDBcDBAYzGdiXKJZQrNzbyXDlfPFa9g8oqPhYGe1lRRmQryb2ccDGOqdiS
5KL/WLsGr5RxrdbGkZo6TSK7EFCJDcVWkXwQsVcyeOBPvQyPKsG/t7F2K++hvkux
XWwGGNPoiDzYerGDqVuvqLZjXzHQ0aNea04O1vVZudFHzDnvx0gYezoyqHA0nS7W
4kddpKfZXcBPpvGTQno0vJBFWzDfmyTya1uBpj6M9mUGKybBDUEUe7Ux3YJ4LEf8
BPJmQM9TRGmaGUFgbjAjJXC7XadM919E7lyjAc67aDVQnQBBcC4pB90IknkMF7Pz
0TzZbCFeQSpASlodQ2SNd5ho0pMyftzHu8YeMUmKbtWGCiB5R8AAWxLKp//TUXPO
RwJau/xbIK4ndiJGGOFuGGwgpaZHDBQom9tnhsOJJfyBT3vzHZOf3yMoEHx4x1iN
xDqU5uX6zbCYLYebpIqHZCXnHObV/65jviqMeVWS9cYbK8/XsLOYlJndo9A/sHQi
sFRUZqLhvAfoUnHxPGEg/DlH18CqIITQuwAAIS6htkmktvhIQsMmf6awr3Kwb5bX
qydH2QIikvB/tI6ZzxR/GJf4xg9FgSd+xFcvWVyWoKnxZ9EDcA1bkxN40B5f7xCb
TA5AobSMQ2IWq+ekq1By+N9fDs8rDt2dn2Bemo53i2NygTu8ouR8Kpd2TUu0S91z
JZWhwxhLCz3C1I85jkZKcI6gserXFF5WiQoPzeewtGGRyuOY4P3gbUn4HKHoA4Hj
q/ZQgmnWLDh0oN6iwz7R0roA4x8pdWiFiMPQ/yWNT+KW/v/RIY/Yl5sg965GOUtg
21LFZngmhMU8/e2pI/cfMQFFYuSsdGbNs7MYxb7TlBFAEjSnbKpffQLkazgCcIud
BWU5jwgScxRYXRGrdMEQKEOMy+AQy3IIRzGHwcxvwNqBv33K2NlpIHNyUX7c895m
CcyJwfgksnIPlYi1YNe+kwGt2OHnQVdRmPdA/XCBmLlvL8SjIE/mcsktj2GCmwwC
CdVnfZJxic6k2mlDWtcOp9ZjnyC+ktABn1+HAlxFcSXITdgghVD2h9ZP/O0obZBv
pHAeVQ4H5iwqa98yXB4jkr6ICxp+KjGDMA2HtrvW99MJ8aTTDSlN7VBrPmRgIvjD
PL+8RdJeBHEdo499K78KOf9+JM5ye8F9XP6QfN7Ib/xAAKhVIsFrx4DWbfzWaK4f
8wDVrkaKfvOc1xwQ1RZXEJ3Pf2cjnrRtHRg013y/JYQ1xNIw7qP0X8VnAOOOwdop
LceTqgLsZ0DxhKDHxjzwMinOkHXb1dwNWgt77iZZRlIfWdtiuDbWwuBqwEMqzuKw
cpw2q7sVU/Lzf94r0Wwq4itGJaS4pilWxnYQiZ7hnyECGa8Zk6W9YWg6rO5kL06b
VOPNR0Ea95rvwZ4Nw44DuHoTxVSTZGmDFSngzfNYv4q1wbuoUZEFxkNTvuKPnSYt
hUBlEqhL2ZBffUUqPX9Lqqnd2UCbLnBqiB/ujartbjnkknIUge1Y55HEo4kSdqAQ
wIQYp3tgeniI89x7rqoXsrEAx7mg/5+2vo9ciDxVVibMQSsOi0au674Be267p2wa
29H1Lu9DffBCLNtRVIu/9VsETcnt76SZ0GCof9BliGY3AxlWbqgXh+Clh+cCYlDv
MADREMv+eC9q0znvoyL+HgwhMbSMMQSR/jFxpNXmp63v6Rpdx9vAHjmNIy1Z7h7W
/oIu0w0xjMjzHZINVCDGV0tvRcJAKni336wXdHntVyxOTdEiZqBrfqPchOEeyKt5
EkN7ogjlCUX9bXgRkjQ3dElQuW4Ms48gYAA/VG2zYkGepT02TZilwuATSzuyiepU
H9Qz1eIa06fLeotXtWc1xu8ulhD/0Zt+zNOZaytm9pAhRgqksKRSUgIshFfeOuqD
d51tzP8bIaXjVCXOJyuwZsRthsUP8ifDuSNJixD56G7nhALS3tTVZioJjStdJmYC
cTjIVmb6Qt1cq0cqV4SK7UrAeKksTfyurgbTztvjvfIDJD+umX8beSRPoLar/qn9
ry3I719uX2S2j/p7SUacRyqh2PNIqPQ3eHKgE2iKGPdRKSnGXVMA2VgM5n5YMljm
gYUbe2MibXpQJKACGUtw5XZivrXjL9YOHu4pQ9DnioxfygaBY9/wjuxQxof6iuIs
MUxORqw2F+k/oZiIXo1aTd5H/YwHivKuxpLwxbMJ33xx6LDEioh5Qk/P+oKbmPZ2
J3fhMoEjtKZZcE8D4AXRPmb4LvKlzcHNq4lEEoI3kLngtNamZwTXl7Jxb1Ackpj5
x7/gK6Vvt6SAtopksF2x3QO6M7ZoH0CJXJc3xUSxSCwoZv4FjVmBd2Px96wPBPEp
C5EV85ejPtTnwFcu47ZeTIPJY0fs3p022ZHk8P5aF6RAXz7+8lQ5x4bJWY4wWm5P
NIdIov5dM117I4O/q7npEhHG87nOzYJJESAE7347ntdQk1C6PCjO1I+ha+TZxKs8
9uNQAtQEFZuPjgdy2009WWxMksrpCdBMe6xxk4T9lsYHvXB/1Fbo+acJfx7IzFbb
RkBn9OPBsrWye52tUVBiugD/REnpkJR7+YbtsV38WmV7/ZQnkEWiUnhiOXTmz2rG
++HxAM7kVRl51gjRW7NR/UlLZ0qpojodJhtTo7c9MGTzdILplbMyPMuOKX72eGnN
hvKiCgVEb0C18vbgTXqDYIvyAxrm9fu6BTGGOrMnWBJqr4Y7Qu8LXYE4/VluzVN/
4FiaBFVSmZxE/E91PrHq6gVlgxToOQx+Xl1uXeu+YWjz5jVLOzw4a66OXSX75djM
uuIiL0jgIBXDvQRNYKyIPe4R68USBx4bp+BRUlBOwIzj7wvY2DrrZUOybVjlaWH0
QOAR9G3k/h102vtHUZ0Moc2pZPT31lbRQ/FqkA9ux+t6/wWJUaqQPiznGmpeggJ5
9zbp3NLqvi/VUWsqHUkgjhdHdQG/IQYlKo4fBG0mbs8=
`protect END_PROTECTED
