`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qrr3KS2WCQ7r7IzX/6XVPbqNCYxsb8djbj1r8RDMWqE02dovqwVxGYWViYCG+FmG
0xwg+pzI+ZAeuLojV4XQe07mJy/EN+mXcoOMPcE9172jHLnUZt9wm8bb33ngAa8O
wta325w3R9nUrLsHU/08u3VqzHtDwnpq4U9idUufekCWc13I0v7IFCq4Iz9zAjJE
KVMT/e+HcxqJR9WZLHKdntx7ERRFZjv/dq8bMFEhXQIAkZO5hmPIADgFRLc67w2q
RPN1j47WCbVAM+vrm83dwFPO+0COKg77wNUnnjia6XmYy8SUjiSj36P5IaRHeh1l
onQxroIyBcyLKbvmMrtV1THAT9kZSqQgiWS1X1C3aCqw/59Bvy6HJz2kaBzb7IPc
zbD6wWSWtuUj4Kffe4wPAVx2EYSLVnhugyzya1BviVrk+AIUexnWK8AYDSFnioAK
rGp5V/G8go2oiuD7ctlBQApabzgQhFdtySil5nk8xos=
`protect END_PROTECTED
