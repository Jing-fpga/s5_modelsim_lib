`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bNYPYcjgxV1FcODs0iGkEpKvn7/UsHmvbAw5jsDvUmFaMc9aDFm721oggIBP25D9
k3Jii9MSzarEMY4CxD7cuPsSPiQK7P25yZay6btjA8uQjrljeAhPUtIA9IDbH9bq
PQ6o4JlX6zCZBBCF3QsmLP1tQu/w5mKMZsYnCusZP9MPHeQtRhS4Tr/6YXkJd6HF
eKV591d+yfNgaiXIfwaEkv/xkFQtX1GFv7xpPsVIha8YKUvpV0h3TKtibEEUz2Dz
UPo416FRwGw8j/bn85Sw0XGw9mDmT/8MGHdiwcQDpIpHdsQSEhKL98s7vPxJuXp4
67UI7L6iRn23mXAY+Fi9dNeSPyHEKm8AhfHqDMXKCd2Ym0ZKZE7LPSSuzyqYxAGJ
6+jATSmWWam2Fy6VXwjUXnhamUb/wRGDtLImhjkl5bDLbpyBEQIh2NR2JTrTGsm8
i+z2e3HATMYVyK5OdmysMWWheABxr33I8mEE9G/tGI4HfGc/e5uX4JmOzh/3LpI0
erID92NrzhVdVfHenWNc0XHHwJwCVsGbY3/cS891kbPidkaIg7P++JxkgfWMnKbM
oUlO32clMriMdb5Jh5BQrls5mMY/FmZqc/vjg1XfIw96jGLy+rv3XqsSokhm6kJv
S9jGOXdtnK80GOqwqvruTQ==
`protect END_PROTECTED
