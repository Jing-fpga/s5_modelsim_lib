`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hoz4RlkHhByMBWnqZcdLXzdG4snUASvNXLpa9JwaJVub1U4Q9iCVgIfzr3EYDMdm
/V6FFidIZIhb+pGftGUdpcwYYuL6vmvoOQu0Jqc14cjqbURgjVUynbOndYwOCenu
TCm7ZI0lVaUSoknNWJv92gwVCA5LloiuGeEJgFdJGn2P+u4C5pRpHUOKHXUQ6sRM
MurVtSGe1fZkk03ctQlMlxAF4OfL7VQ8v1cbvq66SMFWzLqb7l+Gwb7c6zTgv4I4
nhR/JXXsic6sgWCjVixoEFUQ0h9kd2hAK+3Ht1jqwt+RCt1HyQFIn0FYFkVuIAI+
hnKEnqtjuGbi5dBZK8+jVGc39n40/KIcghF4g4LS6MhupPBghtMkd8O40th3NrZ+
rVj8dlDXhJjr6tGsWZHS2KkifllUIcMbKdy4SPkt8P/FSL/w9GnAC+NdNoH+OLMY
kq2nptPM7yyNS+4uwFzKAQEu+AdrnJF8ZIal5OjBOUy2NwVWSmFT9d9pNlbmeqa5
09jp1yrZI8GUeQJmElEs5oxJg1oChq8STaAXhp85b3P58IVf0TZeoYDmyAzcrTF1
8IoSadu1+8xsohXj8lwbJJSyCAI+AbFLSmtPdDUZr4jfWSeR1GfdOgV8x7dMMEpD
4zyn+8+WF0F1huqrQdqVhWw9Mru4ym90FItsS57Cup/Mq7074rLeRAhuDqp58xWu
thoswsqdjMU+OnbL5VtcIutjc5ZSQ+Tjg2y4qrE/+Mf+J+L5T7LJtEvwhNXX7wvD
v5qdmHg7V4FYtwoxR+i0rkTAqUPCdqoldtB9miq5mPzVWymHprT7clNWmmTFBMX/
82UN3pcWtSskkOHOfwAMLsuUF5DgT42m1wVUlTpizVMCf9a2tOxMJA8UAqWUMtbq
+GhCNWwHtnZ7rgXEzS6RWw4tylYBDZS8Nm+QJDYlZiuLrMSdHI83pmQ0FOMk+nsJ
NopeRkWrPoLML4IfYH4yxugYfyV3u/k6GhTr6GIF8GydYgCfT6nEKeku2m28+y5D
trfVda46NByG18g16Uc/uSyWE8bxfjMJC2MdZ/8D07yJCgnfOeE0v0LMqoOmTibx
+P1pKoo3s9ow0WFDWqFnb5z5GcU+iDkGq+46P39R19gwAepKyWFzvxsjbmLYk10y
W/uzpOjPAUFF3nEZ24LQsaG6zwHUMthesI50nk3RQ48WgbeGvkTXVJRh0LQOtu+j
K7BXELlKZWWpYioan+oAj5gTvMBeXm+NAYIQ7Ck2rQHE9C5TtlsDX/JgU0UxqV8h
rS8NCsrH9SuU0Mwpjno0/ah2jZ+gq2YLMWNWtKjW+73WVJjtVeEVx2NAkCPB9ig9
aTM+572Pis5MrU/+4NRWncD0vnaTmIrMq1STxLOP//MgYlgTkMXOU9+NIP2AAOus
RPJyP3nXAKH74Q0bz1a78TX8rXL1+qBDpWFSSWkDe2UbWtkucrdPNgsQrxQ1+Q+j
RQ/roF4WLaq09p3AMD4k3TEjdZP3AB6kt0WxHb1mI+PnEUy0jizIyfA1vyMF8usM
oxfcpae5/l8z2DdOdqWSVu0tCmefcLRbWmijBE7r5VQopSkKeLlDFQUOZCUsCxBc
gQFyGHcj7gp5P7yO2cbO2ycDhET4xQ6qyJ5pZ1RPOxpUTI7geUa2xSGLUJyH320j
n0hwpBxNK39biKWYUNLYgVRZ7U61RMLCQ/JqYz9jgnbnELKkjKRdxLlSEJAcD3QZ
Sq3pzn5wrxV0+/hgPuavSe/9PyliSCwFq4nPmPpUrBhNRBpWcLIEyHQ8b4OcHnuv
k5J9oTMdotS2Ac+5ZEyPAy8jzOW25XqOLZXQu4oPtUmXV+DoOdwgVEOwKKYRdtfp
h+/PH7LiMRK46ptf/zICGDqwddI4fo6VbOAHrrCljMIXVZImlrhm+VOqICeqodGj
pe6hro6Qg8JDiz1n4/cJzrI8vic9OHWVQQ9f97pTP2EPNL1HGRBRUSYAS1put+pK
SI52LEqmUyeIC1ay8IxNzN0KV3GNYsDgcKb9iEuJiNu9FXrPAcUxH4n/AWLp4E1k
d5z0/cBiIJxq3j9EemaIW7Eue39cT1MbdLngV4B4JXRJNljH2BPylUS0F1uw4mso
5zYyu3wbKsbv+WLh4O/KGx4W9jXfuWujBRLktCZztfAE0dILJVDqw1dp8DvqPEGg
W8A3hYsjuNfZQuVqo2N0FiRJKQCx0kK821Ry3r70ME6/cnoc048+FN7nkGZyhRuk
QuW+gXZEHNar+fXTQ9+a8A7Qxowt0oVQ7Ntyj/qXlbKkIUSzgjXlbg2Df6PWplBB
23oigi5SYKt0owyqObGB2mbTG4aM72pCTwBGR3lLzNi4fAfrfkxIpApw1JC60U6F
4zNhoF0Ww8ub8tIYL0ZLVkYyPAJYG7TZTOuntpG6R7UFTK0ZBqtrx6HK3BL8GT2p
IC/b7TkqzShG4o34XN3vVXHA1HKKEt3PcWo4b+PfphL8Xe3wNMRPDDAbtg4Yur92
T0xxttulx42S2uWziY3YLqH7fuSR+7+y7utRSVOq8ddSYt5OJRLqiALJ9P9UKKo9
OmEq9r+2HwVR+5/6mRems3aor2whnZarOgoaG32dxGczTTAEBvVPDkNUI0iqz6PD
swZ0OvGwLRwh0b5PDL/y7+X4cX0XHfUIPM2H9RLk1lrLQXbQsqc3d1RdPYDTMiNl
jGKncOQDo0HKp55Quv6C2NO7FmQVodDTyXAF47OPtWPVBp6B2u64h+lSTs/KIJrE
PxwjV/95pohMMqxOWyIEByomULXsmfqg58ykiqngCfHwCExnzD9IXH+kNAsFgure
BOE1xj2N9RalzrE4BZm1pEyY5U2ucivVaxlBbpe+F/XHvjNGn8gPVM3Bi1Vj52Dd
FT0hMzzwPTduKXNUEodmESvHqXSEOFoVF9J5loYvVgur87qVZ6z1vnJahMM8Sabd
BETVMoX2rEwlyOvyX3AiNHM2We9qkiHW3rJfPiF4mipJSbhLACJGp1m/fDlCKPw2
iiBB/DkISYhxQDsHa22Wf3YgDXQgsDAAt6zV5NnL2n+QcfQfoMGuBSgubwTsJRBO
9V56MyZAQWXS+aQin7H2QG4WGMoO96vvS1VuOMpuFoktd998lo84SKqosYqbGm1p
5LWj/7b2F2/tHalE/lTPLUj75eSJd7Xk6BQratySY9N/1wzuWItsAMG7J7mFT4Ln
90H+wq0tHiO6P+VijP1Ui9xAsa/dMQyZWeK8QLe/U9mMpw3Rcml6D59D8q8TZNYU
xAIGXbx/ZsU6JNcWoz/9510xBQudfXLfW4RZDgg2DXkDhl3hISfQbQsey33Cu1Rz
jXn1RGgFoioyMEJo4Q4e7eUV6XkMkiILbclNxQBI+JUvYc8+1y+SuP0b6dLjIXOZ
g+IjtLZt0ptdBOMzI+q/gHpj5G/Dsb+xNGoG82K/zR6I8gPzIDiuilgF7AN6vgYW
khXJvQUlNcaTIXw5zNpRB3WJLQ6+3htisCIYOIONqIKduai3RS8DWPjNbGAz+Ak5
O4PZxSgYtuLit6yPPGvVPn+NhFS7zZEoGU2bc161e2gHhsDLTFistPg91Aw2q1mn
YXI8gOeM/J19kAIeXWykpJU+dFiCNnohw5SstZvBgfbq7pVT8cKvsz+k4HRtB7M0
R/zk7v8VEiqJED9KEGw4gNpbXGt46Ihhn3aTCFSnxrDpoUd6a1JF0ek6kFyl5QjI
KwHdTSnjzMGxMt6WYvxVoSL3ZrC73SwzkxEAIyoRVvffSx/no4ESuZaVtpTsXfp9
mlFOVtqiq+iv0cE0dgM2QuNxswRcwxD6wb1n+RcioBJzBuwsuA6QyhqyyXjVTEV5
02STcRti0XEv80MwQxAEQX7LB6N9G0FPBU/XuyzxMnP1eGLgga4jB48YpBGnnXOI
l/eHHJ048If9eBCLyH0mUFg4Lh/fajNaMqu5s7CK90y8RMJ6tDe/4nfjxCN+KWnb
5ZwtDo8ne7d2ZYtS/e90uAsOnLyyqF+DZplUIz5jWdS7h6LxZC8Sry7b86YQGOm7
ZU24DWQgQTiYIdslwPAvlgG0x01nInTi/ThMk63FlSwbQKdvbXwcCXxuFoPRawR7
YpFqH4V6jduB3cpUnhRA3FIXMJKyLR3NxhCQ17/xNHoo9TkNuIEDfzeA8SgktwQR
PJj8LlCHKXyy12JsKpAuhYQ2usPCugDrf371hx9Wxana5LiagKoIWi30ob2nfSBp
JNYAIoOg/0q6pmLzQhmUjOARCshVYJHXMKNrW6R1lSN7bYP0mjdtWNo7b9aiyh7z
EDNl2dCFCguixatScygWJB8FtJsTEelrVIGi2yLBSBt4W6y1+ycUY61uVPBpuB2H
epw2tWf+oI3CI5pRM1dLG4h13DPNlP6H6Phbpw4/0HOHVNeqDWVjSg4yG0k550gg
PF3W+XYcmDZ7wqv5spmiIVhXAXIxsg4N1uq3le8FAMxgWb5LMur51Rn0tkE5Mvrx
axG0thMq/PLWrbbWZB+9N/PFbt7b8Ugr0dbbhtjesyqlVUaxU+kl6l8nh57Mj9Gn
Z/tOAAIKxIEZeyzRVdHwNa1hGdD9L7PretFmldYfnX2FGsu+2UlbVy7TGEgOmuW6
OH1K0JfNKVT6A0fnFFHc/QY6P3vq8Llgv6WAacviR7EHypGJPW8LSitC5N79khRj
hU5D5q1x9VqhUrt4czIw7HJnZF8vT+dNeHM2XZnVj/wWsfaiaDnkS+Oa759l5Sy5
tocd3VM4OmENoLl/HCAD81HYKMIAKJ9dc66gmNO70beDMGCl56IRdlw+EQLDl6Wx
z954LyAxx4OoVne1nU/8GEWjME6P8SCsGJD/dfxjje5xCtHUDHkJXzvBdDVCDv3E
YTP6woQJkSxDyiaHhMRzM9ZIfEzNJMntm1VDj/Eb/b6hp+K/V5fjCpuAhUnSAY1j
U2z1vMY4cAat39YCTivaN3zoUVQVKzDYVsUXGvYGVHITkKP4VzWxzUwZafXQi+A8
3cJnhpOk1mShMxhJUEnwglRtOx59J+ocKH/8rr81zb03LaWGGyi4AgU57pJpk6p/
yy7yECSpdLQ6opImsiRv8PlfLxrRUm1FU9Xt26XphcaTaxozAQG7pFZmlcx5ptQN
XwgnRhvNdcIeAeRWzUastfYvYWEv+vcuhdy1iD5GbfKz29Zs2jfnOHaFIKBjS3AR
zTYlt0G3fBVvgGSp0jl8pKR4zTvvD/RDIEaGzCB+s8sxuUkxmtwTWBJ79fX970I0
c1Ml328OiTIqY1dYW0MR35ZeMlx+7qay8ove14IrMBlPy4pudQpj11f2LpkABVI8
gQqYWL6bZjJJGv888zePzr3EmrvcOJ7W3skkKltsErCWsN/d0dbHbR97qADDRC8T
cky5dC/FqDPhwYO8ZflYK+lB07KqXL0XjFzhV3K37Em2t8rEmU/Fup83DCdJ/Zlr
2JM9CAtiljks4YiCwPKTw37vKLfi/sqWnAqBFa+uS+4UATH0uwIVivoOPmGxUook
ZK86uHf9GvV5aP1MXt4L31dKJ/4RKsdZsivxzOhG5pMk0cDg4tTzjmQ00a0+2qVr
PoB9EQEhLoTUdIkvej3WNatW+TLQkeJT504fMkB8Sco9AF2zpTXjmqxTJ8Xu9MKQ
RlGYqpp6ptiFaYVl1Y/7PPTApbxJeQZHY+67Cr8eFSQiiDTzhLFDhjuN6rdtBhbZ
SuHlaXxj6hj86P+RUzrwgzYpHPBgE9tAWOQTQ82Zt1YoAemfJ+YC0bLpOEqoR741
1q8et77uKnhWQ7F0ZxmfFPXlhz/k1eTfegf6PBr/VdWLqAU1Etvfe3Gkc/pcoE+p
whpomtLxAmxAxSNSMxNyPsxoeFAciuaYvpmojnjlgzB1IQcaIWFaF68Ue/QpsmE+
8VHgUmXehqlqZX8A6jXT75gj81wG200m9GTvqjhw7XVI/qWsU2a98HwO94I4s/zj
q+fb9xlULOsDKGU3Hj8pGC8ryvQwXiDYhL/EdkjGwxlPj/lnEAaAQyAF8rAiy7zp
cRJDgNg+JEfj0nh6M4TzBVShf/GKWJXGuvdhqVuTX3IyZGnTVYnFqL2R5a/db5UZ
k/LGhLQVfzRbzUMC2aq+w3XyD2JhNYNvTTL4flcfLPYwM3mWTHPYVE5mhePOB0Qm
qjug/HgCiPAQNuaYs8QFWVvrtz/CWqerpO9fOL9KMv1W4V/1cwSf+ajVGkVRGcXB
ym77HZGgPqfWheRd04n5rPgQNBHU49M9a6HzYn7D83X6ZjOghEXPMxIBFGUGEJSi
pp1FngXg6fI0Sn9sDa/bsBLkqUJ/CE/ymm3cvNVnBIdMCKG4zCVvbN2+n89I5Npb
OgMd6ZMngKeaLpM5yfRGgIFfKiwpGtVN4JX5QDeE8pw=
`protect END_PROTECTED
