`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ot9MpJjT3UiOMMpcIt9CGDj6uNk6iR7KA2JFuLJ64bHN+vPv+bscxyx0HbIf8ygi
DHNYRtU+bD+QY8BUJ+PPz9j6zWcliObj8UcNBkYeN5cog1pCLJEuaq8foB+R407L
N3m6q+23looIoEw+UfhjL83JcB6xdT3WG5+d8NMJfDekJsXARFo5UQP8vR5DkoFq
E6Za9+7Ati+UIUqZrbnr7tZ7UvzsIFKOX+4R6ERMYvVlWAmKT7jgSm+aLVMaeyqQ
Nedm+4IH+s3zrdKaEEx/HEeBxJeCccKOBcRVJUFMBluxeUk01/j525Y1KYoPSYKp
HLxyGXkZ9JxPLgOxajje90qcw7aThHga41YxslzPhNXfa2OlUHhnz8XmzhgmnpCk
wqXC0DTNZlxRRvETljyx/chsjph8rh6EqjH8o3FYavlS936iz/qixJipV1jKyBdu
H9EgN4BSejnY1s8CcZ1H7jpp77ofStO/FiMmowDAvoZkwvASYKbYvTuqXwTqpZck
9F0OtbB6oi4+WTbPDwZhBK4ua6MRIeuzHSUwH1tkM32DH4jCoj6eqv+cVdGsw146
qPcOYRffmT5FRMCM5lFgN3qTLK51CVPqB24vL1BMHvPls/2GMUdUUPXNajk3AhL6
R5wQzYhWkgn4P0ccXNWlT6iwG4MmyuhJWKQCAtL3sAj2AYWYTDp/J+JcDNGPOw8u
YbQHy7gRyX5Htijdb/OqKA6+xa2klt3vTT+let3trwaHV4cJbJRTgEwOorrhRHbg
EhAJux/9e1vfvTsHHeMPHuScd7Pbi71AnQ1xcFAlBfvZGc0rMjkhzcWT/Ys1u+ng
fTKyrp/PljZVKBwuPWl/ZqivvYSELT1wlj6Dqg9u7r4=
`protect END_PROTECTED
