`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b9UvlWgxkO2ummB3nHQjv88HLQFcBwLjgGYMUzxrR6k5wqCM9GSr4ZDi3DwfBuuG
KwxoWEl5DaxFNkZ1Bubwa7Pd5VycRyjTrUnlC+5FGDRuAOmZPCjyZmw2t0ijcqed
PW4VQGexF73TLft2gatxjHs8z2eF9KR7KMUQz0jurJqFs3ItSRRwkiUZ4aUI8fxN
lC2vWGxozDCqJMir3sG8VA3ks0X7mIfISd0nmueE5tUQfno2Z4IiT74HrKkjcCyi
SdKbj6/ccGHPrSWRt1Pf81n6KaGGNFrQGvDtMA++9tXmyeBcBPZ2CJi3yW+kWEZa
AnKl6BT5OlkqN4RWwfgK5L33Dihi0r0EpJFfZ0ySqouySo/386UON45b6fpCsHfd
uUft0phEAS8aE+W8izyEyhzLsHUcpV+a8vNVBlEq6N7iVDMgWco7iMcDQ5dsTxPq
GhhdAEv5An6bY/p4QaZ5cczzAC/YH6sVqKPhDPYDgXvvUo8dW3uMpqdg/W6bcIJ7
mR9jfwcZ46Vxjil3xGCwqwWE90dQEd+5h+SIfnsUdZKO9IeN+R6cjs404SpoY95X
oASJP4XfflYsohsfHatHuimlANQDEYxQ3PT2hlOcwTFzzZ01tWOLbGHFGDY7110c
b+zD8KrURylR0Ebiymai9dFQALhqPOBbRuDQzXvQQHdTDA95p/XYCn3JQPUV2aYW
3nERc4BUE5w86lwGLtEiaoH2jxSZSQCnrJqtHQVdD3eAU8vvoOGOg8HCQrzwIFtd
MH7Y8Hz0xspaxvw0uDtCfCsFrbN+JFiRy+n7/dqSl+owz3BX3f7DsEmoVManIvK3
qkoyANIfIvqoy97t8F9jv/1cZhqAPSCA50FjZq1EIjmwa+jhjZ++NdDPl9nHPjfX
YfAC9lGNYwD2Xm+4KfBbU2zam6M++VpUpPu3sHf7VKSZxVdHnrFqReh2mMHUzktr
UAmzX8qEwNB21+3YoU9TJ6yQZdhWADYXpptUc9khIMZtXEkxH3R1ESs5z8d7Ehka
u9kxOZu/NLg4RonZlRO5EbAwy4T02+GwJKaaH1KFWQfsFyCVncz6dwfeR1AJhnEp
bgVUZJWYoCs83leADywlv76tWrU5pusGQJYNZs+6XJjZcaW4DZxcb6wC99zsJBS+
u8vv1IudWRw2qfL2JFbfShqlBQg0SRZwTa8Bsi2fnV6M62TTYw7lh2sWpuljfFRE
tOQb3ieHGJFaLOlTRYwoFdbT9VyJqq3z0DydTjGn0kEfIRfS4e/kx9pHrz3kZ5D6
UjONmHVHzjXCdIbBZRfbQ2/uh29ZL2wb8GXqMewtPXGGWKTFvK1eosNZE3vbjE/e
xRRbSLdPMebx4HTJzgUoZGrJX9n5dq2tHGhskBFk04KrNVNvPtOdqZ2xwMnEJUgh
Gh7NPbXr9Svs5rjbpcdw7+CiOoLUHAAB3zBdjRwYtC+aurnI61yw4mWa3M1XKWa4
`protect END_PROTECTED
