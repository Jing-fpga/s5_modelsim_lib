`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z/baMk3JPJXHrTGJeG8wRXIRoA/rpyEUPJ2T6Ibeo6KLdbxveNShWonswN3mRNBt
DcYtiCBu6ZvUYOtdbKQmcRuypd720vtIo4nLRUHi7ip6fjROac/i+eZ87s/fcKxj
W2ZrRYALnga2IEBfbC3gdYsfCvBFROqHDJVYDUcjDApdauqmPN8sosjBh5/blpOn
+1e/ZVQbqaov5M2ZL+Zf6cfGscEaPWdBeNavWy8xJ7xLtcKef/jqyoPo9ZOilyHG
u9sknuxMCv2QgkyFSf4GwqMejpJ2niW20CHT/luIqprZY/PnlMDCum6OE0drm/+M
RZ6RtYPSGTxwLNfB1YmA7KoW3bh7rFGDwhKJZmN7DnQdJjbtNvGVMOQGMNceFcI6
hmADvG4oCkHjsriscab+/gw53zI+0kHIl/9K8713wLvqxJIzr+4n1zk3RrzkJt4V
4euItbUtnATwJKIeF/6SbwKqgn7dekQz5GnynK4jLjCNq6BFNPYTCY0dojXR7+3P
uM5PnvWjTxjj39PlNtVS08XcP3qmYWP4cXaHtwk9u+1t3BI+44Bze7NzqkGy6zAc
Z2Co+swmk6bOLszeA7XzF+xJOudhF7cPzdV1kiV9QhM=
`protect END_PROTECTED
