`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xPlo9u4qEouCCZYKyx7XH0tkZXJocYBT7nETD3y1MlEOX4JVnnhmHbgO3ZpU1pD0
TDTYeWwOmi59mz4CqfEf8zI3WS3nmSC3ybXWJzhM2Wq7I2hvZIIiHuUx8mVesDF3
caunje4RiVNVuM+nAviWperwoBf69qnU4ibadrSQVjRUORRQm+9hJ2E9VTvcwtuZ
FeyxrZc1W3iPg5s2WYiX+J3+rqoKY7xzC1oSMqUUPbYabnCCEgU9JEPyK+mbE+He
KRRnxfE0Uh2sbc49lMZ8Gge135zcUqKoPktGTIxCCojOgjIwIdT+ppsuuboAcszW
p202IeayAXQctIHLbF4STYaAbUn2Y2G9RFk0zRPtijLSWw/OZKBgjKMf/DARNJXS
K9qOon5y3UXvsZmc71Xhd4GRq+YVy8dSnnDIZa96hNvJZlAO4jZgG1Z+b3zKxUCM
koJC2BapgO2eu7q4lbqMPVMW5ssVTyD+V808B3GSA+uFOjBKuEad9sDIQpyPmb2d
a4LZUkhRthkvakHeC1Y8XD96yr1E9vyNiB9kIc4+3wUfuokJMDrBZVno07injaCj
Y1M2R4tx4F48hSL7ooWvxBk8eVaPLHje7pugqOE7kQ2ACaUQb69QjF5LbEHH6t2H
hes06egLo/53qz2YkiUPqZpBGjRyd80U3T79u5IoMan6lP5A77O24j22MNk2oc2J
FnSOW8mIVA1C08mfBdtZFDA5sj/KiVCo+QeXngShJfUsqEdO5pYAz1o1aQEfNJhP
J5ClSXGqrjON9LCQJ7WnPmeN4iwjRG75pgpJHQ7H9nJKJ1YUoDuWSN7gJaQgSM8V
2Daj4WwGPLBnnQ3Rel+15MVIPGMLEKMuc2RAFGCAhFYomL+pHlfKG6lwYe0DWANS
uUDFMGyEOoCYFURyzIluv/HHMarZf/WaB2zxp1DyaxOG5TlLGrn7vr5kO2dp1xqZ
YVWBw01dON/DTYstCi4e5xeiYAGrUmGkfOe6XeE8GVx8gqeNMYLq+l2rk1NR4CwN
SWsr08EtinU644skirpdj1/QI9QfLvxaYCulUIfuYGpH4iTWtumPwa0SIxyRbVUO
hD08RbDZqPbfGWcOs4s5y7WmatmQNHZPfpwi/+7UfEC3FKU+8BaoKIZS3gJHBEbK
+2JcsvvbXsZnjtVNEZOq6uHQkeZjV6JePfpcEiTE2sKczOInz8N92P6KvrMpDb87
XrPyj216/WGEajTw7EqN/6+wl4IxMojpeffHYCnBaRwMrmRfV9F8OEgYvOmdizp0
s1VdO5Fl0MiPhBNYHY47htiKS7/2KtSlY3170TwPeitLJ07k6IANwkPMcHaGNQVl
2vlN2t0rtLQxfao7SeBdRROPuUfPSRsvHZYxlfJ785DaHvhxtblfz/vuTwKc3/gG
D66VZF8q6yli565wgRBp4nwSrh0nB8ZjTQefcyqcCxWDvK/THUVxg4PxbiT4pj/9
rFv2tNcBsprqul5gbzx4AIiSjvD64BIPrsEcfsdBT0JWY0iovuYus4cK+OvFGAS+
5ApqkTgoPGmsz8IWYZzlZROLpZswAbmXmRZ2jJJ3rPqYWOPgngJkOC+lYtwHPn1F
Md8oOg3YPTK19p1wxuNyFiu/PklbkfAEBomZms/o01GKLv1ecp2GcA418JU6xviT
PHCPsbN9gegLUMyzsNwFj3VNF1m3cm1/UZp6OAhMbfaXd/lfhUCGGkv4Vq5cp050
IYYgwOb2ezC5D8sZFM3FzdrjJAYp7HJ3WYOC2K7bFu61AwnCvhNMX6IWds67cW9+
WzcifnAXQIpE/fubYcnaQ90Gpdl303iLhnyiZEi+aayQZ16Mlo8oft29TVAcQy29
G1TiM63hrRUrX3zb9KWx7vE+tE0HlAjiRND0G0Q3QxNEV6hUd15qVkIdersND5cl
+9sCB1BTDDiI/cWMCoMAhE1oigLKKmOpi3mN9YXoV11PWclnMxSvZMUOtcGsxKzi
v4QPAOIxaXzhMjVY4pyWh690v5HGcpBci4QtLAH+p1T8fHu78qWCWr8LBIZ4Uhyx
EgU6EVsSjzxKdU84nTwH//H4HLiAdjYRLxSg5bM+jzTRHs7bVAG1LzjItCWL5FSF
iHunSw87UL5kAt/x09PY1P/eYHS6aWRuP0JxkofkRKvgP0R+/4GVpXAYx3pTjeFo
AyftbbQZQeilBaJkmQsenjT3Czy20fTdmqxTWLV8pCLDzZNN0z3JZqR0DbHZUS9i
5IbOXxgYFr7my8ojJktW2bpGGhU5KWUMWKq+CknPFzUfc+wL6YZsxL5KssCnb8/B
j+a5ZV3asj3EfLZ37mOv6dZ7PS3nE2+RRpA9G7S6LcbpNO2CJzs5wG6yIYVqpEzL
XQ3vsIhUONYTefkB6VPvDv28DXITQNehzlSAE9TMnh4VGlO8qjEJKu6EeBgShUzC
/eV5u95XQvSz+m5g9zUsQ8G4A8Bq1ZfcJMBGw/tAGNyZysLnvHF0a9d8av6BeHor
89dsYSeq+JcGplzwoSeROWBA3CH4A0quRZDG6f/GNM/KbPXwTob+B0E5znMA/JYX
zwIz9bCoNuWjPFlnGKek5p7IYPP/OQAKsNE6bT2E5ckypr3CEOTvJ+wByBPYL3N3
/S3bB3wIPH3SvhrJBmUVlavlSmunJaz/MGucxBUwY/Fk2CN6Cd1fVfxSNaa4XQua
o2IoqTx9WbkGt7bgzljTg2y2EVtsJW32ndFMNEx6hR46xltb3xUzUK2TipU6WTMn
p+WbWlHsnhUaynuURHithqe70LjnXGeqq0AOLzib8hUcGu4TbYydwzIxKcPqdDuV
aqk4Dy6fdDZ2ht75TCb1Tnf9WBWT/MlbrOOw+wvLFu5bUWGLXBv8dmzposi1C4UY
Gd1sA8E7Vm3isViqayBKRrcDEKVnwB3vbCeOH+jLZJyB4A1+csM0WfKavxfQRdFb
6jb+MUk37p5NXzoUQvH0gxZurs2N1ySeUdlowtYLb4+D0oL01Lm2Cqa0G9V6JaEE
qfD/dEaHWr8kc9NteZFyHl70C4S7ZJJfmbR07Jpgf+nQnyB/aIZRYvZcuqyvitsQ
uufJLHMFHCKcuw9rM7K/Oa7IKzYljCVX4jivE5W51Hr5ncrKdIcSZcy+mTl7rXbl
fjqZNKIExwEj9o1Srsc2dQQAvP4bqHA4s/rcaTRD7K3wNbYauyau9BscWkNBYues
PaEsmrksMy6DvwZi9OAVcAB4JS85MMWTK4RsESZsG18o5pMEh8v1HzxHr//uKQ4L
eVaHrQi1XzSQO138C+iEgV8S1wdfYDq3Q2CrYjUUHp3yrj3wxjkfnAEBZx1qWzb4
e0Ww2F+bdGpBPTj+szuzIvr1uV6yJ7C44VA0CYS6MVeuxTJ7HpXzlqp9y6TYsxuI
FbtCtVn6QcaDZR8jaU7xE1RYMglMrkq39oTYq8k/maWU+lg6T+KIRfXDiUlsUVVk
MvZftyuyIi+KBaPA+oodi1m+iUxtv62Jgtnq68RDltmh+j9LT2ytGHQ03XQrUMOV
PptayrMwBjk6ZrlNB/siTIMmPB/dUCxGddPPsvVg5OxkalQBoUM9lfzSy2uqiret
yPEtUZ6AuZPvA86nKhVBIquZMkCb1Zenan42P91eNptGHaC/tEHewqeB4shOKDzh
H/rb7gfU51r/9GQ9Y26cnuDyZlnyXvVUmxMD9j0DyZaxcPtz/mFFPC13Vha88Hh+
XdN1mFTXX8kQeqGopHXQ1h9lSwmhoLnON52VwMzq0cx7543LBNgXL1EHGDW3VEwS
3uzLBHyiCRbBQuAWxN48j90OI/MtJs+kQ7nWo8pEuR1TYoU8QLMzS9Mv4LywAXkJ
rqOrfgNMOF5BthzfsQJefQB+0dYqD04zkC8Vah7jpqCugyQqIT0lTdEC6nDHpwt3
q2nv3z3bT//dZ+6RJu17OSdbfuhAHbcpPJofmF1d2APZlJmVDgQDw1BDYHZ6Bzwx
P4PCOcHkkSQ37Z73D6T5xLQRaBiqSNGdQiChTcQZ0uXfzi8APTGp4opyP0Wrg0/A
ZVIIRMNMQFMJqtMGxodJvBZ5u70kxFG1XSL/Uc7q9MSQtIFidLQ6dNBtiLb8Bfq1
w7y87XfKs9SfxHIlPQvR1+1LoxWGXoHrn53BMlF24oh/PJVpXExzQgJMdP/qHj4q
0iuFcTFGoPF3D/xmXJi9ox8KT+L1AxpqlQyWVS4e6aUvz/V4v9JRt285+DSNMzRG
pD5iHDmVIRzdumou8UW3lIqrfBrrBPw8NxPzdbXwb5aTSp7OGc6K+CgPa6z0u5zj
aGjoJc8I4hOmrlukBgo6wkAEaOymkrm1/JJmehZYbgnjVjYqSjFLIWlA6S8Ixt70
awIBjxHTAf2KafkPBZK1VyFn4cgvsOrplBZnMw/tjYnlmfRZbMAO3vIAhDz9nQ8M
+ef3Qq64S1WtwsVbPGkfHExxYAn6PmFPTddawr0hxWNBK+7LPfVYdlBPJ+n/5I8G
xiO38HuGxGIaY1kWRmuMq9EsizQqZWgkvuMN+qd3dEIWtJrRbGOBp+C4bRSyh4TP
QrPji0UMMEw883aUQthf+APeA3G4RdITkv8BwHPUbdH2934GDyAC76fBMS8va1Ve
iUpXb4gRX3rGveRzWditXHyOsDc1cldcexi+dKgYg2engub1tISpV5XwR4ezhRW1
mOzqIeNL7TX1YnC1d1ehBUR2OOFvvmjjEpPilvdU8p1UJGhJ7Vj2IN5JaERiKrXE
rYkKN6fF3TPfXyeq9vcG7UWEcCGJ152yNdJI23cNjB++PRs3qfiJ03MIMwk0Aipe
cK76ZWld6oiOY1lvdWPva9YA2Y6jWhsTO+1Fen2CNazCqVhXYNeO/7xPREEXoKjd
U8LcItTHGLcPv8ogKWz0xBTD/oduWb+4kXzADPxlh8XJ1yeGTyPhtU7y0Hf9ez9E
Hjcd4jP1X1Dwl6TCJHAoHHQBzJpppQlPJzyJPRh919QeaYhadM71pF+2HW9N4zwW
xN+2GpWYKP1p8Nx3MBMdSWqWT60aeekoCJXMfH2tdBK0rXyfUQly+VAWnjO8Djzz
FxiYIk1ra9/JN5K6W9ecB3TTI6sEWkR7Z1RkOhyqVDlHBA+/UogO/BSs8jCe6fll
2M9uBbRFlUf49xYDukOYFWJYBtJXluRWu7eUUTsa6MsH15VgFKmMVqIb1ejR8Tw/
Sz4cw0/aYvO4Wvs8eA02KQ3SuY7UKofEjq8aglHZMcxOcp/hHB+416W110egHwOb
krMceyZGt4nmxkaXgCxS6BOdIE/qqhMbYNfhR1zqbSZvzzvx+X0Era1UgvcI+Umx
Jk5Qwti28YSCAtWCKwkortDzQ8YRmgj+60LQXI32IFhAh6qdZ4bZbnL4BX6BvagS
z+z+N/DS+RQIKu31Q83odkQa9DyQLUk8s7Xhsa0xynfYwLVJ7mTFVC5NED4DcS+Q
Fgyjef/BXmtyNw56O5KVoat5CInlfma3DzJRoQwKRUOaZVYAnGb9PiZ1K6XBCs7h
sZEC8qx3xplc3J9jZ0Ogu4ieY5C3Cuo/CJOIqbGcG5Pa9UZj41qSrU9PWqbu1ZB3
O9ZLQmmtflWWJn/fOvkdh4u3XGUngJBXVjzKK8xvU9Mc7FnTGJFyv2eKONo8rXhM
9dxpyMrdw0QItka+oRbWMYLTkKTC30aqqLkCCRT2PwbffnLfJuSWFvoISrShkqPf
Yib0FAlzbQFTM+UyymfSGlmHnsPQa0WV+QHcSqTFzbRf2TgrquyIbrpAAV5C3COg
q85joLbgIqizvr59mSFTxa2VnjOb5LJ2jI2ZyoWmfe+Mg7v6siiLV9qoG3rPCtcq
IZv0H5ctVHGcL1Apj5uN6e7kw+OR5z97apnDwy1fdoNPY2+eajyVEScIzQ/sI8u6
Yuq2jgmCYjLYp/feFcxCFKQlY8BA2L57yvVln7wzQ9hC3QzwXMnukCdQVa/k+Pdl
HY6jSmB4HkI1TIsLgBa13DV7sR38UJ3BJkummHMMCNetiNhNAQulo+JGMKuwLDQG
3lBtuzk7J7keCdvcEEo8EHA0EUof0qNMRC2/xJKNnoCrEmy6E34poeQRJQKjV4jF
6CCn9cHV8I4R1xwAmQEharW1EzaJdzw/iP+f9XOZSDN/HF+X7qKRlEAklRGuk/IX
JeR/9ocAy0h8XxAuO463p5rixSs+TvXl+Pzdnm/w/yE4L0G8W4IGqEWlGzeLF9ma
JtbiHr0eHFwUBuijbTkoLjCe2orTvz9Muu3lKmKIjdJpJAziZ6L7skrTQ33fM+Tc
N0kn4iyso+Bm8/l2++uAgpKnWJ8rdX5Z7zCKoRU6akgvscXeSHSxdBaAcjPBCfR2
qg8hWE5k0+6mbWHP9RKAoQ4scznYIhVVrBE5Y2flGZwQ/iTmwabK121tfqspnIv2
LIV7DfbiiPxaDJHhwhYVb5i/KrMFsuFkXqRGeEnOdWunTHiq89Lt3umudPVY24yC
fodEuGAxQb7Tip9W5XSkWL+9sOwSMpWJMTBoQ3UrpMOO+9xPs2cnwykdmZEgTE3Y
PjQoOFpazjuFdacp54wwnPcobT6hIfZomS+fgVKJmvTAuJoIePBt/LpM1xwIvz9E
B3+k46jky5UUGEzr07Npb3nuX+qEexgu+0vfqPg8gAbMjMy5+bx2FSNxxXidj1Vh
EeBwmXUZg35L+1TdMAHixxAZHQ9n+Nzl7Dp47Wmgg7nJZufxQKHrbNRn6oPdD3na
fSgGhlZj+ICgS9/o91fopk5sr/I4oQpXnyodJB63SXf+2mwDs3oD5PlcuF1bU7Xv
EKLBhb8jsq1AhQlwi1C0fi2jyvJ4kR1Cegg9x3c0GoiQHAy7OQ83TmOsDPSrWOWB
eRiTR+IhHknnbAQ1ZotTwsVq8lNFJXpQ1KVlT2gaOtVPSf29bDRmZOwIsu/CUS5+
UPHbtupt0d/LYOtKnP6sdmTmg5vNZvZU75iVhtCrtiPZa10E169wywNiM13J6y3Y
EcgDFGZbEfn6gl7qEfyv3w9rbVkf8uhGQORfCEHPKSkg23G6JchKqLuuq8flKGNF
oLZIqkpI/d2mzIGp01sYEZdLQqNOb6IhYXlnXGI6AFapuXrD+zPRqk694BRTAHhE
3V6QUZtsXHelV2nTO2arCvZ7Y2Ms9zDkQpPsD3IucPVc2BQkmaLfJiq92WTgkheT
w0Lk4d9iC1tfp8rGx+AvlAlq+8oyZewOxL5lW9Tgxeg8HjIxEVuRj0NvTu3qnLMi
DNObHnHUbBuWeS3T5QUtlpT75ZzA1ZDTkwAdFQmrH4qLGnjyP/AlOoPybRwj+Yex
3JwG6wstlxgpHOC1B8NjktfUzQNqDlvkEATCxtLO4ZsVliD6GRCb+3IjHpgch+xH
PZEYEKGdf5ZnsDyYN05qJjOho3xv2hE1wmMIpkJtqzpC1zWRLprKHV7OgMtPaAxL
0wrPJq0PTkTe+pQdp5qIFPWG5HtJ+36vhBrk7d54hQbRxJEvHOPtZ/rppmSdA9Yp
7x5trWWWLWln375tpoev4UGI38Xfz2dHPd9wDV/0lvQYUQpoLhQZcSrqzh4hmXsG
TEJ3h9EiWPT8zS9G9aY/l8qV9sEEQxInE7hzm6/A3NS8HsX5B8cv0qMrVAIr0n02
z1Gj/XnNQGNIe9hvMw/bFR/4l8xP59rGYXMvtqxzzqOIiApN+kX7+xKBYk28z9JX
rwTwTA85ApR17FTq42rjMG8jK2UB+CniqadrCauF3W4LburX1UEW6Xs1/ZwiUxRy
PnvwIQTj4RfYUI5B6mwgwVrFT0fG2P+BDIRowPIZmJn/WuBlayhmrZN6al+7XkxN
JzswGdOOz70/LTOPJOj1bQccksKpEPyzSUE7YBtPZEeDBI9a40um5fsWkKimlPfe
XdtDfPQZ7bslbN5ZffrurGldo3GEpG/52NcfxgR/Jcct1KJiFTgfiw1zhl4Gii8M
YOgJFrSUE2S8blHtTMSm697qbw1yTVK+PWde1F9rx+MArog1m+TIp/u2ISb9ttSw
ieMDLVsV8LekLnXvZvKtXKindhSMEHiRfo5oRA2gFTGEtlMMTVjHRPGYvdKlPmKY
dpzO4Zjq72Z4x/OZXTFcFR5Usq46qi8wvGAgLAHlUyG0ZRXqxDCFPquz5H6mQAM4
NM7eRD5AXCGAdZKFgdwY1f7ZWJTR/EesKHZyhIAT2CPVgpZDOJpzfbZ4YM4qs8os
BptB23Z3ge7yeO1qWbQjTnbjLTsdHelpoNuG/r9S7PNpYePkisNhaEFHVsNpjKwf
g+GPN8jGMOKv6LYYLC7mx4nAGMH1xJGIlewljMyKbZwNcGsGHcKXsHv4YYzbZClB
DoqnV9PsnTD3n5cCJUiKEqMMfHgyurK3jCi5jbWXgKxFrR0Q8DIjCs6JwzRLcpMU
JurUj17zMvdZ0r74pxH3Zky9QB1SDffN2J3h4ISV/QPjyBa8x3alWkg/YNwicnOG
AmCJJubMZqt5GgO/dWcQ6wfF23RaWOk7pI6iQrJN9JU3DmoP2D41J0hZ88axZ+UQ
OM5f6yUAUkV6ci7qZhisUig3XqLQdhxdKcRdoFWy7+VWam+D13xo7bcue5Vi34mu
EQDoEl5rwKdbgbPvCXc3NpaCL6Bsd6uqx14jnOwZlUrL9h6nS6FwSFmFiUbykUTT
Wg1UrhManQFfyDiLwUYJFyFHGlkWsW65/uimvuHm1c2kdJn9Hy2eAXHxmlNHjTqo
1poiFUU+8qeRNpS60Egoj1QPrQHkMTTsYqZqEPVQpIcKCNrnInhBzOx37IEJN0/x
Pe2BERK4N95mtizOYhfQiNj//CTlKeCDAOxJMtnBQL/hK77Zi0b3WdJ7ej2NJKTH
FnDxPAKzF3C0FaSAgejnVbBPJ2ztpbItOjZNXA8QGre8BKWKrGOB3LQ2DQb8T5BF
IA9Pa6gDuj8U72VCAuMkjzhwVWxahMJ9K7EKrDpl68T85D6BwSGilJbVriC7RjVS
0IKoxj2pffulETDPxTKYNQCM4Kb3EQOrrV1w954Od6EAStQykzF45EqmnfFaHLtQ
4Nm2EXd1qP8Pj5a5PaRZzeH9SbaHDY/553K324ASJhyhgS1+rykr2WtW5evDTpVo
gJpMlvrei4097TidyUFJ10J4c8oUIYCEZjGtt9SJSX78KgpCgedvHObM6yDrfrOr
9XhFGq5d5qyUQyZTQinJC5ViYpvI93onm0cxHT0z5iUPtBm5Y9fzBApKeslMV1FJ
jpslhIq/V28vz+jMAt8FI2VJm+hkIphzWX4huodeI85dFpnbpm/InC+NZ379I0zB
1CYrllio9iV4IpezBVLNzbDyGzyWnzQhD4Ze4dlTVQkb9zwmQX2aIJCxuL8oftj2
D1jsCVeD/AcKPOWscYYkoY1FwjzSeu6TRVpIo1R4w6lnAiyXvcQ7O5b1P/dTD5N3
LAIGR7lEscRxu+8OrSAtyw/4FN4HpLJOGJOWwM2tbInG68StncEZBvxmITfmwlLa
g0F0t8FfjIokzB8UxRum8tY3gm95CPUHTnNKLoZF7sB4dD0nzJ5lsBz4jRdGj51i
63Utue9HJKY9dgD9rcfl44bSuULO/xwq/I7TU785oeh7cHNRrByR/orJUqr3RaBK
H3hZO1k4WAPvNsD+pRLePLKUtTE3Wj6qsWlTO+jDGMxQzvtFS2+fzKh8+Bkx7NE3
s2Xz/4az/r/1GayAyE9kkmCcPkGpsBIPy17TycrPPVA+16m7AXOoTVfxkTyXQkhD
LSMRzSUH6oiLwBZGWmGcz+8Uu/dhkOhgjI1yAcsbB4K4VD8+Bkwnbg4bDdA8G9nQ
yfbi7/f3VXHrFdOkm2uP9dciD6LMuJUBLOKxMPKlVL7GIbsfgMe7XcAKELnnCtch
n10VlxNNtR78QbU63cjz2UgHo9ROTZ9yo1ykIiP0VMVvrvaOF+GAOwB3ofr7blBS
Roh7kWmDESgEFMkLgnAocWRPsT9DqjpDRGqUrxE1Tq8MseJOkQ77caOk5YWuSSfG
oAD41us0pFCXs62AlscqcO4rtLe5gIjqH6u63YN2ocpnrvrd+JNLYpwW9rSwcF1e
JR76pZnj1G/S+UR5mNMBYXi49xB2jmklNwGlPcrxxFeKj6nY+GrCKyvn6Rrbuxfe
kv6c38pCi+1pdeboU0Bopik/t0BW561ZDy3j6SFNJh6ckuhDmgbbVCv8qhbTJ6L7
oXy6zRIiqOn2oEWYvzfnogjs4cX0zsu8C+X6s9FzJuvHreA4vGOm+fBKimKfKKHe
Q6iqVKNIkIp3fqj2W25h5MnP0kXAhazPYhbxKH0+Kwn8YLaAqgEF5eyJqgiNE/Mj
ibJ44oRoaYr36b137tCjpss2NbHBh1WWeJT0Qk4DMAhogTGY/sW2fSlRqsGw6rmd
IjLRexw7JhGDXQL4jxkSET972u9BOSzVn3u1GRrK3qtrrqc1W0Rv5BUNpedRxBEI
JsyMx7N7JwK1/GtZ+OPX6CfA4inPeCeBQM0F60f2y5K2dr++c+p3XV2IhEX3DTwO
WJ5vcVHLG37Ri9VgRxbLrP8LBMWWiIkIh20/e9kRMR5ak/C9Aw3ziCwjoQfWEjoD
UFgw0sPMbXW8YEkSApobDpKSWWGaByO1noFyMrWAllw8/o8+P4yV4Zn6QFkoVq0W
VRAZ4i3hqSy+jYjWW9kOLsKQo+vy/ewoRcGc1Q6DvPhJ9sDwi7X5ZZ+6EQvDxK3g
zhOvgw1lSY65G9FvgQLWE1whPPTlySmelIDE7ezV1L3W28E8at8nBxBGwYiRXXsQ
l6hyZrqKbticMwhnlTkHxaxeRja3+CfDrVZuvLuHMqdRFkZEXvTzteKPqsV6MOCs
DNtm1O5LNLhNXT2nXz38vKVS4S7H4ekA3hTkWsJ0iKXXjWAJSEQWnZV0zF3J9EBK
m57A58SDbGZf0lT/nVvNJh71d4TMOfC1+THOhBfEUIxevnqR6W0piKCnh7Z6y10i
F56+C54dyYIqfPATVGvrngvFha5PH9h7F6+3QOoKB6HupyXJwTa6Bj2Fpuzp0+Wg
VYtXUE5q2Iv9fXxtbO9bI7wmTt1wZK0sKg/y9YlmixrukkHM5B7QNvytl4cS4XJZ
RifY2JZR5SH40flQ7yi3w+wnpO6oimZD1h5QG1oxAAGuSEyNVxdIdEkmtmDV+an8
aYM2UE94D3Lx7t6sZP6IsHYjhd9xKBHCNeqa8AAUJFp/bf9dtkB01y5miboyAwsN
vD3GdjaPxoSz5crf8XKFH5LlXYb4q1+0wIhMPEocfhshFeZ/uPtE0CRm0kHI63/Q
TfIywxO+daV2KYyWuw39IbLyTsbRo2GBH7M984svftM9dXxkIUsVDNDsDuZ77Zy9
WlB81FS+LHl4+7VFkKtHeZkAjnshWh+llzd8ZSrGkT+MYXHQRJDBHw9e7FQyICDs
NqQd9INiaVlbpPitE3ebF7Gqwut3zboDxm/Bk4p8ESLBCPPak0LShxPh6fBGyg3J
7W7ckT157Y4p4Q7CFuVyHRsPmj0fotVqD0T0zfB2lnknF+u5QTl5tozxwNrczaqB
mjD3GwCRHV7MRVokLbHaBSJg0tZBoG8u64sLqBbunAzBclCv1w+8dTl/K4NtMbzt
DXGQJjS68/qmerOQi9Ft+6HGVG9B9QCm4GxM+Rfjg28910dlbaUyv7YIFq/uSyps
pRdo1nYPiKEsngmd9IXR3Tap0c6HVaKHnM8aY5b054pWNIvbjwdPNS7mtF0RozVk
fubtruNNQiV1yQkSU7UMQc5IIw5ZWgdd3N0ebMsRgf+T0KK9Hota7NeBE0FSdOO5
JQVF0M8ze1aFRY5V1pYH4MJYMQW1MralDPah5clypm3PA6Zik1FzjvkQ2k/XFyce
fsUwtuhLKHo0A7LN2BJtXM/9F7fZ3focIZ693Fsp3CD+yhnL3jkxYnHj7zJVb0YG
kxf1culThsjHlpeZmdu7fYufJegTxZd68nqAouXyjJ9I6xWN946DxkhdhzOPNr6I
qKTrIYOCkfXeJytvtmWLJgwGdLWItsH/9dv+VKjGaMMOhlqzbbYiEiib6GhWhKLO
Re66YusTm1M3OxrYbLAtR9AkcvUyOZggZq5ZFqWAkpPH3Gm4cGWzy8qgOwG/UuE+
oyX+EobhusLnkys5KhUMUOQQ92OnSLN7a33zFQWrzTSKHYX+2XgkAx5lAtHjf2yH
OSGOGkqkzHbOFIsMFbgRQRz1D5D4bDMw3u28ej3GBdqVTVXDouYnsGFwhp2aIv66
oArtBqLoG3q2FFs4N7j3o9Ae8rkouXZkFVnBwyeS68LQMx4VG88YicvTHSQmaL3/
zGvPxfANUXSM9sT8U9AFbxvrh6IX649anCDuC3GENJpN2PV1iREXn4aRpD8ypcWv
i8l0wto+K6lHk9JA7+K6T2gB79k8BPOnRyI/5hqH0KjnG68zZuqvqohGl+8lj8mV
R1Sq+aGytqG+yezsMB80N5CuS/i+zNWpqUWQSXpeMDlc5SYwqPEuZhLEPkbc/sEt
Grhzl0aRc+OB0fEpS8Bg3ZAkJk4pyua58ERxr4D2wR8JIOhqANuBy4/jHCnGRlOl
SlCvWfHSD2pGxdP29n3mJUBWZrDmux5vuKhV0DQDLmx+3UCiYEFNQrpgHle+tfKb
TmECIoeTgTqcP2WIMTTzNTaObFOXWPNen7BKW7+MQNmpIn2T4n4sLxgwsDljmDyl
+je87d53d/csSrWYgKQZbWAEwBgowec5fp9LG2HrZnOC/Y/cB/offX1S5d7jMQI7
XXLYUDNetCKBDHIgtjhOQfOv27gTVddT/zEBgW3fBbEhn2U3+NzPZxoFWPVEzVaB
UF+5QKwbVv1L1MvzlCd9Qb9VpfhI2wqTCaP3raYbALLdzj9PDOSCTmGy2Q+Qh1Aq
vmEvOmZEJXqSXZdVjgHVYrDQLTTriYgN2JlytFUJpnbHB/rJ7bwogBnOf8svJm8+
ZP+q172sZwymWSsGuJwyEnDSq2tYDFzQ0UpOQu4D+FmZHt8FzHYSCUbEA/V5INZm
xbCimI5jVsb8kcwWq6KXvw95vib12xp3LyWya3DzaIyR9PK2rQoZsze8XO/h+HUI
j36+eKH/G0ofkac55MGKHq2pLMAYOmOMdK3FYSwNFjtow1q2zZI7pfn/8PhoUkSa
BGcV3q9KTyAvcp18vMmX0NHrbUf3jVU1DNXO8MwvtVwj52HhUVO7ZPe/h58HvTkQ
YzPfXFuZh4DtU2nthmv5Mv2DNYaY/GSXhL3oKjr2hCgL7R/wG0hnm6z6jpEZ/Xwe
nQSznkoOs905EYCTGthEO+Jx9D/T621CFst6a/GzIPLeub8t4ba1bMopqyvDy1Ng
Jg8P0JKPRmWz6Wc4919uHNp+ISafSmErUpR3bG57QBpLxZQOfV+OzZum+uxKNv6v
/q/+ZGUWs3kIfsTezPjjWxqHZm9wTik9nBV2JUf/qCnYbfv4dItfn2fJmKR4W9Yo
QID1BqIYcstPbS5G0YVNmGkuLwHsMTjIrz0aKRSKt1iQWICTNZlwNeTFTV+/CIBR
RPmMgUPVgNVV/t3PUZ3QCZvmQoCqBdsePg6asQD3fAKmQp2Syv4PYR+P9YA2keDS
6It6B6UR5Naen/2TiTvbKbGW33FpsdkWWzsf5RoOI2O2nNIOAOQk3enjx6GAobkn
AIIfZZhhi0jMVcXlseXWZC3JKGnLFZhWHKO5CkIRjr9ovCvClqHb30PinjS2qT1X
HTvalddQnXoEw8aHyoB3ERUbK5ru1czMQCRHA1zLgvNsgAadQZ/ZJ/0RDBi4w+rf
VJbcbhusVP8ZxL7s9OtmOwPERcaiAdtTFF/NSwgj4wWa4s/AR/lXizw3TsWmEq+J
6Bhr3v+R0t47zb64ayDqOzzjtL1GZDkDmzuUnOgDOACY5pIUrTyadnqCCEGY6hN8
zVftaT5nJD2HyfYLULyW/3QsHvY/E5gLzc7RkGE7LU0I8PpZ6xqgzWtVGvxSumxc
kotNbWoBoI55MYnHxZkpvPsLq+TdCtPp+3TpsdPf3XYZcfKZs6b+OTDakd1YL9E1
8Cka7xaSGb9e8KnhGXG/Jz7SJzRmpan6XQY1TSZ+70nH9fclhawULTot3nX+2xmE
9zsIF3cYKUs6n7NQFutaPlhUJpMGgrTyCnlXl2qXUXZpDHmrwIxOaxZFQWYFPvAQ
W5Oj/2sud/omaHY5cSi/saAKb+2X0SK3NsUSTC24SHeb7BHiAvPgKT3yRJVz40fH
L/Ts8r0tABs6fmshW6rGIPKTQ2EqZVPXOSqk30cLTHfVMLNdpfwLTrr0U7KtABZi
O9B9PCmNGonGjR1JVFUgb5xL21QLj03UxVPpmaTPZZDShZV0f6DjuhNGgjB02kqs
7zSsGow9sjLLWCxqazHqkwb/KWJrMz4o9cjNzyNeX5j/UvsQc0CXc+oYxYchurKR
8vl4zq21YVbOdkBzDN0amgfToff27H0UdaG8d9aDd9PtiXYHuCDnI7pfE8NvQ6yy
LDOlrsQGdbU1MLk6Kx3FdlORSkufy+wPI5fYFIA1MDJm6WjDsl2uvKhG6wPIoFte
6xRe7oO832MJRJq+SxTX7LRMUfr5AkRF0vfjjFGUH3J159ocZGb5ePpXDXK8H2Yv
0pfqwFBY+anHbI66bLRuSDk+F71qVPQM+ER0WymVBmz9CnYD95r0snMaVIexUANh
PZqCAGuAYNOIamVT4jgElxp5Dt0LcBcc3hUX3x24J/UwXFdk/4LBY7lFqjSf+Lr4
fO9gATDYFbSkdnwwkYGj0IiCBCi1byuHpST14AYCPQJ2R/p7IE7JxFTw3/F1FX43
gWQDjTmPcguPWZTJeEuXk7NIvWOCZfxhPzI9Xlr5RRxb4h1WU52WYmvoBGrsHcIC
fb1wilttElMrt/3x9YlFpJ3kM95XAFpIks3FxLmr+xikZ1EcRfHVsHcfKTTVrAHf
gAjmbF8XpFCCnNMIy2ZUWxPA6QsKGal31Y0V8kfBTy00RSXZ4flYAFk3ltqTCANe
Ytqeawdy31+OuG8pLOtHkFjXwUq7OjgIgwzaRax3+/W5XeXWqWUHxolSq7se8cTp
3MdCjOQumfQ04XCoC/1LZkS26QPVmRBtFPnPc9/zPGlhg3w1cado1tLGL/L5Ak0w
ElXEF0nXQ0AI+5FbBabqJGDTRS8Lg6zeZbhN/yF/dZw63aF9eN/EOmKnGtnKWCEv
EutTyxr80IHCSlfKfqFWmQ8PVrv9080RSkxvXJ7BNH5lVG/4cF5uGWXLzbljfDGt
BBOSnNQFEBRvGe2Hw/WUX+t4iWvRzwu7r6RTqogh5TNepzRKDb6WVtgO6LkjbXK/
lu49EK7xcGXSqcgyi663wUuVtys5HtU6iqB8fNaGkYaRyNfQLzYpFu6zdBW1ijh7
5s7vz2ZdyY8VeK7B9DdAcVt3AcDXgx42aYjs6TLC4P8x3T55uYodDOVJbtVe+/j2
8mnboHY261SSr6Q03rQXKjFZnNonga3aXYfIO0WeEL6eIMu4NB8c1uuM5IaNgYnW
gtmBFKLbHqocCaZGVe4z4fB4bWI/7N/8YnSi5kh06ZPVg7Nw0d9t3ThYxg6yZjIk
BJFASHufymgaG8y7mv01/d0ILXSuxE7U7T5eWkQUM8OiBkPzHJA3depgsOE6wi/v
nR80aWB0y04CziXU1EqflJs9VFYqhSyjo50OyPMg45SnC+ixvSKRNoftgqdXxtpU
RS2ehVEOnE/Ze8r3BvLpPBPI0rSowKWoG55fd8VnbmBbj2wL0EtV+oeodEDvdM2B
yM7hvkG9gijr7XD5sBEZjCMdVgcsqnDgFOxc4NJKCF34bhTUAI1i5go3kn87nJF6
2vpoJ7dRCKeLl5JG/NcTTKEv7xQtPZUL7T3yvIL9AtJ21HgjQ1ON8sGazE5mJ6s5
htPc5OQJzmInLBcGWzsPtaaomPadRJyngxrXrYAJx8CXddbv9SigxPNp1HHLmm4L
LFGb/9IAGkPogIOiPMubw1QtOMXu5PGLOsxU8GUaM9lY0z6VwcSAOenfWZNI+BaN
1Jjx6jMPvm4mFaw1hBhstpeuCoHEd6KEeMmwk9pqMhMHb6P+NQQjcFoDkdE6Ktwz
lPPuTp2sn8XiZeDgyMa6NSBpgvni7KuQuH61chqAqulPgo2RWsumQCLkyAx1879P
zPohMO7NNF4WciA07rdsLpdnwlXQDXB392lmTXeGejXIy4IVDB8vnhQkgBrIR6Mb
iKwO/A0OEdZDggeWv1J6gF71pOX3BgPFDf/bGkmppLX/PEmn5nhs6h8xfoFUVxNb
ab0Idnlhu9Lla3E4egsGRGdvfCBgL+NqRMNbIW+8tbD51qa1ad5WWjGAMzCbohfp
0xnudpdbGhtF+TmonLUy6bXuEJ1sO+vVJTuxqUfYpXq4R92nM+GYoq9suQkt7Nw2
3CtoYI1+2lb+IvwjMAV8WQcsMXAx90o8WZmRUO5WxNzCOMO4vfXRStwPDdqIMb/o
GYthJY4d5fxYhRgwWaBVzu+S6EKrjBexTu7FlJ4naiDM0UowvMBCwoMHPYTc1Nj1
qNGBMrrxlQMQi86s49XeUte000FUuUKkr6PdzqMmfcYnMEo7bLe/rU8S2I7KDakA
w+DxB/n2uiTTq/laMjuQOi1IRMvIqroqJZRD15LVS20K1/OF4MnCXC07y5pif0VI
i24UTM6PwnRJds6cZXpbFDOuS1XWb0I87/RAjBlCZDW4W0WFapfghyfPkv0YmYiw
DBSbN+6unve1FKpA21Tw1DjPynMrLgnuMImYCZS4ZuzvQURSlmRRg0Zk1D9hsViB
0r4Y/Vvym8Czig2rgL5O8FVo3X1sKihLPy4YpCM0b+MoQHfzocAOOfYcGIk49Ucp
ak1451mdazyd0+Rs9Oj+FGt5tqnGd2SPZ8nU9g8Tn8kojrLX5XciVdeoatPIAUmC
+1J22TgMBRPkVhHFXiCM4TL+EwcN9ZP7wl4q1MROVf7b1wVkZjdb5JGJvcYrquD2
xrFW4ZZH7X1qDHDoJyb8DcrT3mt2LEggplFpjtent7PJ8+Uu88vDjySOTEZtVATB
zfX0L7t/fvvRkSkf/QJPXrbjJuuUNHBYLwmxsV2EVSG9v8CM0Cu8uNLsxoyk2asy
4pCLDOXFpJ+RiIydWVFPJuE/UU3lp9hfRcYbCbe/MwuOutyrrJGb8zQ7kRl6xUcZ
eBo4GKy+9+zUOXz1LWYibXjB+qBFMWvQZmulhnIBDZH6sNfrvec4HRB1xKKGf7A4
WneRYtyl+K2pPa0TtQL+8KiESFVc2lf1fL7ahFsyYt5xPq882H1UE1Zac9oAHCVf
+ZC5BnfCMlyTvCFKgdOJzOpWEE3R42YjDvxcanDvGWr6IRoKKo3D70Y/MR3w/xbp
xQMzkoN2YA2iuPAM/6YxbGYnP3mFZqYGLG8RiMP/amB6e3jzOXiJb2AXmBF2b+wL
0I2jqa7ENOK1MycMIFELRHSpF+M8v80lI3RrKqHl77W4TI1sVPCUaoREyFNpFEEU
2jYHRrSi1XjOrumIN1QX6xJkLNtL/iBqH5B9qqiu2KRLuC/uOwYqre0Tnb4/3hz8
Gq+QUZ6/6TnWDWq2ZFruHweHvT4qNT3FSOKEw3fvMrQZgSnx2xuJS8g86hpDbDDS
ZwfcAVfMxUzZ+h4zsc9mIBsK5Acad7/Nbh8BX40Hz0PJbOKGX8P4wqWyS2h58XJ2
ek4oRMgR0nHnjEbPJeX0f1RETgJ/nX8p6oaku6qNe1acB06If0eiBFdxgdqZNpzQ
xRK1tQFDmJbv1Sk+vGl4Wz9XyonqvCV8DhgQfGV9GKtm7H+6DQsa+yuoGeGTt5kM
+XAe0dxgVAXM/39frdjnNVA2x3QEfvVparlto0JlOGkvopeeSblRef63uI3Q/N3U
Z4hwpezbbPnhAKdCzNfS8T3dWNU5wzA8aJtp0+BdjIfPexb7ihP+jG5oBuHEal5L
UEztjMzBszoHjQppqaEchltjb8GY3o3wlP6kQmj0VD+4GNYCGBZfkwrG2hLEfjGY
n7aT9cFc4ZjHjwPH3rxLuL8s79DBPTDqE9cUleGyF86GNvEwQSXb/ThPJt7XgjiJ
AlW1t2EyISfzjifMMrQbofjsC8V1TOgWAkYwCsrbrGgM1AYB4ppu7GjFbaGlcwA7
hDy0SIiRfpf56U6cqUMrqMP+yoWNZ9fcvOISZHelx50uQxNCbhfXk3UJCGeVjEAK
nSUinJhTQ+DGm2vDpFJF6jIvMAfKxJAgYeohXJQLImG71Yttgo93X8RSQ8C+d6iA
7avpr58qAJqdFvJ2eFsfeOYVI7AkXalYp7/iflOc3WPHMTWxwxmUGOm8o5swAZOP
z4i73IF2HZmukcRNa1N1fEkG2xXLMPYIda/hwRqutAg+0xWtNiOv/zvSSR91lOB1
Awu+qZZm2twhoZ+3JobBAi4xmEX0vnUIt5c5J35B+hOF9w2e3ecm3gl51NZbzErq
ZZx0Vl8swWc7n9nOT8xoFuEdONWSQnIMYP56o6JUGpaY7m+Xgmysup27fVptv8mf
af5vhxMxeNr43dOm7/yU6V9AhNF2w8kjyjznfsrq7AUeamz9crMLE16S+28RWjra
330h6Fxcal7t9EUJ4Ljt6PTOYqb1OvUkIwelgPeqmlGBlwzukId+juoBDDXJ15qa
idTNdmTohz6Msj9xI47K/KvrJ48UHNbKXZt5HjwIEu0JxxEA6pJUNFwijCqy4PM5
/GXhyxeLR/3QW2DbsKcvLmn65BHPnqCT73wt8CdrvkTZ4bhBE95NGz41NkLBeM7q
ZllIRJp5bjs9mnZU4iowvvvmKr3B5yKQPtRLoZ36v9e9UVihv9nKAhb/pYA/DQ40
12JmujYoaTweaRpKqb4iUGI22Q2Kd8l0MTRZRbL4B09JSWpTDFjYZRzPoe1euskF
EMJkP+G5oGZlqTBYYFQU1bsl4B5cHKJKEwR2lUIIGc0kH62YAl7rexWNiFz5Qh0Z
T8fwH8HeYVrrYf7CVvUoBcIpmQOezZOUS/7FGyHOfQbnvV9UgZRJXuTpYPgYJaSR
xfd4DroRl4UEu4LajbuoFq2a/+pYNF0MxX+7LiZBaRSus9DFEGuloz154dUuORrP
Uxdhb7xZnMYtWEPO+iuYKNqRWgN0wEXFCS/ZpmY1bsjL7qxYcYm4w394h9/lhYeR
0DA8bUidsAsgfKi82KnGFmbXImO/cKAl4LGB79fca5e2nNEH/jUZRU2nnTD+Gv2H
Q9DJlrdshf+cUZvdBmZSP46ZMowUecOUDBqrLA5ufw0=
`protect END_PROTECTED
