`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/L/g3s1wUlRDWShJV2whNXTeM9AdVaomOhaMV/0XBh8NWztI48DqtHMlDicDFjyt
gzZlBZkBn9rxWqhe8SyQkaTvQsAgprolDBZa8m3r9x5WYutsFxGqi7LyQ7yvn9Q8
cvh9AJHqfHW0y+iVp/307iQBAsNKFhWti9VGa82/ZYN0TAWdxDmamQ+EpqcD0Yrc
FiYuw4S1wER9VmR4M7TPr/SDzp60QZvDqvRDQsolKRMVTtGaCZKcL1BTmEYDESdc
2L4Ba5xEhWOdnMNsuRuceQz4hqsO8r808DRgr+btGQiTY+m5dNKykUqCXAKvgPwl
lQGVIEVWajAeGjW3gcf9IYL+FHsVnuvZXzcZ5Au51khP25+mggcxmahpYYUAHlrD
cVgBCccMawmOft4QkMVtIWkaC6xwdszhmJmqj7sy55UaddFox4vjMdXvMfGV4guq
eDxoYB87goPJazOM24ArDj91sq7VQOqQqt6c3WyM5uoIvPIp8ehmrJ0DN++z8km+
co2nKdgT5ZOc4rpuLyf532bb0rJ+5Qd9gm9MRZ6ShwGwfNki5F9ane1dgs6egn6L
9OxSkyty9NSPgrJjF59YMeI0hmpk1QxG8sogGBTF8QUXFJZpZSkoBmkOgDPLNWYB
qfnfrqFEJkhNR5Cq1b5Pjc4GUfjO6ofuw2/s6uqLOM3/D3SZf9w0s4IkVDVqxJCw
23ia2goJmUibTHgDqVNRiL8rATZP44sGPzK0cQSEA5gwiUo97l8sVsHi98BDid5a
VGz+WKYDS1wEWvpAkik0x5B6Tq5oz6QBhc+SYjJuB1P5szbxp0KVNwqaBMwUdLav
5JhWVrO9EPJBWOL/+h+tZ18Q6OZ8tVv1JyqnAnxelpAcu4LgtQKofbHmz4wA2s/F
PVaU0uMdWMirB+tmGs47rGOH4K0KxAPc+vatuWvx6KvBVSzIbN4ngND5tza4aZW2
4hpQLhZqwvCRbWFFT+MhsOHGDzP1+2svi5/ZQFLkS0rTvsYt3XM7xm5eWFw2Lu2D
QQriHbeHI4U7sEvP1u+D6bMGYXZww9/9XYG8EJX9THis94euSQkNe6BHs+h/RIpd
AmoeUbZabood5Eig2mXKQJQBhhb0VH5JtJZucEu0r5JSTca0URVAWNDS0vUV8nA5
z5S6d9dMJnZ13OruoFJQsSBplSkW6+voFEnXm9rNItajeZQCWzhqrVzmEbDx6xYe
WRUIKFMh2L540mC5OwSpbbxa+U09QMQWdiT+8uCSaYZLWfG77tZCkwwwBlfFz0+W
/pvq+nrTK0M+BMFPW2kruWcKHQNM8TD9RhhXh9pXs9pJRwhjB1LrQgZ6raIGuWgB
qY2aKKkKU2JoMthDi4q9KOEQCXg0V/BFB9bsQ0prINfvsNoGKMp/l3yzG/BfGr8y
BUZ3kHHYP/ndBNwPeQ73QdHGbZlkOOr/iXZ8zOVIjslRgqDfOIbtAytHWtJivBWk
aLaSKTGnvOfziG0DPR02bD0yUFdH50XX557Mv0SNoZXPIvs/Ezr+Cay+miYRJJ5I
pwNrs/jpo2IkJTzHijibaRrLWKO+fPAtGPqiSQSVd96uBlSgnLTxBOLiQf8CCDlX
3LYYHzGzg7Zy0T6lsySbM26yiASXuneQCDBi768LCP/eITyEJ9OILOQwnknd5o3f
dVc7j7nQKNlR4Ex4YlYO72qcLwI8lfD228AKwGEKkByCQSUj2aTTjKEtVnC2VZ0L
ybGGthSRC0wTjo5NsHB0wXcThoAKXy0a3CtUgOCyUvU3BYhNzzJevgezfmnp70wz
NME8ldnwyX0sZimFpGhV4IesdIfx/Lyj4xByZRXx8qiqnn9n68KJdHpqIsAkuZc0
B6bLOTwqFUMX9wNisy7em9tEfbyVKeUxWg5cpm81GWAYIIqmoZm21p2WTPHu03Zy
wxDsHx4/V3dpEWvdqUfM+mtpNW9pyfJujOgZYgqo1UPHBaUtUqAmR7/0l/YiGdkG
kVC8u0GgewzgEpXYzD/sMnrL0qosL+NnJpKHoMII3+byhjdpPCu4E/SlhJEEjSbp
LK0tTGR8iAVQOauKSzu+m3a1A9uJ8Rjf61SyaMP7BRm9IpOEialLZ8jX/HE34mpU
ulUsRX3cj4OtWThP+HLMBOxk5NiMiTwkB45idJ4L74dcIzOfw8XLAnPkCmNHaGak
Rmv5paLHm9Z1ft8uISNxUydKutxhbo/P2LsnTuI0Lsi7l+LPjl1hZ4K+C0lU+JnJ
WlBw+Sn+fww8bnBfgS/eYLl8DGvMIOqEnNFXPpAUkaqL2RsrtvNq8YGAcyeZ6TUL
xiY3nBXYLdUfTjjdKxk8/k5FCHxMDutDeRUxTSI/TRUDw5Z5PgHzcye/sbZ3JTUk
LpF3zaGoFrchHbvaX1F73diZqMz1u5B8wa5j+mZ4e5uw4Np9n6dRbg7zFZzQvfbD
/guO9fXqkvkm99tv2dC4G6NPKze+bQOCWYmlscAc2Nq1oCEB11+6DHvTylqQT4SW
Mf4ERRy9tcw2z6l9ZDpPvVvvttFW0xXEjIJZ479kJIs8i4hjOZuq/sitDxUZebUs
XgeKKSt/Behi61F8z6/FZMmpTsP1KHmAC0yh3uSJsHv+NIYfYJR6G+Q4OQsjMRVV
RVh8tB85nnLsopyaWC7wMw8yrWFOHU8N57xuIOJBf/w=
`protect END_PROTECTED
