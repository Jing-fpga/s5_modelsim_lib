`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b1S2+kcnbi2cy+aSRaCbP4fsUY0FuF5A3aoDbNYYz4QSP1IBxDUQourBCEpKB4yP
SJfzZG7QK9c2Ml0Z/V9t+kGTZA6NGvMS3o11MITOKYaElnGRptVg4M/7w9jx6Qev
u0VoWr96UA5UO0t4md0J880vsodWkZ4YMIhj9tk7EqoPlYbpRpjRXBk5u0phcQq7
zQzMH+sTlTNXareJxFdoZQ4QURiJjmH7AoFA71HdU1i91TRy3+Md+it2dFdnfRuq
IJdsQN4os/wrlYY629Ej8ZCF2dHr94a1XsKx0IXB135dyotml/nrnT3SteVmnbi+
K5KfLpGYFPORQ4a4H7pzdG7zlXvkubAA2AiX3j/cMvya9T42EDc407zz15WNGa1s
RqWF/YYalx87jbKi5bDHZ3QcHIeXGeDGZVAOdqgH+Bn6hxlKvu9ZJ1LSdALXYEbe
1Tna3HUZ32fqXQQ/Y4Kp3VH5G+6OvqTQFrToM0Hmfn5gnIf3JTo0ltQSjdImlGDs
DL95QOOnLoVZCQaVKhcL2vWJHog1jSp/FChhQ1a24STPiKqjNxNqPExVxSCTITiC
7wUL13mQsGL0HLESOPJWl1EwqrXR3TcHqJYvTYFvQoy5ad1aYbmGeZ7dedXaTWGG
/rAt8gOT/YFZlvqlRFgo86XEgC1YVu+KZR01D7PI/L0kNVhiKWE2b3wbuMC5Sh81
Agv49ZPBKAuixaHhI1IiDyo91e486nENHPYdO/PCQBuJTizlj6Uac1ClfwVNwSnU
0LVmloJzCn8/BGhwvm1tV2Q4bxKZw1yHgzHQPEB0ux8d3TDh6wwSS4gd3xssxIag
REAF83FoWQw2oqbPG2D+ad7yhXDdYkQ08VSTqXvKIykMD0nLtdJ9LAsba/NiBytr
XnjrgphiwQpCdjco/ubdt19HnUkoP/J67+lGGXUm5Q+TjwR1tVUATNYZnx8o+vbR
ZzYdjEenmhf9G4P1P+vNp7muVVlw8sGjtFvgS8/CMdtXmgHWVuBIq5DAbi8u5ttF
ggBL8bbmMIDq5L/VIMQq/C/w2n8BbsuESFRXaZOcv6siEzM5qwlV8oS1Y8YmS9It
x6dDdvXUmMK22QjKqjdnqagjm95YW/D4NOZp/KVWe7k5aV5AZc+u7DhiqhaDKm4+
4DLAgl/YaoHz77hTd3PVcluBljc3/gV2l8LBnuQF1kSld5PA33pGXMxCtjcPEQUQ
TDIGGTJGW/yxp3QZnX5VglJEtDqDz01DuoWIxUy246RwGtQrIG6+dLpQqBFdX3wb
8EychvqhBhgrMTKtliL6iqGoTeH9btqFyBk2o0urZ/i8NIOep6JcJ+zhzR4ftUvS
Js5PHXTem3gitOuFJ19EF4/FbuVb5JXb3SwGFSHh6XlUry0KvKmonK14MlkCJ06u
9RYhcK0f3d4kp25l5h2efqW34pkd5SPvZVcKkybIfyrnahpFM5TkQS+wiEodX7lu
Qykz6Bi5WJVF0J+KsEonoGd74a+NjF5lQtvdhRG4HlRWBF+p0jld23R8h5fgWHpR
`protect END_PROTECTED
