`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LTcOUt91Ys4wh3u5k1b76AwznemVx69BwMjy8+11Tz6PLkE0QLft5MMFnQs5tpfU
ZFETkCPQswg0iiNvnbGAO0JHfhQ74bprQwn7SrxEqIjt8Q1uw9ZrSZ+ZXeMW1V/N
yMSWpCvnQmD0EGUMv9bKMGgEqSnfUVnwJsd2FbXIVNo4rKAo1SY9P6Vhaf37DFWC
ZpdaSReYXKFCw4xxm3Iz5mmmo9mb/D/+Pc5bUurXoq1kjbR+59e8jGRoEO4yU0fa
HEtp2pPH8UqRPNFyRAvNKOQC7R948FLLQ4AAdHrNQGaT/zR4b3xDhOY0wDkUH+j0
k8pSrI18R4DlGNZSzk/D+ADSWnpLdagWDf2nsgvOnAT5vylt/cG5KkHi1EQy3zgW
Wzd98XZAbEMczsqboF1C458Q9z6rXxzxuxdaJ2xN/5Y5BdhDxOL4zn6l+d1sHu7i
DPTwKZpWbpC9IK/xiVHahxHp3x3enFLypCY/lc9yIzpynSeApdNe0e3TZocvwd9x
rUH09U84qSs8lu3MW/d2Am6UVUsfaIkQ61lvTAeNk9+39JN0K+y7J2F5eqTA9m51
dha8x6FlZu4nWq/ZthM/Ng5B4K84RGSfyAEHlnRw3SbHRO1XMhXNneUZW8j9rCuQ
POLQOuO0gx7HlF6C2Smh/k8vXEPgwGBYkSEpIHBExiRU+LYB10L8j8AU2UXx5yRh
13xCuIN5PjMCfm6oNTZh+JvpRHgTx7zOaSjWi8HnT4jeTtXjjNipFIkWcccg9Jec
UtMuOEkifs/ZZL68/uQbjav4NvLPgbwQRenIEoqi5WX0YXJwl8EE0IaVqz2HQjR8
0yoU/ln8F1q2ihXmUANpBEDp6uz9mMR/uLoiG+zg7GRYA/MC6nfIZ+agu6NH2osR
TFBoU+OZNdqlkXJJ3rTC5NSIlrebdwV5PexPkF4Cro14CACPlMAaYISqWe2N5O4v
GFA26jCyM44sO6hZh2+B+4zP2w7CHBKUi2rcenrXgMcUTA3PgfzTLHduzhT+1mAD
iD8X8FQM9EnMgaqoXsCm2V1EofeVgd6880x4Jwu4XHrB4Oo/QuAimH39dsTj0vE5
Ua0OIKI5F3V/B3tiOsWD19RRseKiooLZWunXK47Ff38SrfDXD4atWBsGPvAnKEZ5
5R0tXzFwJghT1huJCrVFNrX9emHO+yHNu4pQ0zfyQB849VA5sMJprFqblvGTlojW
zQq4Gzfw1H6/kqZJxJ03vUwXGH/OuZC7h3NMAJUK/JkYIn8xrcpwGzXafZVtDpvN
ZGrKTGPw7EIKthg3ZSS1/Ix7RRXWjcz0F7UqvnPwrKwV9FsJMCb4wOY2iG43vLVW
Agf5S+NqWwX/2pQ5f0pRq9g2Ci1TVCE+u2Tu9uNKMdmxBb5lrLPoS+HKfe5LtKdU
RZjgRyVCn9/pUfpbycAOo8VU7FFy21Wi5+RT9LbLDS4g7XobLEPqaYLHEMCI+GNo
`protect END_PROTECTED
