`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qNlfT9dAcVk6f1L1rWBw5m6+n6q0Wumnl/789nEprGWMJazpfvxkfimM/SwqWzfW
CYr2qvelzCrCSI0WRcjY1NUBd4nogo5IWySyjFLq/gmSXGVW1x/VushG/xOZUXp1
f8ueG658Qs0Gf9FJzeKCJteLJKnxUnOUgTyL5lp5G7lui0/B0vAPtUhvaW1yA7yJ
e968AkFNdTNEkdcnXNHBlsdg2rTju5wsS9MBXX01IKvlu0wjx8NY7gk/2d+cOEEg
ptmqPn1S1PYiiZ5xyzyEXz5YWURK0mtWXKWShy4pXzA0Pkvha5PRaMxInB4deIqS
S+Q53ATM/tX3i7hNrfOsWuhvKMcYdFhrYFK601b5nZS/TvWuSxSac2sWSpq0TwZD
vxzduSg9TuMOsjrsOokzThWwALxeOLFy0Nk7m9EsyVx/dvZCNvY1VNCMporU6fBl
PMGcnwwPhBwjoQTmlj1iacryhy+5xfrgxwtRE01E3E71V3/Ela4PT19aWs7gKYL4
gy9iUq7W3MppgfVmJ6w+vt49WsUaT3hoX0UYrsZSrVnvla4AqDSYFQMvtpmJEFwd
BE1vKk8vs/R6ShCVWSYcXfWBQZrn3qD6Wq4VBH2cQVs=
`protect END_PROTECTED
