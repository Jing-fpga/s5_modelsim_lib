`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lKu+ZR2kKHE4qpWI7TWEJQwHVethdr0v4n4pXMXYzZzUpMC66bhNXUapILZCs/3s
Fx3Kcv45P1ZPIEytIxqkGksKIEgAE41AjBGudS98cULpwwFV46U6RPOL+R9qxIHQ
yf9PDjP8lXfmuL4cEw8KLJSSJ584ti/Z1pP3LGms0ccRP0touJOt6cjbk0xH+Scr
GVSG54wv7hHiN4jw3lCRXpnhhxM4iCETz0vgBQGAADnTeFx7J/XCV5uEK5MelomV
QVLz1uLGNceiw8KDd7J3+nvZxcWKBH6IV+xLmiPzoHP/pnbCRpJKQPjpLmZs66RQ
WHbxU6jqNfMEtr5/IyLsCdC2LXOBCXra7qplqU/lAXsx3RRht2ze/Zu7eQU8O7V2
IhdU/ycqXFTVuqAukvxGErbvnjcVwtPEdrg5X4/CmaTpvfy+BJxMOkTKNT/cHVjA
dWNyi2lYB611SZXH1xl6WSNgaxiOfAWFy2jkRjf8Foo=
`protect END_PROTECTED
