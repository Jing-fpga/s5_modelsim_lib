`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dPTBkE0hWakX2/Qcc/veRs0wLa4qbeMOhfN0AYvjH2x1wKf4Zd9J5WXewX0ALF5G
/fNyS5FF7yk2RC5n037uPr2OkCyhk5ghXn/c3xpD/WYFk7vIrudSFsSf9PsExSJa
HEbZeinjmDAdieRX1f03h1uqOaeX3WVbBTlX3GuFZnNiIUyou52izWJ6QXrWg4o5
JUWd1C4wvSp9iCbTaDW9X6iZm+vOnRG782NKGiOJ5KeIhMyRCh1mY7OOv/ryUA16
EGyc9EB3t+Q/+KiMf665pO2cd8x331/1igmxYnYsbklNMmx7S3+uGVX+jkjCyHhz
V5G7ftl7nAvuQYzrEPq5kRG44+CBBi4gQMe2mHpp8f5kNjRxUcbtN9e5s7G4CkjV
QPAjhaQuBpe9fCNhPuJCmhGfD/W14GJCrUFHyG7k35S/yo3s7CK3NgWEE+wLSDh2
TsFTRXquLK/Uzd1l0Orwxx7LtDsBKW1hXVa0Od3pUi0Etks/UkcmX5lieTZTKsjt
d1dMni+JgYWL/s1oZO7w3OiUujJI7Uf0+4HdBQRzyXB3Gw5sm/YBXr1nO0zlc5tw
XvZ3wrLvQ/paiVXAjp6yD5ggU9JjKdgLI+F1isAtiiJ0UHXaaT6xm9u+prFJxBSa
dQd2b1daEO+CuImmyKCK+eIomXUxiOA9Mz3EbBU4Jm8gECvT/7UNbltP3LSttkc5
3j3S2vAZ5bYbSf1uAPsMoAsvXCIm1fFV+cTXkQW3TyQDMcOBjVbgJX+wORXZknof
lVFMs5Qwn4DQa05Npa10+ZnGeMCCPOYYkzgNgWZaMWNVRhVlVbw9gp1toamVM7Dp
XQ3wTL8m0NjKUACX3d1oErHjyFq0rVAhbHGevvgtkpt0YFLi/b6wEDAWWhw6HhVm
+tebV/qVPWfgpBs9cZaZf7GN3hbrkNsUWH7LHI/erAkwuQEINPzO/k8yYxm0iC6m
ErXMUkLzdRsOUd2tSz1/9DMTO5G3JV3L3DFAOYBoelaMwwOE4ZsOCbyS4XRLMDCe
obuICEerID5QtTvR4BZ1KiqDWUU7+eGkUKGOCkrg/gREvCvvbzrxA7ZQqCBJRthC
RwvXnkTHrxEw3CwNM8tu7P8XJu4QFKMh0A0dUGMkIiuoCFWiW++gOKSD0/q6ZQXI
Ue2+TnyIQb7O+65eiqLdvP+NmQ+iQM6cKAboPtRPS7TfydOsBorCvEMnd0cNBhgH
UYh7fQXGOK6J9aDHDR1gz07/TRVxHsBTg0AmQiBrPmaCHgw3E1vLpcLo9t3sPSKP
etgYoofhJpkv0V1B0hj+WhtDp7O3NAFwNPnylilLS5Enzx+EnMjxX4ZigeKmsIIU
bcFwEK16X4oPI5PwYdTnK/TkHr9AO0xdPe86RFmYFczeiqlUpsGBVYOdY4YoQTVg
EV4OmTZubTXJV6XDi2BRVPso3gciQGYxVzujjr5OQDEcKzhjWB/wF9/Eo1PG4Abv
myjccupE8lRO9uCEvSJdChhxH1N2Ec3K+7JUMBOOqsQ=
`protect END_PROTECTED
