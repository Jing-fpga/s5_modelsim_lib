`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Tzit4IKNBWvO73ZcabzJyxfPBRd+YbyWJ3lAwMbik3QsRIJao0e2qvpXEV6aRpU
eD4azrZ2TY83zHh8ibzPHEP9p2bN9p2Ri3SIDize6QT71yIHFtis9inyZ24ZXG/n
+DlzHkXmHvSgn2+aHsvpKB2z5GYQCbEmVvEaHzeg7KpwD7vpDMqw0LO4EiDA6/iS
HVHuDStTKFI1sJzyy6I1r+SopL5NyKSBj26qv9i/Yd7idHr8GNWbcYcpqrVVAnVJ
tb86UHSPQ1I4w2J4HfOS6LGTgqe22SLeBsXC6tYtzvhM9bD8OsGzPkcnpIDf1dP/
ot+bxnbTIO31ZiVyB3Oh9Ca2gARNG9tru9Cf64aQsy4nE+U4ENnlHp2N16CwhF1f
hA0RH7ez2f81HP61bricaRvolA+AhVk2+h5Qh5dXkem4DXHRAxT/I9ZeHanhYCEx
ZiCFDn2CfRNfkYBYXz5zU6pjtVvhiN8y8S2fF1AOaMpoCzOEglFk7p9yVnxkEPTj
5sesvlspOpo+1tz+TjbgMXVtXGJsmM4st7iqhQAN/yFhJl4jA3yd0PFEQi1l3Ks/
Lr5u9ajAzP9lUn0K5fh9CMl7d8RxgfmqVG73RFuBc+PsQ1VF+48/fPK9JXSHUROz
ZfNfELyxb5HCfj+Dmwa3JcSvkRfVyHsiQ9JFW0aKZLX9nIGzzcBlT/sXaob/KxLy
xb7HziLcjndrgx6tDYFWj6GiFmhE7r6+L2180JvfTKUAKz4IiUgO3OTB0Oa0r1pk
mxOcT5tjQiR7vw2fXSG/HzDWha5qyS601iv9Z8RtprLgi/oCYQPiXfS4zWGdoK3l
9C++1a9yhyTKea5qOwxH03zYJ315aMgsUC56zy3XgU0wReoA99x27Qt/GOxXaRkB
p/10htaRq+cg4L9cXhUTylfGDGv/Kp3D9/nqzTMlgOQJenMTYd6yXPjxU4rWV5PA
8ZhMjR405rVgyxVG2/2+EPMjcEx4MUFEXGhbIiOZAIRrwb+nL7vbECt/7mg8NnZE
R7GtCutWiImn2Eyf3aFYKCeIhmFt99vrQfi3k1+gQkryDfWL5b9ccqbMUqUb7w3a
IkfYev4Ul9QvciWYTR/q0IIYUopX/XeKBRWUk24jKUlu1dgtUdMQJg5pHdYmgLA2
TU6CnVbnFDBD+LgKmleU5Bxw1+2Fr/I6NVElse1TdYZ7fKovowMXvUYCy1Y0QEIF
gEvPgQiO3jg1ipxvRkuUWCQY3ElI8UAAOqCT6pxvITObQPVs1NKHTlqfemlareqa
ZNRfJGF99hLmKoilfN2fL57YJdjb0CBGBjv0Qeh/VEbMFzePUimHjv0gz+lagM5g
LcVDHuHmxjI0Z55WAAYIg6p2FRnHckcCmVqNOeWJw3Z3iL0MJ2iIyR0d48BF2/pZ
AFZYrho7oHE+qvofcau2/ojeCAkGJIB8HAL+uctPUOJ14xUzu1RVoAKvFLBYrdqh
dmr9bLzoR3ujUDfM1BWnFnTM5itPr5Vm95Fx3KGMFOJClj9eX2CSp2ZeXCaA8aQr
pizN2eNo0fsZBHtllUscQEKN2xzoQZfhF3Gv0hCCPP31LPCLmb9igpPXoI30MpBV
V6upjSCYqxF6MkM5aqP7KjKjulVgMW8J+4K3/vjNUnOPTz99OTOTk+AjbSbHDMHT
0f2yY+NEjEkfAh+YjdgCoWOWKXrCz0NAQr7vF1tD0um8VaRMSYIa9Qy6eghF3Oz7
RkKkRHMQuYGsXtP8D7cXWwlnmcu7masl+R07eshWOBH5VKHO1aI3i7VEKufRvZv6
/zl3JC+CakQZFxU3KmsAYmhCqnct/5SwgcGAp4A7BNfr2SHEYGdf8XzflrPwWyMt
FXQLCJr4iYqVsCBCW0omf5z1WJlhzD/jTtNo7K5dn7A46RBFSD8hLL4Hp2hH6AsD
FIGM+zEf5Flbq8OOJ66AUL9A7AJTJBYKqgLiHU+eOaBWWINa7NPMCSXpLIv09zKf
NPGrw/omhjs0hWAyzoOHZA4ocbrTKfi8UW9e//alAYksUxdLgxZyGTf+LRpTTp/a
FZo5K+ZtfwhcIcvHsD9IVVuw1mnRGo4gUU4UcI+xxWTEq7VJ46NesHVrqsdVDqw8
bcYDn/Cf2FVSrHPlUGu5pIhWhAw3EHgr6pcu/P8+KQweSnrBb2GYcXyh/TrVIAPh
EqFFar/ZT+egS/ChASgBM1nEb91Fn8ZATiZMD5Pcr82yX6Keg79SS96iK1o9BKRR
aDW4ZBFKoOew4sTe9PJ2HH4mVt8botyNLdqakv648EGd2K07E+c38HRG/zIv49gz
dJyjHww+uP8eSG2OTTbwXXAmLCDuOzHr8vD1CAlfbxo8ayTS+RFlUONGMYgAnTiV
fjVJmqZzcP5ZOctqyHlSdEfzu+ab7rpzE04nNa1gIRLFyWQZf+5HMNB68/d/ekV0
QgGLJP/TGFZrUyyLQ+v2UJHfQd4i9GJxW/y0TFRV73P8zdrzRT6VHMTOn8+FuQCf
NyVXGiHqWGn/tHZ12jp7cmSyVIWqzx/NQgAgSeMGSPKdLnJFGAfb8OOlMfSfdmuF
sf6eHD8rTuqi6clFCThtKfFpsxBjuJueJKTPuZqhuKflPFhPMZHD1OZ5UTnel6de
4dggdwB6QyIRskv2OlYzcUpbPuF0Lmwa7ixZ99NksGfPb5sUjPVJEiZV/h9kGRrj
AfolLH/Kz6NmF+wKC7HZfEy5+JBSuUcuvxGr+caowxRENrNviHlUb7XDpUlmguDv
YxrEMRyGI75iyOzqhwfETpxaZaIww+w/oAEmvbzU+9hZ1/cgvjoJejlthK8ial+M
OCm3dkQiGHVK9o2YnqmbphjQ3dPA6PInKaC9628NHfM+I4u/2pFwYaGWRsgvlC2S
AX0gfUOQLNWplIiwd8a1FedPzpjtF8MXbtFF6/xbn4brvyT4V+QTaK8n5BZg+cvi
Jrnk0qhn/SrY5pJnq4fmie5HkAvCrIR/XzIJlaB+3kwkufONyuVGQKunTIyJGZLq
IadLgbptyMIu/p22otTMq6zue4LeguEamZp/y4XY5JI4BlQaYKFDOcIGwQa5ZMSA
XG8AQfDQuoavILQf3VvcbergOY92wjRUWlqZJUePwZWM//TXMuu0D723cFDRag4R
Zm3yiMlTNAvre7TsrM42hm5dSXaZubYxQZf0kZKQ0bAD8dQjiQv2LAE4YSfpt5Iz
jjI/vNlzn+gtyW8dqpj3+sdamsD4S8903uT7VRZiMm36khqFiB+tCauQ+NuFPVEf
h3KqypG5QKSLmBzKiBarlZHlN5QPCJuDGaNq/JNhGckkot9xETTKX2mBlWunYe0J
iaTNffDP7GGW1bRsu4BxUpEugoz3QTBdCEynniGMNckn8o0GpO9Mcp4yvD+e7eSE
CggrpGIceJyMZnWE0zVX97I5uamUYKtyb+j0pztCXAtG62wyIDR6en+COzSV2G2k
TfKWUYMmQOz/88Owz2hrrFIVHjkvHMjFV/IK2Hq83G0orL/05V4r1CyIkwdX3jmT
`protect END_PROTECTED
