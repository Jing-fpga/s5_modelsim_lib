`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y4sJb2aNzq4jQTRanymKa6X5cSszo4aC2y9tikXfi1FMk8RjNAj6GZvhbSQ5J1lf
uTCip56zEsGjH65WR8rpuh8hs5faoGiJOMFWoochBu6QhDnN/RFvVmzZDPYHCLfh
Davd0nmczEC5diCwlDp5PQxJVCZpb4dq2e0hQ6TkyTjdggj1VleKrpB+6BAA7uoR
Yx5jWbbzqwQ5kS9lr/IlFMV14p9Vhxkcdw1mk7KZkz2ugcoyTDbqGfNBp42tjd8i
QSDAm+CrRBR7MlqpXsq9Ba7JUSVI8B5R7WSSCe8evSn/dL/kQLdA/VvMqu4ELYW8
beM3LaBL5pCtR93i4EtJvkrXFPzctTl/WmLSHmnbKL3FxrXs7rIQrFVOsqQlBmCC
PwINnnSFJEdqb/h2R6swz82CEu+FkzxCH2h5pl80pQzleiqGSkSr8X55HzUlPe4m
pub7dHz3cxCkKy8mVNpx/4ZJeT3kCII+6YplE/s7CS6mLwa6Iv60qHqJWSvo0MEr
5dsHJmLWJwqJI1NAAjnMpO5hzoJP5gIeXEC7AGIwUEbmdu6LaWAHhyhZCfaBrHYR
CLPoqlNl1SaaufHIS795ZIP4JgEkMXGxeVwRjrywIEobPgyXH0cuigrk87JwjyQM
cQv5+ESQW48bZj0LZ/fJ6v28RZXCa7W6Y/TXTcgtCl/tgjp+BMuxFS9N/wB2BFnh
NP0BYHCAyv0C2TWmMM/b8P0cb3gJdts35MAPr8RET6mrA1w4zjO1Am7rwDTu3NQN
UIaKgrXRRHXbjHvQ1UjfRwWodxG25QVGi+CD0Vc9bCo48nKDr7+7vxHybRRhYKcY
dZLliuM05lVu05Jl8DQj3QxhZP7QXyexqLHYS25PiyadkAMc0IPDbaxlMaMHCiJ7
G7FQ0AIfXoUx/b+AIxoZJlXZBTFiG+Lccvt0DKYUBnUqiwdUrRx5becehBENt01u
N1D756RZw7xmCTWojmi4uTZ3oFM+l5QqiKpp7DvAUYI/o9WAEmxxm3WJBrTi401D
6EcBJNs8JeEw3ZiJt0mcR/cgIgq+PmUdNyDYsP5hsMozb0Vk/d+RoV4xuG3oT3xi
mCitPX/pjGjlNsQ8/HsMlsVsUoYYX5T9EOFme1eYMF+7ExcNN42cRHhWgNv44gZk
hve16oWRsvy/W5BI/s5Xp4y0GPEdiK/6IE77TI4HNw+1KjW/TKHsi8jsf1krHDCo
jLwhKmRKpvtbL/4i2URg2VFTjBKnza6ZN45iYxO8aGEmjXsbhQ2mVowypjxh07uj
hjw+SeVeqU98rl0Z/KojoORgHaraxo81/6KwMkcdoRqTzeTNNnnWaWYLpxfD7wIv
rGgiEv6eFz0olZb385uKtXw/HXHGEbu533zdUSIayAcJdWFFtBJfxY6TX5efthzM
FuD96y/XtMAVHSGKhtT3Ti1BvZLIb+5wbMQeI0yOXtRnzkbNzx+Yift+PbiM+/jj
VD2Sic5GY8EJORtX0kklM9TPeT6RbEuDuixqgg8BEQS4iHEfscaOX2L31Mc8/+7d
TrJqSPw6GW6dBgTjV5ZRF10oQ2vD8K3pwlo20G0m/3+Ec2B6qLiSBMiMHJGfjexu
JjaeGw2Aze/fs+elKQrJDOX6MmiagjwldNe9VEFAAuKy8xkAIBG4sCwrvwJaNuLl
h0HtntxEWwjhXZwdLQofKjVpBeskAEi2naoVxtogSrWIxGzM5OosM0nBCElOZ1e0
hwQ05KGUsgL7ryh+XF4IDHv8uzOcnk0pV966uPtO9y4maerVB8h7lfRUvumvtWVg
v5FBW6+beBOH2XMSKNkx6OGbzW85Y+z7punYpF8vBxnEFLj4xli3I555OHy2oo0M
7GpwBxkuv0J+yvM+CZsVW4qBP7LpU8u1SkurZTAcyRHbDY5YM9gXIGe8zLwX8jAF
ZB9nxj7hVfqmZ9k2YLkxq+ztItm1RGaHBZDXNkdPhOa8uRM9+rj25HZoRDp5KIgJ
VvjZZn6+r0aXHcH17ttjXZ7hvzLHCMcjOpqb8J+JziGWYRdezCQZqlDPXRyQAsfo
B/K8GPuYogWqHPScMzNLUn0WJtRMLwa41nqBQkmQcR0TEUVZkiHGEz4jHFzZCkaq
e4swtomSrfzz5Gg/ca3/SyMhUXQSxeHXDuhSp7AKMQc90dEisM4JdSc3khaev7jn
RvEMQYR5lWpQVgFVRC+ucQ9uatOgiMB7DtBg4gbElRoeeBdUJJvLoeUsyRdH/afH
La9FVY+mUQnTIJgvWQVR2P1zT08hxZqHaLjX9u4JVVucN8IoQ0u7p74CrJNQpZjT
v5WpO4Y2HtTTUiVmQ8/PxHn7DiAR1x4IcMF+KFRonA+k4BEW2lrFeLZk4BqG+AEc
tQ8PpA9A9QVaMppxiAj0IIqFxEBnJoMJayusKtp72CSbDfNCJ4wFZrEyXIe69YTr
D0iSH+AQQPFSWyC37cFePBQ6S+r58yQtKV6qnX3aiqhkPsoPU/dsMo/95ivGi3xd
t06WN1VwG1msHUOXBfpBtzqJ7i+aS7uuo+9Mnuwig3aQH2FFZPxFrKGGgQHyCfCZ
Y9iTTa3Fe9uZEtgvGB2WprZ2KWbz9BXhNtSy4to66v+dVEErF1QsAkxY2t8G9M8G
FoR42UBcG/UNOE3opQnJag==
`protect END_PROTECTED
