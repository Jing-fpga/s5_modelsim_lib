`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LpG1bnZm1gKNW6dF7P96J79b57OaeQEf6YF1DAK817saukC89CnJWniY58YSVR1s
31pNO2Og5cXkkpJ6Pr5LxEjQVZiPphNYgBTlza5QGaw5WenX3fjOeQwh6HVEece0
SWojoB6HgxCUJu7re0s3jpPKCw+wn+Kk2O+VBE4LSDyyme/igFvqkpq9dm0ksFrU
5+sqI6vFQ5j5wVbPWQipRHOZt60jcLiwZL0/wWHxj34hhwdkDerzE/7663m5SzZQ
DInwWH/JRTx0nV5h8f2RTuUUinVzvv8BR4uy82z9bX0PAWA3CfpnCXcZinRd8XMt
/ExzElbGch+nbcT8XyA/O+Xne2FL/V8eR9wBUyPWHPUfB8hFiXOHp2beOfBvloWV
1cDdL/ucjzMXUsbXR1AlrTHlsowwNyyFcjujXZH2+qb9zKECrnalB/ASwGtklPyg
ZfbJNdGTT7jgVtIaiM7e4QNw8PzM6POh8XBaqxrJ/9JpgKc2Ce2JFLl39DulXTLH
Y7AsRyjPBdL0QR6dYAqqkZvhien5Xgsp4nUI5QWUctxoJAz5D1Pj3WPTX3U4Kt3W
8K53LPr3qwO8rRdxcfyiqqNbeUcxnzhZ3wVeaFL5+DR86K+Z+yKI9/o4E0rW31up
3pm6wMY3VokxSNPLkCGBbL05YhatMfIMVIZda2aDqvbtJzPLNF7u5b51x6By8Sdg
uY0ckFOaI6NE7497tp4w3AH3k3+UD1T8Tz0R4B2FRBXKoCUMmH/SIlcyftoMYyrT
P5NeiZPJFvx8TrU1KMo79DrbvzqtDJ8AZKkNib2o/1Tc6ITXKh4TVxDDm4cuKZ62
0RhYJ9004fxPIxzGrv36IbkA1XfsC9vngyTxjGiykeeUkm5iMU+L7PUUyJBwLa+a
y401sUWiIxx25WLK/ilk/SdmUTVxnoboB1c7TXxkKo4duOcfJELwujtq7RZHL1h+
6iG/UGPl/vUwZ34UH7t/3owGLN+SlR83Xa6hIBM09qJL3tR5lyXzT0QSa5kzyTDU
nPNI8vF46WduNcV4R0BVV7IJ3h05Ic7iH1uvVUOv/g38WpeFiPjbu1rHO1BxEIEw
gLF7Aq+UqFiCXfhDkd/TjuSpMcN3QKbCuE/QBJi/Yr6dKP12qu9Tc52hnrk0k8+7
J/tI5Nnxr/Pz01VBIeVlWHEaUazWQV9c/XcrqNPwReUkIT6ZNuuSpCAe/UGYbNX5
+PKVMj23irrB+74RNitsLqAPS6cBkEbjKzj2wNbTp5TudDiBK6gcGxht0uH7sRZi
Ki5Bb+3N7olfpyhCe+m5eI6LBFIady3ZOFMPU7SySC1FfT1jcOew4DuTQyrwJYI2
KPrhtyM6A5mb+iYd+vrcniDJOcgynH6EnHg70mDO4Oseh6U8oejV90wlB2w/LtoO
noK+eyhvZa3qhMixxNVMWSAhmvPATmUHAtTeM1Sn4HQ82ilufMw6ygQ3BgmhETtN
KIMtf67YMA0LQ3n8j3xgdjEUmI7tkK+9UT3B46keApVUPStIVI1YH/HghT2EKUwQ
yjBGCgyDG7kWTNlG6mF+VZK2CPKwEN0yvonGXmFLAr8uJsXiKDCcGFkD6ONeG2hC
mFSJ4OJ2PX5dfb9yJdUuU/O/JlZE2rP9VseMnvkdkzYxcHYaMvxcULRdoYXuaFx1
kfKLEbO/8tF7UGNT6eZtBUeEX0V+wMZTjN8pdwiSMz/qsK5BtUgM0uvCaW0TfzgI
u0VYrM86Vf5WkncNmioWXPqbyJqy9b2WmUCUcgI8rVIEOa4W4sLOdVkU5SbJ+eHx
mXuLDIqvqzYnDyOacY4o/TTL8FXX8Zf66BkhEre60KWmiovKqkK3dUa0Tia2378n
S/4oSjTD8NSeBKmfKbzst6qmVhDIty7L70FCw1cCgciBgEugsumMIgvd+vvsRk96
+X2pdPyd0dvRHRJM03Z5QFWbTMO+9U1ybQ1/ATg1QMLuRF/0sAG0jkrP6wP2u2i8
DtqdM92tIvgOPMpNsJgZLYx6f+ND9HHKisNqFmqyGCX6FUGNN5eZJjL+wFTwvYil
37OZdhkpTec35vCuDbzLl/lC+J2FJCHFJwbIp++jvjCz0EX+J6S1AZchvsJV/jFE
3uJWHBiWvbUQ7XZXTqskwWPxPfM5zjydXweGuVi0eNrFPSUFivXsCuhazvgyje5m
7z2R/eDgcrLXLNdE0SiwA7votOq3mltT3u+26PW3e+nfZhAkTQ6WNrFaRwDpBqkX
IKrVV/qoHn1K9eE5pJJBEI6YXMoeg8aV3gxG2GoTHSHr5si+qZqayVDdV6I02bg5
UOKe7iRyjAVS9vD4bxWvPqP3u71sYee6mBzmmtRkMAmXcFOZwf1vUKSRcCc/aSGc
/Ut5vk7zULJLC783nVBw7SKG1HrC5oblUSY2/sxOSgHytq/Kb4LPDXqZvDTRrVTK
VlG9HTPZglXCMWXBZ4TqzBvRsY3mE3yoiPIRHhEf4+fPfXbedBjVOr1YUDU/rwNF
mvLldTfjymUd6yPIp3FoxP7rkxhJTQsHs64+wyE/op/RzgCCWMComx5XcmZ0vzhb
`protect END_PROTECTED
