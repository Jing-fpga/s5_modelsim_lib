`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
41driJXqDfbQtO6lawUNR5VEadxLDHSxpBg30/GsPiE5QrlUcz0SNzvJOshGiqZI
7/UuVgQNH1dHtwE9INxekdxFQK2yZy+gLZDp2EtMqZ+NDiZDNBwj8wGJ21j+ZILk
O9i1R3idE+EXo85gjv5rlg9678BjO6js2Xk05NP4zlphv3/zy1T8UXX2fS8hBoyp
MEAp1fktO4G5Lje1k2MT5boJ24DfOK7ySFCKjfVn5LcILUMVyqdMIjJkCYxH0ecA
THG9cHcUDCDES/BDEaAlns4Z5/x0OeBWYV1G0dSkf19AylCAvpveHKnP/rx4AbgX
MB9DuoGfXy3h2PUgaJNwMXWuQOiATByWWZGo+OXZyV3/O1YWSjY03ewgzF7RVIlI
9F1385uE5Oy8DpNF/hdHngVwrHa2/4vGHL+oPhvA1u7ig9GD1zYYbdipWm/Y0NsY
3uadP0t8UdUg9jjyny8Ygpzsn+GFblj++3KvVwtauB8A71vZ+HgyjmwIDvogNx1M
jSqrBshn4CmGGZjpamgcY/ydiaHP1t29yTwzxZHoPZdpqxzHOxnvdC9QbmkG7R9E
A3CDXjFtxBQG5bltnTyRhXKV8u+HwgD7SPeTjaE8MR904aKR4wejFunZERzpF9Yj
11BhIMz1ThEKQrmp+PXmY2QIbX9jCjOI5qxfziCAwp8R+NXE6PMXpRRUCYT5v1K7
auqVdtNQJ0jaw6Gqmb2rkXjo5oiubA58Lx1KmreM2vt4GYYr2yRdMvoovfvugG0X
/x2pPAP5Dfk4AfYu+ko90bDErWRIgSClL0/TLDqfXpRCxiLAfUnjLfCv8mxqMbUu
Z737jmHjJUmY23hVccnpya5+le/NdgQ9EWU7zoLiv11TQYhBaj7MKkoPmv/oXRf1
GX7epKNQ3sXo8gCQDKqv1cuKpyzQizxsMnlrKhSYbrmx134opyw3vkbEHP4dIHOR
GB9Cv7KGqk7ONAwyeKft6EHTKV/bXNW2AXJc7Uyg25I3M0cCysYGjaCSjLNNm71A
ma7ZnNXr5hood8zTTWYy9LJvulISDuOJVgbl0Heu7NNhyy/RqOSrYdR743YGLR5a
S5Eyp4qoMuNBqx5DSkFpGSWtu9mkActri5OLZoebm9vGNGFLCP8v44yCls2Sy7KQ
3UcfNoBXetjVXK3nUAK/CVX+5yeXKIZM1Y50RbwZ+eKBOSP4UuuDrPIB3CiN1/iS
UxgyQNwNHfv6Ub/67feiVMfQSPfPS7pOxLghAlDbr7wC68FagwnusytcMeJjSLtG
ai+bZ5aQNdvaDWF2AJ4ES8n40W5qtjeCgq2gYn2BXycmgKxr+tajeGMfQFGeQDt3
2snuEZtoEfJZgGyvEpSi17ZNicZ1CCf2sIavpD9epJJH1saavyHeuy+c9pwAjCmj
NrDy1CPCuI6CFH0MoY/jtPrXd7SCCTFEWby8EHHvtoJOfhDj8CfaIy9pJfO2jIGM
2sIz7sC8AIQLrwvv7pbh/cuVFgJ53HYJshOt8MhWCMon7lnsnmMQbV4q3SGKIx+Q
LjzviXQaKSlETv/eyYTlzJj8Fg9GVK12h+pO/gGG4mZdrJWQdjIt4v232+Tz+bZz
aVTfVbvpxh12Szf8vooZ2asmqV8L3rLBGpA2j6njU7MffVZMZp0eXDtC4W7naiHp
elInImg7/0n5exDeU5fxDRvbtetE70KKzIt8IA2qqcyRzJIGpGO2GTZxYV9zsxq6
goslB0GbKvZ1TFsnEZM6Rf6R43pWH8PN+P5M6DAHbT2j3Im5RnOoeIywRq5PRjWR
SVn2L5R2Qr2Wp3uYGoLWc/PxkydPVbQb4oGA4I62xdhE9QQwChI6ihporAU/0gBs
OVoEhc91QAo8Dpw+PGrO1OxDIUI+ShdqcvJ/jcCNFJ811KS9nDIEtfxRN8XIfLE5
vejGicQahPEoWYDWQXXPy9ow4PyHNGTFYZ8VsXh1Xw9rOFzVmSO76KjOXdVT++P5
61Amlsc4TnZSqji4kR8sBTOhUQXwEkBuS3bdDbm9c6tjRVXymKJpDfeb1CYql8xg
OOtw8S/oNmOhvv8G5VHP4/VeCOsZj8P9WbMkB92ynTO52TlDRPhT+f1EG8BO6xOS
DO/Tn8rIpj756fqAMhEc1WaJ55+ucvZag8yOwCmZGFoODCawhgFuHs/dTrC+x8qZ
P5K6aoRDg9YmakYTENIO8r3YR97/RlH4WEdW8aSQ8zd/HRvrCLT5vXXWAXl4Ez1Z
guiAPC7ghBKnPhb4waT79tG2QwqLSuBUIYvwAc1pBK2TTzaNrUytnmcxNegooG04
XZO4No2U7mhI8GhH8GjvXl2kp0dhXC1QWLh3BgvwNFayYWTK+U9IIR1Vdm+0HCVe
msY98xTN4iejfICykyTYOnPwEBkaWGFhQq3zKEBB2bfKf40a3Rv08xtWA/DmNZjK
L7G8ikxr9BH5g2rugzTL04c0d4EHphp7JU/kV5GPevUi+j9eUwEvxAO/aXEwQzy5
FXuY9Iwf7puKAPs0GEOEukfro+ncuGtIqZ2llR1GLWJUM5WGK/6T0caw6fMV3vxV
/+184v1mo/tfAqLo1oQrUMXXBbM6JvhTL+oaF0nlPKo+FKN6zhDtWD0HIEX98Fzy
nx8vvLYFV7alp2aqsMcc92b4i3uSXcs/dCEjZG/Y4J7ML7FRcosAc4PtRx1SjQlA
TwatXK59Akk05UsRPNuBPlqe1YzRQOvCeyRa9XURRbU9I7D8HnGVMGy9CvZtOxtu
xJqEWRfL5ftdc7TORGFBrTBkw87JFA768NlZCLzzGo+8VTN/x/Q8dm5oBOolCBI/
8i4eqt0hTKyjVVEtf4I/GvU2NhykVSYmO9KX64UXVo2a9UMIPG+X3fj8Sfr1HfE3
/E7WaikLwWn+AaceooDo8/9uQSeSFp+xd9A+8Roi0PFD+1j6CLgbvlbY853SjGSk
vdiO1InFecJm4BVYs4ErBAK9p9Y1uyqWXEo56ZDOzqeOCowvSytJ7m79EUXiZWrr
snd+/J2J0VoZk/+k89uk1mfZEdGhHp1tEcBRZykcIxdcB7ucyU2E9zKNSr9LfCFb
SuPl8kv6jib5N81Y+jvc+a8GQex4ipy/PJXnCXEgwyOVHvbgwzZcJcwqwOl9aItd
h1QEU8ZHjIuz2ubGou6igkilpwfO9f1H4FEBdyOBGHNJfZ7Hs5j845d8sM1QwJx0
T3AN+t6korrNKhOUYkNlEfCYBRgJt93WevnAHGrpKxlRA9ClYcz5tQ7ZYF7gjGnR
xd4SjbHhP1yC6TBZ9/docKF88dhbtWSQOrNdU7yiZHQAdaHm4u9hsHM9mNbbw29f
qRpHYTiBQ9Ks5KDC0LUrJB87WI3Au8LdPKOMtXGgP+/j56mEXqzrKmdxhrp6vs69
SqelerzaHRWq0jcz54gbG1WWc8uCrucR0tBYcZzszKCQx9iZ1CQMdtStYwpBay8N
OGZbOvjJEMm7UDXoklOrcd/+8POV+KjBzO45/fFz76FoxznXWa3Q//YCKUe7zpRB
2cBgTD5nEMV5bLk4t+v9CdvcZ959GXMTa+NJcwJEGmRYcDQ4/MkmLQTjz5597jMH
W8PdOrhwXjLJoAlkYobDjDtuUN0ZHFwkbalmKMWfmCvtW0HaP8ZG5KyUaoE0bSYA
nXFU5fffic1Ei8tWIBOS3R9Wsv7+5iJClSMFdI+tivrjLWVaHX5B9zz5gI7wm0Lf
Fv7Xk3/bU285oXr+we/ZDxQ1aK7NKizIbFdq1jaYZwA5miW/CIgpcRQa6S4+/2Fo
Zg+kmNfdHcOINkXiKtvvTs0DFcIZciJh3561k+j9l1HGRf2+i1ENU+WmwnssAYQH
TPm7JaTjVr+H3zWIny1AwisSurqml4ENtIRpmDFFSoryZQFWQR92MBMMq4xFSCfS
yJfomcFQ3OectM9n7IYfr97ZZjh2g1eETX7Bx9Zjk/ZWeljJvkTdHlQcVsQjGV8k
8bg6ucAMfd6WnqM/bgxhrOTeFWmct7gSz1EppgAqwwnZa8J6ulbomnlVTP4zXONq
z+9V4nkftvCgd+Dw0kt70g99FgtOyineNAwSihPAELDF25vYkKZjF+fnJr4JD4U2
y7+EF7/HGiTzCtv607EJ+Ov/vPIwrNpv0Z/sBoxrmEn2csIk1gR2RVK7diCghVn/
bzM4jISBKtPiJCE8PNl2t5plqt9+ikx/r7DsPFm/d9GC9VqSXGJ4yMOeQo4Rs5ud
86Qvl18ZYCoNglsHkZ6caKMe7SxJ8eyiHekepiYr/Qpp9ckciRTKND+e3QTroinD
XmjZuFSYMU+voeMPmwuyqE7ych6DjfbsQqe9uyDEKrMIWoFzSLNhxxwXwils9pnR
f5umlVIf7/DohJf04X+12LL5atJZ06m2V+qrdd6ofCFzGDsRXMMmKP60KMeI3MTL
X8cyu0945cmFFtQxwXsNzq20+RvCmuEQ5+GUq3ElomaAP5ispxBHGzeXmN6pkevB
RUuv/7d5O+t2NZu1uXWvgF6cLEZhYH1fsKRroaXuOEeyUQxa5iDy6ehnrNyzDaJa
wkkErJzRj1jIovczPlySqBM6WMLsL9uFh+5GQ4LaRn9JK6groGLfs6FFNv5+D4Kt
+rAAg3rVL455C511nE6RY7Hu05H/nVrIhlEgrqLdSaNI7blrJpz8uPZSe75sf6xa
shY2I0m/hu9fcPU0qfeTsq2tHWYwDmtHtfISatob913eYRgPebnmp3t9ixNxuayl
8eVA8ReriaI14yBoToou0eX0PW4b4zn0yIJokVWabR9z2kbnt3fQ6nW62O3VV/LP
ryjhAPlFwLIEkORD+rCdsgXr7hc+x4si9Mimu+vGe9n26xEPu21VARbK2atR4gId
aWMlzGyHAW0VyCSVdrAd4BqaSz38fN7KdjfsUXSH3K5hkpCD+8DEAUv7/Lz3pPmC
SivBgcb8v4g/1gFP6XAx1XCTBVh0aZc3jaPKjVzK57PPycdbqlAGMhRfaqWc1QFB
z0XHtCHYgF3JLShu4cZkDb9muVLYXJaLRZus6iSgDhE5KON9G2QicBY0o93cqGlh
cp7lHhd629K/EbqFLNyPq3j3hyokbLzFqqh0FnzbdH7RCRVXgY1LnjBd9yZgMyCp
zkzCo5J3y4Dd7TXhJylkNwVxewmvzRXGwx7gqmgQ0A1AahHgXKPdZIxQGmsiSwzH
+/nkdF2BucD+60d9B7MGFdRNEUcNxFOs3Zn5gzKB4MOdWdf5qd8a28E6SsG6MFeA
N5KhwSgRFmxGnmkHOH1nvcJr6+rCSpL2RpmooNy6CtDkQv/q1V0l9plhN2v6B/lf
eJo7tbCFKok0WOI2SNF2jsUIjtQNNG2FoWDlyYbTjAF//ympqyzY7tGHGsVkeoV3
E9IasEvjuNEybry+OSWhyr5C3ehAHBrvq6dpNNygyb8BZCDAD7IaWALH7+CuaFjV
zechPcEPcqx35F9+U7iJ7Z4ke0crIGMmp1G5i4hC9CeqGO5waYGRG4ol2Rqk7ywm
ys1L2QFvgd8xlEytxu8IHvTLncOgeuTlAibia7p2Kv+KTBVLvaaZs9DFGB1S6zLC
tKUMmHNT2+Nxxlj2me4Jyz8pQJ7pQA0UCEPR04C6WVCZVBho9IRO8eOdFhpLP5Cf
vfBR5dG0gJAR5vWD+SbFz6uMo6+cUMtDEEhjZZ63UNO3XqHtMzzOO+fp+MDZ+Ayt
ugxd2x3Kg9TY1SV0mBZeDj2+nTHnBTggEtVMEEJ3G3Oq6fNg8RnryZ9iRY0nxlUZ
yjOTgmp3DC8utS91lI0PwmMdngHQ3x18U3b3iZpqXKxfprQa5oMcWq/xl0uFYx7B
ly2Y5d8LJcgxhaNwjQ7eM7fE0T3USguS5QIlFu8LcAAJ/9+ZLeMtCsDvrc2HOms2
bRc89euLKWmZhUHEi8tcXO/Nnk6vTeLnLK51YiT6hgZVx/4ZpS6a4+19+9enCy0o
2gBblK0EJF6DO57OY+wzWnvgvqpjf0q1sOf0q8gpEwfYq4H98/FUHm1KmN7ZSGEx
sYDObBaHeQZmGbWQ3egwVGfVRennPiQHh38mGr6Qt287HIv1CksJACJ2yWhi2nNw
u5cJ15r5ZIbCeOeYsHxHG1WgYsyOQ57h/CUQ1JKm5Ue6wFVv/73FLNjZrUYkZMuf
jvRKIGs2I9rIZun+x70ef8j0pStP2ZZ1187IM7wHLjdEZJrmTHIY5hOyAHWIrlXe
PbmlH44M0KPDNIWj7xbeRkNqERBrrdr7BuGRCUivcd5VCZ/UB8V5Yd/tFrPlSbwa
qWsAMbWIivKyBCnR74mJ9D9IoJ0+VWyJ4pSNaqF12XmR4IoEPZu+scIeCjBw1rBS
csKMj5zx2bvyLF2mQT3aZ2PhpJap7hmJYOSkDn6OO825Sj4L2YCkawGLFCO3zb7H
Q1JZQMWqySCfGgjeyzLuirIpGZcg8vdPlKXVVFfmEHTzjlnH74rRfHNotExvnXns
AvT9j4aUlrHCDh2B2z43L/mjkXJ6noxtLtS2hLfDJh2Hh2tguPU/sOjxCQFQ3Ue0
oZRYqHAzsKG6PqRAaxqJAfRquYq7AXt1A+aY/ySioACfEJ/tQOec77sY3Ti6UFVA
0WcXVoRiCB8zzVTsx0aXRmvsNPNorXPJeugNTA9oVyX6fmrqaGiXWOdM7Fe4Nus8
cp+1SJiMyl3gEYnkiI2SG8yzTnJS7K7fOJyftq3GR8odFFer2ZNxr4mgRDvGL3nM
ezwnXNjfOGGHCU31gIQeWwETE/xrDcQ4yA0tCnD/9Z76uGB3YX1UUZwYBvF4yj+l
lyu0x2Rwa4IYYqYQwqHLKWBsX7B32fIW1cpW7HZ3aNPCAhtLiDObVyJT5fL0vVhM
0dvMhAk0Mm6p2qZ+PMtkbhqhXLNcUoq6e93vW8UJxeicJ1s5VZJVUpVz50OgqDpc
gqjmiGsRhj1fmYClA7ZElVFHvjYzND4aswgaBcDh5Ay8hxXhu5ksFIZRfPzJA+q6
gbLAQ4Z2u+GkeGZ5JKnOzs+0hDfb6D1cl2/ztQl9ticrWLMVJGV09ao+uzuu2whz
ErQquPDDDXTltaCtUFq/9wS0ZcRdlUdsA3rfNmtrFmTN/Ht4L8F9U06nd16QFZvr
DXILEoDoIhn1dOsY7iP2JLGBd9O30GGBd3eiWEF7+I+89dGW+ChqXLEKsbvfBttS
webNNYF9+TLWk/ipExBfYW/ejKX3vTyzpt5FOpq3dRype2G8VXxXb2Xz55Qq70qS
zU2plRirqQBtvhJM+bPRdcSmd9mnaq/3CT4QiAgn9gSm5LnQvYVlXggR4evw13GX
J0TO0HaTxX1EldsyzHLUfmM7uBaaoPKN2ZYtdwHIDN6EqOKA2V183P91djrWDo5x
Ph4w6wKDrE7D62LuTnoW+1LiSgz/bWGKEN8noRbctLVSYx8+L8V6PT5M0vF3tMue
92oi9MVPBshYK/4JfxdfKCkxplqiKEVHa6eGeAAodLr8xmgbZa9Xj7RTVL0dlT15
PZWGarytQevkDHc6KP+n1cPXn/ytVfSFDic7miP6HU8h+/NAG0xTgVAWzhmIosBu
DvjAwLDwS7gDqsATcG0lHXtZfvxo8kYtk3IpQJPe7KEHr06B0S/A2Psky46t3eRD
qOvZlUA/lPwIpI1PLQf5NhmYg2ya1uSlw2OPcpskAJ1W0G9ZxRr2CwFPQgaO7y4P
tMOfnaifoXgYO8N2R/SNjwbbW6ElvlOTYPabSe6Nfb4frkLPnK4C7XDKpkQ2L/y+
uHj1Nh694YV9wsWQhvXg88bkSrnN3Kbui/Hl+LVb7p/laHKnTvjPj7neTg1oBk78
w06cP2nndSTrPI1Wj+lFjR5dZ/lenFO3rTlsZB5j6cnXo71vq8UKzkC/UQCe9tvj
uIKoHscUonQCLIivDPoTHCVAjX4O9xiM4Z75LoEj+JADywyVl/9fBrLb2WTwc3oN
frrI2FC0AgudO1zYeE5LydweM6qg9pLv0+DlyfVScSPMYhoI/4QQNlBHbbGjGt/K
A6BZiuQMvtSTI1nPjFItL44kAvksyncQzmvED2Sw0wYNVvIduwIplWXPkN1/kUWi
e3ozYhEnklFhckkcm4k5YcfTJi0/XmxK5aTbmu9ChQJ1b27joOWY9qqwEtM9cX9M
JH6F+QV6lT849TUN2QpCwa1hCJCtsuS5ZhLGsxj7b0Ip4OaVgPbRYsdUY7D2rxqa
FaY3CI2b9dlfxE5TyhbSTDR84YfKZlp0bC7MVLHNml6XndBxOBG+FW8Ofldj5BqP
1iaskMnjgurt1wITfDSKsGT9+fqWnfjSEiM2qEHrowh0GQFe+8yCO+mtOx9kLs2q
lye27g2A1xWOBti1S0f8qRecU5yOeL5IMS+0XBTkMYyMC4zw5+sZEFlxJ8R4yiyr
JArhXD7HLr0Yy/pctqrp/k/vpEDxW/74ONtWS8sQ0wevEY0ERoWaGqFu2aHzaLHx
nqVOBRigHfdiAJZjYVeBytJjyYvlI1VC4clgsfmPzMf5lEB3Aup9Jrooa7WE76Jl
zY0AcKrvngJuNIikMai4lcxWwGiCNtFX5IQBYMgR0HzTmoaIB5r4DxWktMr4Ex+u
F6MEmTyndzoXnqBFkHglxFy46tul8A21xPorEaNX0dniaYThqXKm0BvWIvOCTsZE
6U34viWrb2Sqgz/0iQqVDKUDZCClr66G27sWkRRp+7zFZ2LkEG1hcruY2l9vMTQU
AT+ge9rmSO+1ZF2F8JY0HKenYQwsXSBYk4jdqmKwHZLozCfTsVB6L7t0VRqxo5Px
UCBfoWX8BgKZYfoHdtEgEkiPGlCh+Y2nY5U3h+WjvtSfpbQfoJTT1Nj2sYkaStsC
7YrQO0oOUP/KC1qFSqD2XM0btuINDjsrtY2weuQj6+yp8LL03APxVrvOBppkpfTN
aWo/sM2bPRnxgZoj4c6us5N6pzVBp03jSp1AvDS21I0Zh47o6AIIOBE9AYGYg6/Z
5pQnODS1RYri+kskwv01wvK9wjdUldxXthJo6NMYz/kgnKDGDMjgolGmymZzMv81
XvpeSen2Td0ibXk4jBKuew5QfrWbio0K8hWDX39YDSPiSjy6t79R2oENxR2AEXd6
ydCW2WqBHQ0Was4dcMX/ftpHxD6Z3A5P4flYe9fYVzKMCOqUpH014H7fn2LwJV0Q
dJ6wqrhwVOIYCJw8CaI0bvnv/YO+WTu0rh4NzECUoOYQgkjE+BTA6+FCMuX2yPZX
9cO3VkQwuvEOzo/j4wFnvlr+oVY11CnUxp08UpjwYvih5OvvvVbgGLJoORx9Z9VX
7bbh2wHxl8h9uoZVMBU2LR2GN36OjmGPx7K4OonKvUMFhwr6D2y67DhhoTJ5C/Oy
q2SYs/65RrexdU8aAsAgDvpPaS3T71dxwUWSKvw5R4rg0sIshBrNavBjH4l3l532
t+0XqG5BTl8JUf5zWi+AOW5j4Ld/IcbsvoPZJVaazXjK1xaDz7AoHg1ET7eSil8G
NaNj5KKWuDpnV5OKsm9LeIstmGHWBBGU/7AvaJn6mrjx6JZzQntKitsl3FT1l3xG
tZnNqQ76KW4+x1n300HC/oDUmXPiExt1LhQcIXWdO6fa5sRMFf/oQSfKnSA2ZUff
rZzTqjCykezQZFeSmrYeX7NtbRy0zN7xk1Of+CdncgBqMEH1/JSNBjuI/fbh9vAj
WiwjIA/iPZe3pdmGyjxwptLaTYECBOnE+oEKieSvmuMI7/IGCKbol/Gx99mMX18M
N85nf176QhIoZRzPtXsfIuaIpeeCIYAed8p2y60lWwfgWh/xFvguWPjZkJm66PN2
CncTZ9b6/j9KipRaJam7q+SVC3CQBIFcz0v4CsF2vo/N4I+YK+WybvLb8x5K0Aj3
j4flipPQj0Wzs6wNhYbdnmNMlKbQE3FlzcNhx/v9/nn3mj1RhRCx9VMQ7HCeFvty
jGBcPDbQnesn3ATbRzrtQuBuwr/2xBIE0rhIt7EWZR8zrHbwMK+zo2dhV3J6ylTQ
Z1ZYwfsexj9b/czwDcPB3HoGDGw0J7nz0pJgBKkRhnk/H/0TDUP1XWMI6QLXJznc
IyznPyOMq9CBybTDTlrvY+YQgPaRiBZI1geKXbfRXhX60NMclLZI/mWvU1ovTUNN
UFafWuvqSnkbRXt2A0XsyTfFogUNnLg15tjXIi85UTQ1SVCAAtiwOvIfnM/s9uZj
9ANou/q4npHAlhRr6cbozYtvElr+nGfltWZvRv8JsD9pW5Q9o98zL+Y4/v/V9zDH
Me7ffNa1EWGNi8i/0b/DxyUnrx2DdLkT6BygbjZeBOuBhkZBf7nxiIGWxT0ft2Gl
KQswKRKKPixTjrKhWyhhg1RaICA+873ysvbd7EojbmQNTtGNqCMFZ+ITitMYxUQG
bI1KNzCCY6bGQV6nrd3m4lUvXthXnRHAWcw6wQINff2HMnG+2hsoqvFcpZp5AfEF
69j928SBCKI5h7N+RpGzwEespJaXhNOGlgsKKDfeKfBuIwVLs74WQPhhnfJnE+sI
YlWWQIhX5okxffEYTe2Ab6VqrxxkkspRkGhYdYX2YYeAy7E8FyA2YeW4EYZyrDjy
jxyWQtnRkYNtyI66p+LOAKCltFadV2nvt39TroS1XmBcKBPs+ytOxGz75anrFOBF
9JYQJWWM/Xlcj5GuKUG1eFQQkHUiO/+Jii6AD3LmKQ0ikqRpZXAkNHrk1FreZiJ1
cWjWwYE2zbz12SFoHPBtm7AxoriBxq24GDRgAX9cLXkaQqg2pQvoz39IpvSNBKVN
rvvRQQaaqZthgJp8j+Ql9DUmXs2e0vse1iEwnessZidak0cR2XoRLagclx47imp2
uMyizmf4AmgIcZUSyuUL2Q98va5LD06Rl6/42GrWEDXXjx004S2qvko/le81xdVb
823Us6TEftvlyp7qX5qJMRd7jfKRMU7K6rXZw4Hk6iJyWS6X1XRmwl3S8ki3cOX7
G0fAlVz9xKGLLSyyd8cyLTXbrPoabfRliYjT2472C4Z3E7Gyo3J1F+4jyx1K+YKf
lhM1qXH7qTS+RZ7OvZyk4e3Eu9La9VMQcSK+3vnHDoU95La44zJ22IdLGf54ERH2
yTTVUjrtGHaWbPhrFN76YRgR0z45XoqQf8pMu3QQWQWXs0srWViSYaBVjj68IS/9
99D3m/fJzOEmzouT4huXNxy8VydDgusbhe6a4FEazH93K3gLuLqNwLxmPyi5RIGN
J5T6N8lGbm3uEROExwZ/50wVkFyJ9NYt6WX+FMbaoiqGWpEhIbFA5hnLDyEKSduI
ksGMv7AmqEN403jof9jFJtLGQH6Mthp6X4TNrA2DcOG40EHjqrHfpBXRpq43RYtw
Hdav7trDKOEt4t6z0Y/ADTNt018XdujdtFH7/Gj64IhbFFnK6udgPjPAOeHlprGV
cN4CcQ7scZ/dNizznWULTHXkIbVtNAOh918qA0nVHdCE2UFe6isVV3yeI7NbqBKg
RYu8dECa7ryRK/I6fPzCBGDgh9AFF98Y/U5Xhy3Y4aRbQkoC7e7BIGu4iIfgIS8n
/sGSdt8G9HHxgfHaL5Uc3WAXoMqcexTY9PTReffLRfGCg5QDN1iHpKQUWxyig+t7
8RuS0U6yZpmVYf0xbbwaIf2rTExA0ht9oNXNxaqHFTRv5EolSHWvPrR2XJV8HuzZ
V44F1Rl3Kb7mXUMxtyL2fRn7KGl36YfhUFh9nHd2F/pkdRnxgBMih3PdiD7tKSWa
BPGv8ufhRrGg/mEB/VYwH/jMn7P1OVlc7JxTjQ6cjyfnf3ob7QzNM1A3YbdKtwj6
Iw16wuAvh7vaW5rKFM5XpW2u8tecs8p5a8+Akb2mwkq7wzZ6+5rtEmXrqNGDH7I2
DXSZRwQsBHU1hQX84T4DAs3cPsbtITvwNr9KZEp2kq4rzq0kC1fmFxdvpxy7zSN2
c+dx7dXnC/+vkGYEd/2RUAXFoiBVLuzzgWRSmSel1I9402Nf3hiv6HqTaHkzNrjB
y7UM6ZyJj6L1US5uB8q6LqSkTawkt8jRKw/K8EwkfdFv8bD0Pg02mzSw3HKR/rJt
scgXd0yIK6atfAG148PPP466vZ5Cqjz9czCEG5HEPOwVIp9r2JXk2ZAGjCqNLOxj
M9Hu8n2z60ELCqCfmS4rKnpi2cFHIPu7LWbNUQ/Zou1/gZTercM1CQsoDb1u55kK
nvqpyiPItSa6aG/G8t4pCXhMrTvCUeP32BfaLQnZ4XnE6/sT6kZMTyW4hrfC5D2Z
GiB1fmQBISVt+VnWxDLHpDuN08Fe1Y3DJyhHHa3brG/OJpyyJK3JytbbpNWk7Nlg
5FWsOnsrewlhP5Jyait0qQ/TztzK6n+tEeQ+L6NDXIKqN7qBXOcoALjUL8BYPGuf
6shGTMTxWCittjRA9C0CR2urYxP+xypGTTzsQhFSX4eG72PvhHiuED10yY+24ow5
7EWdCSDjymZej1GWBmYYsAdF/wYS8SX6Lcj4DSwarz5/pixLaLY++gkwiBQZ6ZcA
T7TKofGHP7zAwjQup6TvRBX0fUt7oaJttAu0hYdqWgZv7MWNv8Ax/+RUH+ao6+7J
+ZrmIYcqlpp/ufGg1fYKtHIDvpfGJ12QAbbCO8eApoDQ/QKwuwkA7m1KoGB7ou47
ejK9JGiDBzbDi2vxyJqBxw==
`protect END_PROTECTED
