`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZE4fmSdwXEX6onOP3XVYy9kSHtFIInwEV3Pl3BXWbP3dOVmBYidr+BCCieE+v+CH
pwDsPpZnKrQNr6TnCFzvN0IYNT8Z1hSH9NtUMCNEnZr/JIkqgyNSxYdjwelGSJ4E
ByJcxIvi15ffZnBwmV7nEnOdZ1Cpz9+Ug291DeK/Y+iggAqe1KtnzymtGqRhJ67u
kX7bheUhx2W3OFu2+Yt38Fc/7bLhgRRtacqED2TRW0FTHhzib/sEMHu9YHovODU3
APp0+isU9XoFzWUQVegPXQTxYSVamwWlmM8GmH/o7fSB+yIHufbTKFE9Y13h0up3
kB/L5yi76iZlFam9U6oYd/Uxw2xVUw7YTP2QDSkm5UstBsQFmXhMeQmxUwnXJ8yc
Y5fi3A8iKZW+ZyWytKGJx1ov/HwP31sjB4F20Hnq30bFZ2fQudrTsWJe5elX6KpT
E3KXI7j80IjIeBWf6lpvZCkiDUS9f3aJ7xUoGUtMswuZMy+F2L8AZH94FZW8GvtC
o1Zy3Rjhastq1CcAXWpWhDoN0X7HKTGVfETuVq0c/8txQ49AjmeoG/iIMXugH5BU
1yA1lARROPF00Dm2sn5ZYMD11SlB7r7zQZv7ZhSkDGw2YbsNUAowrbSch8Q30uX1
sO+9uYzDK+Xu1F2Ui8VIY0GitKcpTrNw7sWAL2PprDoUWD5oKFHAPryrPuZJcxpq
yAqy/jJs1fTPKd58UBE2vLj6HxWNaTrPtgas9OHrweoBXHb/eS4qjUptlP050T2I
jigRBarVJ971drMgH+7MYlbBskolHSD9F/ymdYV8WKS4BdWo1DxkbGVlShw3JWjk
+7UJXYZgdl51c+qC9HmdjptArRdnXMSmbpKwYNEOoLEhAdVNZg31xFY8+q+4Y3Xg
Lz5H5WUhoTEcvTeDekhqH0jQ3Q0ofBEBrVpAOINVeulPfN/7xofcNLiPUZOUmOFe
G9b189BylIdYM1sHk1orar2hAf9PSSgP8P4IGTEexz0Nk8q1Jj172GIB8OiY/IZj
tstmcIuaPBQ2M+N7iiFOKWEk2CcbuEIQUQ2k4TP6Q6nWUcfAI8OMT9GeOI/W20Ny
8jLVBbg4/9gq1+WOB6s2t/n+bvGxHBOpPwx5SMdqG/Pxs50NA17ZqxNLY6IYj6dG
gZv3o4bU26ua82kLsJAfgU6bQOrf89AJ1IvNEqmf2D/g3Bjv+bljj1V5XQ1OhHvk
`protect END_PROTECTED
