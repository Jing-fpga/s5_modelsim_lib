`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oTLcuZ53tuXnBAsv7ZWdDgBI5WyvDX1dZ6kOyvL87f9A0U22b8qMtQ4BGfFlM2J3
rVUlOA8of8giI+NvbJeSv+orhGvplRmrmacwTWOGpGOm/7AxfdCDHVRML1KyRGdN
fONM1pSdU1kIdKVVrsHw7i2tjX7clJ3uA9YgxPLMAEJCKouPbbPd8pdxogAZp7Ia
Fu6FRQa/fYbMV+jkrtbjLFw3+Pn1gLZB4wuyRN9+d82V0brgvhefU9IMIVzKVcQ4
nOq9K2VOZB03G6X9jVrl/Y/g71Xg5F74n4u6XlI12dqzY7EuIHfN8AaJ8/muF0C9
PaYhT/hB9QgEHEkiQPeZG+tnerHyn+lSSG8OBGSMkTF2k0MqeU+fK76LZUV2Chdw
1wBFLZwoZnPJnmx7YcDD0mGPtqRW4xEQM5eKEXTH1n/MYQj/qe8RTegVJdB6F9Yg
uhNqjGKlkIRvmvWX9uLlKY8MSJCMogRfSofsnttJlre409ShETsVgWOmxsYWB2ac
sxkHMEVfuwgrxuoIb7PxIGxmcdFUyrkir6/QUDcY25WbA2P8+G8nx6tmsjwuxnM6
nflnCwt5L/Ybm1zUnVel1pdGoAPJkrmQBYdPfYwgtnQU+mnFsBB68kdnWwxo2POS
SkOE5UK0HhPNwfiw893sqF9HSiXbtyl4N3ZQHSWkB4wntUvcTwfQECMG+sxr2HRi
8GTtjk9/2MsiJp/1RsI6PiNM4Zdbee1vMg59lqGXxc+h880dPDM6Rdc+m5Ic7+D5
KrM3ptPL/9Eru0KONiOugxjKXfNcvDiT5Loh6rozWqqLi9Q/jdt8YR4PMPSifl15
MRjcNbKoAiyyx6OC+y5wNSdOwjjqWzCKTv7he6aifkjct8llyFPAhI8XupVJmnhJ
ynjc9AcFcSYkEu6afGFqLnLsVil7zvB4F3yRb7cu2tJWGLcR/5eL9BMVJriMRo0T
VSsPz5019M3++rlLPYYOhWfmr/GGQVa8PkiUwNW/FuVTUhWt7gDX4Jsy2WpOdqC2
RA/AOnjV3787O7up4y5d8NNjA6+GxtPlcSSgkn7wTvXKX0GM+Y1zZgCRHuvqftOO
BTb836botU1NcOVlPiqHtUOGS0SBQuTGm86AEpGu+mZBikXEN4oKIrwN4JcSQGUO
J8sNcigmHiT4KG9+2lou0Ar8Uo151L9At60Z/adUHzj99Ezl/lSk1qQsBYKd+VyN
8Kncl7OkHi3G/cnjHZ3wYsiKaX7EzqRLG87Gacvd0wE2OPOWtKkVR03qnXzUgboq
JGXKyHQLLO3ylIPUB51VITt4BVhgsSDzJvdDoo/U1FezB5DH9ohs0OXjp49ACMhz
zKYU/9l1GmDyyk5eOtmE9ojF/VDYxzGWea5saznfEVjFTW0dZ5K05dOEYpcXoXrw
VwxgrS6mAIrprxYV1kMO60jkivJNyAXG7YbCzAh1N0+f4arYvXYeCw+I6vm7Zcxm
0KyPp3UaNXeC+C44wc4FBs2o3wvHcVoOQsvuPA9k6n1H0UZmZCP27xt/HCpTnYcq
Nh4j/6k+CsTOJh5o3SYfYivMXxYY+/vauVcCG8689gH6vxr/ijRvQ2BlVWg0xNLq
0kD59CZa65sXVT5eWuvO09Nj/GXiTXuqQnYyayiCnOGKuJQMfsleEkvJ3MI0gEuV
q1uwPsfXn03UKJ6/2C5DyXf78Hi4c4DYApGjHH0m6CceOwq8MQDpXstVKQcyqnH8
GwDTegfUZhZBKPGBteeA5BnNypIIQYaqvuPLQaz4UfiaQ/sZQYcL972UdR7l7QsJ
L+RfGhtnYcgHnle13emrEKzWHtpxPI19zDh+XaInJh9vO7EJtPx7eYOq057P92RS
2Ue+IOxgCSMpd4C46kbf4Es9Zpm4XHeFsjdMQo4vUvIbC14kAta1GOFZAho4K3Nt
HD3tSsj+3YhMXVyMt5vt+mEoJjpQWlq4/FQXLx4JI3xuNk1Ov5tZyjM1KJZcXfDZ
RVlwlSbDbNDkO+kdcxN3TFwLyMeZmTpxYdc/heGmBS7ytxU0ViwKs65ZYciIXI3U
07YdM5V1fDxskjvH0UlH3PRubI+Q+f0Qy2UkA6jKeysXub1O+KFzOASi5wFLrNUQ
vaGFd4EyV89UtoweSndpnCXRDNX7g0VezxL5cFGOIbnsS8Ji+dyCMYWkrmn5a9uL
fss30MvrWl0VQ5AnSHhuxxv8qQl6p+q0LxFjQu8oYIoOYJeJS1V7oDKb6es5ObmW
+sPt+Y0V/ogff62Qk2HDPMr6DD3MUpyopR6+y0yANfNIonUh+G0wqKhHwzy1tCWW
KWHWTtYtGsqbrBgapwynqNa6g1dxQXho1vV786p8MfVA0pZwNfhSEM/wXkgNxB7x
LSBomdwe3uffoWX37BC2Gx1SWLkv6ut+r++ggwhuICEE90MlfQG/DXewhRscxnY2
PBQz5TZ5IRpIK8txz8PWMs5Vai0HjHOm9dqw8aqTuka/1UBZybBJ41ErLPOlQhU2
JXKLFc+EQ04TJ91FFZkT5b6k6GEeW4wFuiWz8sEYgtfWJUViG3JIhbCfRhzLeVYG
4Y+wkjWdNGwMgLst68w7q5GTLQjqD1b3rw2JvZlJsYeYJiJJy1nzyk5zCdrpia8j
8fFcmuRMvfJovP2HkNTVpCl6hxkRMkQOwld2gkYfKan6/Vu5dFqYPPjspNo7hndP
AQu1s94eUx6fQmeOs9XJEPBHWDRUtDwyWKL7NK/TEOdjbNxgbXnrhv4WRNihKgE6
oCOUZvulIR5zwz4vDvEspj3EBPCqoKEwxVN2O8Zy/QuXDVi6zo1Qm0HwZYL4A3nw
J81tE2LwMeGeqhavquRhSogRilLyZq0calJxVG+89usIK3lfjKE4fd98Oe9eKqoM
QMIPRBKJPd1BAe03omBLYI0RtRKliDoD7KYfKAHOhW/XxYDzyTrcv4FhfAyMXIkP
nwdpOSAaIX//v5NmmEawlbD/K25eWmbO7rM/SWg13WfUhD+vxDK8AZ3dSXBS4Kl/
nqCScvfyPSJvbONvMuztMQbtFwSrbZwh6wTtxXSeNxJjyw4yIakraHaRkNclzIkM
gx9uOMgBhePla9AI0e01Kgr51sV4O2PEHZJUhbcON4Vu+vIQ8n42HyrS+j5p94S2
jnc9Yb2FmfniLsDXcLmMC1SGg5S1owO31WOBLCMTKHzRNAux1Chh1+H+wrmDbi0P
LuoPbgD6VoByfyUKmpOelwVQ7Q20WmP79OBs/fAWHtQj0ZIATzwuPJeEHK8Tqu1N
MaxOeZZO2fS00apTGNgwG4mrj3jUA9Dq068g5yvmjSUJmM9ggUt06B6sYWvQxDdg
lxx0OelY6FbS+GeCf8os5Fm3ILe8Jo6t8SVyDe3pwJS6gM32rmffDsv3+7o2sTMO
MZHBoX9pK6uFCbCA8jqTH20cm4L/o+8Ta1LAANnhR67wx0aVlrxL7FcIGq0NPurQ
LLC/WEaM454IeRGVki9dMPqNLSgydub/ZXiMy801Q/k1fsDO/1EF60iHX+Ao3w/c
ilWckyED/fIZsD7iZWsfQ79Qd90hpOq5fegdLg9RFg7pr+R4L2b0IvMF4M5iIm3H
8v9TLVHiF7OgDbHNgb+/o6BWX+afn8kS4Au1Tu1H6KqyTUIZHxGZqLmMBNzUDRPp
/NKwgzNuh8emm8r/O3QiadOjy7UxMIaLzG5wXCsIz/us/xbxn0727+oZ0Zc/xP7y
OVpTpR7bruAkn84MYglXJueKBip3jEIo8QUN3zVf7JUxhxHqHO/OKpKxWFdu+a7s
tKy/R+jLCbynmrvBT7zXuPyz56J0Lb85nEdQI1zRMJDaa0LkN0W/SJTmJ8yt8tsj
HBrENuBzD8vpOnt/J57ZXZ5JaE4B0aNQBKEif7S+PvEI7VL02oAgV6MhbujuieUe
+O4o78I2iyDYzL+ml9kAlNlp6nblz6rNG/e4qjl36FXcxA+miLLzvfccDXIE0ojx
lQ4PsNgRMF90Aj3vv3s4d7Q+7k+Oys56rcQtch/wrxPgB3VikKU0h+RgmWV4+/QQ
iR3gtSnu+ZB4tL/fOPB+9+TnooOf3sESAkz60GhWe9TrCHadXxaGiaUhfaF+GBev
7eTE51DphkxXkb24ZcFUbNxA/ZIx+hw2bJmqzqLSypswX/CutwzlwQt2CkbtrNpV
+CQpgFuQdHBGOSdZ7Hg754vycvYZZjLsXtg+bjd64HbDGbqsVswNX90Wn/EZhgIC
nuVnDYt7N7isvwoBds3bcFEv/MvvRqj5cwOlXCKMImmHhhj1Ealq5atVdS/xs/1k
P29mEpRWfiuczekgi6sZKB6Nid+WZN1goNyM/6GL4XoWv3G1sHTnI1GmMgBHJ90X
Arqv3eN1Gme/+PwTwYMGvOIgHMUEg5CLg6p9tw70hc0MMD8i1nKHjD9jn3q2YzxN
2ZbzZv37NDL5yj3EFNFskJec4wzQ80YgZ6rWDr2MOZ8zCPoUJpnViDf0r28DOIkM
CaZrZ9zlTEoUUxhfVhgmruXRcY5mF6fHtY/WilBr5T/7qAawKvEm8CwCXsDbwJnD
If9I8aFVFvL3sL1C7PWfL7J6KkXoc/Twma4HGdjgJ4qc3YtYVXuAYKeRHezDRQmL
RTyCBopMXBuqvKx/iqVCtZqVKRLdEX67DKAQnqn2vBvLqcKGtT1ib6PhXDXaIZrI
g2FHK5OOil9kN5b+Jkv6qwYkUid74PVa6gJI8YjlKBQ++oMC3Jan/G8B2IONrYRo
xReln6qm15Y7d1a98mf2HHzp72zI0akPyWEolOyAqANGvz0VkZP2XliU8EJodi3k
7R7CftprV5Wnx6N+wrlMAemL4UwnG/n0qFHuCKnPzQopriMj/3d68XUFwhOSvLzo
vsg5jdvAWHvtBb33RYZNQEPpLpzI4IkJYUG9i+xjYljrKXRp+r2RNEPwjTk33I6F
nMVJSQxdCP24FoY3x20Futa0GHqLBmgQGtqo7E2ZklUm6hO2Y8g+t1yNDKoJWTQN
EGGyghYeFToLp6gGAzdt879QIT2/bVzLMvKmLAgbFtoLSdBtFzznq83dnvG9nvTV
0kvUcgTjQ4BI2Wv/u7c6sQtoGKmgL8BFGrBDaCS5vM8cNwo5huYCpaZZtcs+LLSg
DtMqH1MnMrqhO9qgnE5iefdlwxvPZSCnTBC+bXEyT3/rs7cBQgUBAspykILtzxkP
rLoVl92ydJKOI/EJ+Xnryb6rfZIhgnFzL2zWgjF8TkYHDVRC0N0QGQOGzBN1hoet
6mnnkBc8JVq1oo807FwU9na6FR0kuR26fUdC4XhIjfo22yuMwMelceiKCKgwgMZh
a9Vs/sToNLzIO/hGHlS8dgPRUullLUL4Ruv/XAlJC/3qTOtn2+GP2NXYnR75HjUL
rHA0CrdsbaWjmo1oFkh3EvHPpxNBi5fn9zVGihvp5eFZxUrZgE6i4UqGVz7xPnCv
X1AMDJR2J2Bbbb7VGoJ0S0OLVfv5E3d8gNXF8932X3CrZv2Yybdv69cTUmymNZk2
alc0fjlz0iewtLs8k630M9aY5Sa02uPeNJfyLbd2wPquTnTictg7TbeFkvMfKgUa
f4cbF21QXRqNThCd9q7NJPPRkd+hkZBVPoGFdOTtRjKhPzan/lzpth1e9149Csad
81lioZj4Hoi5NIeNL2Zf7ufMaPCzWbgLjWfgY7cb7V7KbRMgDOJBT5KtpsuE20NE
6BxSuIY8KGYgfLzqt7iqhuwL6ScqMkodnQmxk2PXHroMXzbXYbjuQqnKkehFl7ey
2exY4RCtjiR60esEZFb0OUJnW6d5R3LhD6enu7w9WgBJBMy7CDgjjA/0ywf41fnm
hPyO+4vVoVwu5e+aCtmPbj+1/I6Xeyae6j7GOjMrQFHoyE+2PwEBWQGNS3BdGnu5
bqZ3c5Qt5wdDEYMgZiIcfzuIyn+ZUXTGVnu9+eW0SCQYhgmsv5pQRaQYsylWU8y2
cI3r6Pz2sKRX9Eus1CGBy2q0zC427MRyaFsfUX2dLukqIx5RBoTN2dGYoDFGJTnm
EY4uZsIjVcpa0rqK1i3K3B7CNrEI15QjI1CN/ADJ5/y3ybE0QG7Z8+LZ9wAYwwd1
r61+9HH+rRSzxsAfcloWkQjkIj/r4tMNfvbfeFURWuU7E+gF+OJHpp4MooQXxv8X
BdscJrqarWm831xK8WKjAfMznSXa7OuxUGB9Fwkh1FOxeYv1ls9cfK9jKQ9EgpXn
AsXBj4sTdR+qGFosUlr3WxGtaa++xpJshxbqnjbsPupo02XJgNvstkPrFpeHa/Na
qf53npUf8ah88F3IepwwOPWv4ogYQ0b1T0OdLH358VJs6bhMHrnn9Z1YaVbpY9By
bzHFIeXeutekwLFkuJYXvNluoXCy2NN6d0bT4eabtJzKyHBt0XMyjDWuOo34DY2z
EIxM4sW6n5ta5T4/328iS9nRfsHwxiewJ3dB9s0mSKP0EgsAthLBrLiLM8uf9ULi
CBHwNKmAfKikmXD+YP7F4zQCLnvj30kPZXVzLFzixZcOhBRz8g12mMj6vBL+tRme
hJ7mqg/Thr3jdCYs5z7zMBEaEUmfPMZ7mIozMr/eEqI2RhwRHOXvugKteNx9UVnP
LM/p6JZm/zPhZ4AIekWI0zdFFL5X8ENHQ6a2nekT5/8PZ3Z4cZlhDkyah+YrLJx+
9su4QebwdZvrKjEIkR2tj+pJJXETqbs1QHPXRN+GmGt1wROldAUvPAj6g5Ii9+MZ
Kmh1IUWbENPZ9Zu3iLL0JFFgIXrj+YKM/bx14zW87zXaL1q+upga3kvwum/+uq8n
VbFzcOJDIDHs/PvmDCF6UJaliR3JK31socAkNqQ6YJZXIxs40IkNS3attWWysTSt
EqbglEHYMOr0seC8SJxqRqfIBZCzSkCOmmQEJlHZL+cinFtJOc8ahw1URYMTFBKk
K6o236w4rmIzH+bo5dQ7OChOYJMo1qmCPx24T2P+Ry8gkZzNiFSw0JcFw69YJx1e
d0AEi5SfzrSvc8RX4gTPncPAomaiifbBCkd4USE+njH42fziqspHNd/AoKsrKcAO
OvK4IsXuRcuKmsP5qQO/MwfMCMpL8amuNRTO1gU5zKigdaULoQOEdQPiwNjdo2Sx
7bWF+p5o4wBZEHoCLvCLmdofsbQ9wdI0cA08iS3+mooBNjSz+WHod5lUXP3xa5WA
lE5aKFUu9Ygy9f2AYuYoGkBpQuulbfYXjTA/b2r2LxwMN3bheWWThD+SJkNRfIO9
Csf4kTO+H2ahJgXC5RGCpBlbcUW3LewfADQwNH0bdz7oe5IL2gb7q6TywcLfRVjF
+SKCrdhwJkXheb4iIr0oU9Pp+fXcTW2b43fNUGTs2TTe4hLnEw/Mxa5rfDUvtdkJ
NSpsZ1clpZ4OZw1gB0TDLhj0bo4KJpXtooc34g0847CiLnOfbvs3nvERviC/qmJR
8unu44ED1Q/bltIywWQ2EDe3zi8mCPE4rQheFQw8FodjG+VTaHWIOGF7jmnICBKk
CnKu0JHEA5/V7Ggv/LH9l4QXzrFqvikFIW0UodQ45UPmNkDQ2khL+qP1XufjaVuJ
xdv3GOvUFPmDMMTTr2pKhysnnMRuqvEwu+7/jlfTONs1qHagz6ABGK+4GoLlQpLu
XvD+OE8GcVhY0nrQcTBTZMT0hqRTG8CMpiIZ93p9I7AYtQYqC+fuw8oSWljOuMQc
HNcpD84O1O0Mp3i9pQX4vySxKpgvznd0ybzMGY/SWFJ2ysKmJDZM3Ks+yebOVclP
SJ1FKUIKho1gd+kiND9hHJ1ygYedDBo9IXftteIkV83vaEgy/nJWHnDI3vIRsfWm
voj+2o9Y0e3/NIUin60cn255sLMJURMm60WhNJ0brNvEoV3oWbk8/6J+Ldr26JDh
jCXb3WNktjwe7/5SpHPOHqMS6FR2Z6U3EYoF6ua3l59XlBMpP2y+m0WQYH6qLjwp
L7ebkQcDG7mAsx1dR+4n8/Kb0yc8jFceCaVz+YuAaqyGwUSEip0s37hQeT9g1MTp
43NWgeE84YU3mYyvZpvXBdAqLZPrasksxLZ/MITZR17udjkYtlDFbLLOIf+LMJcj
y83LEYFwc8jwFmDdX/1mThNqU7qcU/aPpGF3lZJd9u9IwcCtBdmxbEzYA06yS+7J
TG3oTr+2h2/dzo/lH8QnxcKdt2hxcwVXv4XN0QOTiuE9O5/nF2Sd0E37a+YfsWW7
DNw3J9T95MgmUMY0TzLz6MjfhNIupiCZp1BBQU8cVQAEyw8S9j7jFWE8bVGMEPKZ
6tUT4RNFhq7eNf+eCC3G8WicoJzcv4U8TtZw9NoUx9cZSfsuEWgupUZoSdNBxESX
x2jKoLPRcSqGcMdCwssna13roPtACuxW8qqxFxXLMH0o4db/FFBOEFlTusiJ04n/
SvAPTuzmNlOMBGXnmhMnsUciLVcg8yqb7p8IWJpKOMWU0gRGUZwidcEbNQAqye4O
tAaisFXHOMgtORYBdQ001SZPAD53m3qovUeh3XjaOy69lvR7jNpYVnNNeWVSzZnp
GXSMuj6ERkRTnweBlAmVvHsfqhyNR4CA7FSQQ0J2uUgaFIKBtnp/TuGpZmYYv9PH
L+A/QPltMCEvLLK4pzYAv+o7Si3KoauNdbJlaSSFA+osHApoOSmIQLZ+Axe1w0sL
ij38mS73kWsAKTvVBV24WESGh//UpJUpcLHyhhJGska6RQsfuMqX6KSQ6yt4GeoQ
cAjOq6yQB7BpHTCPGuabx4os5S3Vq5zyy/zUJrFv6AWHU85TnubDCwoWfKkyZAkA
EeE6H3XArO1ed2iHToVuoCRyOGfyFIWIU90ZnqTN4i7ZjqZAzp6PoLuPri0JEN+6
3J8M1bVfBNWhpcggL4Tao+2rfq98S+wt3CbIZU2EFmwHAGE0vZkhzKVG7TjQxeiZ
iOt44wkJsiqLoRFLF0vY121l30B6JbD9bdKsejlvbVIZDnXHEQTdtuoKbHcueI5+
7ZfB3y0o01Gw2U6Ol1ApzOqpgMG2KumR3tcG/hQFht1CR3WcQ6SWo9EmgVjLmX+y
/ujYOMMRds/8Mytg/YLVx1r9msOLJEKNHaevoXm/K9IMIa7znq/nP+N2a+XwHovn
VGdj5D5nlRstnQF4Cf5MXdIFPx2NvQTvmDanHleb3NAvX0scCNW+0fSk7cCWYA5K
LN8Gtp/3dH0168SQV67am6YqhYGgCV51DG9uwJrAOPHqaGM0qu0GgVjHJ/7EDrsh
gqEB/HyN6sGZoepj8OviVB/Mt/bd2yFdKgDgr0Xo9N3UIRYPuPEh3vwsu03k8j3M
4zSxF2AInDFQ1NszRISUweF8s57RySMgrTwsxLbn3uQz7NsdvTMwUgcRYO79U+G0
DHJtYth4LL/BI/Hn8bxPNohlIgNtriJbOR+VSoNePDb7PyxyDU0KEKSO37qmDOBd
KwbWQyqwOp67lBU8uYZHXXpJ8P24bdl5YYJZ/KomcKbjEPmYhCeoXY1KhOZY9dV3
I1WIAeqzDwqJIq8oVFr5Q8Ulqo/p2u0S9OeE08Nni5yt/pmpHPAw4MGDHBQvxLev
tPqs/gX6T7XHj9vvyP5M8/UKXqTuJFIqHRY0DYh6ioTMMBSaKMLRJWl61fvw2Hqy
8MYqarcCVXOtzHu2VNcHYtKcIeCTIdJw4yoxEzTs2DmoKT2xqS++zMa73VU+vNFk
MXO4Nc7hqbQ+M0o6q8ITAa3tT4AKOchjCIjizih11YP5wxIsDvVvn7g0TXBUTszm
gwXnmCAaZ5pSU9L6x9rvvyWqqH05upQnLnG5+EDhRiqFBc44XeXJNFpw66FF8kWL
10wJejzbCFKMrh3hKaowx9qzEB9DDrxiG85xg6jgJjzX1Yu74HotPb6E8SMCNQNd
CaQ0gJ/vn5xtFJPo3aYqFce/L2HOluBiAhLRtXsoQCdj47Q2yIUfx/3UjsOXGo2r
/QcngwFb7h7hG1vdJlZGs3/nmhlzZdG5l9YfsEvueKZEAw1/IIbY15AHmjQIHzB1
w5MNE5U82nV56Jtj9+ob8g6t8t/4+pH5ENAJnCIuo3CrLHNmdIY+WjUVk10cbQNq
IgGC9Jru6t6XWColcyl+8boVc6jxOwryqVjIsX7dEjK67X1SMQhtU+oUksbqGacZ
FOPqKI1UdAROJ9xgbcNHoz5n2S92OKhwArUuogxgf+Hwy09bgcLFOSN5nBXVUUcU
y4ZVSMWkCjL4Q6YPFbCZfFzDyLXXLLAr7qnmWG7DVsjYO5EGuId7XBhg7T0Md6mc
Ov4Jt17xP3xPokk0tMbMGGeIprVDRtFlZ4O5I/Td5oPixX42To8zl9aIJ0DpyBeC
IC0xh+5onQl/3TnucOwQQxVCe2uRfrUpKUe0bOweVpXdkshFZE/45sJlQOs7VyWR
FOm7/0lXj8WnMhNGG2B+U7MIQxsS9EYcOeVyijJcrt5UVrTPk+QaWNAPADhfnCCy
+FZeu4ph8xYM0haO7Nhdz5vcyQdkda9e2/vYhQcgF16phc9NJYUuR+CYjytXnqyo
FaYE5+6Zqz6491BwLojMrpzQsEt/qXRwy7E2Q5cU6U1RPdkpdDwFvzigNPnZ8eP0
f5osxSJWu+E4pByleLhhIwh330N8pmwAePmtRxSgKEnlM9WeCzUqJZ3Iz+x2B0Hb
HN5bHhz0qMn3laxffQztqpJItDIb0T3ATAg28Lf2oXgxwkKmZrVpzMtMSbIXCIE2
f/BJN/istI8QvyPysvJSCnO5DdFImHnNF6MslIuVJXmIs0pj0CL++1x1V/6skRxT
3d0fzbINsHLVkrwFK3qYcYdHSiK/NNXGSpqZe8lMekaqj4uQ5LhWRr9t0KpeJ5VI
Wly2XCoSi8yw+Z3Xy7+J8U94lZZSQOtfpdsZZ5t8HbD+lah6/OXJF8hzRiqO+kQ5
MmsC7Fk3jj1GZtdZajbOtAQ//xq4Mmx7EyQ440aGwZJShJENhypetzNoS3o2YFww
zEosYavQCHMHtZM2AQqeQMWsfvIU2P7/lqIGe+7syMplBuGwcJGIosYBZ+EwTOeL
xoIEzK0bZA/rno+OkcitwkV/HfpT7AdYKGZLY0VKtvzWYXfwlbE4qbXxzSAIiHxr
3vxi3We8yUL2viZFp+r7ctM4HfhiQifQqZXWlKOBMfQjNkgINi5LoBeYlIy8rz7h
pL3s30VWtNPPJ7Es4rO9foSqc9KnIWYuCdaplQ/yRyKbVqUwaOOUzr9WUPoUnXUy
kRrmhKjVCEG2kuhOM0YgsRGnB9nenMM42bzcZiXDCxzPVZyfS9M4kwJa8PSrgTmO
tiVVwYjrWwER9PSW7RMApkxS8rLWd1VRCHOkDbZlX50q6uVxT9IWZcatdzHV/kko
KFKTnytdVZ5WW79+ncsR85hNSPmzDxVDDotXDHqX/q2Y1QI60MtoQ4anZe4t0iM+
O0oZ+OM5MJBRNPxtEGzCO4zAhlHRVK86UfsAG3P5x5+iSiGms81MCQsWeK7dbT6o
nw1frRvEavOTZn1lU3JLUQzPerUZ/0vvp4HcwunHAa/6ojmNldO1Kl2FYoSGcDJE
TtMOu0eZMXT0/njfB8cfI8lOMVqWLI3vDYSsjq0wqWFV6mLehpSt1bnE8LAi2zVT
U0bbAnz3CBr3KDR9Kne8c7BnSTF9/0NLFtfw7gouQA90uYfV2jWVfYLomJXkqDt5
P9SktmblCiiOPXR7LJfaYGzlbLQx0MIaLAZmci4/luYezMZtrjyzp0y74GazCcfb
CmdOSf9KPXkJhy261eHsnq8twqhfXQ9AQNlINPBGqzCux6n2ctGAmL6XvXXD376y
Yq6tbS6eSBxmQLY5F6iL8zZkwyRPnrTS/qogEM7P7wKOQb2sfEFOHjqHmtHv/y1a
EUWQ63qcob6To0QdwUjmT4Pr75N5aX2PpsaFL7+Tv/7f+dldXBnZ0IVQlM4T8ZVy
G2ytEIqy5gc6xtzJ7CrRbVMglevhRxMSTeiak/37q2eCg3zA9JwYI+3sKm4L+ZfJ
4jXw28m3CcuRU2/lKAnzI1KK4eHJxBg/szvg8W1Hmj2d9D2R3F++6CxzeHw/NX6t
Dg9yBJ66vOQneeN1YPgCpLEdlQb6r5V8C6DbE5qWDGomQg+3R1SjI0JmEhZL19SH
kuYfDQPrkIvfljpg3czAshkJ8J/LDMFf9xp3D++gJAy9HwwEzjdCDOLpxwiuzJLx
SSJrhXJ/4ucWPa96ow51SlZb49RuaQYwA/RhNMq0Fq60CZgydnIZzd+7H5gQQAKr
TozjubjfLtCzZXwJFuHodhft0hJcOiPz6YpW20/OJCQoJFnXTtGvhMg0cDaKgc7W
xfDK2v0x7FjqHiPG6RIhAG3m1EnMP4TDsZWd5m5rVGi1uIZAdf5OC5Rn6OFqsj0/
HbwRpejRrHm+cpeyHFiiimxuP6NDDwZbDLg+LS/AodC1+6By7vLnFuvpFIgkiGlE
9TUKgsnppU4XEiofrdjxYkj+1o6WcSDlOgXcdATkIfpmipBsXkKZWq6sEoPlHsYo
voSz5eQq6bha/Wrv5u8+TY5zQKI5sse+fMKSqbF7LhctrIrS+rkIidgJ5PPjTTvk
L+3mDMxPKMA2gx1tgEcX6GpJ/yEq4g4YzsEJObmS/Y4arxTeHmDy74RhAGqIVD75
gkdZdtKmEM5cGlFthR89MgPpH1eh91eb6ZVstukyT7j7QuxspGRUv0oElAHUtwtq
T+xwelPDhhCaEafbaBZq9SKzmuwvnFVzedrYFAJJk//dfJyc/+z4ihMlWHpHpq2l
W8efSpfBhIBDb1VZ9Xa85IBYgnA0k2a2VW5oT0YUaMhvdwVeLfP28Cr4G0KG4yLl
`protect END_PROTECTED
