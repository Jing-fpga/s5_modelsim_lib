`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KwOUKe8h4eVJ9cA4Lpx5M9Dvwh5pt0u5r7eeMdG3Uey45GJKLHcTMZFLD2ITuk5a
xXb5+0atirXpvNPhRlXcXvJpHzN7GTJSCN498vUx1T9FCTmr9U06KCPcHIQgbLxC
vyCnFdrmPvYoVfXpENWhbB/By+v2PldXdJBbOhfuI0dh9lqQljJE0Y2c3EwEn0dL
rZYCDTwR9fi5b9pwr6vt1oa0OOkQr6evsXq4xGgZxyumOzovVq/UH3GE1YHK9iH8
QYpVS42S1EXV3z3+x6n8/stJX7ZWndtY4XfSNClhSSuXu0Mwvvv+npqdLQ7sEd46
PsFsfW8ErAleIm0HBeLGm3P7eKMx36WUShcwM6n7J3ro6PPf6/H7uvUjl4Zt7Auc
uXH2dKBFOdYKeVKQtQg/RST1Eex8B7nJGT9j9waEOTpNlYsXK7T4Wl73mSx/WXgR
VLwgVS2bkQxS087+JsNEMN+ynGIo017eNKHVhcNmwx4Yq1MLjwM1oGrn4N4DuwMM
DGg5dhk9A4TCkadfYJWjuPgd+j6aILTE36OfF0wq2xxNLMoKAJjdDN0G+UwyYVzo
cb7rvRCChp73Ukdhx0yy8/mlWgIJixvrzqCmA6DUgDmUlVne23NQLLEJKBg0o8pz
ALls9vIPrFruoNdFZ85VywZMZO26y8X+9pfRuzFs85y/6dyb2lfgs81JyZcl7qX5
1DDcKQygifZKaGXmMQ2CVX2PcU4Ush5BXaf24JYUo8IegvB4rnGsoT6zesXMTnLe
bZ3GFTc6pGWDIEqlrcT5L6xbJe32rG2TOp+KYZh2e+VGYEbB5zOQk6Npq+ApYsYY
unF1q7VC8tAByM4hyNcjVSgGnz1FH02hkRLjML3FswUj6VID7lMHWzco1XPSNyNz
6nFwObBJsz1gub8ZadUhxXzXfV1zpEKYadk42VK5kRAoO5vYtp+AxZ3di9yzMzlW
SMSZWs/WcwqvMjjn7CfKmvL/NR2VShOsFpWVtmIZeV3GZ2O10TsIIDEUFlpblof1
O2R3dtaO54eQC7XBEp9Xzs3i/PoQTSaQgWYBqDUWEdoiJyEg9Ezdl4UaWbl1hiIE
/AINXaNW4snUkfjnEZa6u2B06tgqqR8y/FCPT3OrWrLOML7BhLjhRGk/aPsEwHj5
okfpkFcKUvlVXoDUnqpltwoj9T0gPwJzHl6G522ia44AzQo76Zzwi4wrhc14/kbk
lStCpFbjC9IKr2Aj+vGE78KAWiWb1Ecc0GiUB2eslm9inIh7dTzhd61DCGXvXa76
PDTilIm82zf28YHyLYmnnflOV/lO6blpqUQ5CJi1Uxj6YPqZmiMN6tpVJP40aR6c
DrTJEuBMwjI2Z8VHlPS0vCYGnUbnTxhbH1BRFw83EduY22vsee3NeqsnuwRrkA2n
W4Myisvrd5c7E8UlRxfU0iK4ascTGqxTub3bLXTXY4K5mHVtY1nnGoNzLHzDD0cH
ANKpPzHcocXNFYH+wM/L3GrBR1LSEAOPeXQD2v54AQgIqgBiP6IzmGX0abNqB0oS
c19v//r3vDzsZDaRHBFqJ7d4w7GbkgDZRjye2/Q8vPcInZVQtyZMFsE1F3gdgCLo
e1Zu5CoCSLu1xPrVg2yuQIQCMjMORzaiTNUrJpk4l9DLFmwJOXt0qOHBGiyLKQLK
qAolYz4QMEa0R1pMvO7/QFf3kwgwEy6zpyjzI0qyyr8as3zw7k33gN6avpcvNgW0
Ot9XPcDzIuPsasBdpXy9epe6gxE6hdvnSoyz8uWZ3qIsOKHQIt7parRmMN5eyMvX
o6XMElOTOJiFIyJ96P6o4zNO9Zxb8AnFWdBb9M66Y8cR69mE2TGaGWynvMta+2i+
44LoMJdcEk/yDCY/BV+i8rVaiYN7ynZDitjwcK4yfXoeK8wegb4L88da3Hp7/9/M
NO7uB7RaJRDyM5xXCNkY0MgVai88gL6pF97FeHDymsSm4l3dDPutZp/0yrgqPPdA
TWn9Ekx57JKGEUJxnZQUS/CALWiu1KYg5paYYS/VDRSJkVvpzjB0xnjrSeLzDI74
wMyK8UWt2vU/FHrTxpJoNt24DozFBDuT2bXE73V9aL7mk+1ENNsqOyOUIvGHcRRI
lqnnA9PwZkPMAklhGwXlIhVc6N9Efu4KXWZuX+PLCaM=
`protect END_PROTECTED
