`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ik1zxnYB76m7CpFJAOOrozz2D2CASM3NYt68iORHKIv1ZHB6eUU4yhcyOIEFX79E
TmLVKnfDdkPLsjwqCGwVXQNtApGrIPAjsXnEs7/jqAjIivsqnu2Z39Lr7Jvhndt9
6fnA/V/MBFLSMnbJiLJBenwWJUezs1U9bMmpUTGM6aIfvNW9/vpO9JomMUxhOLEj
nUWGRyGFLUjOXcCI7Glk5g2y9FrlLNSAIZC8x49Ii6zA5eYqzrfHMtbgdLZuVYhW
7LO7vavTuxiKmU/YT9QLBwXyeE8b/B6EmqFg0pbC4JLHbFw0tIeVGQWBe8Z7JOQL
wNQ3P8xHY5kCWEUs8nuLhaTkqMqcNqkappMMpdrpTkxi62/ECKjcuXT0NzmXHdnC
NMiasbusvZJUnnt6Oo+JSA==
`protect END_PROTECTED
