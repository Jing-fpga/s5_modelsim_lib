`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8tiGbMdfFDEO7PytvhUDSzBJzYY3yY4txX7ovvJObCJb4bpO0825HGZZKzNogeYK
thPMqMZnrycgEjPCfkCHGNhlgZ9VA8MckB+fUkZSGllEHp2ItCDo424L+roB/0S6
EYoVxe0bj1dmmXiJnqWuK9zQiRlDwUB2J55zXdvG3TrY7XTWVUm/d3YKzpxieGyN
8/xwQ7yyUBIuTXiU4YeKLc9Mz9vhI/GFI23HhNbF/z1Cdh+oRkqcBR5PGDy55Fov
+55PumI6QefiXZkPiKYlzqCG+Stv6XbLfTx4Vo6cg+YKYKd3/olWZAexUzqiCzrJ
vAu2dmXwf6k5yS7VALHkOhUEQBna70vTo2F0/XbhuZKwsppvS7cfBrkc2D1fwX0x
6uSy+JmhSvieXaMHKCxpNS/7teY8RislvavsGVkOpX2BSmDrhIv7jZPLicId9Xge
V8Bybaiw86dLs401vw0Qp6/C/KHfTuEfIdIWvCd6et5x9bsJseb0QQwR6QHT83be
xQHBmxA0KfLA949KXhzOC7BSHzh082ap7uV00m7Fz0pmS2m79F3wF2qpA9CxrKAM
NFmIBp/b4i+IBlNPTVMuoS/GF/VR3faIqcTNszX59gawfbKEE6XDBYWJTLQrlkg3
rIeF4l3lSZE4Lw8NPBx4GvAnNIiCRChUvq/kczU+cV7wtXCZcikhuoEnguqFUVr9
o/sJxNSo5i2lGmKwp6ge1o7uubD8j1H3GaAcAnu45fQTuTP4faEqhGIQQJtTSmGi
`protect END_PROTECTED
