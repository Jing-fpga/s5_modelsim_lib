`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EuZTaQAu0gABLlSEkwL2OiEZcn+2m+qXx4ly6GlozDtdDXXUW13pLmFVMKcfLFZk
DkW9hPFeXKbP4pkF4VP/NbOVCgjTMebYWWMoFQ1iv015c107zAU3l79rfatG33m1
IqsmeDpBYSxtEw0y8eh33WFQNFczw3BvIT7Uub4OqbGgVPuNHjxk/pw9nrip3Mwx
TrMabsXxQMOySeUgE87B0J6ethrvgFU4c46i5WsV7deG8F8zSLQWDYPcXEGYX1g2
ZnpLV1rjC+11WbJ0F/VE31JVl71EO915xy0747mGjmes/eedxWZEqnoauvCrq6TE
U6E4Tu+D6q1IRMC0bAFaiPm5V3o9A6B8Xez49+ZYOzv/UsZ+tbBXiUrNUFY8hqcM
5IvUYrZWZHDZtm8LRdL2bye7FelY3UOs7nYpvX6l2W71wBKTb3pWvHjl2iDCqd55
Aq1ihBAf5chF61eLIzFFrDAM9h5+xztIBp4WoBtllozqty6GBeBCpAWGOnFX4nB7
8/2PyhtPSGKlT/PMKdwlTz7oYWLYHOFhj57EAiDqtYcyeeoN/sMkOci5giUaxl4L
gve+kssQQGwX5SXFvEXVc8wKb7xDxMJGpTP2/FtI568u0tFHndv6w9iU3r0DxOH9
/WUjBPnUMjRuhHmPfY8uA6sXXnels3phwniHmdHmfzqyZ+Vo3HRCJrBijKlDV126
Ip8p1o/W9q/ufh7Cea9nuLxfIvB1Nygr2RoQPWOwrAx1uFo9Je7hk2WafqK39m64
Av4gbdsRxaNLGyucX80c+GvuS3Xi2/9FlCLU3LIuCvWvVnRd/QlwK4OWK1rHB5rg
TNDh2AH86/Z+zRMuNnphA1pZSLG6EMaavK57mE8jGQw2agGgwyBspFYoyXf3J5Sy
36zGz8MDnxBvU8zrNhayszNFYeg9Q85q8McNpyw1hJPF2juwsguNpDLhpvWsTAjp
YwznyrUhlckBzwc6Y02/LCyP4SJsRSaINFW+ncuWpSSMeCEugmqlqOX/PENHhraY
JH59bh5f1CRFV35Yo7ujXDoN6Wq8YgB0Kfc8tW/jjLirbsd4JDMXCfTbMWCn/duT
0Z++tZ9jDWXj/XspfIQTzcexQT1njsEW/grXX+wC7wuug3uh2Y4/CPkPLEg+A2/m
xuQ5rr+sl5zZB+7ZZRKehV+PpzkEBU72YrLGhP8jVy539wfqgS7k+QOwG8sFyTc4
09hh+tKmYihLfMeTGFQQWRoRoSmMybMZl/FoWZgOiKX9KgZOq7oYjAXkYKpEh39K
h7Oh2Hzg5HjChH5pp8P0zqfKpJ9G2sqSMdIFTUTPaxzlQ3W4ANQaHfdZyVQFQoSz
Mor7mcwouY0dqqPNR3ZmdiwB03Wzxd8OMgZ/JirlsjyyIBV9BB68Tr3ecnz2G71J
CoyNHpoxv4HmpBLEbTN8NFUq1FSuInLx+I4NpYep204sU8HWh6aKimODVhrT59Qv
4PGt54ID9FcKRkUVzDKfJGuK0//qXWLnx9Scqd0jn9dFrC7Wmd7zKLdYudO27Xna
nGi9SzeTcsjY2wgYCKSb+aWCt3CumqjzBlTN4cVgRlgOiq94m9wVUhlxOSsTkHxZ
i+kaF0+PmFDf3jXr0eT+EGErG1Lt7cxC0F+UJfePEJLSGJ304M2GTW5WhpY5lKI2
BI26BD0bZyFfy3z5MVi6omN4oRE8DJpYP4mEvj9roHJkx7BTTZWFl94xGjxiI0Ev
1TXnEHP8XCic/F/Johoq+PpZzzDNsvPGqAiFCq2Liav+7txatmpFiEse7foIBqGM
/vHSPKNLg/ApMfIMgvm0CsLB0iZL/2pEGTKL7C0szH3Ztm8KP1oNZLht29PZvGNo
jkTepIXZIn6k+3/A0zAzPbgAztzfH/3QdUgZIUX+HJUGUXfwzWa0hbVemjBj+/Z4
KurL44+MdXWCzBB4pA8+o6EKjK7WR9Y+3/IruXxCxm6VR+7Ap25ERcut6jc3Ovs+
LPoKM0kKXfZsvhSdYErryQr1naUoT9agk+P0DzMg0RV5ttft2FaDDVh/5dAMKEjN
Y2AqOJ6Ro04OIC9/66fkGb6IifMlt7B8NasvdzV3l4+GomAwxLIX5lzR8JB/2RWX
8nmq4ADmY+Lx/ZLZVUzIzEzlBXKqgJ4vXsd7hPNTtXPdUw1GW32DPq2FaY0kth5J
11K/SXeNMmaT4dRYKCBWo5GMhjKqB20OZx4wSozdMaFTDoK8+Au+wdwZzlcYxQrL
O9S31WoNJ3hMni6TaFnJ53ZIC95zSQg3Hgk6Bq6oMcInI9fJ0kJ4yZ/aVytl+dzc
yQ+K77IJCSZjnBsdAwuZ8mLmi5nfxeHB0KWpUh/rKiD0pGBe5nuM2kmNpFFl+x8Y
bRhZPDKLJTRpjslc26cTmkTlP7mFWkwg8Y5AdNKKHS66/EOWkLIsYelclS3/HGB2
BzxcLMHfjDALF85rMIdzq7ejTfRdGb/1GYu1v4SjPECiXj6P1X6ZldF1iZ/u87A5
ALy4aERespvWaTbJJ5EFGLycRW8Kv6FmfKqUyQfNvv38cPKMtIa0tb2PkLFRYJI5
QRxF+bXGdADQBwGwkzpnGgY+oRpomtNAefxuYYW5xiqhwwu30tCRxnICcTZPzPqA
nGHhWs34CMJyPjJEw9u//WXXzEQq2Vo0i66eWKQBYbxCXu6FBNxMnEf7VkNaERVD
WE5x8g0Q/t7Ae5H+wGoaDDd/F4WeGZkEpvJbA8rcIu1pHRBu5qagboKTBjNEv6dv
GJbyqYK339cI+ymNovWanCoLAPbuqgel8Ve57PLGC6VJ49ggXgPec7z8QrkZ76QV
pXyRba1C8HqUNI/2KpXLfCUpZwuJh5vmPwGCLcnU5NcAaBCowv9Zrbr9vpvu/FSa
MUg+usP31Sy/xpGxeP8Ea7lRk1dOjNUM5tk3cE+XPpbhhnQDKMFZNz7h3AluBLIM
`protect END_PROTECTED
