`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eSMofb7rrjuXQz8QuwB2+1MjAjndWEEhy6GfkdPof5nrDtq+AShPb89bYFYPqaGZ
mF6oTwzWYbOmpTcKnGH1PBlMSyFoWt4Sjo51owW03e7M7crNMzkn5VrOvr79LrDF
6GcK4H5NyISdSmIvuXe8NXVulPLyHV5052gk7AAlT0DXqAWKz1md4qlxcPgzJ1vF
MaLq/oKFvptXZefxYNuUajjn16TX+M3GW62VmWmEwh3WqS2WZmqpEe1Eif6SGoSk
banE0hjLl1lQUup+bdSd+v81edeiEnKOMmGmoqHvHGtxDL8gJfMMECL4id6CsnCM
3kR3kH8M8XNi4t7FSiBL5frXcTwLhVnKln3UXOsnDDc8Y3JkJ2t1XZhPQm2aSIcT
Xf2ACjgclUnGENtVEJteCb9i8DbLnhFk3nLOznhu8sEniBGpWGXvUGbrbgNaHJ+8
9w76Q4VbIpXC8vm2VC64NOYZDpZlwR8rLktWmjmFt660gdl4uW+342bj05T1xVDM
n6H7b6cN3VtqPV8flWKtQRQr2UQJ6lpckpsfb3ynshHeQJsfctGCOAg+qKqcgCVi
sipOdWu1FdE5VT++h6TAcZT4WLi2rKhf4V6/Hz8bvfP9a41Il0umqrMjG45yJnFS
QIttuiQln4uUQgUibwZN48X+aZi0PeB28I6Uv0ea6vSD39iSvVIveWCjX5cxvEKn
P4q9xWyCC2Cl2XL6Fid1vSGNrWmEtStCpetbuAq25va1HfDEtK4OPibbb47AT4pW
AY07/6CJUJWyUHnQ6uKn2yPd0G0+jmXkBwNXS4XY30SiC+jUHTg/59HbDNJwufvS
HMRzML/Q4iPF2lbEbk85xI3ROu/D22dSOaTIZhe7fGJ5lUgzWB5bq8CNalG6I1+Q
QfvkUgRdNJfsgtJM/CtwYJ24BTdHjaPJQHI95GycQTcYOj43ABug1XiPScnNqbxS
m15JGzvrcmpEaHflXGJRD460wpxjFJCyQG03OhexzXOgeN4OIEOTiHUB2pRuPVEK
7NbSMsnIde89XFcBgyI0VzXTaaQZWxSsCoec8R/39kzuBgmpuw5hp7vct8VqXhmv
Eq2ks8hIYGN2OJYN8eKPs7pKr4rgoPAYAe75HuQ3b9xXumkZA5Y4ZV2RKV5aEUZQ
JuWmybU9j0heHirlpxqoGZlbpGDH+NJTBA69o7oXn9Z1CmOEFuBAlxs06EPwuYPP
zhnTH16VCwZ2comGI8g/WpGB9dmRIpSkaWm6G7WaLEiidEYR0Q/chuKCNfIuIOzW
bgIYa+HL/pkrMroFeWHuhBCIZqiXW/l1mBhmEgZyd/g7ud/dTqLWFuKrOVa7ibig
wXIYJJMNFQZhf2Apt/Kj8IfNfnezlf0ajeqLcecQ5yXsAhEm8rSu1dAUjh0xdZAF
ZLGR5Y/B75ctVxPN+/WMRB8bZqlDeaCt6j3hBaNL6HzrHZt/QFNxq8aixA3hS0KL
sRBnb12bUDg220W/5Tr/HUr8Nlepk01REKr7wEPVQkgIKNhKjplgnsPuVQu/Ubpm
klCnd442/CGgJ2AgzfR81QKDYwPz5kxSnhPofUrGtZQaEwIcrWy2eIu8fWQ11mHv
CWROs61+GDzl3pngwyLp4VAw3U+0eEzIIdeBywwOfkpc326uLXq/8hu9YXOB2e+t
7kEdubQfmp6BBCwINvQcU/XUmJW3TJtQKN7PpzHi9Rsfo6/3QFOb2FsXz0FhxIh9
mGn2KqvvBN+zUxWPcF5749ME+i3khZvcFzgja9F7ru0x5WzmH2ZfHe1y8gPFKADC
DupOiveqluaEPPFjPmUHnUPRVqStbKK5d75sK57IPFCEwHKUO6LisWfvzBJ9WBl5
qJgFZc2G5v3emVNewqbaeLf1Jkrm++eQO9PqbjBMyTMP764ky5eVDmxO97O2pPto
I1EiOM/WF931P3+Mr3Opb/dBrqBz3+Qyld42/NHEbO1Bg15CjJ9mt84KkBcf08RT
5cXbJGb1fUiwy/7avv7mRnvKUaGpXA55DdBLzqzLoEEsJcWWAIaGFjtYzKMuojIH
hZqXrzElsuIRWXr4UeyANWON87axG3eYfk7eG+EPMN7VnmC1UI81vDJD6e5Uj4vb
k1ivDBcuO+lVEsdg68n9T8/ERwLpSDwess1dS71f31X7qR01aVNHoLZfWZBTulMR
ndGF69DPR184eDDFGZj1iIOZj4zCXAsFlLDL7Y3BHZ2UGccDJmEA4gpC8ujvvM3M
45g1Il5KscthlyeusVJKHQ74NSYm/0iNC1ZYhC1h9+rL5nSajhCs/gh+5Foh7/tq
uRrvaXFcfRc499l19XZ+bka0UvE3lLrzLAOySqb1rRTsC+RFAlmnGeIAMu86dIc2
UX3w2H33POCyZ7chuGkXKScyl97WoZAle5EUGxyNYFZQNAvw632Iyi/HLaWzki9D
dZmoXUgp2Yi3hjjl/AnRV78dTU2E906CvFRpVcvbtjRPj4vD3pWn/HVsbOKXICu0
5E7gviXCHDTyulpG0jYSVYyIAVsJv9tM3eHQsa6gK8Q+M3Q2aKcorhrJ6mrBMjju
mrNohu6BqcCCeFEU0nl2pXIq7HAqdHFA/1Fy2IgXlDktIw+xojHWPWPmBbtDb41i
iQZPSzVpXQawfFsKxE+/mhL0NGnz2TEMec7dS1uyrPLiA5bcnsgDmjAFiENB1IHH
ZaPBlf0rfLiew3fRXIrJdhQE6JgyPFPdw67JNbxLhYSZ0VMEB3eQdRnhxB0OpLGG
AlW8kx0F9Yc0CQw8sQDzEH5EQ6YXROnPgo5C73+fEOpFu4kRoS5H7xt3VaIuSUD8
ALiO7rte++hXHXc/yOGyedykxOXhafGq8b5fpA5jfW1BDCkt8BaF2TbaCfgBi/2a
XTh6WDZeoy7c0MNIhCSaiZfAzjJRBEevCX2SqrmIdf1N7jsirlgNVrcw0XCojKpy
5TImzBBOTHWIxYuwph1KEBFU+ZPSiKr6slTrtFP3mX8reAT8PetQ2qCFlffCjyca
2T4tuFPz+DJ/Op1IjngdC4tvDNev8fbVRUKdGBf7ED3I+JfFjueXEJw+alskw9CK
q3f20GK1tI+ajaQhHI+aRh6CdQMXK5sbfC8A/kZ4WoDfAHTrwn0T7ZL1mubPH3fe
QwFMlMU9ym68iFI8qZ4YXgevKvDxqTHjO2HGMAW8r5LcUxkmCeW+t3ix89mpEI4V
8GoWnBqedz/rAktl80fwGfFCAqX2FEV1Xs1wte1vItTaa6LsO6m5y3Pstp2QkWs2
kXolAizlyghEsqXC1iZ2x0PIUTQa3KE4mJT5TtfpKLddpzuTalAehven2jhOs7vm
EHxSPZogjYztY/Z3J21DFtrHfKhW3B/EthdFM52hPhxk4nwgaj+uWgOKlPMvRWvz
xPyLxarF0y3sSklKfWFjUGpPRaX46dnRcmDed7er5aaqeFxC68Rnb8seqy4TeeeB
r3grWGSK7k2iF5t314wZ+SytsTYXw0L+TizjehKl0L2UNt9qesn1sp739d0Y3dFf
Wkgk7ZiVJdn3xBGKAvJlvh2g1lOMwkV3n1PQc8qnZRuir/bS0B+dvGdWS54zv9FY
QguRaixyp7dqpNTO06SfwEG8G3yIYLTwVDHOHLmo9Ofum/iM21UJlMs36QEdwbJX
HyntQoXQBU2TmBNM2Ny0YQFx0t6M4B0Z43fDr8xzN7gHtm18Y5iPPSWk7ApMSToB
WRKbcM60jgm4cq75Nx/fMMnzRfllobgVaNLu+FEAX/mxYdCEGzuW/O/NHhR/ojk1
LmjwmYhdtRM7PhGgpK760RqATtV1kR3vND5Lz/YOVYqhV768pUP61QKmPJ6V76Ef
YChtOiJOXmz8BDiskwwJF++XOoGoit+YCEO94WEQCGjy9bsgpX6DMqwrxnUa+xAR
l7DHJYj5ujgmRN+CLhBkinlGdbUskAEF+8ve509LTsAfb9cOqhaFstiDOHULBd4L
I7WPbVUJWtGpxap0KuRi4rPbK7vQqvDUbcqjTiHaaL7xN4WsXXixweUHtonBZLhy
PwwPAImIMKPUDk4qoZTUczBv6a6+L2Q3FDIThErEARj4xkXeh3mr1VvWAQqxoevx
UYlP3tDjILP5ojFPe3spSzSpQWHuoRgNXnXQwiMrZMkOTRkKk+F4y58eEpjzCcfQ
6HYxSHAR3V8o3W+7AF7rWqD6eJJE0kcsKvzDN7AhmDYytdsMIvFePRpkRCT4tWDs
ODFQ/N9ZleT+G2GtNLV9hiJ6xh4CPwHemGX6fykTVHj4LEpcFdtOUcNDWXSmlSjO
GmQiy91neFF+i6THr2XPFcBQaR9d5s0ttalVh/5/LULHDqZSBp9GBrlFsYLtRseK
eNj0LGy74ff9IqKvn2jAW9dPyF1kMXBCPGamqqsiLK4xEeju6SiXksGzu9B/JuE6
FRL+icqtw0xKk3evgazxDhVSXUQLCKVClhSK9CjGH6/e1VJrdf0xrBbGQXtpV07q
wyHl6oWW3y+Vw0kaeCBGuS2swmggr331Vs7Aw1nA2QPOoAyCbRpI+7nQu7GymrS7
D2Cav4OKDdn5udm242lYpt7qJpFgJ9e8ntffZghHG3+8yjMNLWYyu/jEgGi2qawq
WkO6kovAWD9AYdHWsmMvabzz9SmUCdVG+X2olczgE5rVuV/lhHHd8lqAIhEtKHK2
eN9j7UD8gBxe/fm13wAnl0fZ+3oScuu6Q/3Hlj4taXukcmmtbu47kp59UP23XPRA
etu/RPT6BIgepofIU4cbEI6yhFqfNJfwpgv5HO77T9qf17swBzPi3D9+AOikIgvs
CzVC5WiD5aPi/ooC38hlOLtKeCMfGtP27ADveoGodXoZGud4NFC1qQTF5UL0i7Cg
kRcmedB61Vbsw4UOTgxA/+jINpQKxfOce96YAyxevP5tquLjUD1fU6VMpV6ICdtF
e8IbnPLeFMVOjxcRWnQ5JN8m9Ade9fcWpEozfyFBW9hJl/bvzJeSzSD8PQmE7b5B
Lo9TjYt2ivHMY6bdXz5XMszfo4oXvTSEy+mIK71R8pAYLn2u4W9C2g48Pe0g7cua
L67Xz6Euo050HU3XcDuGwFZ0f4XpXEMs6NHhvfndkIFCRPpk32GnI087x/PwPh9p
TWqMH9AWULZXv3XGYVK9U6X8gcGAwWLXaxqHrSCJwPDfxMnFZQyIKMu1meB0b9Fi
qwxz/pFceMneWPvgP5m9ogxnszudx5ucCxqMvrmbHzck37H4TYanH1Eamhl6RE0a
GHK14JrLNSlUs2PuAySc4xDBTSDr7J9ZHFbGvTpw6mfzjqf+GpGTFs4gTx5MbN8c
9vKUXf6SmJoOBbHiMECxI0EWO2dWoEcQRBqzsiEppYz+fq/wLV/aVUOiifmMjouH
EIgD3FCXEIWLdhySJyZ+xpkQlZr456kSf3HlDjv71LBWFgEu3IjFZuKwBAUgucEN
NbpbK/bql1D+i1+1nvfJ8GeDmyxhDrgNPTF3Dnr2XOfEK2aZm0Xzili5H++rln6D
vZzMykHPlhre0dgatJ3AEuLMt6S5SXT1Xz/9HZs+eeNLkbVpeGFDzMX5RT1StO2U
mzVlKy7ZJH33ucgWduhAuIl6EwMP0tR0KPkvdX2gCNGis6HWOQK8xsX+hL3CGkg0
1hnqVwtL9+OFIyNLe6cRIUMx5fzK8oSBBnGyMnUEGPDMsDSgwcnT3Bnki4zw2HrU
ZJ4pDSHxr6+YLAGaK9pSFdHO/HCMWHiF9zKmsFITg0cFFpaFCjMRL5zFX+yyXnqZ
OYfX1xwTFr576kn2qc9eC9l+9f5iiwdDju+8atxug6JRoNb1Uzt143DRKLvmTw04
1JLVXX8XNkZxiD4wygdUMzRBx7y5zIGCX2TW/oDmeZznq1F5ewby3z+yQW2YCJSm
SPeUE5F/B/i9ByI0h+YVl5COVFyH2HzGcIXvXizSsRYyZxzm7ISrqhi9zMMko4IS
TNQ9ej8kHPnGhu2BE87Tf51lzCUz5/zeVTPHN1Qlj6z7zr8Wc8C9ygjb9RAKZsvp
5SdcTArKbs3U/LXb53a+//HgNGyvMdNiIXv//mKJF3Bd0Ft80t8L91NiyOHmxW8L
wwcWQD4aq1Dvb6i/S27CnrHQWvv2aWdtKcbJ1LSb3bYJXVfS3GGAUye48inMjQke
JVC8hFKflEOHCyn6HiE9qltSyrhfApi9ijH79FallT47H4ItfANvbiisuPesUB/n
UrJYkG3AVWDeOv3y7OvB2shnzj7nbKvDAeiC9Zl162Xfzju07AnSPs9QUxXwWhph
4krl3HtI246QN5nmMfpfKGWdpgfQmx7BJjXxjh3F/GfTe2C1PfTq0gYUbVd3RXCa
ZfxeVetpStCxEdLiTG2am80Zsg34/9YTZvVOpNHIBYK8ZPrNN7GSWmPrFPG/lHfJ
zyN+tPVH22fbZVfOk9Ct2hKwlQFqXh5xHn5OPAoYaGqafCHxHzc5lFQcPVNwlUFI
gzKV86kqcsFtr2gDp+2z7n8r+tEUHn0CNBIbhOEumI4a87Il22KZCi9N3Ehs0ba9
pw6dSTB3sJHRHgDvop487t8Ly9STqieOpUTK8fcM8UqH58N182zusmcS/Z2tF3qn
t49a0u4MXN9z1pTCgQe/ixDzbwBh0isAFrHC0CrNC90hdCsZdxCRg2/xwPmE5M8U
MTz2lF0AIu28PREQoatkORvLdCE6QYYkJ3Z+mjE75rrx6wEAoqBRez9tOwgEaQqj
kZI6+J2fnxkPztzt/PeYdk7l+LV8HOy49S4QYVHO5i58Lui8a6s7pG81ZaItOJXh
U1xa9+EiAC0f5pWgAKKVjBL2B2GQ9bsmBlSZUTTgQ6Z0xt6X773evXokdhfZy2BD
zvaJysN4cvcoBmK9+On8nOJWrit1vjNIZybfKLovNU4WG7T5KXXdoavETA2oYbLj
iuOJazAa7VKK+eFHC1uutnNAoYS0UKVH4HXG6K9DRLhmlcEUPShdwLpb8N+63xr+
5i9dX+r6ABpaglvy72OMi7GvSP6g4QJYDCXVW87aOZRs1AiDgn5G0TTpElh+zz/g
dIk6Xqa5pH+Z/1RSTeR0X9iP9TkdzFMv/r4GxwsE+tLujjWOh8nqyaHPuk1y0Yup
sX4dmYISRD2dKfiV/0bn2JCQWrk4oU9DYKsPu2xRJxITJ4dRirmgbe4DQ0MzANT7
j10qgd6S8WLxj8rRl7EWQSrcdPRDwNmBoBQLTOm0EXD8VlYHTSbl7baKHUDc4bf0
LEfPEUaSEa4PCJou4JXW7LFappZ2raksHA2PwwmtWnku3v9cyXqCtImufrzPOOx5
leBwsNu3I81nqpHPvvxmn96sNzPeFVwn6S6UAxwKCXntzgGxpreherd7BBqgsCRC
xEtVU9EHEwxuhF1x6ZJHKhpJRdndwb2vSXhOhTHKBbCjfyjGGinr9RawZb20hkpk
Pict/xwQL+mDbX/FzY2HRvbZUj9TIu4e110HGNQDCU2PHN3W2fv9sIhy0yXZnm2G
UP4VjmT8tAxPBTngRjt3ISd3jbDYRPT9S3QVxa4Exmaw9DvhoWCCZ/s8zMcvVJ3b
0VY57EbAxMeI7oLgLR3YvzDeYEhjvNwSpwODHyShMQUn1RI0SAkvvoGIq1J25y5i
4TcJMvH+1uqLSdcXKurUee9Ro5/csS/TV7rmlfNSrfpBpN1xxmr11xkFL8bcjvsL
GUS0hJ+XDM2NqeKPeXipDY3h5UZ9RsGDdQddrO96FykhLC3vV4ueb3TlIOJMfw+f
Qpey7gkmHEqxmsjTsr6cYqSSgAK7unljTb1fk0aEy3GECxkteOvP0r764cSCi7fQ
Y0kPIqJSAf0z5CCDUWsestheTI//EJ+zVHz69GpN/n4wLXWCYLih2DeNg+YWLnDf
oNp/NUTP/ZvgZcKR6+kWsKazIJBa26XrjeyL9/FGrLgvakMYIo+/Sg9seBGWZd3r
wv+JWQIOj7b3eaeK/mOf8YayrLZSTUjYMP0ponANWhE8pG1kxdnqjY9O9kLWg8yU
bcALjkm1QfPRZbh8g9L/9u9mSWDlEYry9+k2Xt8c51RsRH6XP45cj01i74kQ2Tod
CNjIvBnbKZqlsD6nB3nOJqxJ2eBgos2Nlj4linxqL5lGEPiMWyYITtQxUD2olCDC
S1w0N+I8dbAzf/BOhABtAnbaDxqcTVV+gENiDTjTzPp5tWcNeiXG4bzJlUP9W0d8
A56U2MhP/zu1t220DHeEyT4bYX+uHgQkKlvy/mYEjpaUpxUBfD4usGCvlcrwvOKL
FCqagvv6bbA6m6CtOKYt3hOX4Lvp3ezQL82pACxku7qSeXhHCPFe9XN3QYT1mt/5
IrBDvrSmJhkSMixduKCErXlE8faIn6X/kSe32iFKuTtK7TETQca51cq0iH1Ls51o
4vXULMb5UmhY0qhpEzKy3Tb1IKHw4Djp1G4QtUUzKkAvpQoBTOntQcUISbCYan6p
rzYS++RIUGLASd60dRJt27g6sOsYdCRBU1EFI2/YyhxW6f52Ncxv2XB6nv6Ch3MK
WYrzuDF/Ju6F+EEX2maUmlOsT4urTcsObQpRxv7qWBOShi+N+oy4dMWIXr0vWa9R
YSsdTAuIydSZ2xoftwpRYiJZe7826kMSDz1+n2m70YLjsi88H/Ok+in1nDZtZdiL
LzUvJTUuSyZzqRrKc9gM3jVh8gSsssY5FKvIYQ2zUzPowh5T4MUHPO6G4D4WYiUq
LuyktLhGwrNJKUxODmARx9RTSYcbyCDP74sa4ZDt4r4DunPlEZb7qjl2fxTZLgwU
pgBPhlhO6aAFO9bp/iBKkUz+12L8F0t2AFt4+9PmdCOcfMOWeAEgIYl0+vP51ljE
+MJZdubjoG8i7l6IH/1K6OQmyEv9l+nvGgenDO9NRhOH7HJcmMvFw9i2ZloxLe0l
/HVCm6S/oTp82KJHMCbhuHrxrYRZYSJO2Q5iDlHScgR+5QaWkny/DlrruuGi2PP8
3WgerlYnbCRGILX3WyCb8JQP9Hei2kCjoY8JddfS7/m9LLEfo6RRcpBC/mf4uRNR
M/UvylgKMzwVxhBHvCKD1HTvybTJOc9WgL2r+hdZyhAy9ltA2j/uHyAOF5CZJi8p
u8jmqYErahz0R+zxWK2yWZbkGHfkYtKSmR+HC9jlHilG09NEySfFfHSVPweBsTDu
qefyFig8fu/ZEmUmQ7mtJrZvlFW+VxT9fKGoNJdsnU4lyrJJPAdDSpJTAljd62W4
WAFjx9RiiVkYfBsVIXNRAQxWFy+endGRFetuhj0mn6rcZ/c5S6ajUebvOr9pidcf
ngAoq8FkIYJwQ3x8WtD5YYl+dTjJlODEDBm+aENe2TxsrSRKv6/LaijBPMVtgh0z
3Kvmlnu7C/dnDfGFXqJmbWhaiqFjx0zhU2G1NygfSEn8YsFRuBcr5LR8kOod4x10
Rahmr8Ty3Vn0TtALrl3SfF0FOsQCQ9RnmWDVKb0O7RU/1zST2Ws4TwO9aic0/Qzz
xN+XSe6MLrzkw37QnWuHp8Q4x9TEVTJNLEdNEEdBfzxIKgZUj2iMZXcFkWEV0DiZ
aMNZh0rJ+Ann6s9xuSFkazsUDvRq5mmM3YaSQDKMItm54ASVOzoL5EzDNKiib+IH
QENEQJXTSsm7ERlf4/y6KlkLlDPRGkGRImHMwxION2zrg0YiGOHxt/+7f/+xvVkS
7L3igFO2WPEIraND8ZmfWhyQMflzm0lNl7P6Ug9JiOo5MASrCsKLBSPnepocxHYU
2rfs6pvWqjAK/eipcNlGe/nFxd1+hWky3ZEkkWo7YyEkVVspsSdrh9S2Kyg/XdUX
ii1hqCU+LoQidhu1ckiNNnPNtTGT+rfe+fs5y+itYsr3yGeL+d71rh3b0OvY3hKs
WRGy/HfCF5Bqo5IoBg0IgcNwD1s6a7McYowNHJD7UGnyKnJ3TSre6n1IAgnlT4wn
hmj5dlCXactlTTDo9T5U2qlJL/3VEWclVVZA6YWA2PPz5KHOYiw8siIioMGUUK+f
bPFa7LgkjqbyVpaorrEuKTpQfuRjbjnpn2Zd3PKbtkuaT72UXeeIBjByZJNAVJUS
H/JrE8dS/01Gdy4T+pqwwVrYLzHCcnNTvFNFV78FdsdL9rKSLlZeLInGTnOzNyP5
hfcumaXiaCsrSW01oNpv2Aj1ij0MDyOEy4YXYJCvixt2tWe/2eii4f7vovO1ibR1
ar2sJ03XRpp7p/RCdqdB4DM6BiJBspM2I5X0QdVWSmqMAnKlo42sx2tLtJRB9P0H
OEazBOQgA73G5pp10NP/aRrYCn5qQpXt4zzG1OXII8TaE/uYiIlZ9NGOjk3ZzN8H
iv9INbMq1IghaY96OsPkwUJyKOH2FuaDvS9rER8gYeb+dkhZEMAMCGB+MahuFzbX
Ult00++bhrRowIoDSe0G7z9Fcd94b/keu1QmEw1HWm7hdmJECsw6PJU4/7FrfdBO
+w2Er5ETGM2I9NCkDdhJwIm3wZEk7yl89mjfs+FMpe4b67JXiUoxQP+k5R+SC6tG
grw8X1zbW3ObTsTbYcQoGZTrAA2jA9zcEBpC5/0TRHMuY+rfmPHkKweYzTY0U2oT
folf7GY+8sSgyuh+LraRuZxmuehL3Il7Q7Nz9lOQOz82k9+GDgVx5VPduqbDF2w5
4ZQXlE6f2+LDv7X9TZykNfUL6cpuCFO4yuzGtu0/leaR6DpjPxkMJGJ1aNpidnrj
cWs9OWmRIJv/3OCo0nFmmZh9wrCiujiV09AuG9St8SrWvsHOk+bQcLAFKYXyzyav
WaxFMPM3669AwaMmvh+JAvfyaQy4NPbYkdudIPgk2S0XvzwTwzxzDIu2T17OFEDk
dCWjtpecVhTkgtHNBuyzbrxU9ET4UWvIx3D03sa0aWi5aHEVUtZNym8q+tr9HAag
azCjHtlck9tLifL2AMmLT0hw4E0sRFq3/QlGnBBSdcDst0z9YUlAlFmogLx/g/AV
Ih4Zz3CnT3H3ba4MMDosUE3ufyBjU28bWjLrwe1Mu6Pw0lVohohklLsBtxhtevNq
U7tc6OmUmOe1HYOJWQzSbEZzovx+s4BbWYBjPtNSyMF5zR5hiUi0HPAFODLYeyjm
ZNXlqm2nL/KPXTVxY89QaT+uVORmcqkyY/NZKANL9dh1NGK/ywDFOFy7NgG1VJB/
9HMIjkF7PBPWpDaQRbxAWylxwWNpeBRtTW57pEBnltILfQTW/zPUtJaPxYouGiLK
p2WtztJIZXiNXSB2BAwtOXwQiqbusvKpGn3wKVualcP9t+KlVOFsg/EnJ1lrqeGb
iWI1uOV7Sa9lMBX0HelfZWa7LXt8BcacTT2z7lfYSXAfoOkZ1S8ZHCZlZ1yI/WCt
mLTxwGT4ECLbzBN/69414jxMszVQVE0Ufg3ZQuC3Sg6z0Mzj4ZrARtSNg1l3vLKb
6RXWxxxwfNnUZT0E+orUXBnuh2P0ikMQnE4n2y2dJeUNV0bT3615ZkkhexfP1wx3
tN2VPmlCeWMkqAhNCPzv3Nk/zWQgUHAxBt9kD9vDrYg57csLVHAdnfWrPTMtG2MS
J32z7DTija5zlJJhDwYz9fnHWrRbLxWN0uv0erozuSV5fiMsfjrGuNcXArVwclvO
zSsET+yowJX4D6qRRPmiNxcWm/rgPWz9gZQvvksEuiCL1yuDTooF482Ir/EvJW8X
O0c+f+T+nz66lFBSOyRWy73LC+KpUC2hWXLXeqiU7cmapVuhK+XAFaAE9JQKlnzM
FtrgtNW3jyvBRtKmnpf2EPnj0HT9oHS8Gz2O6oFpDVd8ZpsalB5/oRlLn1E+t3BK
Iqf2Xq9YKzAwHmnHYKCPeg91jgFIDOEw4YBAD9lPecn+1bnQEJemU5e0mtUw5NcW
ZtUuklE0c1VI4usCa35pWRtwuJbCDmF9Fy7g6aJAP0Qxb31G1I4UU2H4I8OnQYL/
aK45teMWmnfflV319HI58e8KfoxrCvBsznjmQPhSsuB+CsI0LTe98WZih0xQMXFU
hC/ArPJeCghlb6d8dR0yz/MRoNi6P3rVbh4q69+QvTtYG5LWfA+FFDKSmo6vHYz5
X0ZPPBbkKFDW5pOnkTcSGZUdK6isUnCynTqnf98dQy9mEh/Aoddz7kJSKO6r1jjK
jXque+xPmePnxYYIEML5unI68pxLVPCb87iGcPhHw+aez8BtB/SWu65iPqVBEAYt
cWy3M5l35oVPEpduumVtLef2ILG7bus96eeXF5SmwQeC1pou4BVXfLYkFockj9Vv
n+j1iHD4wOCEfxDsq+2aCutMaK5D4lpGWwBCjSW4NPIeerrOSt4thl2yuNPXosE/
wbrXsw6zqDneorYi5YGkUB0+Z44wNOAkIbOK+eAoc+Ls0M36vqy7HZTb5ULsdrMX
BpkziPkT3lxGxA49f0huY7TI6lUA+gUyYZV0y6QEqZ4zkmTE+3KPc8HaGxN/tEIn
xtFS995txEFHUMq2GLH5TtvsuE/lIcBQx24789fGY6e+5pnT/asl7/sxOdyYPhqr
AgMcujaZ28MyVt5Pp5NoJuUaetVyXT7KJVHaGi/7gmAJZbkI4QL+8HwLwmxvQyg/
AKwmpEr9HevYfnUxUU+3wm3alCcc3FWEV2RrHXLyDzjcEZPg9kIdEm7dgb48fYiC
VFBbvpzVwraiWnNDQ2gaNe09oG8O5Xeg5/f1nMeQlwOiz1I+5D+A0OBwDPaVP/gu
MrcR9zt80QfO3f+HIk66jqBsNGPBLoGCK+vJNs04ymc6Tifv6zVhFQuwlt5QjiWq
UCytRmmR+blDxFF4w6kDFZ5TwSAnI8ZFVS+EXrVMoJu9Z1bReJubjeVqfqmqNRu+
4ggtiYiJVpStuDD3X19tjg1QjrdZGKzasUrCwxhtNIsEAwAtNkCBe6pvkTBld7BN
e8LPcyAXNHOr3wPJgZ0hoESs0CviwEeO2vhgoERDO8sMJnOCCSepioo/o+OPN5yO
C0rq6FP9LUeF+k2fKgrOr5E+uPvSAKE/7laIQbwsImaVwSiCyRM4dZWKulO6O9GE
hUaNDqD4muqTC985oKbHjZt1raUMyBqpTO9/m8+qczgtUCsELWyVAr9OVT+aS1cc
WHjqTDX4a2xFwXyTDxaYXSTFTi88WEjyZsxWV++NWt6Wh1AP/GbCXWb+hoZYzpLL
XRaMil7ZsxgVnRJDfg5vCEXiJLhApykSOCqmqFHTS+e9ms9qCR/kH9nNuf5xvcww
c6avvovM3c/czSI797SSECpZINNjhykwvgza7MlSStW6jNoPJaa0bqGU7wswVA/s
wtXzYNLiTr3LKN7/Iaf2k1+C+Id4awaY9CxEesHz80ziZFLHdL57tiFRHf+7/bFO
o8PFm3bLXe/dktVlYTMe4pFzq/UQPAMfYEQ05CvQhEpKEwdvmotwP0vlUISNOc25
1gypUTnX+lYtawhoqlwqr3Ku5iPSXoiSnZVSCIq4kFw955o08ZVwBch/jgnBp+4F
VM0BYNoOIwZyu/iriskzKiMpCApN4osMR57vWZKLmoDLXREx0A9Uecf7FVXF8mI1
TCSpaUV35oc/MkKkP0EiTTZ2BCtdeubQ2UrgrdYAIAMrlwIhYITozLw6x4VJFPJW
lD2JwLVNPB6u3TOtC00tdmWLhbdJRP1VWqIlNNN8kgAB/S2ZXgrsBu7eXCzY/bc0
bMIlVraGItV3Il3Enpfn3zcxuSW9Q7InQaM80aRjB/9vuH0pP1SYCCiUXf57GZT0
V/HAXkfuncENufYJejos+fSVV1tUUWZzST6fUgHi6vTUqh/iVwH2zoudal585fCW
H4obshY1UHpxfQwRYDm6yumZvFe1WMAwGqtIsq+2sqoCE3nG7skLAbBrLd5oilx3
DhF6M4eui3O08n/WLL/dIlndufJh6b+gZaDVd8WH866m4AzCzIO95RCOViup6Mgy
8b0R1ypi8xIjcWrgCa6SnltJSFZLrI4aG5nbRZf+k1Aqur2jukBlQeDKXdbV7ASY
ZyOpoH8Ti7VBrg4gEPM/+WUKDcJGeUandeqiEtFdhGjtZyIOUNCl9/EEw1UuibBX
8T3PzPPLT6S27f0HC73HpnrSMxm+endSMIaBTuY1vMQ8uMN0FMRxKWHgYTimlu8F
OpKVicK0c1seqLIvqSspE6MO6lZ6VrlHIl87Z5cskGl1hmX7MwsDuu9NrdSyhFpb
5jL4f0ssx8oEAxcrIamgGeV0OAsSjKNTcnbx8IXWzPCN6tIHeJ56OQpyB08SZOD7
V2nMs9/CMhN5jOD/b6KJl4w4WQwre5TYRt+8xdLsGD5haV8OcteftweZksMRXTNS
KT3GMf7NH8xn3aNIkf1j2DOeS9i/Xy0tV5ATyouu1qvoQ9ztlHAKNBjP796C4ib6
2zH5t3cw3g8eE21tW0nPCWpezaU/AXBbu9lbhU62rs8c/674q4qdIwDfsUdydfgo
zmtEKkwSfybR97tRkYaHwgl96ywdD5TUa1SZv5jdVl7QCA7oPk0IO4XEDBi7RSEy
tkygpCcHHT/9/MIqv2IPYaqfCeZFWyMYXj3JsUDsRNQTvuI+4sSdIdbO7sKYl/fI
rVo2PxvTeMofnE9W00RzLE4YUTYugYLjDEXvNyWBN5++S839VUqRkTGxQ/4izSMS
zmI73oaLg8pqTHQBwwQGD00rkqvsb0WT1Ylz95cdqG2JnjvVCj1DVpsS3LTVz4B0
sPJwfHx7BewxtTzLqqYZCNBsrs/equFRHKBHIaD9VbEcvfu+tdYoQb+HIHzJjoUH
zjikGTIGSlcH3BY01glxuLJv4NVzU+qhZnr1+VQkChJIAq8i5VlNrqk8TQ64e5eN
Q882f56oHD7q0m2VKwRsUCauSS8wdaFzTN5iVko2rq1vb8V8IHrP6IiXeEIA0Jyo
RJba+Yb7do9rz7B8/PDnKqvYgya/AaOMeawtD3iEphmxaEW+8I7KOOxojljpYBg0
RGXjeve51zEmfHYIfech4l26aYhooHAW2hiFAeqU/1GK/NeRVEt7i4lDu+Cv7go+
/Pe0nmCXbcn4JlIVPojYfp9Wx6BRstbLxJSCQEvqX0iTxKHQE3tmGf/E5+4MJqXz
mZwPV7LkI+wmAA+5d6bakRXH+LMdpNpWtLHWjCzvSenrOwHjKVy7B5m/IXhAXKMM
rrjFl+vtvMCLf7Mn1bRhCzinLCoX1k9YYcOFSxeTJN/+EWID2wDyr6EBrTvogaSO
rVr9J7VPdzAnljXv2f9cPzqnMtRLZ+YpOceD6DKUNpwi4ZdKI0/AhnOU5D/Wrvn2
SUpibKhvDZalLvcf/xbmLiG10Fma3BJFaE8TU4SqHr7PPiQ82+QwNtCsKUw+x+th
Ra94vds0rBZJZqZTi6PHe7E4upDaxV4uBD/+1S0osoSS6c2v8S3D2xPoYqXvifsC
rPXPyUHRKPKODHiiEcccx/SOVNKblFZyt21CVrHmIE9+NzX9e0ho84EQZAocmS8Q
HBxpgrzge018pXKrKywuYuexjPJB/dVVfn3FCXRxxBf9g4nR4lVJ0S8bS5seWBF3
KXpfZ4KoEOz97VahdiM/vTxvRwZTAo1Mc/1IkrJCkbjeanooBHhFWmX7dFyIgnwR
CpdV2k+KIlGpXzCR+gXFaxJnnlQAijsVD+cooS53X+K+Bp+pqhnu8U7z8ke4qB9Q
wBGwjViBNJingL6psUcBtG/8BZ8c+FaedmO3hDMM+/PFhYOaXitrcLZMEgV6ke0O
HWcRwonK09ICO6SghBPg5SrwexEZNlTIYn6iy10iDvyg2uIaA6XV3libXGdeNtK+
JX4bjW6uji3VWAxXd4IrWSFyykemuTxmJ1bgL3J+h3AVt5dlzg7ow1Nto7ShAP/O
8CkqUb4c7z2N/k9N7Vqs2bp4eZY4TSxo6otioM4rHBbOit6ryrpAwlXuqfgFNHKp
ydgs/XKIh5F6ARQQyi8HSvabnBu6e7CbcBHgu8etULUNapXu+oYxnIAEHMo5gDBZ
T7Nx95ipBcuq9iI3YOVT2tAwdHa+eqVVLZZaMQMZqLQkPtR/AzfZBwR6mG0K75At
pkPseEcFBpf9Jyll6T7tt7e7esSJ/HJRf9SC+a7DjrqEBk5zIRaqtCEhMg0IFY92
+Qj4ay634SsoIZMBToNfhlB41Ib4/mQXzEjyCXpkn9M8e8ir7TGSCugMk1ENUKke
Eq/FVrVFgCxAtPUqfL5mTPwJpdGGoZ5iDRaF6VRUaQjk2RU8NVhSaHVoaWK+Wx8/
LjijZkPt9Bp5ieDm8RQy9bOiBMClGhoB9aLGPhR4iJKpGt4dMMIUJon3ztzy53iK
K0xcm2jTDTNNn8z8KORIhNW+Ij/GwICF5RDa7vzfo8xkQYv/cqS4JCSQT5xeBVw6
sZRfNe40eDKMY238WFYjqAFS5iUxi1VDMvP8xTqCOCG5aN5cxoFFHHZUmPb5fVEw
c1QwHR8ZlXDdO/8sGWXc5RE0PqAjPob0Xy0LgU9vB2dc9RDEuilE6771saOuU+ap
P6Pcw31nm6Ct5H4P1iWjjd7kU8JFGaWiaw0+JGaOgDdsUlG0GP/mIFs23DtKuLhJ
5BiNBIx9qdI+pSyTEMVMraP0Wua72yiIkzsHsvjeOGygH6z3buh/Mnl75MvB3Q5I
k4CZOahIFjIptoEvyA9Ixgh27SX5ZpYZx3mlsFxSgexjh7vypZ+fdrD4Gybw+pNj
wRjzZwYXI8TPq1Ad4ZzJZ22nRGLdyVLoLHMOFi0TDmF1rswSHAzjl5Be7rJ/nCoo
68vvb9D1Vt2paksjhnJ9CxudI9qHSeaB4Xs6ngKLdkf4d59X1toK5rZ+yWBqbnGy
tGKgc3WPZ77J6DH9G5eOS4d6gLxb+SgFQ7a53szuKf7MNDfZXeVcAjEJeLiRLrw6
rlq+WBFTKkWS3L15J+ghTZo8rcin2gq8wC3xl6WkwC95LQlV8a0ZZO/+zYjovSYn
BwIgnzcEdBB9VG10MhFu7fXuTObELWCZ2Nb6ur9x+9OBiH2SLvgtycPDfKVjXfzg
UHT6Tc8PzEh3gmbHwgTsRwMViH1A6tftHN4Ti0WXtR7DYr7bdj2L2+6XjpaJATV5
BgffmcCp7akklB+YSJkjK3RsOxF+5gUjngSpHHUBXBlaENG8Un1vprfzzP/Mqi2Z
CuZUXij+QLpLBY+4RAxdLzRkbIb4cfB4IhI/6rG0x13QelDTPUDXCK3Rx+jObEHQ
qjsTWFdzXX5h7YBiT9lFcPPbxgcQqe8NIBU0+YAUOStR3Lh2XfKSROQVHQWQkc5t
OR5unXnD4KG7+sKmlyQVb91XobzU0rq2GPDsZXdzNVJri4SOqhfvZsdQBiFWVIV9
M/3vvZmwtP4WUtsNfqqdh/QCcS/ESwqtr3ZTAaRJabryVPFkSU8QZUKas70kyI3F
N/cDDUsmC110zNcwWN6KxcjTBfg3iCSt1KNNGM6YMffiYM5eOwuzhxQmjy3UZ8D8
e0qYNAs0mXaxYY3iuEADkMQeTU8BOL88kpSKmaB99gEFPwKPKpLsO2Hz87QUGwjm
2kXh8AOuUyRftPva1D2GmGY3pZv/BBD9OE2P+njmA+3AMpk/dFmGoJ/K+HnisN4X
4ub9SXndH9R8sr9XpmhYqXPhMVjnjeARzQzsoj00jYUcLg4Lt2wApGATOUrSy4pJ
7Lq9yafJmH+0J5ZbqFFa7ExfLlwmk7zI0ctU8YN82d/cg/MCQG9hIZGJ+jdtPvFo
FtH3hlDjocp5Qf1pr175zVSSeHvpnWJyBqJumHCY4yWVSr6pYSInco/iSnLLzcL6
35zLdMNEWaojpqWDFhp9/Fd0QbtxDVaCZ3FPPDtNOHrgllqK7jtmTnJpqAx0DL05
ga6pmPNkaMeTltpZBWsWQc2joc6Vqaj5TDpxX6vvFjjI74qMRt6oiXwtxVBjT1JB
PwIJN2EQd6+E3kEB2ihkLCyKzMv6QZAlQGRe0AgxWHJaw4qnnSDNlQsS7dxOOSHO
4rEl7x0ci4spB+skQHeng7YEBOb/E7IsUycO7iZUP7HZ6OOrTVXdn28tIdjrPiX1
Eiv5zOPxuu7oG7NllEO8mflGZQme3Q39SV3CGQypIgprEAlBwMl5fnoQJjCWFq+g
NVCTtqT/sQgtmbJh353l3+ubBFSLVH64bbOYCcLBDwiS+NIoUwa+LcyCN7dp8SgY
ffeBQivFSOjlrUdLYTMWtu83wd3hsgljL9Gv1kXi1sGdHIklVWE4fi+1Nr8PLmqY
3bldWquBBOptQJydL/KuphHkcCl/Uc6X8S86LAsGb2mEwRJnbHiwtUTcDizAwq79
96GXRseZdsxp11qea8mWE4RCboZbE2zTCu/BnKfSfv8XjPnLynTVEvh9qmnSGCy7
PiWXj3rgOfNrrB+rAEa6ybhFErVtkg3pi2s6ZnMfb7D30hH7CT8deMPQrF9YXChS
DUiBBFcPRxg8IrBHfRNaDoMISb1+xSNyB692m9vzZyVgJ0mfDlzFg+DDn1rWLhfj
GAtdivgUkPwFMV3TnBrEamsBQg7UuEmjBQh/BJQNSFzcQkcwKzek1woQyaZpX7Td
jb4xxp0Rxki9cie9q8YHq4gv4wsasuN0ybomEf0Lumi3QZ/BTXUjfSeUUrOtux+y
YGHD9N9lRTTkGxJdIT+WLREBgvW0nsV6XkImNAkWFhahug2sPuM+BQGoWIbe4ukh
AxwOTB3U6SPi852OKd0pQfSoKH7HFU1mwxvk1fDkagA5EP/WGK5d5k5yaJ/i5b7P
WgqAOyYWP5dh2qJCHI7Yy09uHD849njcixQBWf/PKu8M95KHp2XMnESc1UkhfRhL
2sGpNOXnnaAdJDT669CC+a8f5eMsM68b0A3qPj9x9ZsDxEsRfKdtbzTX+nF2sH/8
yMeS5IHosj5ls4ddmRggEpeePgqjvcG8ACKtN6N5SIPYbsm5Q237gV+/aDOie+Pu
Aodl+NC3CJJSIOLz4668IoKw+7Y9ML9madx20oTBnU1ozDsa1wxtY0w/mrUbMb0o
wXE4C10KOaLI5YWmePGe3UwKvBOPPgjiiOvFgZcjJoUc+ZzVgo6ObJ9SMv7qNS6l
DftFJWgeOc+S1uRubn3rZ6c8lVgHGmQc5QbgbexYA5lxL4AsjMlEotb/HUllPMqo
OkhwflkYRh/p0Dbha5dml7qcG0ZMUDxlXzT0BJnmpYpAh9FJEkEoZHupb2U7WAZP
5JMkPrBOSCoLEJjyUINk/9gFhAjV5yNTdO327C482iFM2NGT/CCNq5wKbaU6o1xP
ySB8J0hWb016XPRuXfDhGcg1Q99zmbntv7rId+sMeQ1U5z9OZrwcXcc/XS7ID8xq
eDXh83rxXOF5rsu9lczKqL3s5rsjgyiY2l248Sh2Ipus1DeVudfvr4685I0P0GtQ
HhYGhvf70oW+mRZjwRCkpcVOMYU2OITuqiIuGlny0NW7AAGVjlRbnyQGFlbRIta1
ZuVPlk4sgAjN6KTxYl4H7T2OJsmX+DVOP64pGsua0TlwWOaigcODmS0dIb/A8Uap
wMbtoKBKiEO2Hx1z6hcJF971hEs9nvQQrkYcWvOYGGD0CZ3rta+X3jljpm0PxfOy
NAF1+aobR8juEfRO9LimhUxoFDFlJeiYbUUfAVTJIMA425BbptbEJmRxR3zQqqjd
R9D+tN0NPvlS5r9oENep+lDBvQxXgtOitOFmMYzH3ROK+ckj6INxl6p6GI5aLqof
OhdUZtR+qO05ecc8IuR/97SPCmC3m+1krzhfkvIwu0ayaim/p2s4vC4HTgzSCAy0
hzMfUb0UVrVVEylmXBKwEF43T/D4nePuvk5ydURuLXHr7CY7CC8ovfZh1R59G8hY
SDIPVRS+BDpZQqfvwYtHwN7dkEaM5wN+K5FRQP1uyIAJexH95GGJl6CaW+Ul3WfH
yLLHahZF06/YkWCZDvvrpepM+fSxSD6/kfYajXADC/Sx2Qprc9keRt55+qiZD7CT
W1ElZYqOa3VgYgA9VQ8Ems0FkK8RunC6vX2z8nNG8CJkLaNvYo644ofvtwDWdKDI
hVXos69Jy4oPiLD65ncf/WuajQIc9yzVrGuhuBFMvnvXcobOhTNdlI2o/7I/LES4
ZIgAJOzhlzrEW7dMmB47BJar4bKBQ45S3atefG+RbXc2hHcwmMD0pddi5OJRCwNV
bi3xUIKNUhXZV93qnB72VQfjW+rkZLZWvWnsDmfFiNvjvitUoKdnVk7ndg22Ovbm
r9eDypqJwQ6M0gGE9gWFFcI+fytCocMojjeKBwXzKF1dnlYWN6d8hOBnIc75aArb
Zb1KDbQcTSTo6l8L4W+vimhKU7XOfpN3MHOp7/UCV8AQanqq1OJ4z3WATYqef+fX
7gMzrW+byIYO2NTfvwrr/ORfle5+lhjS+cJZX9fABjRNbh7575HURgl7fPXLEHWp
jmBBFdzLvm6bhFI5FMbUV57TJYrWyuBbO1FjlbCllAoSyV6gXOgpyvE3Pfr0PnWN
7hWopU+qiihIUGSEc9/58hojXWkBuR+2/hxQgw8HyJb3R2yDkl3pwnup5sKB5Lq5
YaVb2hvAIL5U+ys9gVm/ODqw0fMFqMkwvY+8a5/SZFC21h4XVIeDGUGnqzbX2ZaZ
3Eq/+uGTWgfub68q5y3P+wqabhQ+kvBVBcNDZ7AmpwSKnG+qbnieXCtbbGfsrnmk
mnYqsNDVNf7ZvxShbJgYALwfX8BN8hUWZRL77k8+di1qqd/0OhEvRQ6DGaak4BEf
xhtvDxyI4NnFBXi/mqmx3cV10X4M92f6DinAxWWO5GFBXOM+LSjorkLmHHqYiLRC
jnDqbmjcd4XGeM7VqSzOETf6Txu2O1J3qS523d+FMQyEwA7y6dVwZEGXM9NN6t3e
/kfKPZeObC8JU6Z+5ZQpIJUa/K970PTG9kXKz4ttbkwK9hl3S44AFCSB5Qfsa2XZ
XqWiITQxgDfG8i3c9ElUMNyq8dMkCNeL6YiZDV8BY7vgA41kGinKmefGpRm74Z+L
iAswW6DZEsBhhiL+IXwVN7beREnHWeQdFUS4gXdGmgwQNZ62YP2NaSH4YcUF4DiB
6dwfowryVuophAzzCebXdF/H5tPXSHhJxuKgn7vJdEl1eIYnVIOJdaMXAhQmYfWW
Yfwdda/CWUR5wjAys5CqZAkyx7b7hPe3FFuGY21xE3ie2EIFsbh006LC7VaPGO0C
Z1uQ3TQ0r9dUYsSRe94hpYgKjs44aKcnHxT47Au72fe/aLk/6v+VGi7FPOdHAhfA
L7TQ065LUJLf7L9iLpZ60zGNpaRhvy42lPjXYdFCiMHVP8Azma5KDptvw5O0v6Px
Q36QlVR+X2cz1HHXTP4xsECFIwn1gTmlgGxQmC1VkvXuI2ZLmdK9cgeHDe6ssooY
QupL6Hg56y22H6XW78CzaoRPiZ6PGD9AjIF2xd8QBXyzCHT4H5jKUgqMmHxoUfPX
fddq7aiSstjs+fF5gmiUs/3RvjFnJ3b9Q+3BM3ppGGCIqCmRUD105ZktTosdJ0Pm
SSfg7Vnp2z7zaABDLeNdiETNK6I7sdgwqM43ewnY1C/gOUS4J6CqjK88lj6rBQNh
C6nEIOl61t4irdPGGiJozOBgmErar0xQI9rCy9RdvzBZaSw5htsPaotF2B6zLwyZ
Jdi+ccYdYILkI5p/B4XFcjsKP+jPF/FpGe2BnEfzixJWNMmh3sHob0dU/jtdN9fE
gS/geuxZ8W/iJ4Nk8oNi+1mI+YeI/sDuG9fuBEfCDv8GelSnmt9GqUSJpMMvMrsV
/JS1lActL3JvYbZCdEVNZFfYd8IjGRAkZKl1ZYayg/fsdgXOHqBbhcFLE42ezeYf
38vLzWKAc9kbemDG6j7Eqfnkhc0IIkdJ08lpQhAIprVIHVrPA/y0oONSWg0Y6RpZ
DODo7CIvUdfNYvN1C5cSA8XevWnCuUgZjcgNxSmWj/A1w8GTAc5eCvW0YZjnVzyl
DlZkGDkKDmZiotCyIo1YGJNwwtOe6I9E5qPtPhShvcKBZLcVc54nufab7/0uwYcX
JIQf0903j2Ynw8w/PWEMubHZuprYAO6Iwrg4kfjQfIwEcgWovHq7Z7ItLsuHsIRL
j4ouImQy3aVvOeZVpTSCAogcwEEZjRY1fQZiMmTO33DHiUOqorhp6YNiukqIHgPh
FtVE95dxfxtjQ/5vvk8VcHWBt5GGNCWKtvPUBMbUyWxqDzoYVB3mqAmT6LBq99Xz
7tww+FZbMJD9viw8EhNd23AhObYAoWkls2OIw+DhQ4RRMHi6sB5phUnst9sEH1OY
1t/HcAqgq8w+kzPmfzXRpAithm6/G8919RdwYRlLAvd66MiDPgo8ANbkbVQemDKZ
PPNcz2U+Yx27Bi2nd+azGFWWQ7jyOsBvUPjAZTz1/Z0k/Mj25bcU8NZmV786cIr1
gFEiHbEu5Y7pV6SVuiCQ5lA0lBJ4CCbq7ONI2N65E3g/94tmDwj2wF/JN9/ILXqO
b6ppJ3wyg0viEAdN8Jqq7k4ka0PAcDBJTDhxeeXxGk9YaoU13sg1mq11a4r+1190
rJfs0BzXoUKRZ3bZ4SrdR3KflO9DIuVKIRPCjW/IHk/SoY4Zrqti0zDobVImr0Bt
BpksFuaqNbE7hwMvpBASPY0Nu1GDFMzNLXXn5mR35Lga9BPjgiYwwHuuOjOJWoas
PgWBnJEl9nkZxDv2iUZrW92fCWZQhfip9zp5CaMFiSH8NMJqjaEoqThovwJlrQqH
Cw/R7hgz+FuFj/vbW0oqEuVv2+jBW5LPQwl5P9m9CH8HQcqlT+UXiSaSymeV74Ve
zlfVUq/vTz+cW4fEqBrfHZ7F3QAAvWBhm0HvtfkJ90xdNzCK4xxDSU3UiUe90Zls
bEl2NtjVQpmVqmQ8EM4mU3xs6yn+Egruv7UotCXVVo1pPxpuuBWb0IE6bIi+nkNW
ap8WpY1MWUeQ57B6ZLreKYvOuX3h4tcEiTPEeY9B4MquCSaD+j5DccvWtA9kZ/S7
gqHpLXjaOQWW7XYtu2Nd4KmJ98ut/ZSH4KGwZgtG9W1R0rRzcnRhJdXEdvtZgA8/
O8dYZJnBX/QzLHNCg+6KRFLDefuDaS1AF14KGs0LOlqjwCDAEs2az1wSIRFNUoNN
pjjHVsvP3nsOT/uGPUlFKQEYbWVcVAvOP9tbKBsVxEdB9Qrqqazhwp+qtHeCR6JH
LweE+ahmBmK+gHh5eKQWYXnlvxD8lMNLcWqBAFLDyt4/A8BFcdvTQWP4HSYrgnM0
m/nqg3yhaE0JMJTT4Ggdwkl1aqfKQahwO5uSf02vI/Z9uV7OB15rf/dF17ATYIxR
brnSQXqkCiGDBX00E437v2ZN67h1qn7wWoa4ZHdCsubPuH4oxfl5Uv6sRYBheiFb
0gNWKdQQ5SoNm1H1j1w+i0hDsEXTpvYf7iNH6eHTssVte3rBNEWL1vKbzLfMad8k
qW5niBSd9ffVT60JSIN4Fwee0IidYt1RLpi2xlgVXjM+HbgoNOvmtSy5+RiSwBmz
RA9mJxlp2evcsMdIQ0TDNdvXZk2gwXYTq8qyU2Jo6rlM3hIJrx1apxzBmZQJVH5Z
mLXfoLZcaGP6Z4LMGe+gxYmstBDggwvQVfeqTrejoyoROrMP0Bte2a8toRWXQB5m
ipk5JyAs6lHSg3FIOBTZnzncdR7hSUNu8VfG3+wMERWGUuohcmxnCEjWtWw730zR
C+1NokRz4rxkTWzt5i6NxgHDZidgKe1t9RaR0wjszCnAWEpI2Y63AKDs3i68/tQO
Ml2yX9Wos/s0GeAcQselcHjfQaeOliD56o0gEKaiF/Spjjp/oJffBGUeDK8q38OI
otjDYx79PVN4bpc1gFwXHPCEGXcEJOco2rA628VX5Okx6Cttl+9PKaUiMY/23qmu
g6smmX3BrA8Ov8oahtfCasiNOJ5SdF5SgRTt1xPaW9SX++mikqEwHHtLZ6dM+9FU
xpa7huEmwiUOmf9k+XPpqzvRcPrpDg4SZXRmvlBde27CeH0Qk1gzzdUhSaRzvrF0
lqjH4zKjYg+vfaLs7j1c17jKl3AUGqFJMdZ1jOJ2Nqo4tD9ywiu3oqBK/j9/5ADI
W6Lem14xFUJHfzrNtVFrAmR5I8Nwnehv7yfmP2CsAGEuQBKR7eXa9PIS4eotuhIE
NiSmqn9j/7SkH2WdyMszS0vrjevIWtYSBuYv68yy869S5CkPGJsejV9ckIR7ZeJ3
rg9EEcpIkV+MVS9Rnu+wOASdbPEAk0+ENOIM0nIk0nmn1qx1cZO6mtYifNeIOAKh
ACEnWxfVOvoQfYRHDImpLk977qQbBZnDkgt2Jamv+f9UQhtAcgxqth3YXMkV8nuj
zHzEI9kXtMymCP684/R00OntPUhMdfd3ZNiWKMjW47DhFlwM4/uSHWpY0k5a3bHy
xvyFDBoiTKru9kG3HODKHx28SI6qY5hdXrm7QSszFGig8V8CLDGvWir98z9u5gZr
B+fgCTjNy/lzrt972uN8g6rtlB2BZVKk+U6GqQTiwtN1llC6WloXxBqc1O30GCy4
Z9MimlY2r0qg4W8yhNSMJg62XB9kZCb8vCOZrapisTmfp/eKjYwWUgiYEzazmJ03
g5LKlV0fUoY2acN8bCnTHL0XIIpKifb6zH51ose0C2N0UsfclianL0ffmpmtpMpT
6oJ5pkz38rG39P5pBnqSnbLs1ZrWk+J5V8bfA+C4LddWfHNfX28E59QOhNI7EBux
vSNHvA6rQWVoOcYvYv8h8NIsLe68Mx5tnOauhwd2SEyJTySdrhuco3mAiJrEBkJx
36uxxHlzhauE1lKAP6MkBjaPzsyrt4rtYv47N/JUUruL/E4LgZQqTu2aWX3RCNiE
Vzjq82Agv0hkhM+/BpdzW83apB7xaD7xPim2BN0kG0L7H5Ycrv4G/2wza/TGsVS2
g2bPGMzgZ2PaqB7/ku3h0l0kTxBClM9SNHKAUiEucKIttVURBGQ1Yy5fnKa4paTy
p44/E/nsetQREp5y2/x8E6BOzIr6tPtOtDWgiV+YeuE9CgHhfh+Vc21ll1k6JmLN
2Z3isXwqZ8PBZKL8qh6EBl2WK9VgLdFrWN/EhKr5xQpZER3InlC8rHTjJBh6LNHK
+UQtRo5Vdogx6LMJ8Tax3xkhYRP3J/OAQiVqmVIo7/U+738DE24UMNUh3iT54CpO
sY9C+yK0SatwYWtflCOt4u21GZUSpGKDy1kjuMLOJoCn1df2lOL4dXpGidP/HzHk
qEybFnhTTNOg1FDLAf4fmeb37PyxZBdYZEKxOBhntcihCFn/TQTOADMQb+7yFKc0
w+vhkzi/xnyC5I1ZSgXIeGkf0qm+IBel8wdky9dCrxzzecz6fWoPXn7tfUpWgTqn
0kbYct6iUw74Mt1+Mz96eQFAlh9iux2lV96z8kLISL6a2pzuwgi0DSJUVsOupcu9
2ha4VXOXeEF5CchJRxpGbijAnNleYNvn53683+ff+HUC6Aon4SoDUCfxY4D56i28
GqX55AteH+2V91EdasIIgEeLeRpFDHyauj68qmBBjIEsB3aiBspBLLTCUczOUXa/
Yx2hygvsR843UyPNZKVReH1ZuREh8PyaqpJvEm9QJVZwZUdGeLPuwLqIofFZKq/N
HMXORGy0uTf19T9pHzRighkT9+iqRhOA+tte8jP/1konPyRgabmOWI/9LFqDLIy0
3bgMB28dF4ePYam9UhVEzvWbFPtsaGXxH9CCSKfbg78MDS2+0ZbldJ7D1fB1C085
w85J0DB+TItkS2CTHn7M4pxd0k1eY757LwLSSFmw8ey/IQKUfsCy8bC5G3a1aS5R
R9XHTJ33lR5NLOd06K94OpCRzqhm71VJp/PlxiELe8qM2dZBj1fBWOYvZv/i0xTm
0+sMsEfZP88uj2+EG/fuo31pwV3COALNFsAsDFp9YoHPGnNUU2AaouGCLm/gWNxs
t6gRnv8DKn6kCA3ADvOKzPVNk4noXdN1HsTOWXE/5NTAn5aVlTCDszgQCfjI5KGo
0Q9bbBVA+DsKaYNWbmNjqN1VG4MhobcKFtF/J8SeSL24k87IC51TTqIa/eZGev7d
onLKbc0MVpG1xUY3cBnhcvLbkJ/ObcSkDipo6iJpZ7RbWgrDIcmjNFUowE7QfOIM
N2o+Hp3HF8seVM6KSYYM2YlM2IUwHjfnydoQj49AwlcPO/xTaSLVQl4iK+g6vYwa
iOeUtHoFDcPplPeE9pqzav9T/ohuBayn672ftKpXlT5MVRQpAaYhUF3mfayJ3SHy
RKGAI3rS8oWySyhTAb0FA5gllwJowB0Xfxwk6vBwKQn7SO69AHRshIEXDeTY5IKw
5AlVT4kUx7e3wk4YKkz0EhX90X69eZDdFwQsm1rvNW/JgpWAhA0MFULvgtVFCCy/
p+jn5grESUGnD/ew2/JttWo412yi9WT1RE5B6HDI/hF8D2xZ/+vOxGwReSEoAKwa
ir2aoHn3EXqkHJA2FyHs58Ee5tRSAUgIBsrxZ1IjwlUKKk6Bbre4To2ZsXjMhZya
kbBiDSCOSIdlOkdVa1KT1oS2pET3Kub9Q9oEhjmEql5kg7beuobzN4X41r/lF4ns
6hY7j59Z34Irom/IORNuqNwR9qVyD3f37xYXJrw7qLmGat1NAAGCXLcYV+Kl5N4E
EKvqEXPFl9iHn5CrQOPrYyq92/n6oJ3feYK+QyXoP21n2OT2ecXa/sf1+B5G4M7y
tbV+KeLRIY+1MtxItq0N5iqPpe3GoEMh9bJfUfhVPEEx3owD7sBbYKCSZTWlrw5X
GKokhMY687welPJEJNVWM5qCg+hkx2lAnZv47JVv+SLXCyo26XIikIXJSd+jnuAU
b91aw7GpVilsFTEM7Gr/cjA9TlbqEEf9hyZCIIq8+XVAgnvh+ZoOKMosyw5EZ63+
TI0jqp7zGwMkdWHm00kakB9/hVFUU3Gl7F2Ax381pV32xP3Nc7hp/TZCB8x84vTD
cdeROe2gjc9ID1PTLTeeO64QBP6s9CSmUKAW2lbCilYzyx02LE7TLl9NYerNUP/C
ddXOkKmNVx9LdxWNT/X1nFaHR+UjxuzGEoOoyjrm1N4KIcNGZiO4lu6WC02JcJRY
oF5BP3Cb9gAKCg9Cyy1kI8AU5iHVldSV+q2PZXJNpzmIt6PfgqAA3jLHlpxdeYFe
m9IhQOOLUUbTVYGX4fWuPgdgqOCiZ8LKzdT9aEMEc90qSbL/dZxwWHDpUfCWfcTC
GA0s0sppbRYvZfYmzqqVRW9/UmPI+6locrxCG3VbmW92275dKD22UpaUjv4NatX5
08ayd2cH/b+IUXOlrouOw6dQ+q04hfqbmjZevgUAwQUsXMCfGIYTUUu6I3XGdORk
nrWijyT0HJIKnPHCRiyzos3MlZ7HRcEXIOcBTRK5DUhX5eIDFGhDiJzAVRv+TplR
zm26lz28wD4+I8zSsEmfc10tY9lV0h1ef75TysfGvQsXd1haszr1X19I+sRlR34M
3ER8WqQU2Ivsjo1B63urISv9+O6DV6tk9n5o0gOgpKkv/r4K5Ep9OAWNtWuPOa6h
NdCAP6Ck9Xq2DnGo5rE6VJEQT8uf+oQ9ap3dscI9R4Xp6/d0FGgz7WWO0L0MGFwC
vzdvHwDFyi2u52trRwnrRhZNWnkQ+xc7MY5KUYBs6fyon9jPhdFC+/JDgYGAMtRC
LKNem7BtIINrwk9qG4OwhStXHhtKqazRSQpDID5sGSuYGthgG7RXec//r0TS3Cuz
ScvacUmClmGHIGW8Yg9WnX/U8dH9x8hiClCWzknXCDbzDWkSTaNr15I0ymwBct5y
3TrHna9G7SiXqzgxLo9W6zP/GzQ5Z1My/klzMi+FcrFiH++CPSXnmxi7ZztNnGeh
17XJcf6oK9zVWRnhitXTC8SIDs/cLlQw592E0Xry+Kpl5qUigaInE2ZUCHA/vE5E
wbyCxLTWqVRLe+7+DbSGs6tCGloI2W4WOfFB+386q8rDTaOUXy1RocDUwsy1xp5d
slwBkfpF78zNhgfDl6SYhsgJZ0LaZtAF5sYHDEkpgf1sJc8ecl2eZ2k5BGvkX6/T
EeaxqvXufrFgCA2daVfQNOD5aWYuscdd76YGKtizYH+VjUpocEdJiVqc5Lx6s+9t
TfVGWXeCnWGRXw7hpRU5/7PCDzf9BYwBHPcu0GARkFUPRsy7mzb1+mxxaCKOnTK/
tx2xsY6a05WQ/cSHNNSVswLJ9/8CbLF/wiIekYRhA33g/k5HbflhoCm0nJS6GUwN
EhsxToiEN5J7E1JYmhEijvrddVamjK8OWWx3weJGb/YKBcefNOOhVWn49nWhzy1n
/BbJvXpDnVKzb4EcoIFPkRCDt04EkU4PNxrI+jJP8zZ+S5Q2OZl9n+dZn/nLZWpr
ksQJrMWw7wkM3ezTBSVxiLmI6rbpPUUyooZ7VcUE7c6FXfro7cpOX/OII7edhlS8
Vz3nbcWE/8ch6OBfwfTpa9e6HBi+quq3sp2T7segzBFWAjWTUXTGKppmbuNI7Y/5
RO2No9sWj0Xbeqx+VNzQzKYsR+cxNJA3Ukp+cpPR0XURCmVfbRPZ4fZ2YexW9uPa
y1YBaf9vifpjq+qD6scOUxHWLXrxsgNmD95Tl4UtaAbi8rjZWv1hSw+ddJc1qQKW
AYvrGvFc5tSEwoINJ1mX3FMc3YtlTQVqzjmHHwWvF9oJ5TfSC6MywTK1Gb6ML3oC
g4RGNnCwMy/6Z8On/vsqP6Z+c5yAYyN09akGCtXo/8LnGwLI7sYlOOWn8nkoPdsE
OlhKgueeIncXppkqD1aN6pRCC9epxfmP98xT+c7QnixF2y8aE5taWBdRRaJr4fKP
a10yi/vdcSBzH4ZsdnJKtfUnuHujIWKWvzz3Hvok2yYs5Tf44Koq9UL3MYqQXYJw
0PHY8f6EuDj94FOrtjaSa993KbPfaPbTH+hRzOe/Qdbym0iG3W+wMyWjTsCYdeaj
MVyID7GRbGAwG6r/GATiJHz+AU4Q6uVDv87GXAGaG6EF2lJePWmTNhxfJNRUeNHw
F8C3QqaJUhk1IV7zRy5tq+0mGqMzIURJ8A7D7T4zRZtqqdajQrP1eGEA7bNOR3tP
sD5SrwFeZiWYs+m0yEnnnGfVYdfE4yUz3oejDBBqN93fwJizpvieB7DhRxLwpduf
259Hj4+MRXPTAXM6PuvW5HEopkMV24rR67nWZDUcnd1I0BHAqjEfPBFJhwqorQix
iiFD9jv+0Gue5iff0JNa72tf1PyPfqXYxzp14OGcwV6FqmBjmzTlw4+u3gzGRPv4
o4DF0stFvw5kcDUGl8fbK+PYvcp9vzwP4fz/y4bm+EnDaGQyuuBZux/O36aFTucj
7K35WPXz+BmGlUAmAukBrJFac2fIGriNekzQMy4hKftO7eAkUFcYGhw07iPf4D1y
U7Kq1JkmukPqvczu5UoezLJYLteOC8lCscehN80btEo7vlI+MwzrcSqqGE55ADiE
amegj4D+KyGTYVHv32ewWrZltyVa/IASKftS/LbznS899VtNcwtydtPMJS49IWNB
4ow0L5aeqx37DifzpQuI/nc4xfZI6rcEDjigQZFMzoGVYldAIucMQDUTtD/0coj1
HUqhMqQQJ0JiTV/EKTldc39/VIYnkRVu0VLhaKQkmeCQfmofEuFYAvU80Qtq6FZM
ejIlmjQ/PLxewZ0xzLp8OLRhhx1Nzm/5C5sDeG/PVBMFVfr0dgph9EIykv9DdCS2
2VMae66dZuX0POx+t1vkWZFrbBNXZPwYnNfGG8FgFafl6OljVJNNr0RgHcQ8/Y4V
XHu8DxqvzHyRx5kG2Q+gemMs2Ci1RttQwMmMR7e9XCe4yvmFK855uyAcqvHkBHbH
b0NNyPhj6EvMXL9yA8RcgilWXDouELOEqbtpo4ziMX6FtCdzjh7LcMC1wQbS8Yy/
Q0Tyy5e8YktJO/sd+JNd0nlXbT221vSUakFgvKn5TYJ/IcpUJ1YnsDMMJ5dLNl+K
S2tER/fILwnX7QANbVCOjAiL+xmoakbKkh2wP/JdXzbmd8ouG+o2SVFGZCLKP9md
bQfeMqStVxiHg5lHtIEwlbgoSF7rgkx0Nea91o8uSuKRR6jWKZBNZ9S5yv8hMOpE
U0oRrFIOpOUYgJp3b4gtLfC5BlL0Nh6dq7CHxO54oD50E+tWmfIyLc10O5/quHud
b7oZ2/KM2di77Ds66JqpjCN6i9CE4beZYFbeZWz6YrTlYT9Hm/WViHPzyBaKHs1Y
Sz6DHaEclLMCKWbTsdU2NnbaGxCqMG3PRUf0hNw5KAny3pnPcvcb0Xh0k4TaEiUh
akwfjwtDPdDC0wISsIsoVBLB5rPNdT8dStVEFxB8jFM42iJQ7l5oU132RY3pNGI9
LKslJ5ebK+GEvz2mGjB1SMiwkvlzNGjwQZ6Hg3qSnsXRtMNulLCb2d1fZ/VXL0h/
x2Wp8hGyX9v8Bleq/wN5koyQa51dhIWYZhbD1paQ/x445DcyaKanWcXBV1igZ/FN
MRL55LvUg8I/t1ze58mqf2QPu7p9MkYOZHOyiO2rC689b4biGzspYgmc/221312H
9QVQZ0JPR18EdZ6i7gzCl3XJQIFkfUtTaQmPWzbVcy/+vxrzRQE3HLrQs62OnSmv
saGrbv9u8qbVISVJqSFVvz3Z4f4Lqrw3hNyptj9aDau+SxS3GwS3e1ba9q8JJ58n
hBLcTNkX+dSrpzSF9uVyK+ydz00XfHa9HHxHWJdwHgP+yGJ5R9tFYba5AowpdqyJ
5nryCTIcKrTRgwveDQlcJ0QfmyNN4gHyGEPN74wL/1dH88uDBgw+F4nknjyq4nli
xkvJYLpLiVbpIzb7DKUQAUboFlbf2eFWIwA/JuqD28pH6aM5pCKiZIF2ZYbJETT4
h8Gy5pWQPHDSzayp36DOhHOk0HXZyYuTwX0g9zjVhoCD99DVZPMagHiUB74YTeIo
wZeE50Hk9XbrzlPo1z/YIWowyWbZ6d+JbavyqMh+aPBTnMVtms9RXnyOcgmVLWxV
M8VUARmfNdLJtFXyZ96OT22mo7O+rxkUPaxKricuvfrQ2sbDAbaYHvDHSaANHubj
gWX+FPxEWmWZHzhXRML0WLuKLQMhuyM14LPIlk7bfg7qJzsXvk8EIEFfJK6PceRO
vVlzuSyvVa5t1N+cwrV4HnPL/4XLaTvVKUjsAP6fwT0uOwALWeFtcboq0v/x18Eg
2C8kGpkoZ58vdm1SmuJzCcR9jBPxhIxZDTodrRY7zAjIQ7r05dVD5GvVmkZ51noO
TVYXvwBx3rCL+qVA76RFVl7j8L9pOjbFktWvysKg8kdww5bk412zuJNU+IrVBxCS
QlhCNOQwMB7WKElLeJBznhxa3ELL354jhId1CNU6krs/9eNakYRwfwcTVt3p42u4
BHpYJTCePkvrzeKi2S4a3nflU0YYazNcV5Gc6lekrfqr2OqIHyBpV7ZyN3sRsntR
40hB885GJnc7PJ4ZPRo+6Fjv20m3DnlcATpmCKkxrdkMHLhdp3n8LwSLV/2FV5cB
S8VSJRQNYUeNGOkFp9bHEsrerBbq8bVDp8Sbmbb5GuFNddWAQMT5wVEeZvyTLLLF
5PUpVbx23k3sXJY0MVJUZw0vMrop4AaPt2gREJKJC0aQq9vp0HSzp0gfDfxE9VgZ
2PoboqL/nFSPJXrt4ISKVdjH9TkXG6CcoyAffwVVoJdNvfFxP8rGEvELYIyUDkh6
WuB4MmALDH50oJADiMzKp5lbf2aJnGg5AQ4J0evsTRcGcMFDsF/ZgoEryzMhASMG
3d9B6SBuA4OiwEbYHarRGXgwqhSUr6U+js4AXlGO2EekET24V1TXxbQIWnQguHNl
rmtNWQ2hgxDQ0RaetUzN13rQiK9iON/DuJQOt0zFA9kdIBqgbhmpJLGdK+ohBuhJ
uU/kLVGs4X7IE43Dn7hA7J4OqRbpntm00AlIIg9KydQYaXnnYA2MIYdudZzA0cUb
njxShhBrk74v8eoHMu+FU2jODqkXWo0Rk6TsUOTjmElcLyr8fVMFotJoAT+rNV66
SHTVNaHeUqKPFLIU/sgkK5H8QPOv2oMhGdh8afmzALuCz7AwuKMxQmxQvWLdC4/w
dZZSgl5bNReK4Way2+qR0qE9m5sTRN6236dlR1yXE1LVlHAEFN5RCesYQa9Z9FLs
s+SwgBcwTMfRDXA8dTLhutW368c0HZjBcKINttVrRTUbOcc79NP09CoxCC4hDyqe
yDyRT2FcJRU9kk2PnIbcbmDNlxJO+sz0P74yxPiKD4vs8SXnmbZvvEjSsyzn00qh
5VXGPdebjkcj97691oMYEk9tsyQkVX8NyMA3ZxmvF1vIGsA8fveboWAoWqAs7M+n
hWnQGfJrawFQ35ZttcY5TlE+zpr2j73Thq42Y141JvI/+jTcT8U6lvAAwgZosDrH
jFxGUnYiKTCZQOVMLP87EANDKXvo3yDKXKpoDUYvNhpSFPCyQIS5uyqYRFzfz23t
KAkkL/Na5SIcgpXRywzkbyHniIN0p3KofKTgvjLCXcKFpOOjlKab8es2cxc9GSjT
YSSB1AX5cGWJSPqG4fJb3qmYuCF6curd0f1k7dpLL0CVEdHrMSPIGQRNEqSOgkW4
KAYa6EQF7dT7Sd05s/folEG1h0datozvcZ1L8kOw7apoKfWDP2keiB7x8kwL1gjo
u0n3uIq+vt6XFluPmEm590iyLON3mhVNtcKk+7osNRwOMCV9ijgtFP06vuFgOgSa
Fj2znn6rd4QD65WEZorFVJ/ilRMO4EIcZ0GrFlxzAmtx/CT6ZM2Xc2i698Xpttw3
zN9+l8haF0nF37jakypY81wDWDH8t8UWP4gIJKiTDSaeMyOtxXe5rjgU1MWHrZ2n
ERbM1IKThkPTrXzGdA75haRblzJa7va2qY9wUKDLUfOfhyrP+SuN3D63WFVWg7II
MUv1mmF5KFCLB8iIOxxZiIriHvUYeytGj6KAg9rHnKPC0UBoEgOEaw+ooILBaIv2
a3lezRGGJV0GPbyGRQMh0uQSEWyw7EKm79S0tpCaTviJogS7O8B25DmQ+chAcKVA
cmXkLG8SnYY1e+bgY4GdewCOqt6rd3cZXVUKCQrIS+WKvhGXNixjuERBrO+sQZJ8
9AsERHI8ZZpD6u+uHlQPGaKaOyKAClNKl0lIQzpLfzvnpdbzeAZUQKinn1U5hm3S
IRdRthZg7pfOtm+93rguIhw2jsWZPVS6ItxoMUP5jUKTrgq/oJHyUZ4kjKOonPVf
WiLIoRxlS8jdZ3HLoMR3e4zmkXW8V7Ph2iOOQUluGjI=
`protect END_PROTECTED
