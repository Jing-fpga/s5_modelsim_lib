`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r2khB3SmNXoGuelHHTP0Qh7CHsx5pza/ajMcHLrDj4IF1ZWPkwO1fD4C1AMdYuIo
B9IXc9ZB2jUi2Z5+99UzplFkCsygzkaxHf8xvHU/4XlsLf6hb1iCrNxTQtwsaD/W
ozCIPZ332OmexRdog4Y1Pqgm8BHSmrA9x+2jy65nh7S6XRKafFQ34mqb4QJxeMQF
fPDXcymJVB7abCb7pk6dIr7jabtARI8hylpAHAoVU00J5H582ARASW0ayXbRR6r/
mkSLfmfn3zPaNPtAhk2MDQYt0ixDZRYgGHOgv1AsTrsugPqkHwPokZUqYACLCm6F
L8/WaFT1KZXJwFOmpsHVhnpQBLNjcja2NG/UwWm7BRMPipf1BpLrBcH19ZtjpHYT
NGlrBi8sHEl5yKt+C0S347L8PvVbjPN0605UAWeteVGHeGZoc4Mq2k9SGgh7c/Mg
y8c3TJDDA1lfW7gEEubfT4sWe8G+knRuq9VJfe9hrf9g9IFI1FgxBJM21xNoViKF
u7ijVSjIADifPmOajB5rz3JAejGmsnobGmzGdxGsoxBS5SpODUAo/D6bElrmvHNI
hZJU1GypjfytR1u13Ls2Fv2nY8NTsH0WjKd++8qI4Q0jpIvFesOJ3oKHHsVbkguJ
nHclpCKitYBMdwuJwi3CjYHMh5wmyJ5RheR5DV78BLU0DVzSETinB2hbs60zreF+
hijhCn8RZJpBlHdHqR/aGRaBdRN6tjM5bqN9QrK6/2xbo+2ZSh+MWpRuKR7ujbJT
Jfphg4gDxmBlRNdzGiTWUowNZF5oTAcG837Zk+zeclrmIqg8Z4z5zJMem8iGW6g8
LBLTE/KNQ2K9rgEG752lSSVifA+NNZ4MJEknBqtSajWWobJ3vccOrZC9zbwXYO8Z
a45uLQj4NCxbqQVNTuqBo5R5OGVRjeiyzWH8atLjs9d0glnMmVA3OWsrmvrWJ4g4
S87n+BqjF0zNIy2LxoqqGRLy0eyG60e/rsBgY80Mz2inYwgitu8G2+fMuSbW5Ge9
KoeTIlT05U8rhWPGhBmy6eMCrnRRAv7JL7bTQ6QsesbCXHgG/mO0XUGHbgASCPu6
Z0dd4HMaQLQ46P7tuhtWzsUnlK/oszfJ25qtC3c/ryB5xrfehffW+s3fmlXzO8Kd
/AHKhfaHDiJI4G33sO9b1tgESIQDnB2bthnZRoIsGhsVBhW14yAUPxkkBxZHcVB7
EWHIlqqiFuwlYzvnmzCyrwx8WXek7IJNH7j8zBcO1e/GIY5StkEaCRx10De+9lee
2T/gCDDREx5HwQ853y7GYIvlKw5ihN5cT0JySq8Ea6GDC5pY8dxze2v/qCMe0lIF
ACaylgXIHAEBS6mCGe78DaboHbxUCfa1IdDZlsr+rnz9CIJegRxFs9t7SJxIw6m6
g9wXIKra/5yn3F4fa7ieJuereKIMMyRm0SHFzmR3XuppnSKoW56r+F6o4G8tqQS4
yc6QaPozCSePJN3EST95TOhrFkqivgw41jG16olQSF7St4am7UQs8n53HJpHb0sH
ofzolMow6ZwkX9NfnmSD2KUD8D2ZmB4T3MW4s9k1MDvM+wsUkTTh8Cb4bsrDt4fw
cYY/2S0vZB9t6mq/JlN5TahvSNviev9NkVwwDBISDBCEnmKJOebzjqyHpFk8ImgY
ulhvd7bVSNo7jIqXqfPUrd/rvZLLQxUPGS6WmqVLbaDOoRGVpIcOr246Fpq798/r
MNyBI8vkuf8wC5PLCDwJGuYva5cMF/JQr21e9nllx8Y2bVDYtmSJTRvSD9L/tx/B
mQvTjl9mHexzphJcFMtmvN3VxFWDm+xQEQ0W64WKfFfTwQW8oSqm4zZOU/G/hDu1
ExaUiV9Tb0mnjoN7TN2K3Abt2uV6Qz6FxnJLaqVLxDEb5lXjp9iPvShdGnYtiQwQ
RWt33fwZs+NmtqVzGzMAVMqWWsd8rzfl2cqNRNMeHrOhI11xW6NG7SSaZTxcxrJs
p41d2O/n9o9du2Ayjp4ymolPrx1Xq2sHlmv0C1AraTgSwoxJgj1pafr3I+vBMYEW
2I7Y8jB7OHfmLV5IfPl13SNzBoz+GhKFqlmr6ndQGZAYfWLyW2RAakdhFfi2BBIx
1jnYnY01UxLwtIobK65d+qvGjrn+BuATvxwPaWH8iJYgmrfUf8tCY3QTKYLVTpp2
s7HgovEs08ZHsEkOtIDfg7dDAY/P4ENDkLcRfqP+yp49yz3Q+6/W1fEW3HS5zsWV
g3/sTNgP37OawtjogldDxn7eIKYn9bQqANLUpb4Dcia4GNTtvVPOk42Ctzav42A0
evYHlKV445bIakPQMid6TTCpWm4VeEcBDsbsKL2Tf/0MNxeMhamNLQoTSU8sVsZs
RWsrCAUR7lMNKi3p5KfiA1ogIE7OMSpOd6WZMFYZQRIlBa6mWNYilis9SzGGWiD2
pExuK8EixX8LquqQYPO9JgAqaovaCkmRwwkrJ6128FXOI+IyDf4xv7/ZIS0yNJEx
f4YaCF07WluTpWeXbjYt9jYWpdB6ltBZCGCvn6gIxwMbBT6N49xQq1rGcZ5C0tYX
jFx0yxSCmiYtwzHHP04Grt7KOJl/dGLlKJFb1QAb/i2Y09FN+ri+/vIr3fA5Qx9y
AaWuBUgN9G0CUS1rJdACBVVff1Z/3Nex/vl7AVrH1gS7CsnrCUJ3F6F+sqhFnrI1
pxMTw9NE7CTMWY7SKfbZ7baaYxqP32EtvaQRO+HXzNFxM5VZ+hAZIU/lHDRyYYk2
LwHoOqqjy2mY16bQQG11DlOLbO4PjjwK9wENlu9MNN+zOxr16707BxAiWZGOqVLp
3S55tDBhSVjwDi4Cz7a4mdqvZJ7l5gIXGKqytN+vCaLqS8UijvhHZ2cu1nMbUXhA
61iY4cZo2CvdetBC2j0EQ7UH3X9gi4ZT+B9UzdQakBgtXIhLC4Rdcqr3AwJoeCfN
vlXSm1xjVOkgALT7wM+dquLQE2/YiBj+i4ounKjRI93dXTb5MKO4iZobSwortbGW
z52unwlHcS801v8LEXs+TtQLPgWqUjgRec/Kf4PSZ5hF2BEZrtJz/SB+orOJ8xtf
ca5GBHQSOqmrurEpZmU8H8/MXUVQJ/B7kUwBNhVkNmMtDeoZW3eCHK/xN/L94Tjm
2WJZWdYiPfAf4qZRuXuqGpDYgUSKahFkG9FW+UD+iYbX50mmnZ18mKPbOFz2JGnZ
`protect END_PROTECTED
