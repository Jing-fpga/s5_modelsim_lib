`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cq4ZGD+c4ZGFaqISPSQo6p71iheYk/b+RY6mkuXF89CNgnhA146vdygGiuz0AI97
QBFJ8/Mvfxm3CQdQNtDPsPxDCZyDxWHC18ovADhFdq14VplqexkuU8TNv/+oUnYd
Vnt6B3d51VU2LyTppuvNwEYXe7YDzNbH+CT12zlFp23os6XDVWRprVoeCCs6owbu
xFHRigUfUabN7D4VkOB0GTiSwiAX0wbDVC8u+AxZBKuDYnQYOHLMVYYTxnL2sMbn
4+HQbZDuFV0fVBO51MiAyNqjDmQcuKMaYAy7wpMWPx0XAhkLivx+m/pT782bPgTh
GzN9m2ad78wmlDNIUzYC3axCAc0aepQy/zKeRS8IIHvF2tbPHzHqHwKOFAgUzv7M
PVnz7+Nev0jRosjgNIMCdqCQ6odg3QXlvCUjW1UZzLNSQNuEMqAMOmHJbg5fwRuQ
mXa4uVyJ6j7otgliKV8SumgJSbGy9ClgDOeh6iBTPKXXZV9FUd4laiWB8pyIjk9L
TU3FzfoPUyQG786V6/CsvpJ5k453MXsaPhKkfS8BZ54=
`protect END_PROTECTED
