`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yg36kn9W4dvTMagS6ABbwOGB33FP7niiw0B3GK4h5RFTiDnATzVl8BetdAqKP5oO
zAkU4n+Q3SDtwlwxycmm5vkmUKaXStvsVLSB0/n5ZGCi3vFgyNF8vN5Gb753U90L
aT9GFx8aALvwbVLJQREODZQk0aS0xXBMqG2wXo0Zal0rsxdRSdDBk8zfYPsX0yoB
tmR4EUaFzFd0nvS+WTAG+zcYhGkLY/eomgdRwctLYxL+Z+/zrU3PvilSCUwXX9H/
PCksErjsrQJ1MZFazEC4GJpNi+PT1v15C2gqnLJUVvL0+3NiNrew3GApg+R1XQkH
HtdY0933w0CaetsA4H8moBlgUkT4XtcwKUQVE1okrQtskIuTuh14BAPdEEdLdPNT
opfsJik1z9X/mOESxYFol4IaenZMZpRJT3IlSsiPSm7Tebo0+kuXO6WVa24wMZTR
twGQk4BYv87pTICslgBp4RxbrTwkxRRrp0eLwuhojog5LcvZIeuCkeDySUQytsaI
YMJBu8btlLEm92gXqI5ErAwkVDgWjroJ/AwqkeamD59XLVZxmuCBWNIBPgGR4ihy
bnnnOmVNI3mlz7ynPfqRNq22Z1IP9MiJVJI6b2vljIiI5cp1KRQYLKnnfwBviqzu
JCAwgwCZEHvXWM8fU5qzN/QfagZ2uLrgLXQytlgtj720PXaC3EPoecgnn4gaIrqu
OfylbmWVbjXPW8jxzhCxviabx3WUSuywd3EkPENT7p3jGawqv3soy5sAmnfvToI7
g1s6Sh+hx00bOz0dELTyfInrrbjkHzgCq+YKGstrrKYkRgYbWQIilmzSfCYyiBlC
lOs8KNwkMbnLaq9URnXaXdkALnbxu5/7lKqiW89RXEXLBt+hhSCIWXhjA0FEyQzg
3HAqoZXobricvmV2UgHJCoclm4hYO8tRbIaLp3Edot0YRq/6P0UReiCr8VXoQe4C
B7TzI2DXjzJ/YOwSF4j943YskgjOtRKeFOmeg9bvKZY2pZAVAWPTcDWEck+1AYAO
7pF5hkfvBNXDJjVI8UoSx9Me/HqRiTPln7T1//Clj37vz3i4eVQh0Mg4nnp/kmyD
zwUmUAq7eNty1PGYmzTGRzSkP5tGfag39L4+oYI5SvTMQxOMls5fL5k1kzV95rNF
n4WOScn+lYUezrVvR/BU51vuVllWxQ4xoc1HXMYZnb9jH45iyHVcIiffL1Qus+tz
YejaEzUZVX6kHuwa5iLLaFWdbF65p19KebAH4BRHD47aQFZAwF7f/oP9H7yzzetX
KZOOoXww1vdyQSCBIZA8cYXJn+K6x0RcKxccqaHW1Q9U6Zhuih09DYcCWnT4sXdU
et0qmYryoEaEKBF4Q+sslOL702ulB1aCf5tR/grZFFV9b9pDJsq8PfzQcCWx7AOM
Jc5iE3z6xEKEXz0IBAi2SreOTUd9xyIoBCkrHqNHSO+8dFJKI10F4tt4nr2jC08K
lFII6+eStoB7deFM7Zdd2ayrZXJ2FMilObj9Bpdq1OZdjZ4O9pAwQ9EC4Gi5Dvmn
G98U9ywzyWz+vh6h+Oi3M6OT+zewLodGSdF7ze6j/RA=
`protect END_PROTECTED
