`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rCXLt3JkfWMHjrS0b1TXWQYSxa40kwehn+qBzwoMOTUtaZx0X/m7P/AxTJMbYx5d
aPaf34HZO16XpjP9P21qdNkfQTtphCtWZPqRoZPq9aVKb5c9d6VvIExu+8UeiowT
Arw2l3V9ffBP2WirGi7c65bcEefFdqRrP9poqjLtCksrqrENq8dPuRdEnbnSRspk
EnNn3rNL/g1b5KsH2ggPgzAiJ/eWqftqyi31ASAX1liNPdRhG7ZkaZMebJN4T5t4
ITA9S7Spnnh5Iv/hR6/580nIYxBHYmSw9yhFHump7aE0oDI7rs+O8WLdoi75IXgA
IIARyO4hWI1G4Q/pb6Ddxrz5LCVizJ0VBiCGWPbKGmIT4UgmyUr1NwZg7gRX0oMm
vnUjirQ2HTuia50i7HTRpZnM6V/GIx67Nh8SxRrGCl2ZBHIEMhFngSflRupte8yX
yoAFGyxrogiIKer8dwuw5QaYi455y8UJY7XsDFU8Qk/cgGpPkRhP0JNl55/+YY4I
19u78sTdEuzu7uS1ULGowGFCK4fdLOYXbbT3AiiccFYGmjNP9h5+eJryp6CcjssF
DlVvcmD+u1ddRGCYIk3tjv7MAvoRE/npm+SBIslTfDLe6WV59rV2tLfGnAEn1Nme
CVumSaNqzJcJbW0jvpbrMKt3kjVaI3Guc6lN/XLw07Szr/IieCS+//auIpKMnWy5
aziO/8iPAslb0iktgqP7W3DFSrOvsix7j12hFQmddWNO+JuhICEBWuJU+ieYhF+D
m8irrMZuT18QBeRIXh19gfeX/9WiGZ93pt6n6dFhvO/UjHU/5EEjsbliFgOo6Bi/
lrNBNBQ4SgllrIuRfu7UZbfG9BGT5xhKiUehU6RHs+JPF3L+p2UPnhqdCCRtQ/Jh
vASPDj5xdJdACUMAeMyQzApdjCDMliLsk9WwtWdhxyPIzGbYhmd3/kuQyKeaUhjd
KXGQN1/+tfKmWD2v+t5GaGJjGPHawkKzVxae3mE1yRUvNSJCWgjbI2OmReOdMhII
WDg758Ck94RxFxJycbRG4vhG4pYr5W9xuEyLcjxSPdN0yArSVYEKE9TGnG0+wmqn
ptuqJUbRrHkJJCXTBd17gHQOgSkPYkLPlxoVz4KJhOY4+UPKbaLQIDKsaEN7YPt1
ZQwMr9b3cgMoiwcEUkjhX01hltd+lLVX/Ntk+rCz5WJdJ3n9GO1eE3OISrCyWSZm
PB76VHl39pmUZCOajtCaMNbJFr93P90o/UZGKQquq32hllfiIcZPcIUB6nq8mB4L
WgVUJWqG+CuFbob31HD+H8Sh5ATzNU3j7v5TRbnsIiBhfoHMZSoGsrGlSxup1Kl/
giInV8umxkkGvMaxXBhzwcXJg1lchFixa+pXiF9zrlIUdbrhCWw0DCW6vwFdjUYN
QQunWOBCjqz+6lylDoPh/ebAS+KPR1zdgL3sofbv7ubijX9ciKeqT8ZOOplGOAra
mf9gVHFxnzCZeCDupz6olRoav5+JPEKrUIuLwoj7xCCNxQ0myHOwJSPDQ/G85cjW
A9mxNe5MOMvRyq/EdDJ9yLy0/A4xWwZi5ZZhCfWHGDgUZwiST3DLYTmj5ogrIFmZ
8rofmCtqDK6x8ZuR7918dJRhpQ5vUV4Onvf4T6B1ghsdDS32Y+iVXJ+sbUnFh0w9
si34lkDLYHYYh4Baq+QdHL/4b/HLaWOZgvW+YW8HAxzLrJPZbDLLMR70kZs23MfU
oQR29Rwm9iPiUfbKp0TV+aiEp6l94LlWbi83KEpRFuYANsSvgSCwg5cYegxf1S46
Bp5IuiO2XmzL6ZIPIxMadpfA85CnbEp8Y2ijUhxfI1w+CeOY4lJ1CBBZqHr+Zs+b
gIeBTVWiL/LW0nAZyJE7Hw==
`protect END_PROTECTED
