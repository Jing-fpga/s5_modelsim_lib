`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6KGIMR8Spf4Lbd+elhVFIdYceUpd7qxBcZXpVE4/JHak5pgS5z0/9vI/TCd5+XQQ
TFI+EFoDlqliF4kqYdPfxVB+yyQ7W2D3IG/fEpE5H4AGDbiOpgzFTUirdMCZVJTY
Duym4JrgWLiHv+OVTtnKGXmWV4eKvFk+ExtWtqdLsemPUTbtNTZoXuKWfX2KfZWn
zjVmRc0tN4IVa1drhuPTdUKP+pjpDjKha0fcxed3m6soXZRp8Q45ZIY3Wuxl2jSo
a7bVsR90Ou014uWd71vn8R1EcENQaVfgqrqzTtjYISmjrlkocMdenppWYBFa2+nf
Nf4E6lowpuirPiTVvKOzh/frnNpflycNlqf80xLpo1ocX/8EwzOplQEq4fQrDbJS
ZcfeYmq+ITNNtT1TgfXyZdauhoFvPgPfc0+UENC6pTdC8R/+QV7zQuSkgE9ycd9F
EoObWflxgt+3nT5swZpPRIR5dvpPIHTGCi/nQCy9LkkfFKsR0yY046gsBb6RpyNk
paUqKvMIeYmIYwtEL5QUKcujfTASVgm4TkH1RJXLDXQWpPAnZLi8TTRAs7PRyORv
1XlOMkzfwtEGAo7rb/9U7BvKzCbXCB3fK6rKko3wyAe+HI034aCv1zGzU7PW7ly1
jR4Hq4Ix6AEIlpgQ/AgxWboLdnKTDDFx8d7+hKaf2t4EoezAT1GwPqU887hkX71j
m+5RQvTZY0FHqJmV03NcA3LPOK3lbnjXJUS9HgUKs0BxZygDz6CFHy9kYKtC2fD8
zoXvOZqwRVWQ0X0QNbX27jP/0iEUXd3FigTANVwJaZC5HURBtlDM/ybbJBcmjqei
n9sclMR3VoqfLNrGWrcTTVALlQufkjhEd5eAGoynCnIo1uaHL1KiBOvNa2Gy3hjg
Zkh/+AkdrmdZ6zVxU1/jvMKLa0rLUIivfRpBl3CviT2bWTy9VNx5D6414+hrkqBd
bSIvADjo3JW8W0SCvFgDoTibllQv33z+QnNWYO9Dg0mB4G81bNZs7FG/BQLnfaLs
qDgrLt6Ffssdit06RLdui4mqJcrREWldXZ2B61Ytopyk0TS8XFsvXojjgIfGlhuB
61w6H010vPAnsi8fMYBDLIhjn5lZkeUq8rXThfRE8BZ7Rs6eWho/97Zds7ouVVpX
gWZXLt4gkw3zGMFlw8PWVs7mHOnjbz3ceuZ3wWLusiZjGEozN6Je89Emao9Gjm+6
0derLGbb8wVIH7p5dpyxpHVcu7h6PuspKykQN++x3TYm1P27/uqhhWlQFj69YyZe
MHidM90nAE/GOB4SYrfnXmYLGWFuBjden+XBWUAojBmLuVe+nzV3ujA7UvR4Pu2X
JFLuDcRqLJ4Y1GguIL8RLF+lG75ycJqSBVp5qFtKe9o=
`protect END_PROTECTED
