`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/9tN1IrVh8IaD5uyCbyGeCDQoKk70IU3WbOiWUjhhuZtER3brxTQYZA6qM4aX+PI
SS+lRNvRVkhmfsp32SCY1q3KIhsUuO6CuOEd9mnGMUdGwXQmX3WyhllVmNbKDgQ3
mtNnY1Ps74WCMELOgLsfRnVfV7azF8txhFy739EwWS8NKJEwWmOGOHBKZJfhhXQ7
CyoZsvBTjUZjJF2Tk3ZDpSLqUNYY+dU7xoeBbmM+5HzI7/IDiZGVPTYwWyW6ciS/
5EbCyrc4bAu39GioQClgtw0MzdDhvBxeboBNUXgQDnnfb1Pno5FMNs86hMU9YKx8
BwODtDYTLDZthgEBF6VMDFisJ8Z4MBthNNog/Pv7jXhU5lG739rZRAcNxdv8a6nK
1dUMPuA8xU0HCIGk7Fp1yxEG+xuWq23quOCX5iZ726hS5GPYIHAhngozUSBpqUTB
kHDmC6150qohUwRs2NNzlZDmdOFJ17ZFqLvflmE1KB/AG/cpTgWESGyA1UgTL+sg
ptYwBCwuHWg4LIJa4lS3EJdp6/qFjYXAv4jlwBzjWwIJnYWlPtE83PAp6qyKaJ63
y0c7yUt4bC4oMd905tJf9T9Ira5i4BxkiJN29he9xdFSGYr+c5EH7NhS99ec4g27
duVF0lrvmxTUyNfOdcYyTjlWv/bd4B6R+sFcnFGhCsxkospu2jyaYPtoJRmlL+As
StULxky/wqkpKRIXYlbqow98BpyfW8zjoqJg1io8HEo=
`protect END_PROTECTED
