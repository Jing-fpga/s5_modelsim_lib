`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s1DS9I6VbkxxQIE/qFz9ADtv9x1UQiG9EHlS/gDd8rwdtK4z9E3Kmqv9kJHILMlK
u+8afu+cJIfzuHZnh1Dfn+9M94WE/h3QrSZxs+a2tUtgpFE2NCEPtwXe6ezRvwX1
JMjqvHvMPJgr/LrRg9K/GzBIrjVGYe0+pjuSGXLCkiBRJb4vPjE1YfEsLauNNhBV
ZQzMH6R0dsbhu9sOfT7+HDjgWDhWIfm7qdiL7BEmzfJpg5xPL2Tpe1iHbLqNO9r+
P8A7YX5kSXmdq8OD6eHiUghfZ5kHiW0vFQ6WbmRumzEhayZTz6JaQS8psvAMaLn+
U5DYfvtUB2F7a9nFb57viCzVXHV6L09PYXNbKF55BpUV46VHlTrWVah1sXV5ZIhj
8fpqlnzGQ0J0P5Dz92kE2AtEYeo2Qvn46Xrv9EVvxitkfq/i9J2OpjIDs+oIE9s0
ScSOEeFjItJp91ybs2MFn3j9EjkWSiPYSP9A4RdbaAOhu3FWq5tPACjUdYl8s2R+
Jpv+ATb/sY29Zgfg2FDaAXvRMqs2WOhjm7UqZrxATvksc9WYuFmLCq8i8YnQGVbn
5jnYIrjed9JqrC74B59EqNxZEcI8gixWB5mW/74Nk2dWwcK9GrEb730MzvspQqmo
Eg4pDz9ouIrg1YOrUy3hyk1zVXVVpGa10fVXheu10jUwSBsHJU4eWa5HOPJflGZG
Q/5DVyn+VwJLdACKa49f4w22dYTXxXBISPT8EORmYUuQuCTU8OO2vACol0QetwY/
KRtVuxk0tc5A0H29DZhOfIk/+2vvfrprRpUApctSDnoJcWfh6yFVBQE+bXbXjPcZ
Jv7M1WP9MndLWNk8vsmJsq4DhC65Jf+mPq7rW7lcqNH3hE9yISQOsHwHGlLPe2lL
WtOso7zwIfOSEzElTJfR3bYt3lS/BzTKfZkAyVvRMAZK6JC2v02MNdo0+XaXg7OS
ze9gRqErbS8uJgy5GdcO6dnRszfDYESgxiVCjmUSVas2ith929BBe8P38MA52uNZ
ckoaKe2c1ekxtvshA84+fQFclEgrpVeR3wS9k7iavhhErfX9QQlpdeniTpSYxyOM
KQ1Ib6oUZlD5cWMT88iBwuJ8RgwSxrahsmY6NPDqr++rJDUicQQY39qnJm463Wfw
6dzAOx2ACCeoGOcMyrDmPnOFShVE2OeSCF0saqvKP5F7HEQ1VEq11DO+a+Ihimjw
d5ZQc7Lxy73gDGUV8vhbCVnUMHvYRh7uttpxHwGAAO3fR2DXDpkvPMANUOsNaKnq
oSpFHjF+6DwOkSA+nH2EbH3/aeiUp60dxW9FuZDIebg7uJaT4ltkNszdmiIGDtZi
uvO5ufVh2pXZGSkbxyw9Xu13RsR7f7UjJJbJjp0ypR6HmZOaNDFnbfUy1ACf5EqX
BtrIgYev6s4fCojHqs08/iNzRy6ryBLBIYJVTdIDOBarmQvBytAivwaFV7RNtiim
ecFy+EkZbF1kl8/sS08bwkteJQ8d8TvAkSktrgkUBCsiJynRUKKuNSN11f/Xyn7r
xomzHzM9QzSbkHXwhZiFVJHEzVZBxHdHtuX0j06P7TJDatDwKGIBeLD1buZfg1V8
J+Vczrm0unMncBjsp0jmhbTv1JZkz4B9NoipUsfONHvYXO7n8qVZWmJiTcWXE33v
7bOtWR5iV2S4jwC1z3yD/+5XvnP5MSIrt+itjeXgtZxeUutNPHzKX9yjz5c6pfzz
pO9l7aD3IWm6SyxU+IL7BZi4aMXV++hb+JADQqOvy34gXqIvevnx+V7nhGKBZjFd
m7azwNcuHVUxD7AlyamT8HTQ26k2YnwSEZOn7tql4PwfXLVNFsY9+Qo8XFo7VWrE
tbz7rMUBJgqlb349W09QLdPzzCQlJtpea2sfyPO0rV84lfImTojhGICd3ik2ohen
8Xk5p5f3mhAT/Oia1hQCVcu55cK2Kpc3M+ood48HkMfYlsfEfxZGZ0Iu0wfI+Eii
S732VIjkHDshlFYEgTvYsro2/X7mrRUytId7AZ0JtYEJcaJWfLRwrgiQwQdegE7a
XxsUV6SQZ+sakqrf4gXxp9bXNB8HQGAhORTQ7SHIaZSt1MDKyCpXqcLhtA/i3opB
eZlCQ8FqOfHhUshSEjS3qxYnxjxOHfQ3lmxaiAnbm2EOG2bvQf1yJwOV5WneHk1u
x9cswQmEnVPLWB5uZDrcdZqAENV6E9FXZa3ieviv6FS42JnWSlsjhTZWjsd1ctcF
Q1KW9tZ6G05tQlY2d80SMYjICV9w5QTJDlvn4hcwI8o1PwNP9/ghgIwnHVT7H6eF
3J5ieZIvjjwJLG7G14iTXz42oHW044YHsJLdEb5h2Z306Zk1FtHnY4GcbzIWCI9c
mpqfxW5bKk6iYAW6INLanlxSpNCpH4eHBNHhnS8z+CYKoiH45hSSzktmf7ZdGcx2
ylwroq1f4F2WaU+HCvEw+HFOgR0C4XWY3Mrzpr+afsOUe357G0XCNe7b4yJ+pb4M
PBPgmw9LY3KrTGB4xOA/+SV9iKHD6wQ/VLAG4eJDdpMeKN7yKwaC05Aryn/e9mQP
/PRgUk69YS/G9hjiG3AAFQ==
`protect END_PROTECTED
