`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
92bkNqyDQI7K2oWredqYvPHNeAU7mLp1+fLbiB+ytPex20X1N913B4Y2DUHaSR7K
7JbpfN9Rmx5HhmU4KmX5Z/hYmCzxyHaHJBe7g4r+tZbz9p8wMsEMEkZ8xKXtBuWr
NTmzOpUFfv9ugIRxn/pIbCovLI4m85pCLKHWrTBM5xVc2oB5uiKyzYrgUS/iX9QA
886AEtbRSqpNn6o6TfhvAeVC343A/r74ZRVbHHxULRabjoqrwFjPG10VUInbWH1Y
G8rCs8ukulPhm5T1uFivurmT9Aj6OxgIgmmGrFD4XDq0RzZ+ZpSpTsCZpo+uBVfw
4Yw2yxqTqRmn8yU/S2UpwN6n7LLS2v1fW7uwNDe8kWNsbrtlz0QSeVbygYJhHmSQ
P9vceC/jSSV0AF7GKI2/Kai/LQbAkJJCB1Y/mHBajoffCsGFHs3MyW0lsrrWkduZ
iYPhDUg8sXqzLvXUYcTJpCV3R5tJMVYbhucaIoQJBQlfYo8cKBbsl/JoQheV3FZ4
YnLQxUzIiBIIvJEAfNfRaITuLW5YOppw/DR5NyH6N4ufuVlxsqUpQpIlRnE7slat
oth77wvtAzIyEbXXnS9YBVkCh7Y38UM9j8m3z3c0cqI3Xfq+7XJAZjXK5WXxChc8
CqM3RbTbfEJwIbUAaOyMqx2RTglDNZQbvuVK/oYxayIdssxyB38B4roN5ZhCNkyQ
Vd8LVJLRBaj1RktygezrI+mJc2bnrAh1F2r0PzZUcfzszYiol5LAXt+jqc7E3ltL
+/aGj6ttxtf5R6mBck7dLXZ2XvGNJHCkFFhS60PWohiahBCHm5LWrcICybxdur3t
dtp+N0hvcyx8+PSBS3yjQj5w3AYEJDD7Syt+3M6VOIrU+28HNi1cVvI6y7es7xBf
Ni/aXbu27NLcqTWsADZ0ctRG9YpiOo9RokBOfojjXt7HezxoMd4sf44ndjT+0Keo
rzkjDhUgDeMwgAHwZ5WT29C/i7TJWda93d3/eoTthJz6D0qNmlS8D6N0YrLlGtbe
mkKhWXpqY6yRM9HdIGBRclKnvrPGhYuYW1C2/6we9o8aOHzphtSNy2qkiT7jBeMg
3F+PH+pdYsdxNo/Y3SF9yzWGunSyXUxMV4ZI6GkvGYi1PgCtJSAarg/3vjxOFDnm
1s232rRdxwaBB5oz9gGut+pGSrDkxNLKumWERch+xtKDAs9/i+ybhelHy8wIBzk+
gKfc9MC/yQQA4lRQLy7pLoQK2vHcISjrqDi1AnHIP5J+LRAyEZ7kw4dv2p3QuY6c
CTSRpZth2DvsdoJARpkCn/zBkeFHBB/BEpE8zyofaTPftbhUA5Ob2B6aSkt/G4iL
6e9ML0ylv+sfL15zsv3dPAS5J5pb89TFeUpEbjurPjGu9/ZnDF7oKGa5BgDFUD7d
n3/4RGgthcAbbBnkT0rf/OJEuebRPH0v4KNPY5owuDsSru+/qkuLnNQeOGoagK2p
WvqxD+Oxbg8maw2FT+6nwcWM/rtyKiiaYLCO/RcKTZzwESjYlQQEXRUBo6Rf8UT/
rmnxBHh+ynKG+DtMaU8Tz7WgUHer1JB57k/nMpSYGZWQEf0rIFxbG42Ej8kIXnLa
MNebPw20UdFit2H8TMWXs3TlPNmIVveT4gMmAoUgCqX7zQsfmwaSCc56jZnhdKEG
fadWy5LObmF11SKb9tYEpp2l7KA87LeN4c4auL0VF5Qouke/i1RWVKBTYc3DkfFV
abHYlHkJJZ9TCsjvU3OaQfK4NlzRBJWV5i7TSKE6M2sfwbiSAtUAsr0xu1hv++BB
btycY/qXISbR4Tm7ociqs98oM2wEpTClJd8LuzLgo5Zh8O9WpKzAegZpCifN3u0E
zqxeulwlFbYgQ28JiCIyqa5wsSS2oLNMotZx1ZjAfSUxCXwSh68UA6Pv3vKV4wWX
bLIa3MHw7G7ddiHiWBNL+gGSiagfnAWkdoqca8td6ybqtO5x9xcGw6YhbPQeWXCI
pgyDv1fhkV1KteHg2k21oXDcA3JbxohQF5BEg4XSQr4gbcDxiyg9HGE3mAUFnKNm
5omilZKj1yG+K/gqlzwz2ujT7VwbmRu0hrlQP15/gCHXqWJn6sdkNUI1PaHd5Ism
i13RK7wYo+G1JwkH7h7WC/iDbm/Q04q856/QQrhmaVXTFw5eRREHFuKIHFiWPXAE
jVpyIb3dBFKJx8RLVU3WLLyu8X6cXoIaWIJgRfpMToJ9o2ZpuBgQqGhkwK014/KP
GkItcPpqfAfhobzqgKzJgW786PeCJxO6eFQBSaKSUlh8moRJ4l/fgP3HwtXayoMY
pd7IlSpdtiHabigWYGAVcK59tnuYce0xgQrnlmOfsmM3t3GLyc9UJpxHOz2C+vvX
C5m+4JZ1jS7oyU5Vu/btVoaI0dV3CZZfclWm2TvuibpmDtPA3dgRn9Hn306q/i0t
LXcuARCAO/pT10Y4Xl9zUDBACbKTEUX3AcodSJHYWIhXSbd9h2SxUCasn7Up21Hh
NI1Mb5XCPQzaySzGaRLD1B+h/Q3m/insMRumhGuXs3QGmGbc7PMhbsDiCj6V9vZa
WBXlJRB7BPWh7G/GOdI14cZae9I7mnT5JgBKQuzlDXyuJojVwypNwO0d0yhi5cj8
/fpf5gmdZSPL0OqU3fJn2G5aoogziM73VzhEpJ9fHtV3M6QIzH+GmhsMzlbXbonf
EQvm/KyiBJ1cOrv7zPZpAqxyqU4EbbsRzmsKUBimZQFew09izdR3FcqKX1DRY3ES
ddoqwRCPgueLIDq3SbDQ+oZMNiRzDGj3oT2y2xWGDaEAVt3eP0CP6sR8Jca2D6tI
6cIsnbNKUwLsJVyLGHDgJb2ZWHeupSIkbI6/ijADpXd5i9d9EDN0+Y7il+818ihH
t+IxooRU0MV1bGiZ+/pIODP6XhzVJjOrX4NVOTW4Ft4cyqj82SlKrkwo4P+7Pq8s
H9NdHgccdyxz064EMGpXgYhWbQYf62z0UObrtORA/XC7Xsk0kjlI4EJGMErJnnr5
NAqVvPit2lgErwyqs+sMQr8yIkil8HxyrsIsgLxkLrOFm/fwfK2SEt/KKPrXKkez
UfUTFNVCyJ+vIlCjGFI2JgqfZhauj1GyYgGbYWG//5hifWVwCMXuN5NrT4YToVRf
u5tqlrte8K8OAIHWdF9pCMc09F7obKONMc888cW8zeMzXWUSSvc9vf/noSpZqHEP
V8Q6o8o6QEGf8CuC+dtt2egEQ8didogp6uj8Y+/uLC/DE63JUatOpEkQyOyjUsu8
vt6+p4EAB8MNwz0i7XVUE4c8pkqdG2DjKFrs+PweT0iT0YZwarNH+c5J0jFDZco/
fK2jOxCM5zVvENlmKYy6TeNZsf4W1TpICnrqjfmP225ac3Mhsff1KMNT/awoy0xY
A6r1VM8kV65vxhbvJ6MDgzjvse+yK6nzK4L7q1r74uhZ00Dm2gEp/rDVwZAC3A5q
+GXyOdkYoUJkWWc5GMB+mlwgt3u/MyXIhvyaMceOSU70NiAPmbmPUlZQgWEGf6fU
fuFZeSLyk/wtWfsvqZSGKD2KB7Let1tbWODjr0b8vsrd6cbsbezSlQMZflnxYgqS
vqERPI10a4+36Rl2cuhnJ2AHahboXLpeI6bDYMU5jo/qp3vzCenHDVD/8vBO/8fy
C4ewqDo4LZk3kUczhIjClJiEysVQixry2QyYOAjE45JGXG0uzVeHc6x0bdthciWY
UXh93p9Kgmun4UC8hC/UTH8aVKDK/ix5WJHDlRHCeUg=
`protect END_PROTECTED
