`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ntOKu5HAur9MWVlD/1uKfP/FvWHX+LVdBjWvXJQH0JHl2p/V0ahwOqhtvxyMF4wV
j6mPDQXibUv7EdSILz4M1HIcgYH95bJp3kFRAtNR0L52/1Q1GJJ89BbeHvUDTw9B
eB3+P4g71CDap/CLZmdIpkpY/WfIH4W+cJ/o2ihKDuMFVB+bWyt8EieQow93jg3N
1I7kkqKXxWslucnD5ziJ20F90taHxveV4SDEUKNAbsN6lPsLYdg3yWWBUuhT1cCe
fQtEnkfVGYbpC22/x+494fSmCcAlnJO7cKnbcuiz9vtv3hpk9x3u7tX/z52vSmv7
grarS6tWJWCxLG3Q2jBlASTG8fpaqwFJhAXrjRyrN/y5IehfhDZmmUFeUSz2tB/+
2bi10/9YDAZLr/r8e3yFzi2n5MzPDNKNJdTDlOdAkQsG7H3CF3ibWSKV+EIWgM0t
3Ld9O6FpFmMVJNaRZz0OnVTWHflGeRbf7DH+7qPAmzevqrMvY0btf+kWG0iz3OzZ
m6qx57k1HrBS+VIoULYM9NMO6umXpx9j14Nd1mmQzaKuKBozUNH0i9NstmRh9Hdj
iQlsOfTJj9DIR8tR2fpLb31IZ12vN3DPCAQz/rRGPt8LdT3nUxMU0Mn4CVqMmyrK
noHMyjGJy3W5zDDb6kmtsmMTaVSVZnm+ECrnfXjrZWSFirUJoi6i5Rk91hUUyF1e
HRTDLvNTJ86Q/E3OPfW0hRB+5CrobVh3mP4Hj/YlbqdJY/oPY7CWvQLJN3h2grxi
wk3gQB4PEitpXSvX5FAMNsM0eEws/Gma/M/uNpaNULNOgHCYJ+3pqi5mjMCZam/Q
fQKqYvPqKsgHF3bdRIu2Qk/edfi7hQM8vKtH6UOl2r2lXPZdmsIM9LZkmYEVkjKH
TV6L4t8HtZN5pO0JTcf3zUvnXXAXX/MdSRmKwmOv9cYC8+2EPxQsbnaQGBoAJtcK
LZcxABB2h6veX8Sg8qCvXbjWfeW/5ABsh0XACJVb6U0KgAktpglpjFcRwPofK4V4
ANXIPSjSY7IQnnc0rKCipRqDSG1x9rqrfG/swk5mQ62vp7EXuaTRA1ef96ki6Iqp
4lmGCkFGuv2GBA+hA5+ov8RFtwGVjkeAU7mhWn6t1UVBVNTqA/BIx/9FEImUkWXa
kB3hHVvKO1IiBzRJ4rk2KO5SHTvCFDjQovCL9IGsc6c8127UAilidBb2WdjZdlTI
A57d/21XYC8vsAq1+Yngx00/SxO26LwTueYfh/A/fOcHHUHLfVax7wuo7JYIUyON
JD+S7l3uncNG7zC6AByT8mE1ULKE39KTjvTTi2S1FaOG5QhKD1nZfKr1BaCkzkSu
G9pQVnmrm2UV4rxRbzrabRK5fTphIiCQazKZTfw8PMiMO9MozvNVxM+6QpnJs0g4
QdCO1IWkdP7GHjxEBGjv/L79ysbb9YMCyriaUnWWS3Dz960Rx+BX59OlYutHOXp2
wRHVUpOd7iM2h5Ki0Uqg/jCzZ7t1+2pcK9l52SJNE1J4CVJkRYUkbByrZCk/0Ist
stdtQpkc3MfQIAEKFByYRzUP1CfUVXc0ph4ECDJdai4xBrSmK/5aTAVTxXEB0tSS
t3HCP2BzbM2efNlXU3C6zUwsdVoNOnmFawEUuUONjVO4Bq+0vsn/OO1n3zwxKtWU
0LxpbfE+NkEJMo1QDoa45iefRHPC6M8p3kjVMmwqvMtZ/uWBr9AUapjOOrn+ViUu
cu94vt9j9nnhKua1zqBEWOzz3juQKMHE/jihiiOza8xLsrW4oQepA325oaZCCjhh
qL9uE9GvN1HBFK2yhsXsJfn4hyB2Lskd1/0nghrrjVax3e3n/rfuHzUp0rxzvIxz
5fu3/Yz3+PGaQPLNGmVoqwBuNYt4ElO/T3L6LmBjvWBs5nrN4qIoGIwoxi3DQC6l
xQx62YOgHMJKmRnBnYYSGW1UJo0CkZtuokONXRxICDtHWsDWJ0kd8B2c28kOdK/w
iMgeHnc5Aj75EK/uxvZlPIWw52swFYeMJ7ARzqW8x3EKLOJM5LgFmhgbDLLT58xr
zd5QJDHHZaFKDfq7wg4Aa+2V3/gdH8130CE4aTpqM6RQds8tM640Teb59Le8sWs2
V9d6B4M13d8OLQGE7T/LOW277/jXsLLdLk5Fs/mL/RQ6GP72LibKYqKg+tvWAxAl
Q9F15ROYdI5pEwbZg+lyQtHQ3QXY6XHL8nm9ohx+Fo5jggNWOf6loNlvlGRmbgS4
4S7Pc9sCyx9QcfF/FHx0JaTdd/TU1EHBhyTVVlwgbf0eryhfwz2buO941nYdi/iV
uEPMXGxS8h9AFV2HJACv1uKc8F0btSvsR60Y3XMIwFco59CNrpmR4Xh1kAzYqQcx
VyHaZSbvGihlP8tIsNfeko8/EtWkwoGDHO6IRL25dO2zslMMlnSsx/e2Tc4/xA1R
60RyxQccSyHviYyD2c4Dyn0fMT3wwDC9jKDG69NxKSR8H6KG0Eaw5V0ltn3q78TF
QUGvXudmKOSO5ysrJe7Qw6H9RwQ34DvNUfm4WQGMQzY=
`protect END_PROTECTED
