`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pdSrrfNWAuZuAh01qkMCmRcutJbCl05ASULDaC9RWARfMSvwZee3hXoAMSwdSJW0
gOSADAulPYG1QLZcegFDOZVPuK6vY6mULYfNFSFFmZjKUdf6mGqoXvgNNe6WdmSJ
u9OQf9IwbxO2CT87KgTyiMtBbEYHt686FAf23NQnQYqGUNMlpJpILvh2hEzEEbrL
5wRPH0K45Twc0RpOhqlUolC0iT212EBgIFTryXe2YoJ8hE8UvqRHkUUmwrMzlBH4
KbsJmwi9SZ7xUD03ex2seC8LVD08PeJCAYqBFDDjAvYOO4EFFMW/8Hr8Ar76U8y/
5lXxm0AP+TgPJ1PKw0y3xSFM7JfiwLinzGRr6a7+CDxolbR5TBU7M0/2ZaGleSUX
HdzXLTEizYlmpef9jN9tjFYcGfj8tnLQ8Guk7cwek4u6q+0v+kxLRrc9rj/ms+4O
wjS2QMtTRmHTzr1/9ULeeBGcfyjB7MvG9i2IY/DXBwsyQJ5jsxsXU+TnA0gHJqa4
2aBrtMlLyd8301knMrhIsHIEEjNPvnoRmzZArviOBuKEWOvZ3G/n3y1RaYiVizAC
9oPIMPg4C3XTnbklJbrJ5QHxkhGgwyzZPHroYEdsdWhB4UgjJcCVytDjPltsLkah
k71PjGGKc6KpscQRDSXQ6IlG4dqufTqRnF/86gg8qqgrMmYW1yYnaeM5pmLwkW1V
4srdhO6Le60gnh8Zs5lC9LIEP2jYNiKVVUYyqwLvhclnEPnyr/PyCjztPtCiNGBU
F+7ER48ch5+peLoa4RtpGAN1hr0rgtENP38AIC0FmQw0N4fmrRS7wj+E+Ug9+DTf
zDx4foweIIjfeg7C/DVJ4VxyuMYoAWiRik0J9JJY5nvnGr+5x4bBGvHiQMEbfo0K
3RRaAe4H6c93fFo5br1YSt08t/1ay1KwgGdo4KkkYBSg7F4hsWAH3vJgjQCCyULf
vLIqiYu8Yp4Nf3MRJtLvEa+b1lKjlaxs1JGzI9GzsyzXAX9r6+0/B30iKpOYY8gq
+ITKKirD9u2cSZrPx2a0cY6Uiy/nm8eoulZn84heNxKE4q5dezKfLm12iHrQemYo
TFCWPYj7yOqZfAfli3MtwqsVXO3fk+f5GZB6BAd4depryclxDXA0t7dMSIjCYoFa
oM6tqaWIaYzQ3MJxEoyUQBy8n2Kn4RSwX/eh+CX9mIut4pLLD1Pw6YGuixwC9m0d
t1/ajHuJ6YIzOInSH3kYbEVJTB96rl31Pv30fH/ko5ASS5NMXfKJrvuo1Xq5QzA7
4eJ/TNjze6riT+yJ6RwvtPuerO8R3+4jVdt9SurOlEDIvRQcdgm9br0BqMr+2wzy
J8/gDidykcIjrFBK70N1uYZA0UAarboZ0FvVOp4Wcj+Bd0WIVIqXqUASxwXuctv2
b9QyqtfxoZoBood/LdBpFNfkL3R9ynTPrdM6MhlsRF6s+0O2eQMUtw4cFIde2vTm
oNqFY1d6Ujo4JPSzNMBPmh3exm0vfK4X0A5dztD/m9H4eL1buy4cPSJfw35QLLEz
yyNDo0h+iPTFF1OeJ/t6H8n1Dm/PVSQ3EcnNbGqfYokOMXtq8qFH+gvMwFnEL6an
b8kooJlIlMErf/foLzHVfNXDulk8z186X//R9JU1GIpQ3HAJFL7f1N5s0YiHAlWa
gDad9wRT1AWSDMiNP3YI4ljNnQQUP3nX7bdwD/9uy1taOxM7C3HbFhwbZ5IOwYcF
FRqQ8LeMPyKDUUs13swPhj/kw7AEUFru/HNMjGn1t23rUKK5aby5UuqyJK8SgYvk
l2mx+Ct6B20ZZ3mt9A6bbwXHdgAxyd+vm1uVxFMEjFRwJ992tfoaDSUZG1j5d+pV
JcmFdNMem8x2XrS2yDfBR7gwtR4PSJk2eUcwL3xCtL2HyhKZ7YqE+1OstabpVw0M
fXEGSQuq05dwNSiWSpTT+n4Si5QxZlGgp7B2Q+kdm7+AABuKcvzfI3NoVDXmtaKm
LsQqU29RzLOdxEboXi9IGdUgBIgkCoNsT0oTCbIHnW3bkDJFIvofycvZw7z7bLfq
VmTmnhzaiHwM4nStj1T5KbDljei2do/fx0zICgWMXJ9t0fmbyE3uVK2/PG7xC2ra
d1RD2TfMRvw2+kkqxCSKZAEKKGlPACpWtFcHBT9zkbXTI1zFCxN9/kv9PD/dNepC
riCMb8huuedG7oZHPuQKdgRQBv8keefGHktHvJzFF0u2S0XJ7OhHx6rRpVAOUeqE
g5d93dUFsi8xtd9scC31FN7RtA8+RJxkB+iB7qmEtj9tymGaPxPmWOMUUNExOkDF
HzgCVHuvWFzhWO5db79Fn0P/S7M7slsUOaV1bgoG7oIMnJ9AXO2Dcltfc48QkycT
zQuUvH7wbxNvuAGOzVVLKrCDpvDhF7Bea01deUoowCXQ06B/AeKZGCwUZlAYAg4D
IujzLpx5uhGYkHttDWauGAng+tKOBY6EPX6KV1u1Ozv+jqBVFk1hiwEOwZKGH3g0
6okXasHAZCx2k2LN0Yem9K40HBS19CqwTEuV/xNwuEA72QBqHzZSOGaSZA2Hfm9n
b75kc7f/vvVqgcB2avOX289bAI0dyzZtdyXZkBuNU/ORDNf2KuFKsO4Mb0tj5z8x
UqDaz5iKtW9ZoLqZZb0zDOEqNMlqBnMu203D7yyNImQx150r6tWl6lWdBPjR8ZXM
pI7uZ4sYUEFYCXXoQYqickvgVX6Aige4WBKwDCuxm0r3BD6Z5KB+Te34ix0BBBwG
0dfJOLVH1fQB+SQzrPpmiEk/nOlI1i0yNE20+nVHHRlM9mXPL04hZCTekQw6TQef
6WoFmIv4WC4mIXywMig6QiGoNv86h8/7a6mKiS1T8NnQmap9iQkaH9A4ZQFKTFBI
y9TIciujVIQ4CXHK+9U+PY/0KVrAvsVPFXRE1qYVMjfWH9EOcDuONpANDuJEIC0H
jQib0cFgcE77c1jOxe8EOmqV9+JoeHwv88gfbPrwAc309BkP+pe84cjsGKhYK93+
EoF0Fk8mI0TwVaUAcOgkipBXoLddOM9/+8I02FFmCte4DZk7MS2ovlPVeOHW3iG4
2GNx2gOcVR2VbKxE42qARwn4u9eW3CASxzA5sHbkneLKMP+6oM9Wd2ck3LnEtnCC
I52wAnci7aE/VFG0IesXLR9TljtCqB90QgA8fBcDAKsVq7QJ44oHUN7S7BTj22w/
ng6/kFNB4ZlHM/PqjKcijHZu0BseEtgjFkubqCPrsOCHunWEV9eo0XTLP5MKdNov
n7rN6soX6FRSJW64afirC8O559ooE7gLyovKgXhnNv/hfU7uMv7kwL4wh2s1KuSU
VgTXGboP1xUVbKf5sl46bOb3reS/QKrXo60ulAB5YFkHf8O7kwq4j/D1V1Jii+no
Cuja7rkpvaWOK73Kq1gfBNCSg8fF0PJLbALzeD07BN9s+HImjvpraIKay0PQ0Za9
DQJqGZuNLvfKRUWFkjzUG+Bj8GVk++9qv/jzwKdtF90JL8lWplsSwMP0gwxv7Hj4
Sg8PNyyu3Xl6vv2ix7P4/TTe0a+mi+ObHO+SowG4lF6S/dM9lWEtMWZnfkE231Q6
fATGhZsNYOu/MfgxWo8dnp3cDzueIGVXhvAOHMiFfZchJotBYEF6I9UVdvFc0KnL
lNGZlx/1bbjJpgoJk0T/F602Uk7zN1Mu+UhjBLEkfXNYwhL13DuYt0O/YlCrfObA
XjA2l+0V8FOlJDLvobB6+vsfiqO/rvoRiq9lpDtg5gu6UziWyK37UsqHZa+QGffK
v0LT2slfyXs9p85eEG4x9slS2fftfjM51K7lPkAJOUaaSBze48b5W52DVNNKeWA2
mElC5ZUiTD4R5bPgx4niq6gLSA9kZDgnBhSueJC+d0yBQUETaX5fn4WfSdXbfYqS
NO5ZDSEnxseYGdtFqPqRxMCyQ1Fa3bq3MpyOY+hd8ue/xMPOtlPkL2C6PccIhw7o
kXBIMlPTiYWeQT1XnX9LS8cy3uZVU0nSKEmK2FRKAqycZyJ+bJXqJdIfTtIKtWwZ
7uZzccESIGIc6udKHy/EF8XN2yBm4UfEWClHtn3IlW7PoortzUbarCcIJr4zJcpw
q64Y7blyYp9Utf4VcnGzqkH2eQG3Tq9dP6U8ivQASsTv75C4+K/+ffB/rnuzh/oF
rLw1jsgT47tZQz7V/XhfkdgKfdM29cVUMthdix5aCfzjYM1px3J9NUzTsTmMwclU
zP+fyEWRzMuWxcnBFfAk1k9EQqll4l3JGF+lB4vgZbbqWiW3NprqkJMogx4M2zod
X3fChNo4HYcTk36SM8dzNs6W7SvRIoOCVsYeV4k0pqg=
`protect END_PROTECTED
