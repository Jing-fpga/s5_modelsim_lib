`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UxWgSNYwp+1ohtCdjnMVgDtGpGEy11VkfrRzqPirVFTSqkcM98QyJv0Fj9X1lf6Z
CE2d0/ImfQQCz7Y7gUMvlBKPqsGe9vMqkrcn0QApw3bX4DbbJFX2D/6hspI4mcxw
dmYbdz51ZsRf1csIGUkThrtdA+9tauNEhy8/kXSKvB8gXJZ6aev+n73JmFOjbqJ4
cBNGdKWh5Aofn+WnLuny33g2C+Qk+6H6u5/v4LOHleNownbfNa0tq28v/EoY7OV1
4UWWFSn5CkbTDoCznxePL3EcQsMESW//Vq//iLeJAhlYrEA3PgNUzcOVPIjW/WOw
gn8RTRtQDmVf6jn29xUnSVaXxKHQoeFtQ6xsrkThSwvgbXA1PK9f1tqn2O2FsuJi
+VgvWxC+iNA8XZT5aMDioxB+YTBz/1xLlqmMuqG3oj2W0Yky5XZuSgAhKdY4g/j9
QTLJcBe4zMjxRcaOBnP5E2w5OtVPbp6X2ug7uctO/Tj4Qa/xhKNdTmpkRZopiIBj
QfwI2u5kzriuA2Jqs9tymEeILdszLpb+GdwFknShctQub0Yi+uuXdfMr+nWY5kad
HV5VU35oStg8bpBfFSNbn4PQ8wqBzO5sH5xs7b/X9rMd7sIHKZFEgP6l4vvglbtp
+3VMa4R04O8FPxCbTHHzcV1cI/ndvr41tQ9bg/eQAGYt0RphHJe1sgTJ8wEj0o/p
LngS7DXaZQiFlQrwSWn2BERSaAuPScKIuolbzHMuEVXmDKZcZqfXO3H1y1LaN3JM
NKFkXZR5BH7tQ3HSs7i1GSNXgRy2eWLi3TY26s6ZLFOSqcMZ7yQWcvqJ8yNbKgvG
HdVvbuqeF4l83QSvwSBVGcW3Am0imefS3Cr4cu/6ylJ0Utm0JG24vpeXWmjYdCZe
u7rC6EnCTIC3hs2x4/AZbFvPUlIbYCVL7U2GEO2gI34AjNgda9/ZYsypqig3N9L9
6NjKVAjkKnGiJAMFl2tZGiJi1BetxkGyd++gc2Pavv0hYKYL+INF3S+n76gXHfvW
8K7zL/ygBtsI+g6SvgV60/uVGJMpXcDB2SN1/vn3qopmRj0fBENDI36HtchSYYaw
vVvVZvLb2JNj7eqC8d4NRHIJZ+mAxGwy5anq3j4xnW8gcUyiIR0ofoeJgtJWgz25
uvqM9sABEWHe11hf85+tqe1QuVhk10RSUtPT53yTUvfFAagZxkZGqKFxl9UgtcTe
N0nLYpNpwSuUo1FO82tQMbAENqExOW7J3saUDjd9yYkEQrLmJ5ZE5FKfIqfLy5rW
iitdm2Xiz8nGj4VD/2EW7PKkT19YzRth3s44/fdm+ooo/Lh1AAv2L8bV20J/7qEg
54s11CEess/FAhh1KPg0wp2AgdnoZs11dCh7Unx0enVEsfaila4B3uSGssR4zieE
95AEkeIdwexCh+grbdSLJG4Dtv/x926xWXh5whogr+tIoWvrveRrBbToY3zW6IGc
vJ8ttcxjn33X/9SuaQI+DhbDxgmZfurH6buas9MN5LVF/52V8gBzWsV9n0dfqDVe
XrseajdNVEe3R0hrXygD07nxdeEVD8nPz1HQgLwWz3UWHndcC1vVvd4QHNS1FSQf
ptMBSXj+x8PKDlFUAWoI5pfB5otR2kHplC0FOOEK86EAMXU1/uTnfvCYNjsGCRBT
zgUVqi62x+m8Q0/JdWJVgSZiA7AF46HaKpG6Fo2WnrPzErSQrNCixYWdlR+TAJKd
uUeF6Lpr4jYeD0TmzE3267BXz+esaqganLs0+n7j7pg8CI7LZb1v5CB/rYdoBuAE
qXPbTPykVioeCrCkrHj4BDY3KSQp2Va8M0wgnygaqOlakLuoZhKXd10PpPdY/RWY
vF5Wehiv88dL9qdfPdLu5g2YxLvz23s6Ia6zbOZbaAkBhOapVnmkrqa9kK9BNjXs
nhEFX82SkPa4XNvdwZAiLuxQmGTqQ/z0lEbYqdEaYDvDuA8PyK3jc1Jar1sAp23Q
2j6duiVmnGkjm7jWaCEhIMLOKoOWlm3FAStmSWAWs4urLbFV6pzC+dauB+dBEpqC
mf6q2aA7BYJqnmizCyHqLXB9W0u2P7uN7ZaiUi/DEqfnOuY+zYszxUlK9bAZJHHM
NhF5QFpU+uh6O00357v1mg==
`protect END_PROTECTED
