`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o0vllSGj5a1Q0tZXpgfS5QthZYphoO3bpuMbfuQtNvSPwIJxYgQPcXcAw6JQozvl
4AWiBN1NgIYi3BPn1xw83AG9itGC3HxoOHKbDS2fzQI348tYq82iPGFE2VXpIaY0
kcpk0BTpMFWaT079DDe+DE7RyBRuwvXgKusD1Mwj68MvzQTFti1yYsblU89pqobH
bMWVnBn0FZvMEJa8uEyEtSHNxwEY9cXT6eYBlNRIx1joyst0NZFHJMohGKoLMftl
TZwOmx2V1V5LETBtnTJo4D0+eSclZ6bcBcLj5u0Zxdvtzw44iIX3RholczvFX9pI
QpRkQ/jbDO5Xv5j2dmEi5JXgV9xxZLxmH/Y9LmW2FaC9la2FNdJmEjuKCA5HPDND
cZSP5yKHuItUbBNQdXT4hjaJ32HZMI/u7M/Be2OP6Vft69ZGwcJkqwUmspuzu8Ui
Ay6xOn4k55962wvVBxjuThYNMBiGEfgNttluzSmWQzmN7PNuP2tqV14TNyabpHE3
YlEfxeOGOQjBCPi3bYQOfw==
`protect END_PROTECTED
