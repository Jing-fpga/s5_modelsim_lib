`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/IlKvB1ArWTjPq+xLLeeK0Jg4Bq/A1m1Qi8jdRvjfupOpXo+M0jp6ldb6R5oFAnh
RID4wdF3CH0rH8cDGiyMT8HCRvDc9d65Njk8iPkS/zJwbpPmajHTNzRxD1J5qqdr
mxiK34AnAjF0h0vi/0QNCCXEQfayeql2lsjPJcAmvxpaVT4Muhwa/52mqKkOyoub
3E6ApMvS+RqZWSE991/e0FAblIXMtkv3NTR6t5MtDeteAEWAQkZcv9NaNtN/hmGA
x6akkUbd5eopg8mksX2rq4vN+tyMEeCCmureQ0JwatVPZpWt8lmdHOcV2lv2LUgS
67muaOqbLhPBI4r2JTCKa2uN3ybVWKVOA5lja/DMJRErndjFqxnVPorJlfl8AvHi
cfd2k+02BqmdxCYJI17DzuVQBuQawr5b0ti1EpUawsJHvPMLNUfF4Eut0YTmDF37
tUHPjCHeoKGCDiNs3KYduYu0SVL9167CAFAv6lHT3hfN82gKAAxFyE3gKGdKdcaX
zpTJP+LsHwIWfnn3UtgxxWiwnjOqTswlMLplBg+lPF6PM3AKMct1h2sWaWloRhxh
w17GNGjl5Gv8jS31rx5GpbZhmGBWJ5rjoaY1H9m/kConEfOy4KywesLdUzDgGy81
umg0d9Vd6VSgAwqdPsWi1w==
`protect END_PROTECTED
