`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/4JGwV1XQ9bSZVt+PDsbfm5G1hwiUVq385f38rjWeMjk0qY8I3EbHuLUOjQlPs/0
qHLumE9b7f2+Mu6Eh1kt0vCSeD30ds6eNbRMak+fkFqUdIaMmYcf8rVAAQ9Pba2w
TAWlThzJsZlpGNcDM4CoK/YhM+x2QIeVMPDBRDvyC0k0vNt6mp6WBoAM8HSVlwbA
E3we9wWn5Og6N3B3LL9pQAJnD2d/7BvQf14y83/RZPbktLjnCNoBbeS7CTWquTzD
+p45gR21FWh0KPG1ylkkOKxVQ8LYUxgBkT3U7a9aJ6ZEx1t2RdU3rMMmyrQ6Mtaq
u7G2486pSgR7cpkxI8Obi34gNCoR368O16vGzucBRiC9Lqjl1ton3x7ACDf5E2+X
MlP7yTjCBJqeQ7UU7U6o6ZOg3eUt0tv1FmHnWNYzK+CL0tns3UoGHrZG5zxPDydc
s8gecyf8qSoEzhzIt2Kx0jSsBaQzDIJ5sZ2r+0n/isREk5aTS5/jIQmjtk4Nq5Fz
f0WjCotcnrsWIrZomlkhO0CwSjwyk4tRgtZa0kGg66mTzAWRRD9277m+w64YOfI1
nCFtdhlg1NDojwoaCdfHo/T9SBffHHqnRJm/nYW8ScCD65Q6KB/lAPfFSfvXTIvB
zZal7VKnMnHOaQwtYn7tLpgO4eh5BEwJ75tZN3CnacGeKwEav3IDfE80p/V9XnIC
4X4GLnxpww//7isWAApHuEJ4KeHNKHxployNo6Ma87HCLDaWZhbGNv/UpcIH1p1w
f/tyF8hMQcYb4t4E5xh4SLWjZ2kBBX+v7fQkubSpVAkTRV4Tu1MYLixS5bj3KlsM
GAOFaWTciCIel4wCp62DbswAFWhHBbpiZJoTrhyHHujX6fFJ4okbfPRKMXHqk5me
l0J99TFisopBt45PtDsW7xKLiKVhta/MydgQVKgJcxNciEwfoE5HSkjF7I+pl2Ph
nc7UjFKl2+DvUqmWyu+i4A==
`protect END_PROTECTED
