`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+/r8q+rR3GkFygIxTjWqw8hQuvqnoDPoy4n3BmvHjBoob9Kjn3C+z1VZMdPBCK6G
PwHO4XxgR/56wHtnPFN7Sd4pry8XkSx86bAETCk4UxbD2JfBeJEszzMRhfDc+zQn
r9+XDkryPlqlO2RRWb/RB3aBie+PNlMGA1FuvIOTuj9mOajkHvSnmMbX++IPk/Yh
szwflH1n5VsgF1hjPiWgAoBeAEKBQwaRE/95XIifnIdGsnVwyaginoa2IXZAXm9i
jGE1lVxyaTTT4lHiaKUauvzAy2RlOY4UWIyHJcBSn/ljZ0Rhzi2GkSwjj1bJ9Ife
j3PZZWRDh9VyHcPIix5a0CqciQ8BLQaeEmRHyHp6dRzrUWgimb2JKgfi5RgfDzf+
8o8UQYofNr2BS7GWQ1isDhSUwD3AFjMvckzPCi/bVhIZNkuhwcr82v2IAbmAEI3/
jIrRUIveB7OtVIAWwkIWt39wKGdD8xe9S9o8VRpu+IYL3A7fR7T6GyIHO4vycq2+
GXORd0EkXrsQ+wI6Oi3/VTYvPbPZ0L9HjUOOhAjWuQvBs/HKbsXCNWO9JdjgclQg
UjzLvNvP16KvbZXbyS/rnKxOzZgB4weI3INazcMqixTDhditjRGUr4IYgNZyIEgh
05/KaNO1rtR5KG9CYXCr0g==
`protect END_PROTECTED
