`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jzJGoIMBRnxvowU7quc2a+yfLARKzeRVTCbb5n14cMoYBCZnvCDLQT1pv9WHrHXi
Sxlgd4IakPLCG9/z8GxJw3lL5TcpA6B9L8DggxAR7AR5REqcSZW1sgO2D9B9+nn0
Xtj5mpEN18nNJM2QxETtChRDIHoPAjrVfrTZfvqj1AsLK4NSJOUUz/KavMZinJko
Pkgg3aCtSoMjWyRaY5f4bIoNK0vzH+GYn8sRHvnW438gKfRjUbl5qUGF3XrrqiYM
fShnAAmfzkMh2ieG3TcWPK7wK9DGiaxWBIJfIctpe11Qcjp9x5nmJFFKFr4a9s/u
XaTvO3FB3gvY8dvdeutzKN7idoyctKUSsNpQmymrR6BI/TBlYBlhEtn/VbiTaKB3
lWcHoiva30++CbDdRM5KPhIq2WTHQFxI0UpVowlEnZDezF2eXvYmbpdAxJEoh9eV
tUqTOIif/oYH1HnTl2oANL4Nt9qhj+ekK8ELToVmbD16MWEzhwGofjj2aLin3c36
QUauVz+6wKVQ5rejj1lL1dWia8rmwyOBixR4QIJWUUP/yQsdIXnAgB6CmaGPSVDm
0LwaJfvXG3r+3WM4V5H/xnfFpxQF2AZ+RJnlgFcrS+/q8A5CjT82NbP9V1AvHUAo
epy4o/6jH/229xxAT9SCPWiBj1kSWcxZEPx/0QmEYX4Nb/O8+sAUoko46O+Z+I/9
UVj3mvyg23uyFP1tuv2c+OrI9Xsw90aR36D2G7NOljHD55u/xGFUK3egyGzPyl5Q
SJO3QtUGX+w9ADzxi09SYA==
`protect END_PROTECTED
