`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Rn6AhjekX4qNBgTSRvkUpcj1/g2iTBHshPgqi6GQ35EkQP+2UJOy2Poh643HtHM
DOlqhukZFPX+J5hBIr3ys0DGmoCVk5xZCSWhMVl63tEI/23Hb/KHf+wqUu1C1qAw
onx0GVn+Nq+IVY7mWtXCVuSYnnGZ9O2TARBZpm+r6/+ZKPSxDjO5iv1ORM4tBpPU
t/C0tPl+WZ0MWTg3GNVZ/hZWBVoNwPeQspF1goMNQoLeK2ZGcbWQZJTPEZ8GP5eO
so8FuNB3VKaMzkXFdW2eOiB7i/VoAKvcI8ev5F9CQ5DXiOnCOpyodyfMTVKH2iY8
r+85KO1wH5yDM87znBe+Eglsb8hddKpFoQV/haeZFVAtrHZfrfI6KBD/SojqHO+L
+guAfRQt9edAphLInaXwy6OdZjBRBSrbeMCnu7eZ8QdL1DGFRupAI/6D0C85VA0k
HH7TvD+rpEHAZKBh9mkpcNst8ZoR2rW9NsZROoYWit4bQdhQp+qmqjOEKMkPz93N
hyukmpCPeluY0Kox5ZON2PkcQ56rodgv9j9Dxpk4EZrCUu1jb4igMCPin5JS5r8H
WMsL9+rXoMZGdl+EN8Bz+p41H9h4+/yuU92TpSCZeNmh3Sgt1ecGm4KdzVQhq8Ra
BX6onxGfEKKzWRqKLBv306WDTEf28df6a39FMbVS8QSPo8m1aP8ucf9s+lSQS5+h
RFM6Z/kPIW/SC8WbTpb57DH/yI7zyUfX0QVXsNlu9MJcYIYE5VpzlMAVN0RkOQLu
4ApLGopTmBB9pdAeULuvgQ5WdllVMtD32Y0Pv/xaj+i8vTlbBEa+HdvITyD0oALx
gN1Gir/dVP/MIcvlTK3ndASGOrMv17219xO9EcfbPFxjIrahgH2Jh10n052iyp9j
Ir0DswA1UnfiKCdoo3v23JpMToLSOqxE3wV/Md2R+A43MoLNcPYvZKbGJqBnJY4z
4qKyD96MV94xy2/20bK/BjN8Af1zVsKD9/A1ORYVHbCLHsOYsegyHzgZbmDYwF9F
RLo75JzHkGRaqDaibNt064piMutG07Z6LRUDTER1FxOBIbfTXIBeERh3ckIb0FZQ
2DTiRbyklNIdr27R65rOJeevUPxdbanP67gjUVwoPpaisx+elmQawZ0Xk6X7Q3MQ
KZFCrfMR21IB6YZKoFtGJClbvYVeaRBGUOdlN3NZSHAsqjfAYU9SXGiaLk/M9A9s
IaKMKJpFutVPJVnfDnrAGFqvsydM2sjrScONQPbsWrv80izw70SBeRJ6bIbItd89
FlEEnCn5IW0EYQNz8oO8rnFXZiQ1drl1eFG3G/HfwFuUbu63ZIaOx3LMRJiET7Vk
RA1in5AYMkywvCH1cKfTYN+umFTEM1heHqPr4sn6N5T84Jk1/ppDn8cZqCVFpotw
7ewrJLz5UzItS2JIbe+VZcLSMdKvmBXwX/p40IEN61vCNshLdnS8DRE0/+1/1e/c
y8JTGvtYYpwVKsO++mK5n8rOaOJyeKHXnpvzOGcwC1o2E9h3wKxXmi7BEwF8aDqk
HnouljWK3z8Scb7hq4EPmqiB6BskKX1HxY3xl3ayomKDBo+YBJ1CXCKUw3HTB4d8
6vd2diV4dXmLsCCucjbWp8lAsAIBAiNHew/XgVEhAUQk+QCKfA/Y1kxXfIjL52wj
3LvCv0rHZ67S8oai9MxE57+91E2tl1PNV+G79l6d1wrRgodxNzdTJqmXq6M9LmNE
NexxSrpWbKodLS96I5rfqCw8UOc6RtGo31a8uyhRc4r/sMd91gB5AfYN+AtEw/c2
e6MtfLym9iAyG3WESfmWWn8j1cjQbi0txVNyWxoWXjFRPPdtrXDvpTIC8JDbCTEp
/JR/FgfnJ2RVZW6pCZVHbkt3Op8/omYSZGKJ8Q9YSNGT24vzUJPZ4GX2kQzqq3+M
o5WCOm6I6NLc+HBwm0LpH9riaR5sZmreBv0RxA8PsRNrjxOPeXPqloJTqAZ3VCYn
NfJla0yJ39jguFKeC6gDIOfz0EcfsYlbQKgKH0t/U1uMCGk9VhJbujgua5V/3MoE
XFbgjo3x+UGH66XbK5YDv7EDdcQ2mpNyfCHDlAw2MXwhVbx8RUPNlr2nbH4RirdL
mnG13rXAAI6mgb2l92xs/CRFnLAsd7Ng9BD6NOw4OWhYDLHDZE4hYr91U+eS9kWk
CGu3SnP2KcIJ+l/2Ngn+eXeig/oKOQlRge7BL2m6DF8bZFtnGzwFOCLCVkfeLPo7
+fZnpe+V6mYQGsHfhOHxLpVFUehpUJo32rXU1b7+PLViREq6/OjMUZXfQKajy/yJ
`protect END_PROTECTED
