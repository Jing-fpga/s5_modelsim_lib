`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pR3loVcXEHco+SDFzIFdZsU1iFMuOUk7aNhWRvswivuYKBIQNc0l7Hg96qYPOPY/
+fP2Y5AZekmR9fi7zFLn85dy3AXemVmKfANOHpN5UrHhnzaGSzi4OrIshurtZpGA
SkF4TtnIC+a+snVYLed1Scmd2MCsZr6PlDlb6SUnCCbZVWUvmii5hhY3x4WniMVe
KbZNS2+5pni+Ef0NYAfI3AaQ3mzLQ6iljtGFutyEkCPCSKiKJanWUuOsf4+U9mHI
kGmt+StS2gacJG7YpyW7hAdffVLjj4Q18bXhk/prUvCvOS1Ws3p/fAXS2JMGcdQg
6E8W0mIfCvFzXWk+ZPjYOdkfde67MVfaQpn+E1eQhzckNAjjAs0v3LS5h8Xspvoi
NJf5/oI+7MfnHRpoGdF9N4smtkA1WLxCbkKpabncP2/fDqDH6ShaoDucHWQQsbQQ
D916lsTyflQSkAYKIoG8AqhS1KOIBXznpuTsIKwbCxGFkSw11gig3YfjCy2sd2Cn
aq0uji5fcM2NUfvXyYTy1tZsAvt0EzoEf5vAHi4NtF9/VAPLPL27LG9WJs74RLSp
ClHUu+aVMOlsLMCTyq+yfPGoufKzmVyAyxN80khndbbTeFdeoL+GXPViiikqbFY/
bu925aY/MJWYaskyUq7/AT+wxVIs+oNRcyzSex6eeQR+enm1lDXTlZzI/drZ6ORL
gUvoiit3fhAUnDuYoGZdgMQ7yBn8PsYuD1tYL00fECvngefMNsptmTfpAWMOlgHp
G5sMmPJILI3GhN4VACu58jJ+ehsnwQaY0xIBmzY5bZ5sWNy5FYeQH685eks9CKgB
rPcOZMYJFZeqIZvJXrwqRhiH03i6N3u/4xI6qEi95E2gJrFBIWSzOw+sO6P8afrK
vqk1FPC99zQ52qzS0rhpll5cuT8n93u2LxBrjOJ6x+hgLprEDAF5DnZKfTE9Y5XJ
CB7Bi0KxktluF6PjvCRVJ58Yx5G/ohDENm2tBHNzWvNxFmvpNgLQS1l9/S0fJxMn
/D+cAo+bHPGfglrmWPmJUn2n8eMZp+2cctM4uk21eXzgzu+/KL4/Z1ApAF3ds/Sw
HRlBeLNzQWr0OObTTTRHVFCV36XasXYb6jw4ow/7LSBsDGFpdKu43g5GXfBb+Ow3
EvMHLLCQq1kD/g6KXKQfLt+KD2CsSCpX80+aS9TzLj07dvGIERao/K6Ilp7iOzBP
xoiejjZat1XRXcJXpy1bV4+rLmO/B+xL8RPUo6gngR2B4JS7qhWUpLpjOByhVGtf
+gUneZCOvm0vw+vR3MKgGjapx1M4H3SA6bskeFvt4pCZEmnokHsWwmRanVsPMt9D
IFCxedK3ADzqizmIABP07ao3u9lK+rXj8HK2XGh8IQOuvv9j2ufKrFlh/33Kixqi
FmzFqyZ/jY5gwF1VBv6harHX8ewjaurGMcuQUzQsQLl9qBgDny69GimPHcDZlndu
oMHkz6u/SZs2JsWh749ow0ct9SPe6fTbgWUWaPsoiJCa08ACQW21r7nPAYimCrgy
MrRfku86iW7bSy46DbAJrpt/LnVTOf+JomerQeVzjMxqMtA7hwtm5i2kbehBwX+7
UjPRHiM+XQjri1vEu5Dv/kBE2petCqbVHd754UOGBogqZmek5jQcOfC3kLQBUjyX
Svfgf2QeXo78aR8TPvZMvrfIQOfzwuYB78UHFFWsqobJ+L+ynbnSmo/kMR2VjbVF
XygGU8RuDzpdfLMNth6lD0+GwLgPXff0FJfL6j6b67K8lVEasT3374Z+VU0x8Z6s
rM+2gKyzreDiAPnbaG5joaDf2be8MUe7LiQKL1i/qlhcb4UTfw7yzdJ53MlqUNFw
dEV6Zn7pxZ7ZflXGNj6hnJvypqDET3wnHlTUorZm+YUspunOGpyi24KsqghCu/Sq
1YWnA8cYVnEohMQYlfhdRSbIw9MfYvodn/D3dIPmtC/+ijGWQHUOysqG9KwzsiCq
z1y+HFkz0pANpzNPyQ9FGfG/Owk/m1WqoBYylJmKpHTSHg+EOpRmn2x5RLSg//dW
ZgQ9Fx08sLVgr0fjlWziyuB0aHB4fngtSDc9MWmIJhU7rlWw+tML+f3UpWZRnVph
hZ/0fVA2vJz3U4DZZ16fWLGx86BilhzRMQ79/bHKkdwEUMCfBZYiivsEnGbIIt26
aIeB752bzl+SfyQ6oeegvgRSRwzhs2GolScX7Yakg24+pxQzmvv/foIj3xAlgscL
jX2+oynadYHVfLDWEZxihZjAEAtjWlsEWKMx+j5dMrNiGhk3ZOMANpbx65Wz52pV
8r4ggrQGg5efWGKYmEDxpAQM5LqybMSC4V3+mRfxujVHGxkyMHJc0AlzINGeODxv
UISTdoGH21e8naJUY0gIHHYmLHSXZazdtsczcy2+BgIotLML9nHxGCOz4bot+Zfr
4kf7C0Qs/uStz+b9za1tdOJzqAlfHgthRfCWm5+NHMrh0xZ6x+nAE8ruXl4xnM4f
pewcorNPr+1HKKZYVTPDrXzge1a290O2weqR4wYiq9arTN5j0MOLS3nDtYwWJ1OZ
lyN8xrGYlEkpYslljzXcpcytWqPqiWbOm5Dcvela6rFUDK8Oa4F/eIJUbYHpzRGG
CcIb7SlpflKzBpxdzMM3ER5r2UVM5gi+CPIfUxxC7bYTQemtjeCqTpYGqyPMz+OC
hoXhGnZgiAA2XpWsi+rJXO5LHQ/r26lTRDwfJOOAVHP9FEOcTynISir/DHU74wzo
HkpVsZzAKyku3JnyeveVrrAVoFK0+/n+wqnlP+vBbaU9tvMuslbaRoDhtVINkKyZ
PXLQktUJt+J6rgU4gUsm53GOieYRmoLngZHSsmGCoBpqmKTVvO4w4W+lOkGF7bph
LQpGKGSU49FTuO4yGWAp319iPGJSu7iiaqUgCe3tU/PYWlE+xI+p26E/oj0kiArl
exXPsYrCiVM/WWjXYY+GNezFcqqCIROF1gQdG8vdel1f0c8kKssPXF+ySIX0pbVj
n8/sC/jlYZehFRPhf+J184tjO26z7Os+q7oF3id//tv+MtzF9zXKbr4TNyvtf7ou
QRt/CMtTXeK56LAKKhRfwQuEj423bYGWIrepKo7qePBcVa6L0pRpOIRDozYkDjA8
dIgKl9co5OULJYSs8lx8UDV37GfK5kllK5SFwuXFhtG8KVDtVdEZOfjFdojTAhjw
PVXWxogMRNteqYpcoU/2VN7QVmP34aZ1y2218OwJU0Iq6b5E6O4/U/xiATrzwBhc
ojMgC2Ne/zHokALnS5YPshxtrthHzKBnKJDVWO0oGKM0JT7GepuNesP/tdV7AroM
TyN38drZ4hJ9n7oRez0f72XmfOmYOIdZDgl0nXs9b6K5dC8YBtIaDywt2g3imAzJ
14qFHJfbjDfZWUVFz+BgiL/HxNaUieLoWcp8lmP/KMnGOqMwHnunJ0jd/YVWrJMU
bSpNqAxf4BUTwn2WLa9oCnBSEXRysjKzc3yxBzRsvdATLHkNHq+FL4Pb4MY8jBaG
pjbyTgX9c72uNZfwA1E0WeqK3lUAbAS2eyo7t5ZAEFkbEuzqfqBw+gubZPMDDuQQ
/OCNDr8Kz2cTt68k4eMbiSTfmPNPVFl/y08n+0UGiicu6pXqGZRzdSLnE90OVRYF
z38NywNgkVSWV4FO4Tf9GJQM7+kqzg2HeErXAkqUz/pEdNfnzPPiJpiT3UrQy3ls
0Kgs4RBl52u01G0lT5ieJvw8vZfyLKGbPNLPVAM31JKOlNPlHAfDG6c+F/GZMflU
rQmBcA0K+FxaUByD1VhLiedRzVpmPVk7wEho197sq0Q6rf8bBhuQGrYwwAm2Llgq
GSgj88KM8Mho0RNVNU+TccgaIAs+aw+l6fB0SRxdnGt6eXZxCTF5azNXhUJ0z8Wc
AgAars5cINpEqzX3L+2TLXXVx3UZfM/A1vuarH1gpIy9inZ59U7tThiugWyZlZSA
JKN/26nsglF/WaHR+8eUTyPntWPzfMSjBXrCZ6/8vdYuV7VNIRc1sexfP8Bnk53E
8uN6kDNczgeTcFMYS5bHoZDm6uwjW1dRFvRWFT+zHhMIyhjsmC8NF7QDmRTwKfLB
eA7O18rCNPS1MKP7Z1YDq6RqUYXKJygoBp/31yEdqqUg1Vkkl/gDCMuuYfwkZYtz
bkstV/CJzrsNMGQ7a1jRJUC+SPUfSSgu/GckldlE2s5e+lwIRpqeRrkxqnuwlHNc
LCxGZcUGY3Xhnn7Wh5sbgs1vcFyv5Kit/tBUwVuPdNjpm/aFUohoQnJRd9+xxdoj
yggJcYbwtUvH51x/BtgiY4MrbZzUWHdDc0FJCwu3AvTW+RFUbi/gC3VvqIU6QJFx
eDg7xNoCFV+TfYUCVib1WA4scbUK0jkjRiizBN3S92iQfD0MXCMXNsSOVBmv0zO9
aPixlBibndHqb1Px6QIcVEWmcEaHwENXYtcRARVVTuZJb8qfGAcepc4auiUUmELS
bDX3qyXFv/8lYDOJFslxKPPnKH87jqT/PWHpJVo/CH3nC3brR4lTrdK4W6TyfJtQ
KqQd0JE85kRnmRqUmCvldI5EFHLuppWC4KhAiL/nVtfT0SPKBwycaSBxynuPrFPf
iwQPN/IYhASMfOOe9X6WTV29Fc2WDUud77uEqe8BLg7XGtwEa782Jj1v1yOvY/GU
yDBKP9lOMnsANFIKH9TymEcB7E8OIn+TcPG48ljY69L8lEmoggWXP8i5wy5EBPBp
Y8nqMe0GuAt0AOIpeARQJ5KZPD/XD5huUfyspe3WJB5obBKSknUH6eixNm0mv2sb
7eD4ASwwhhA3/vrinkr0LH04J7x2ec0ezgPYDGhId3DseUozPfEFDQ6nAaap9jwM
yrdAMeNlL++cRdySwPte2V8FlyP3y+rwludAzqTh0KJvzSM5nOgR78SwCS2SUUQZ
THahFA6GynI/WHwlGHCEbS1M+VHWqLCZH3ARh4GorQ6vN9RCb1CdU78Xus8nYOJ4
CuTMnQ0UgTSbMFW400Zl4Z02RK2ncvBw1ErmvAA6QzIFWKl9w/UsswvStKrBq67u
pu5ze1L3Cwoc8Pik520cHdcw9M36wd4/VYAjCuVlZH5Zf0n6fjc8NMrkn4CgIcH9
IH/gM5O7gGapEzG5fpGDQwiBjJfR0iBs8x0Ib4kB1lYkuT4A/AYRDMbXH5MrJCBB
1VTmzGGje1+kXs8spZK+Rp5FSqE/t+YF1tjO+AylGo0F/rJ2SJNanDrAQX1fnTAh
83t+YakrIT1HZWJiAzUrye8vehpmoQK8o+Sd7zZzR+cRRu3GOSY9/eRNHsHWe9G9
5KWJsYZD8ed09BzmffoEOsay+3Jyo0N9DwffFx/pbRtTA6U2CkogTEOr6vfTKml1
/uA/WkuPUvFc5gF7UTbMYfRtIuGGNG3ZStVJtjo0fTP0KIGGtU7XidAOb7pLYbFJ
Jlrsz5IvuOzwtokwRfzx0wplrEqL7XWmS0wNX5/y1FLElDJOgKk9siDuDEdyk9/J
cgZrgaWHjjmOtWMkZrLyWufez+NJ+AqxzfvoCPcj2QImKZ74fWnycLEEsQhIGq9K
6CF0bXdFetYnrqEQcUhiwXhvDhZCY76lUuZ8mjaVaRZSzaGg58hP4rPr5r2hVhiG
MpAIDxD0f5GfEcOix8VWdFp0zaCHbcSFq4JzuZA1JeSdFftWHYjmYITxIZKloRpP
Y7yYRPsaAqJtqOj+UC+gcoFlA4LmoInl28MZ7mhgGBL+T1EwWZpKpWzRUPyoPQp2
kW4lnckVWo0lZqkriqvyx9oZGX8SOAiEDScFOUM4nIA=
`protect END_PROTECTED
