`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5DUXI/4UQxiIo/JDOi6qtRooDpWpWrdzVGlvMOZSF2UB87O8W2/sx0wD0EsEFlv2
cR0TJcZig2Folk/8cSd3HLLhMdfXxO43jP4WIlaMBZvkH0wV8Ef+ANpy/58p2WuL
dx0XzGalmFJlVwrNjySrbAghPOq7DXpopTug7iz+2NO90FSvksIO4Na8oP5hP4kk
m1ESfuoe6M9QEbcSlgli1J71kJ6ev4nFHBfXCWfNmV9p1LxhcQ2UtYQlytHzN72B
GPlA7mTkytvFaz2YxTOMkBnlE55CGIYER/U03EynPrn3j6KkQ/UtSDBEfCip+QtU
u5b6Ersp15p+xSljrtRKaFvZfkip5OLCWtMXvbAzvfdk+Dr8pXkMyDInDoJER7qK
P0DtslWKCgjOKYLu23dtHCind137gQwFYZsTHHmlF0lOl9tz9fTz88VXTK2tkeu7
99HgcYTtyTSLYsaX70irtMftdeYJKzEhp1eqm+bcb+D8KEviOLN+S0dB1ciWAUex
Pyh5nCrG0AJIxlPM7uJZUkaEMAeAXuWJZ+I5ymvaWasBjuu1ydnu2y9GZ6Zp49tP
8pR+NrrvG3BS50nrPETBmzpwvWzqH9ceiwx08QvejhXqJQdrPnsZZiLGqJMHUky0
tEr/WmY9UnJS0nCWtSDXx7e3fsYc20Oe6beVihr9J/TmyX7XzipjAo91qvrPBUyA
jpqbg/AZIop8InsIwzV60IPy36A3odwdR7GM9s2ftgJuCt7fkJhEPfP5RK8FyiJi
2kCsssN8NnFfMFutSF2EcXn5XyUK0zJ87hINRjXJs64Sc/7xyBaUQ2ZN/72ZQwAw
i6D4rU/FFzkx+fYFnNa4SKdLJOdyplCss3600ZEE5CDmFcGWBzixDcbUNp/60vWk
hkk4GjssMtvZ87p2UfAe460arrwEqEDkzWsRgUAezCZTkp2DMqxyINBCKhgIqMKh
cZgwxlJhWeZgXCMGuuJftkCBLLpiBpr7z/n+HCgEw565pURSkr915xubi8ySi9NY
+Ulw6ZF32e8gERZg4RHhVpi42C146yhKKUvuWzgt18xqOzmy/kPh2uBVfkGuFvwb
i6O6jqUQH+dgXUdZUS0JkRVOiegMUBf4LsWZDAcUHO0Goe1OVchDrRM4MRN4gCdv
6mL+6eNijrnhKkPsfOlUfWmHoY3rf30LdTEc0PnjxVSDbvi7ya6jgG898CielGMC
smqH8yyDKVltgSHiadjYIg==
`protect END_PROTECTED
