`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kIYNbHk9+2zNDmuoOPO9x+ET0rB9TD8crS85kRZb11dAt9uYB1EE0/JPO6Y0dJbI
Dj9YSKNSywb1ZN8pbiX546fBK6+yVIVnJxX1ppfrUle/Tc1uLUbi2pecsFK9KPX7
LRSwELJh3C3MdoDzkX65ozJZi0t3ybM17zN3XQAZjN9HXbwOF/Kr368nMscpnDay
g4IeFjmbBmLyzQYHUqLgY08jotfaudt4QRVVZafxtP8MT47EQfbOMNJ0LQvo/NOw
uKy1C41TlEF7jYv+15L+nV3xzQWI6MxT+YtaS4FO1t4nr/SyfTLZMrW0y65pyzcT
nVKMhblJ77opzx23pUK7bt/MjxIhTiD6moi96Bfaa49EGuCoa/vj8lR/l5Z+lnmX
1TWqVmf4aDkIS/zzzeMTcUdYpBHUC4AAnM2c/fJhtz+qS6H5XjPB/5EBqo/AsXNK
ArThQw3W85og6EOj9AORtclCUivg7owDOfxloBsOV+35nnt09gRzgY90+rU4aGQJ
00F3raSURg8z0mODzyOd4WXHhRZaKYUlyYRfR4jDyDDrgFLG6TkMBYHFqZf1Mf1Y
xNsCba6iLeG55aGUcJwUWvHekt+RfuO5yWYo3b5zfKylQRNF67i7bPbsTAd+Qcir
vzfLXLvtmV9iYU2pQpxUU3Ny+CWSSFXyUQVZ3ilMq+FCE6fznQvWwfoipfEX8uxd
KXZ0eHCHFJ2WBFdb594DPcDmbKgBEzAscHlg/bde9wDxoOEt6y5Gl3Cmfbgj3n00
H7P+Yoejbvqjz4KequZk33jKWPGFh/HLiy+R+opwTKUjIHJpLTEEpH6harYtcVFD
GpGi2bMGwQsHMI1YC/EIUKUFHCZR2AWRBHh4GbGUOr9aqunbAxosViD32qm4iN2e
fBWntjppzyoNPA23aYp4cO0PlXLvDgPKdqrycUQ+xjQTypM5hMgR7YOVoF5bVZr3
VdI0tl22Xp/54owm46Bc5773D4334Wauuvn7IuhzKN81G/t+85pX5nj4LPl3K3Od
jP5vzHXeD2PaUc7n30P/eo/gmDP4Y0qCFlfdkzrDpYuk5CbTaLEuYsSe0hxJmp9V
ruAfKXtKADPTH6jyJqyh8r7IVd4jZPbT3REGjcw+XwI+5CxgqPCm8dt5wWRk5OUb
s7fLxzsV7k3Zq29mYsqcr/0MwbARgqoOE2ZJD/yzMZ/ODbCBzY5iunj29lu8Mq+C
KWcUjzS7wWr5ygusEuOCY/HL+emeiULz7jVsEz7zhC3eN40kTsIGHOp5WQ6eUIok
GbZlez+4TDIfmlDMfh3yrqHNfFP+eBLoxWOM8vH/NYjvVcbWYXhF2W5DlgSYxu56
dDOpbDs91yc38xAuabcTEJE3GiIxrXoZwh6PzmxLPoPIy0ArFSONsPLksrqOsfL2
aj4bwdoFs78i+XuLlpn5Vx8NGKvlekHycL6LklARdqk8W9/mlFXwr3hMPJOjylzZ
Vft41uaHxiy8sJhJfiTkmeTOn9zsTY+Qzj8o+deyhUyy8hQv7FJNGm0hzn/QSApw
Ws4SBJAvVLI8rvXLPGQwcMW4zFZYg9MLWsqoYVxcHcyppI0untl5PZElc3enhR/m
skvSd6ReEIiThH1bQtlaYyZEcZ6AVGV5ooYSPHWOInlEJLgIFkHSvLNi7inA41UA
XzFkffSHidsMurKGJDkHcLb8Uh/CuaodfYs7rx2BF7ato4Rm5U8uMLnYQ1QCFa1h
rv0ZcZfMG1J9I3/NWJIUyDIg1owcZk3xfc3508BuRNfVu5qQxPg64TwEM1r3au6L
ptynCPrBQ908RB8pjVstufZK/0hQNvTi/69H1HwkURJ3g/9mRMKF+oIHIfpdm3I3
4XE485xF09fbTPZvnxGYsa3Df4uciKWUCaDBGiBpx3quLW4I/hn0Mk2DQUvhdn/C
MBcK+nGYmzZ+YuIIDJetvw==
`protect END_PROTECTED
