`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o5ah09fnevosPXciDjcWcuEvDlz+frXVcEWu/ngabWhmA130nDF2Po6rmFjyUVyQ
f6Zv+bV5hUJvoG5A55xRqf+oSetB93XhriqaIIrnXfUsGUnKCEgt5Eze2dU0ddmQ
m6m1tOlaYoD7Ru3ktjR795Tou59BvKAxe6r/UkN758pq60jgiD4r6DXrmSub28AT
LA2iA5ietagRRSZ+b2Fq4/+XX8+a0n3YeM+1otPwJAaEyahhKb6f2I9E9xquJYq7
0pWH9AutG3xk6Gjzabow02Y+eL8T9c6DXsd3DRLz8/e8PcMHRZKeDF7eSLjsoN7/
NBb3KkdVuBgu9/wfMG32wPu5gsrHC8JHv5x9o96GErfaa8wHalbT6bYIJ40dNZ7E
N2uupYNLk9YZyRNrZwcJbjDO6HVCfeFdX2ndotGg3qGXP0B0/qS+7VOJGBiDx+kt
AVWs7oe/x7tGmXLD/KYRwvb4YOED3IrusIbUZiC0w1ERBNqugr4QcoZJzwVtvDBx
HNpr0RUWy/XAInfKgvc7WREuQaO1Fz3v+OMfNWktOxlGc5SCHQIpXowrAwjBkom/
yBYGnsztwYHob6A3My9GTAev0AHbmkvGCOlEQ/x7gVZdSlhDfFF4j5tXid7XuI4V
Uokays0m7eb3MXF2c1MoV74ovcW2TIpvf6D5+Cpx/Hoq2S/jfU8+G7KJ0FyUNJMt
x1EXXbzvbEOk89zvhJYTOgwvjnpMk9tJxBx7vVBT8NV3dMseK34NbTVRNsKfb7az
PFeUoAQkcPgXobZYmOM2nd/m3IsWZJDO8dFZMEMiFO4Of/T6YxvtjvpqYD3dtoYs
`protect END_PROTECTED
