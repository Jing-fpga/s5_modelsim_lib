`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cGlaNG2eDR5pmJ1Jp/kXXLwY+l/TZ2Vd2IiYWyQTjjxPAyb9XK3WF5PVXG8RV6Kg
PszcvCEOiKUrSCb8x8rjrUnvy4X7BON1CJ/+8hyZc7G2JkkwQzQe7Y4p8JKH3Iyi
zZm69DM5iTo3oNV8YDfHccqcZu9P97cM+diM0Fqd7gzfhI1Oc11CLiWaL/PSkLMO
7GmKwLaqOO6CiEDFWr8CReJ4i4O9/6Ree+wZvcKSWmjXGoIyv5PAS6yo7QIDOPN8
fnRsdMro6YMA4qojmu0+gfmkwVYZNyYtO7YFaa6REMif/0i1H6yW7uu2HiDsXM8H
9FecN8jnweQvXFQxvrJALrum1xLH+FlIfqJp1wRWzZBAja1fMXaOLjp+i/m0A0Jy
tAinnfq73qM2um3FKgc7OQRb6aUWUHdMEsXGgvAcsoorYeikb4pXknALjRIZugDg
7ObXUPgtky8MxUJQLdbIOLeZAMYH/y0RMAICUuz/QwXjJ2HTxNC2BXqXK1snqSVi
h0kRsEhoDlrkU2RLV2/wVERefWMxrXXBANs5j/bnxlIbgvPidD1zbYTiZkQeTqVR
2TzBp/qsjo/CzzpyZyMziidp9w8idkUH7KZkbZ3Dg5o1O5r3urgCpJwRHipU5UPb
0LrhaFD26P+DYxmfvrixcJYk+BM/HBbethMsEDAa3vtuevFVfjwKwty2VMN/4mD0
M33cbF1PiqccbJU4h0nTvmgENpIn+57Oe25YA5KiPa3XM5LD3oLbCFFImzhelzg4
dIrzU7mQL2XJ73/fWCwWjAZDk8Jaszd18NNn0QfE2cMjkV+FKVc0xhCRmE/kZmLa
xa/+mCH1nKOOxiLdhYuxiqQj9q5KzrJ0x5fhIaYh53VRUvf3qFxviLojjOKll+0a
lLaCiFdRF9XoyDaCcfbE8/fqZVKCrSpUKn/JhqoXVuYfwVaJDsL6Jq3G3wrU0sDy
G1vwRyZ9noOdsoqwvad2hrTH6DD5DtsEQBgLuAHA77FgiN/HBl6UA0n7M7ACDXXQ
+wxp8Z5KifpvQEFCPjT8Arn0UikRv03It9F07tF85mnnh9ZVvta4+8JRsQbrcjYt
Cb6kXbdh73L4vCz691V6QmCoGfr3QOMv6kSYmFQOoAAtW88lchaxqVw46GcnHaiW
Gfr+Z9JIbUeYKT0wvWtye0k2HAJu9CVUX93gWgSsr7UHCj1P5CqPWB1t95WrMGpP
r83WMLxiTTYSAgffKabWcUDbB6xvEBZ5ZQ/JNq/EY9E7LlJGvTUhbQi3AKvnG44T
1X9FajePd9RHubtP2xJUW9aIZVD+nxGP1MD+dKLTczDoSfQr6JFDDra8l89f2ZjW
jV2RJVdP0LClIEv5WY5Rov2Y6B1y93yLJMxRdMcNkxMhNxrI3tLxfA8172UvejwP
Ard0slc4kahEY/80yo+shkGmMrg26ehlm8tcxpQbtZlCG5J1Xme6AJ/O9IV9AhGr
GXm/6XuBf0/gh7U4ypzFGwqmHSJH+WVPVTTAkd17YylTeNAMkohVd4+msTrgUOL8
Sh4wmuHFAKqhA4IiBB8WYoyRhcdZYLwxJITbrLX58CynSZWTP2gW5WlieExFgzha
3P5JqabTOU+pffPT8ChD68hXPAwqvG9f65e6MhbFUeDltoockeZegM02KLOLEbvL
awGmriuHnQWvLDhtUYvU4HSNyRsiqAZjB3MyHiBw4O21cWStbMgLUhUqKN3dGirO
wgmbiTLQunmbyKpVooMrw7iqM2gnp3+kaswRV+HQpB3ZO4R1BLuw5gX/6/UU6QEI
CTFKE7XXQiC04Q5dCJDmBOe3Bn3k8uSZeyLJtyeuc3GMBaTeTgbyLSYd0tjbfn1s
SbxEX1e5BROVQxLfAtJIR1FqNEkgW4Y0WfE+NV0zzNGEMDUwSyyWHFIQmy86QW0Y
XNAAqrggcL0w3iMDNIvv5qPQ3NEOociv7ABBZ/OVoDhjps4Eddxb2yk4tvFIdRGR
j5ygZRotojJXN161gyU0a3MKtZ2asUOt3Ctub6fyWDv9qiaIoknER4nSXawAeW1k
ZAASxFdemsXafx63X3yHQSZkr7e4jbJ9rbGMpSrhRYjg5qzXiOxMbsS38bK5spYe
PtyoOwdqxkYDRgt0r6hfg/1Cw7lSOBW2us7GS49O1K5yAQ5ojivjhlpLABx54erd
3DhZ7CMwzaQbHHJ6MAayvKHAE8Xi/V//e68Wwyi91GpH6pS5xtPgew2xZbSFWIfD
JyN7SxSuAhWHz7OGqvRYp15HrG1lqbcVr2GVKU1UaFca3CrUbzWr/9cISJYtsctj
My4XTqhRkBCESVEb0JuiXKpi4nOny3NrrwpMNq9rrap+pdNnW5tIVUkz/m6tD+oq
RfO3csxGo5560GCsBZCmsa5RPwXiyBhj9MMsXb5rkteg87pmS7xluAeBICKXz1cR
cGYApF/6QFvNYqHO8+gMnMQXyeqdDx2XbJMSVfAnhXhtDoJZJcX0trMl1MeiyCqu
AHL0uMcOgYLoXYxaTN4/YkJzsHCS3PsbLSKOMh3Jove+X1HxE6AexTkG0gSv0U3P
d2cQJdXf0oAygFOXKdZhe4L42pz0IIawWcjNmMQ6XsFthh2HYZLzsXBxLoT3FiOR
4mZrMoprzaqEXxZgGhN0AzgqFpEC7LM4yV4Vjz78nRg7hyFPTdWgemqex8xfsiO2
Di9lG8b1Ya3uH0RILQBInL1d2nF0UlhNfi8QVzBUAFYVUSFmA3rt8944FuFAUkOr
Pl6pHBAAbKPVaW1tHmeuAaDNY+XiJmkNvf76Ipdhu5osF/EJIUkYYeQYq12kE+Tl
9RFdRo6cU2pQflys4VKZqkII8vynH3ez+7DhlcQ+Cn5+iv3ASxeVYJRAj5FI2MgL
RXNs6jzSOTZ6gwzX5+ttmHrBdt4T5l0M+rWz+MwCjcWphl6rTO5g1rvmRX2LLbZq
zJiHTvj+MjWwqlQ1o5j8xTjHnTba2OQdhSyEv1MmlsCe8pHHaQZuQajqrs6D4mpe
5hc2i0oTCX1Q6OskbadZqXD6/qwf4sB4YRvhFwSgAJpfpmOAnulMj65c66MnNKiZ
P+Pu6FUv/kNGkVwnbeRvhNcGek/BVyMPG87rrK4gia3W70HwbDEr93KEwDLySR3x
+NAMvR9mQnPYWoywmA2AMLGBG0ZiM9kEy9Sfg9qyvGdrX4dd0B9AUrJSfnmzdPQF
heaI9U00EKvLKgZV1PsvVescQe+pI9AQ6Tdr9SWZJiMu6PQPC9nKSqGJUcjXMsbR
xsO2RzYOALgGmZliQiRgurYi8Xqp3XxzFPPB1gAUykAIMPXkjmxYsbqG784vkTom
bJnkP7QOLc8iMXJ1690elN6YHg7Zdk+L0cfH46/bydPnNaf3qWAsTfJqsTsg9slJ
X1rvM1PRfpx2t2CSTa0hQG9AC4y94YW0RDBHSd82GbjwQ3Pjy6iDZzSzTSaWP/dy
gCEBAlMlU4JluT7bNY+Hd2rAV0GkzrZK9qpC2gkI0E7LEbSPsG5HGuclvVXGMnv0
/f3zCs+dq4pS1xw/9huMobPgx6cqAZFmQil60HkQhmT411aoBMSvkBUEqC5WcqYx
XofVRR669+v14EOGDmgRKVgGRGnH+Nfj/h14tVdBq3w7UtV0kewXfnPeQhE1+gDJ
99Rua9wTzkGV0oS/ZKS8v130KPiW8sLqPwrJptO/29p3a5jRQzKm2SlsUx+aiBLO
P+edttxsCKZP+R8xZEGn2l19cLThNyxKrzooDfXIo99F0QsnXIOUl7z4aFz/u+Tt
ZIgUP3C186gr5UdQNdXv4+ZkqNKi7M+TMP7xjdxSTufeMmh0ZWoVGfEN/X3UOYKW
WWZKh3gK0zDocuYfa+SHe8gPmeBdkYpHW5soQ0g9wjmfCnVCMh3vhGnkqMLY0ubT
hN6rrZOIC1T7VF+1Z2Zl08yZZfCbg3AjeTqKi5t7+tZbLxbUxdG6xs7PHgWQnEHw
d5GIaRy1bA8fDmizwZLRMHVAGxC8x4btb9ioRnxve9lH5Jtx+mhR/9PDWhnGbr4+
LzWWFf9wu4UAnfLL6vcQcbZeATV1U1GDx5VNoEBPPfKbPpwJtyGXKOoHjN5mLjrP
CFmR1S3NYyRTT+UVibDNT/+cnnq3MvR/RlEw2aBafcc4JaMHGl8rWYTC3REtwdNq
yhRxY7d/LStJo1cZClhfZyn6vfP+s8/u9GPhhI+f+lLXzRSgcFT0A9L3rUTI0hcX
ZtnvFI7bu8AapGafzJonT+IPbGL307RfMdmKacFFJOn+f8Xp120kYCSV/foRQuDS
LA3OIvH9MQsD0gMM1Gea9rypddHJObvr9TjlSt7y+/dZuZG+OnOg2UELhHYpjNc3
wiMRsRF8zl4bOHxyyWE9+i4O/Ttje8ujGrJLp8WW0TdpOG04vqtkhiWUQZ8peEbD
pw/RWsRwglgVbBwJ9247mA5mDLvSWG6gKxUnci4LM++YP3C3jKTUeLb0N+zhK+lR
BjJ3Y6Rr2RKLYXkk7CJpc97RWTAIEv5LyTXiGZ64Ll/+ZJd31qH2r7RCW7hIKboL
IQzsSpfJ/pT2yuld9M9KH798u+HmelCWI9UNEpk4sr/rYfZMr11pTeFD5t0vwYQH
ShpIXCNKSg3n5aoMhPncgA8RnKv3v1eVsnC44oiJUxU6Cpjl9M2skl6iLeFmCGuT
CcGnkPHuHy51VBqiCKhTVn1TOdf5DVxJsP5tgwQnWzUJqKXXMKiPpktq7Nna6CFR
5WrsYzntVTqr0S/pzOFJJytBgDIl5yOVJU/9BWspAOGfVcVBtDjYj65/clW8sT6p
vVlFiMuMpdOklUQ8lZ6zLnjRLPtoARk9rBtqXOZCaQCmyIhQckbwcOUvunLgpKDD
Aw/qNltUqLxs9IFb5AQbtCTHqfPWwl3PBxHEfS4LNCLjVKZpp54FACISyiOXRBdE
lvSP898aFxAbkgA6djpVPrO080+bdD+wL6EbUHUWM/V+2B0hVExKapMjI6kxzQdq
EeoHKWkz3fks+9Q67RMJ67nLnbmWj5OSDlvK5+otTzBwg7hh8vGuRI70/A91UzAd
tSg2mIn5NyisOPsdGSFtUVK2QgeV5uRzr4wXk5uOR7B7P8qmpm+YfAvR2OxjFhrb
xuzwjoXpvS6TZrBpwjtfH0XT4lC3xXO9rZXtyRYU6/wmPyrJgYxIanCpP41KtrGX
AEhbARPszPMNq9yplLsZovS3gLQgBM5D1/EgkLgkIfhs1mA4WM0TvG7+Ly6I+SQb
jnySnsk6w3Eybj38+U5ukt9JayH4pKOzK/RBA8ETojyMGDl6a0cd8m2WNvLGunsy
0vvyVdcYspjEUi6/VE4Vvc9NOEcgrdo3CZHBtRmptA8wldxQv3nMD1kuo9TYTIMt
83LYE3JYVYC0kHBpjRR4ZerXoq5aUfflkIpnLHAiTZhSClE2aAjTKyNzZtYKQH2s
l4PTGrYq0aWD5OV1XufTovxoz1kshbknGee8/dRG0i8Y3B2ZNn//RG7T1R9Rs2IB
Qu2sRn9sCHVuIjS4J0ibCJjnuKPukvD7AhjBECy9TwPaE5NxwS8tLPIi4jEic2c1
uDVScdzSPFLvfGIbZ+xsIMFOQEyOR86cZR9eNcXlFsSpV6ne8+0AkiieF75r6YWS
zInjbYGMw/jHrkydiB3vYnXLpeN07chkJ7/27FnTaJQ3TXMfRdYwqUfw9DV4nKLl
doJq2JljY+xfRky0iNBhXYcngRhr8avgF1AAiAQ1kgXUpsdYDmbZbO36VunFx8sh
LUIdLgO+f9Ub4k7it1vrxvAB2fEulq6T8OjFu5H9fTJ6YPf+l+4V8TAp6YwirNvU
FNrSio78iq7TJua1DYm2OJjDyEdnOd7zWUL5WSNehwKPGCsMzyaOS1Eeq0NDb5ls
YAi8UyVX9b0LoXnkGBPXAvjhvAQnOSkupbxEIzI+QhdP3tyH8qfz5tL+sFz7jp18
+GxJv3byn1yihMcEIxoGtGOzICeeOl+WiN4Q6iBgG7ljlRIaoPIF3QYhqOL6msf7
ih5Q9c2hviHsKXtRIW1bXtgy8ik9LL5ghQjlDBlZ3BCChavtC4nwm1VyGRmUaGI7
teygyCq8K8FEyAMJVtKyTeggPp/DlhuRA55OqIk2fo+la6QaNU0sjEhFx4lxvhbY
+T520ZzlTUDtz2r6Ti+aikHKflyZQd9VaD83lOoHs2y2krk0Is5T3An1BMDds/IM
WguSMXxjX5IEianXketzDpB2LTuBzkr6mZp1Pr9uvtSpy62/ULNvOcuOAi74JIIf
VEu2rNEWpnDmpnjiFXHx+vmdTtDIMdibjMs6KNkkHULwEWi54F1FUYvnXjIcHK9w
0kFcGX0xytAoY1EgiwaiBxrsy6yFfbT80U/p82xH3KMdzzweESom1j6aK085MCRa
IszPjaKsUqo4BURYUuOK7Y2zdHo2f1s8UNwTMt29yKTggmyz65/lnvpZpjxk7tA4
xyMSuwaQm+/rHnRLYkKTjk+p5XAk5rxfW4+HYJZnA1cep2LDmPXWUQMDWthbYkoK
i/uKkYUO/cqpJgmNErEkr6Wq111aNPxQ0V2Yyc9JM/c4opPkNvdn2+cIDI6DwHy0
sI20fWEPHUSWglhr7r+9fS+2GEk3DuLy/WFeJvkivlUyBumvOUA5zbYb2x2h2HNF
hE7lM0d1JK/kbK8jtEsiVNQQaaSaSjmsJMBlJCm0/6zyTP3WDdyO5iWCu1DIYcW2
6KaxzmGGydL+7a7R7NmvqLWAG8vk01Qvp/z+JYv3Kfp/8ucx9KWp0uuw8B9EJrwc
LmzD60/ZQjM0Wr9yepkrVJ40A48vCBCn+z954BdEBE525kjdRen+F7Bc8o3pBG4Y
k/bB/W9lZSrmfAneTFpJEAbZKUzJ5GpJNVy1ikgMpbb/fyLb/WCMjvM5JwrG4HB8
mnVbSuPhgeSgOSWOo3zaioLqrcixtBM3tIYQISxUE/98ti1Tp2E+/VfuukVgoDAw
0RaOLdYbNqma8syDH0UdEdJ+iHBhmOdikyEHsXW9eEOl/jkjHkLMqagrFeIuOT2e
u8meeQZcz+KYUPe2uTbFwPkP7dKrFKPY9Gi7A6qbE9JRmJJKXCDtgzA3hOJU/79f
x9GY0siNKg8uYAwDoJOamlu6Jr32p5HYpAin7BM4UQ0bLrbnvgcgKFdhzTpV4vzT
8Vo95c0xC35I95NUSvBzH5tTzejC2C4ljkQt5s3CPf/5/55eACQa34JUjGcsJO6G
iC8kl0WtXyy96vF3xLNZOaOvSx8XVkA3RmYVAXVG+P79WmUNB0aCaFCKLeWXWpF+
mjJrtlpkCG6JLcJTl6zeFjNaDqzTBjZvijXYCfxIfH3/vll3jiNh08G55oqiMdtf
63Y50h2ynnXahVfKq/NfLt78GxIDfRcZJ3IfagY+4hMxb3wjXcmHzBPYCjA96Day
84d4BtRJ2hgScnNKPFNV3Krnd7S+n0pq1DFsG/ntTKucGkhtc5RiTaErtDdxhjpw
y1CZIB4pkyB5k46hlvllsF9F/NGueIlZIMftEFgRxw33XYaqhCd6PQ3dv1oQcdIb
VP8XPE8fC/mL0YsX8B5cixd4qYEVTRRDD8C3+asiD0iARhaH49PyZbe4OhYhskA4
NKZF/p1E+x/xagpciv/hKnnn2GFBQpkmwtcNe14Jrnl+A1jngu+isOZWiHzcNddS
p3FjgQKwpjvXo1Bp7+ao0V0NOdX7UVlq9ElQFmRVG3T7/ZRlj5lTRujd9ltshef/
BbTteCBUIEFtkNLx44ACBSWHHtCyUprOUHHScOb2bng7cGPRg52AURQdQKiJNyMe
+ov2Hz2lfLUyuBPZZv9ewYie8x0k8NclwO/yVP8Bmsx41bG4N9nzQ5nvIeIalXu+
gsCLaeSgGSJYv7bZR0h2Vbtk9AGm6jGcoQRt29uJoI+zHQBLbnqMTV96J/A7hz7N
THTC/gTOJD4lMJq6qLuM2SlzShcSqGBlzXqYcDS0W9IVLRii54kJGyLUGA/X55Yn
NIkNPzxaL2oliStP8GOWxujplBTn6Jd8agWm4o64ABNQT0TEeds2tkQDJcE87DEc
Hv2ucJfBhzokgXSBq/4MaRjjjq9EPgxfvFeFwpSRnei/NbniVS1kb8pme7XqC2zZ
FtATmAEmY+yaLkdktLy0pW1TWk1KVzaoY12YCMZkuQ7xuCab8XGWYvrYdQAbdVt0
AuyJ8XMbzIn1xskJUjhFAHJLZbe9F2wWDJChFhrSFat2u5lIC0os9MU0BTPemimx
2+67Fl/rfZpHeA10miTUJDO+MMDBQ1IwgTKaZIJsZ5l036HgFhOyJHrqXsS+ZO/7
+eQRx/S3weXFYtCR5kgZz/9oDAGRdpopcSvWdaNC/Abh0kvk8mefunAVB1FGgsxC
V0ZchsOJTH8ktYMgKr3/a4EzvVVU1I2emmWatv8VXQ+yJk8or60ErGD1uBUhYLMN
zvGmYWsQmDNRQbHoXoGdt7vAn/vArKPGT6SteQT/0i9QiM+pEFI7KCheVS20MIbA
rEgv1Mh0K3yzYacy0mbPpW7th2/hhZfdlX8oFqkjCHEx48UwEkesYijcN3OAvqYn
RSLYPCuT8IgqCLhmi2kiF0/9kHsWyO0jZAfHTA75lgWxW/AUdNL0gZhT2gX54Kre
i4LILSUPwpexa9yQdIX1SJWbhl+4YiYxSakt/9rGniC7mB/D2nV/xp0ay44/u6Cz
27lTl+IlGvxe4F6wSbCOyCoDJqRKowIS0/a8ExXSF6uebQ1uT9iVKcOpKY9lKX1O
trnodGW7CK7XlzgTVxQDhq9wm7/5iFHAfV6mqmADSZ7KzmXXiLOrTenk2mqOtLhd
m64g5m/0MzMp19Fs+db84Hui39gDEbDDPK/iolggP+YNfhCHend89IvV5CQ4TLQn
+9A596sMicJwmvvrmHx3BnAi5dzebNzRHKe2JDyClj7FBlBWQfoea+3mbsYvhSHn
BlCtNQi2Hq5ZdYyjUcU6YPE2T49d6uX6HD9kVHQuBf2+1U3+IbUv1ioVJrYZ0w6f
DW5MLrlHiiGm9KtvDdtkFP49+d/1PuGZb05/I6e9zpvtpBpQhGluvrS9M3uAko4B
9TZP6nrRZcDL3j1WO0j1GkjQVfSeT+pjcdaHoyJcho2SLeMsKuPx9Plj/YieCoU+
zjDoOt9sojwioVPuM1/yToQu9gBzGzwBSsNQasLC0CQc+BTnNA4OjIVybSEI1/Wb
Bh4d5RGny1N8fOUIItpuMGHT6168hnZi5NwzfijjEfGujotw1UKA8WbxTX/Rqhdg
Qd+VKNe0UmUXvNMSZghtEv4/4ngHJlBXU5TZ/FWBRbpcUeoVnYNC4Ut4kgyIucWj
YQ8mdG9ktyNj1BZRaSrL4rm7Yda3ZJQFlUQWY/AFycj64I8ubal9DWiks5xHkPSQ
9K+3qnsP9xKSyvv/RrPOuoqS45J8uMLBlEphelHO9p1AcrKwZthnza1+ECzXORKZ
eACMu9BSe3YL/CR/XXDurZBro+Etmh7Mr4hcZIrsHQHzLx59a82Gr22ABy4TBSnd
aP80D92Px3kF1HtGT6iJN9MxZnh3i82UW2/STU5Ad8RDHwgsSe3UvpJMg3enNZ0o
usydJltOy6MU3G7XA7Lpg+J32GYZn/hBvwiBvwZigkzLYMKhS9r87UJfeWo2XxIQ
Qpqf8IxirZIC+bL65OUZsMuaUfhMvcofPc4fPzos9hzp49yUvCiwGUjUGpjY5aO8
kSSH2oMWGlrsDFtZqqswkw==
`protect END_PROTECTED
