`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EHXg6zLwDEEb6AADtGPux83KSZ7f1ywc6b32e6B0THy38e4YL02ZFgKRrdtbmGuh
O9KQE/MiGIfERstU0a1iu3WjG0BOtEUpzEJ322wOlczOxCB1xeSXvAku+SHHXMvM
hNje7K/B3NSWK+23KcE9bmaJFZ888tKsuvIIpF4dLDfQVoeFOplTcgGtPMp2BsHR
efqevmy5d4FVT2jJOxUhmUodpuM4Lvas5CTjrpRHdozWDc3l63odXyzQm17TT9Ao
IBKREY6vzuu63IgxEzAKdd+KOA8MescYNza1EahZ3zJDFJnFtbgZpqlEUa4pnDsr
Ce9NYJwr0kPg3FGUD3W0njddfg9wYn5YyOxbJXWe7pwKxNy5ojAoWoi37WVjTNyv
inVFR1+4wzq6fpCAHqa01oF3Qbfx3QtJ4EECMymdP9VADMmbGoT20C4wYFhBfqt3
otB4+4WOUYJUll/op5UO6USB5krMvAbmBTQPBBEgPVRh86xTqoRN+2oSSqnKxCeJ
Np0qWqa7wvuz4mF1ZLh06Luk0w/k3Ufmnbu8zFJ84NyxxwsjAlCFBheavn10WGHz
QP+aB4u6dmMkGlY96LI29GKTc/E+q52EAnPekbFGEXR/s5nh8fV8U/B3uJKzqE0+
ORIrbS7btJXtjlrD6WOCuVB4ccQ5ez45t0oU5j4HLeJV7I5GQaFwJR+HOJ4/kkee
2bktQWB8Y9+Z6iFs+LO5u3362NlgurknUS3PcgakKvugHykYFWuKemofCXnm3NIV
7QRU7K16ojApmnKA+3lQjIKSyE41nYuRltkOf6DV38xEpQiTcLA2O8aaPFeNnCvN
lOJ74SChBws2FEbmmu1Mp8VkOZgOsIR7HvLpdDW1oOaQsFsrnRlaawFJSHJvnigR
99o6XYxfSvvyJe4a1Fox2yWZ3khMgZgWdsJxSocWOXH24JHSI4Ry65Tb38hwSrMy
ZykIMATQNfIn4b7paktquMnBQoxoMjzbCQa+hB3NSlvBEXP8n15X7I8U3Z/DAZPd
SK8aHnRksnphz8n+RmKi8KoggEVueuo3cjDI5PVOLjJnhaaGAGxdyB8v59I18zZ4
xP8GJIVBDLyrpet9PyirRsl36UqC5VZ3/K3WkGwbJj0J2qSXMFeQHbBAJhDmXFz/
7a7zQLyF+Ivp4TUWantW7dU+Ncvf7wG4rEP2vTNufQvLoKzy+BrMX7PKhD7+4kei
21dx9/5iVGV3SWh2ECLMX1R38oejcGCuQp21WWhVQFMLQif1WZKevPg4JxgVfgQj
1UTRMjkJAgrssQecbKjtdzUawDb3vp+nUASH39dtx24ldVLEZJ6z6ZDVj2fIjS5K
srZBQMJNI5uyemvH1fxF4XfA3oYSVP2JyOvCu9gZ5HnHzlq1edVfuNQNFQhLMxsO
15sjTeEoNYtF9biY2FGfqWbwxlZAKGDCs6L9oW7m2O5IXo1zqU2LkWlEFwarTn7o
1kXP6TBzypN15URopfZNmmokvd6rpHFIPen+oNK7b3bj5rqvcTrQTnL4pd9lT450
4b5ncIReFwxdvNR8lFsOrSzpUhEGP83U4z3LNE5WETckh1VhrsUoo4MlvNsbIE6l
8hmoCwMIHfwwIWc7hTIppJvekN3aJML3LAvhABvbSQ1r6sRU4CDbWXG6Qoto8zmB
R+SUGb47+P4cPXJHe8fTKMBb1aVvfANXbolGvAAuNsCqtNsDImSqcLNSHD7TJHfB
kzHJjRhDEIl0H/mGiCibelOvQ4QzJocwmoE3ODGq8F1RVpuJG+skwHbhksQTtv6b
K+oSIBGKHzS41wdN1+D4nS+OcEpDU73WLdCDTDDHlu6HY4qDxcUtGROIioNH2kv+
JY8LoOSQ3AZVs+1AXg2LDIppgQE0wF11UGOyGlpe5M1GjQZG6zBvXc5ovf+W6PJQ
6EB8y0LAwnAKneyaiIQkfhcQ6HkAMbgejmWFRMN8zJp+pkZ/FFJQE365P2iu0oDT
wLDoRU85f0P8apzQouLaaSVhIWoY8XMrUSTH+cV1LnBFwOF4vFxyPHxg5iFFTI/h
jkKZp+LlYSibWSmByalUF7oFf5Zul8iYsBG10Cncc6J7w+hUhL8nwrJ5wMSjFV+e
KMJ3hxBcuZmJTmPQ3VO7Gw9hu6ulyax/q9H25Al+FlHLv9PYjQ3P40V2bPIdglrF
HrlO5fY2B4+nGEr4Cw/XwreUEfHpE8JqrCw6ssCmkgh7VjamvbKhiYV+6PWo0142
vcYwTgtO9BdF+4FiaparuRx6zFftCfuBKbQWmjPuxPLA2iGYJhAHE5wXM27x5WK0
Mq2nUaxavZ5NABxmVwMpqnNpOwPWetz0CSa/7Ach9qCkp1J7T3s3jMsCMLCYyyWB
0kLI+Em6SrN/9mtVAaf+nudoLXcZtb0rb5KxbJqifj+aaP5hO1NcMmWWhoc4LmYS
YtnGMynwjsY0h77Vx2yzryU2IRAe8w4eg8DMr3+GchJzhzTUVgiTBvfSLjk1MEtz
57OiROAMV4GvNyXAfEB8Iqv6AkscSOS/MTxiGGlsln9zZTVnxwQr2eX6uUSB1jhB
GwiQQ/2ikO5wWFGpElCq3Wh+eri4XJeJ/KrUrKKNVsdtOFxwGhC2kpO/+/s2o52G
KqvVg1Or9r9Llo/d/tuOYl5MU3eSvN/3FfFFjuJse6+fou6rp1lZkQmL9syBsVZG
Vsw3ay5epMDm9YPRTD/vFcDK3/FcxolDLBHhDOf976StTaNytISY4nw4PIJrEx/G
MtEa0jVBLYfVW+qmhk70QhcC5jGh6oFPD/BJ8ryv2us0luAUl0axoYEQTd4A55hS
NCRepR9n3yCJFW+jYLVBySltbVWPbZQZ+g0pWDyNUkCdRBopCLYRzVFDls88g0Ix
z1VXPex6o5opsWgZCmmDUmVFtMj7EtqS/uiH5+D6/yCKdrDbZp2mn7/8u9q0O87E
/nB3Pm41DmHMfp3NfdOwf6Lb2tDArVCg2Kc9d9c0AxbHmPo8NyrN3SFTR5NMfJe3
NXBBmsSAnARBwbTvx1aplhKmYvt6bIzLs7+i6Z9PisED/bG2zofce0HwfeYTr987
Lf6zU0lmTEin79fnDI0/qMCPCdJ77hBC3KD7XiBRo5O6KqeSpFptbuts9cmKx6ec
Gv4DBB+RMcK5ct3OdLcuhrqT+AeF3q41oZv1qUOZ0vemrCy5J6pw+ayWa/uJQeXX
pQMbI8r6HHgLd3Yo8zdOjvkkCBaOhSu+Jphm6kf53DlKWwoAPjFJt0SMm8NTnL+Q
NMT3IMxLcXDmuJi0ZqnafQ==
`protect END_PROTECTED
