`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EN7a+EG87M1U7qLwaRLFkE5Jq3/SgwdabyrE8hOUqmGoxT6PkNso2EY3fR2CdYD9
EJcZwMJbeBk3CmfClJTUi2S1UU4IM82YoDpHya41oGqRpUAwgSyKRYyPQdbk46KT
2DP/UXWlfjuCaA8gOxxgFg/VJYMCX839AAURA+b2i29z+dK1zW3pDyKQ5ir+jfC9
IHQQor4WzYkdPMeIXryQo3r8IfOclYWaP2u4mMx5LRzzm5cFdFWz4C9DL60rdkA+
QxRK6H8xOKSBLafzBy6kGmw4CiIgrquoccvwiDDqMdRh23eI7Z5jErrpT4j7H+E+
hMykG5h/csmswaFh+Nlf4Qp6NSltLNN/JkTs2HfLweMc+WZyZOxLy+FMvJO2pFMZ
nJtF2BGNNlINztArTYyqahGLPZju7cgGAit74S4v9jNTdkVVcLLj0Ef/q0qjXn5t
JQldagUVdcTwEeML6tna82/ircF5gGJQ7sGPR9jH54E3QQGZEnzV6l69Wd2J+3Q9
tASzUH1CEMav6CDFW4bRizZv/yK5k+emgESpM+q5vIsznxYOVWIgtJt+SOLWHxJO
TsfLD7+7C4pYpBdj9ekDezA7lrAwj2IKjU2s+4Fhgj5PHsfBMW3NPuQkQKJ5PKlq
76/uAFQGdpHWNSUkzrQZXXNYiIi1h8XO0FY+j3ReQyoC455DL0/7apyZrXqAKGkH
bR1LkqRzLCNgdVMu24f4A5r8Xu8gdkBXr0ngQ49q9Bk=
`protect END_PROTECTED
