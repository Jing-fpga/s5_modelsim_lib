`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7JWMEwMkn9N4Fvei6uzIVT/AbJZD/zjZKTE7Ppq3WwS+K/EZ+h7g1LXRNK4s/k6J
rk6PfdHYTk9LH1AnMTqKgu9KNv9QV8FwcDGA2ukicrbl8FZ4Bix0FuG83f1iuS0b
IA6r44INxfzBV/Amk4pOYQitQAIrdonDhp36vSNmC3T4yI4T4oqZDw0bW1UAI9WC
zoyhSgk0z9zmXcnVYObOzPKEAF3hKePn0Olwpwm7KJIvqQ4opatMd8j6rIGNQ3qt
Bw20QRhnNnsNlabP8BozCJjvuYi0hlsXgTlS6+54UqqAZybXU+4FhHHOmNVRAM+K
TVql7Xu4lYFoqQKMr9HoPnAPK3an5IOXMoFEV47uMOM5/CgQ1tPC/ALqfJszCXkw
Fl/tbwO02WiRfEgilluCw29vrnC6hY8f36GyMtc30OobMIOuJrUHQa024wRhPMtn
sRTtrUaRHWBQjENhdIN/0H23OLpzJ4u63pwn3oH4S3I9JgpSqtX4NUlTVdbZsoGX
wUO8EBWok4raLJNGVdAS68mlw9ZcC4lbU3+ImSgBLpc2KFtZYT7G0yZCiVNRwiBp
VjC4fVtoffMe9II5sRzXth1vuIjRAXSEyb4cxVNytTqRH4RERaVfhUTqCkFG9+C2
n3ycV+zPzUR6PbdqkOyHqFajYu0wXp8hNWn6HgXSamNsq40LDufKnwvz1ieGD8ty
BgmxIgaJRKDIswisDLMZd3ScPocU5XWQ5jpfqMANxiyuMYpj5c5bcopSjCA75rVv
JP13zMIY9CGW1qTmx4kyGvc1il05qf4QjJLwd6Na2v8=
`protect END_PROTECTED
