`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
si2YVzOdbF/d3vRtwpTfjt9H1xE16aOlT4URLo1GXhedirR9b5IxbtssUIuTC+2d
py/nou5TZHlA7YdK55K2N18SOkoB3qbaxCOS6tf1C9i4wTHIGb8IuOg4+pZyLi53
qwaW6LX+wyukNxcgSfb/pyXBqmI+bS3PlyM4L9FmavHeHhjB+gD4ypdVjTtU9JU4
2piq8fmSwDuZMKsfnFN8op+7yp3lKBcypZ7Mm+AkahE9SjM6WTVkYVxrC7dR6mmz
pmWW8Aq4lKHIy0IF37J7Eqh83M69CmluO9A7WGIGy8f9D7kLGKZg1XrMo+Oquj86
mUKjMis1/m4ajHFpJRp+mqgZHuuBT/fEPSTk1pEgzLvWJG49y7wM/nntguw6LE8S
IEnXyydlwKcT4N86WT5AWUUqNdXD+g3oPw7ion7txCI3pvOoG6rEqf2ZzkOiu/9x
n/4aUs9Sy9hMYa4I9Lp+3gszkX8evpQ/sRy0rZyJlDWb7oWUzwisYk4DccDOPtoz
xA+OjEwrw3QhBYW62T/KGt556rp68EGsKJZVg3QOtQ+KRV2FEBZpxeCtxgAh/Vvc
EMoJh/AH8Sza+OZp6YkG4KtzaZw6RpXhPwcbEu4GVfOqYKYmCgT2GShFv4Lbxk7b
gX2cbmzxTw4GDCtIMKfz4kOM+PNvNpFiCke9ObLsNq5EnQavF2v49nJOa+7EEgIk
F9ejnYzQPmwNu3BKgKHVCIWJld02uKI+MSNOzqarW2uVajNFydKmdV0ysQF586Al
QMYXg65NEYztVsFxynyBLmw0xYKDA9EkKtSZniobp/tgpN3/1vdneo9lGOARbdp+
K9FRHOFD4rxYVijjlOTkDdZUuTucCwu1PXvCGqRxAnGlAMASl371wyt9RGR1BIpl
ZdkTHoN6vENa0L/UsNw2TydvNCe6aPdzfiXBDBOqjSy4gs5QM0WqKv8aDa7B46t8
P2a0L+rrQTczsCT6t0iE4wwB4Ohf9m2CbKfjD6HhWSir8HFZbpzbgV8MZYTWeE2d
ISyVzbHJYXzRag5P4L08KtCuaXKOq4o57n7GZvDXumtcJcb8bRloPJSrMtxuBhVz
U06Qz67M6Lv6njgfoeIDV82WAsA+DoQGDFRlITG5z88hDkU4jHrZjCZTBIpAbg23
5+q0ioYUXHkh/hLxFmrei7ppQn5NxhelCQ91nVORkh04m1Wq7+ogT6uWMn5DeLoF
3PA3dNOqBRUv9FqQdT2ov49GJ6tayz1+KhtwcccoEckmWcNHmwxnRV5VjDnVoYMr
qMyiSrlU+HOm2JHRsHyc1pHg96zyv87lizgQfml5OtBgmJE0MvN+degfhIqxMGOX
/vqrBxtL1VX96+wjsf7HPvwofpahWtSG76DfNahCXjhLWHMfAOgRlelI69up3ea8
jcm3X8bjFT/tkDJRsWCWuPY54KNQNVW6VvrFlYEQJeCnpmDd93OidKzZFe5tN6RW
t+1EqAkmJ62M/IcEBLTDchvJkh5diXMrqjqcosMWXhTxeOv4ai5lfPiztBUD2/Ao
QTArIctiF+X/aXWM3B3Tl13RMzGYfL2YYWFrJrm/J9gq119LMaaxpN2ENtWnt4t+
Lyr+y4506K/KJ426UM5fVYdTOoSL8EGe6/ljpONeDZJ2cXfmWVm/J+LROB0zMQC/
Fzl1P5GHwTKGtix3vCHT608tSH+dj71ffTMEB/a6tTfG4QVwuowAOxLrhY+dEx5p
r+quZqArmFK+wBai358PMGCKCrlnGkeeJcf77Ua6Tb9+bXqIMxq9h0kfaTfhl9Q+
Ef9Oa/Z+kAeHbKo/NtceV4uH2RvOMk4oGj7PRqaJ0yGjZ/C4qth0YS332Mcm3mu/
DCPT47OJTw/UJj+VjgWlf7229Nv7r8ng3cNwP5SvLfBAJ+H6Ui+V6o1z554oJk4G
R3fuY9eb+d0+XxOcWOfrmTM4Ba+igRJnJ9UxxjrZzo+Jk6Xez6kdRzAiqTN/SkEz
XVGRmQw8UFE8NyOY2qCDeci5gb5mofmNm7rOF1/i89eyfGWOrJG9HnrjL+qpp7Tq
Oa0c2SyfmE5dRkOJOl7cV7JMBZm5SrG2veC/KSaNth5hMgvVosek+QVuYY3ri2cz
kRGnuKOlM+6oFBrunDodWzI2taz30hExPFtQt5qdgQdVcpyHnwLelbR6OxF4xZGQ
unex8skPqdiHHydmIbkrCAaYW2cFvpQ3YNWvoQr5wmJfVn1mM6+XAHTS46QPjoJ+
6OSffxfaZ/M+qQtp49I2WG6Ba5cry2rWaa7i7FrRnCoWox57Wcz3mb5MrRM4aRtw
20nj6mLubMmjm8pnPB33dQ==
`protect END_PROTECTED
