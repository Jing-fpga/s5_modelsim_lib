`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a4K6b5R1Ojs5QMV6SnD0n+nFis2nTwZ/qnR8GKIIgwFcndliufmmePoSlJxwYI8N
9AMCZrsVt5MJZPFUw8kxLh/KVDNVi0DGDe2E/pcUKjZibaMQYrFXHyMbq+55g6dK
GdH5phd/ZRtFgjPW+SHl9BaNDgkRuI/DAot2DUK9qdYTLaBC+f3t4rqinBOhvknQ
bHxxEUbec9T/+tYsxPVLEGHjKsp/5wNHG9uQnexZwh2QmYxHYba70C0Sm213Af5Y
+DGr/yjqqbDvb8bJTaQwAU5C6GXaRIZ1MrWYIH+eLr+1C7wec6yiVr0qNUzRVT6D
yqYr/STcUCTYQcSqFwRRotLJ92e4lylX1+0hMzVRMNna8ywqMUGtOAmOYPwtALbM
/hYP51019MSHP6hLPtiox/snIHdH81I3GL6rhXJqVM3cEUcppnE5l2VSkx2N6juT
QCVZjtQ+vlYx2RCh3YNWARFw1ngrjDUlU5X8rLBd5yQaKASiX5ntMcVbpX2GF0+g
s5ZQCIMkq9/J79d63mtJBjvQ7XOKdZcfd/HVcUc8tQFRZpCAUt9tr3U430TRqPnG
GPsYC9vyKii7KdObml+YIAKUq57tknBYWvbikOmx39Yxu6E+SR0WSaFoSEPCe5fn
C5y5oKi8ix4vYvJUvIHan0Hz+DYmQzrddkJbE9k+gbMVe5DuHyr70T8jLYdSUAch
VIyhFLdGz5/Fc9QGW2tWapoQOnhtMZoG3GBs/GVhGmsDy8YwJaR5vBYe5LPdgwwv
LyUSfMpCCU58TM5l4lp6kDv91TssQTnYZwg39wyLPZlrPuBdJcD2IFokzvd7PXBO
U/V+HyBS1vzC2Ip+kER51Gu9bAwz4QvIznOmEoXu5VZF+45/aYQzf7vkASADitg5
hNyKciS8LuD7m+OgmTRPHv2mJcUbx+UDx2X36WIXbuW8bUxd0+/GDjpay7KekNjP
rjbtiRTIY0y6q1WbJUIB8fmexSCVjgUrLT5ryoc5C7GzdKN+Hdv8N/W2e20BX8lS
J60Hpz7+J3rrvWm9gGf+pB/i81T8pCmwP8u0ouWDWtM2Q82sGO6QYvJgpSSYVG08
kBZJzBNrXJY4itI/MoLS+/BrZfaoBkfAXbPryUUEh4Khd2CkSwYQBUF9BkGGgvjL
ULxhM5PPzA3iH37DDGzG9wzBqSIZkbiRYhpshsfuvfAqis2zUPBZbdF3G5ATc7Ye
BQLbOQkGfD/EnjIeAr08pIB3yJ3PzO3tPs0nNF97f7/J75esFGZ7XsYjMsyvB3Pr
FUUD11QiMN3u3+IAE3pyAjZL1SclDflYhaGVikgpALqZfjHZkIPKqu1GB8if9CZ1
nznnohMeYBEU1IlyASUC71hDmK/yVdd0DmP81q+vbLXUjxWaO1Y2CIloiTu+98M7
Doef4WRg9gcmKMilB/WJohoyOzD0GqoXV8qdQqduSEGwQ86z3wpSofUp+Gdm5G3L
CVXppZMSy8vANOpxfvvhUzbhKif00A3cUDOz5HlK8BLT+eRW0oeWO9dexltMGxdH
zC1kFhWjKIxEe2BoN1/XiCSPTZmYPx99TAfS5ebyki0LSDYn3ZSyeWgSH1oV7qgq
ZRS6QS4rIsEAQv1epSmcqVcebrOIzyIZnNnNlP9LCsc3272QdGXOz0eMJjR0RNIr
TVFaE/tXMMSp+SOOh1rgvLRVS70/mbicDLtr36ZGcDYNfZeyb8YdG3Jy7oAHL3PU
Nkm9Pz+ebJV3PU159BGaBkB0LeVVgeDETwbcA0IL06Q5YmW2w93tOtZWUSJW6xc2
5h2kj3CbpJiEAI6G5WpspfYJwu2sM3UZzfpSMMENLeLj7oOoNS/jcMfAoNGHmVAo
U0VpEnEmWBif5lyOQzkyCTg6RUQGwSqloJA4huNngvDUE0SZ4PoH6/CUGwLQcuA3
uBSdqNPdUOPabrHsP9wg4xz0R7hZtgAGKWLHlw4dka9hnc8LKprb+uaXRwMjl3A+
00t8gvJtTkBe2ixxy+4DPIfs6NIOrE/7oB+NaWfIsvpItzmKK9IrQrupEPgIwyMq
g2sa/rNM5yU0UeGXhR+kkgdWNNgQT5hsErP6c7SC5shIMEv/a1cMT/j7gm8bM89J
PXSDSsXb9wzcyus3Nwfqn0wdk0EJElndXuT4qK+0psstp2kNPR8hzdU6rnHcRfFx
gbvAN/497C7kVHec6R4h1V+mt8HxSSJFwBlxNMvCv6NoPVZn9zb6A/9remepRyPi
e9WIEyD/+YxG5RBatLUtgMmMoVcDx/ZYersplNYMzXiJiQqvpzNTlyYJUYb+Sz4I
FaEW1NpxgD9XQTdw8uHFV5b1sT5DC2bHiuIOd9orhBa4/ab3PdI6Bv5Lzn6ccvzu
+0H9ndpN9R5aTnCia84ZryBU2XtdUSRFpOnR/V8ykEku6UX9CCIdaTJXD0o4L3Lr
4OY45QHNgXtdk+Y+0FXK9tUZAcvPzVbyOpauVbh9JxH0uF6HM29YgKgbDNkEMVpl
5s+f896w3nyIHwrXNZAXg/8r43JfPgzUj4qqfGTEsD2NxGp2Bt5TGPMmvM7XrnjF
WJf2lmsKkD9flp6AXsW3VjdCy1LglEwuJimgrCPB4sIYhcFV/AyKm3U2INCwRBZ0
K6rfJVif2Fmx9ew53ISxkSu1m3fZPjGMi3H8GUmI/dkACvVGs7gYDDQFxzE0hRnW
cOLk336irjwt7Vi2rvdx4HGAdqmjE1JpVT68+4O4WDKSeyqbGOK1chAyYcG9hs0N
dZAy7UqiQwYATnrKECUZUm8NJXpZ9h9zedTFpfl9uuFAJX4v4YwiHK5c30zZcu5E
LuxQfyjeXqTL08iPqI56Y5LB3Ph6VRxYKzMrxRtgXHGOTelqXgLsrSubyV7/wtS3
bv7PXOW3WOu/RahntBH22N8S8yoYbW30RefuNsyjudW24GvZcQdSdiOG3OYmFSa3
4NLapVmmcrt+W+mpokAVqaj3RdThePINJoPKmY6Ebtl1++piBzO8i8DhBHa67xkT
maCyeRELX05BGZfP5H3XUcSu9m4iZD3oCmHzwx+boeAa3oaBGs6LlNf3i3gICUtT
2CdMIbVkPqcUVFKduN5yNfRUQ7cRiRV+3dJdib7XzszVmB5FjAaRnJKOemFmaCQl
pF6/S3dslRfYUzLb97cXs/Gtlf3dQnBYCsskQ8CA81L0DXfYUGbC5GQt7ofqQ0q5
FWtyuXR8MX24yujVNY4Zw6f3NDWHlRqK4VtKAg7/w1CEsi98WQN6zVtdiJwj9NJw
WgV9p4F4Kd1Bq/ynRc8YRh8EK/Ixdvgv6hCfoTjLetDUN3nLL/33zyi2VNukUoHF
BQJVV7yxMfj2Jd9yIuiOikuMAouX88fu9fMLHoTW2jE09aKZFt1c/xnUAa+3z5DK
34udkUfHRo+G0UuHLuPn1RaUC2UeFVXWGyzw2+IA9xhKT2jIutlFPn5vFCCq0Yql
H4l8sVqHNEFzllo23t0yteHlReTtkuCswcdrXvEzjlbJZ9id8/NJjOqz6nXDAoOT
+mqmUF8aTNN6nH4InAJVXvJodpRe4SyuahIN8Yi4rMNVxptbfma8J6mR0fMC4y62
yb6PLgWyNHkKdgR3A1LhLzC8a3kjA7gXodiv+pPixLc7scNLxeNyK0cFFJXTRTIN
nC79BHu24Vq4GRiTJwHMmneTu5XaJpeZVpyEqj222ATXeYilUKKDkUjRcTzIh74z
Aa01Sof4iEQr8aD2y5jv+aD8U6Tut+Ub5auwSJcXPh0N4WTrd8C/enls54SvRX27
ezh3X6o+TxcJm2mcueTZmy2+MS4a5jBeaZ0uDJakY8dtsfWFgkgyUel6nqU4SRv1
9XEunHVUQtOF9OlKolRyMJfZD8ALbVGy0JzZ8IxHggkAWjfa0wS9Xt4mY1MGobv+
Ul+yU2C9fYIr0S/Zlx4/Rhf1rkAo5xxMeW5z0EFbgOH18CRNwZ7eebZWzBrodLqI
gfwheq7fgRl+w8pT+yRoEdlmoI1NNNywVrFDPYznsjuIN9Gr6Q8oDm7Ym6dMfb/1
mF40nmSpNYH7XP//6KR/2ZS+X4VU9WTNCitHVikl7xNjQTqytzBIKpKWl0JMP3A9
eYC5HPRATNG3grqNdRJyZvU2jgXc0NiGC4HVd4DTvZuyL9tcYM1GIlC55zBMxY+5
SZ54WPyJQLqvn+AYjscHk7eV5tnpJpxmQ4QZ0I1KnQiStbJcLmbpLdzMTKftEusE
BwbSbLYumGvt43sUesTtZNfx0Oii2MavjizBzlDk45kLxecICOGgmXRtX6aVvzBi
frXFR8i9y0yYap/47yxwbY9W4YF6YcjuH1+SeoIJR7zslOMt3whii7UWcY40H7Rj
Kmgub0kua266WXcdVdd2SeZCuOjV+O3uGm1J65NQQjKroFzIQWQaFphfp4wRVw6V
ySWAmptXJUr3NGZXyEBHGenjaLjr6Kzt9Mmyo6OihAjGv8XeiAZozXtCVMAklqha
Sl0WdpK628yzq5ziB+ZgablhfjWCRXJtbXfr5J0vn66WbgPCvW50QABhEPOiLRCD
2zq3t1o+YqIAsa80QQWrnfJW4824jFJAVcEloVv3HANWOG5v0w5SCLiLAHDSZQJ1
sXd9EU44TTp5t3CC4WabntVLxXyTx4FWHp9t4MCtCpedT/LFHVJtpvLghHBiuFS4
AMbgR0vPZet1TT2ORchWP89P0DDM76P5P8K1oTWFdFY8x+99Hm8QgndLCx0zYEZ2
gcFC7BFSO7gxIJA/zZsmhldTqavSLiQLI9tE+J39j8nO+RNNu9mlIeh9DfB2ayxx
WV+mrAOVAL0oNOhZgMalT48lrzfgM+q3LGPLprHmxrkGnkmdPS0vSugXShkAptoT
63xj/pLDiScxXbCSvWwZXKYKxk9PMXHOVcesXtcGowc9p1IsKEMGJSperG1H2JW1
jZxrx78V47KmM2XJs6i+HoBKZciCfIOINQSSQkVDyrxmgwBQC6zRq0GsB2zoMPgj
40Zh5//OSxBO4BAmoqJfHth5Ch1utYzwM77/Bn1WeDutJUs4defgnlTgKLncle/p
FOZG5bIYfELS8dLGycUPH+wL7ppa518f3jOS1WOtWP/toAI/ANVhUNwknpPOuWBi
cvSUwvZ4C7yvIQCsOYZqmcqL7DW0zs6VnDrFOCYUNd3Lvtcrlu5qOhO5DupkVuQ+
F6nJGDzQhWT/0KKt/B5wl2ESPQwH+YHPaDiiJo46CWMYU4Ti1naySPcoV7EOE9rv
pH6XCBX0vPj5AuSnYqcDF3J2pwtitDAIBIFvVCidJ2q6ShmXi6RTPfEEtG0HDVP+
HdDIDW4g50WV8uv3TfZemhSNe6z/s5tLt2eUhXaMfHUwZlBqusael4oOPIp/+E+y
dsdQp6MiA+MYycW9jlYjGiuw8MSYKgfqkL42lvmjkOtSEDqk9u015jrfFTP+gG04
lFiFU+lrTDOI1qWBfNXwV8j7On39jNAvHXUorM254uXZULm6GKULhG+lBEa7Bk1f
nT2+3cCjxYac51DBMtAtxNX5UtIZY63n4atXwNYHO1pnd6E1TFqgUpeJPe3u0zn4
mzvOvYgZbTpk28pAMcEcBhtz1FZ7QqyFcyKYX1XzURu/0yvI77co/hUzzSQdS8NG
qZ4z6XXHhYrIov6Iter8ShU6d/Ivfr6Loh0Bi/Th6ZLAqVyoaCBNG2sdAxSn1fcQ
R1tprRhsEf2/my9sACUexNpFZfUoxXbc/A0UP58FcIL9BRnrr5UH4mZyVUp9LwY/
JGnNDh7JCKuecpywBMjHYqGBzv4Iq5KAMhTUVXEujvRQHSetCbIKr/LAFy+tVdvk
jIhN+WndxpxEkV4anM1mf/ydfXR2gTJVLqL4h7Jauj7p989pI4MqgJwZnvHp+tON
BvFg278+Hns8H//K8DRg+i2DYtRd3l0ll+GRmt8vdqtFpZRrpXnMeZirc2YdwVAg
734zKKuBr66U1kApaslJwwOK2Dmwprrc94bp4HreGSVaJ9cH+0mtMKRnnOVHR3Jc
JOsnqWV4BafZR2nlcNR+XTgYOUKyMKQcNiYk79GFrfDgwPN40vjH1ptlxL24KqPR
OpT6R8pwke5KdXywkAi3IxccAz6vmEVJ1ieooNPOfsjhRVKPMi/bCXDkKwd2Y4H2
BmQOlAkVfqwhndugIOdJHS5Yg7WXiOPedw5Fs5qcDtafH7me+ptfg/PGY6nBfAu0
XUwhc1in0jnk3o6B0Om+JIRmF7N2B4Fgf/pITLrYBJvI+ynibWDKdTJhwbRHoqs0
SbzzEVw8GoYYCzh9NJJKQ4aZxayXAaRuxjY3hgUTDt34tJTwSiozoN7qSjbjVHvn
rq4v0cX2CL3gszAAjKBOWy5pWHFH5BljDfsCS3FA/+qyEKTQb8Qo/p3bgqa/oHVz
WCVau+fLl9XwgfVCl8RSSMT7OmUfVhCMm6ii4QrN9+54FRnXqqVn2fEfWFSuIPiE
JRf5LuN/9FPISQ2JI3Om0ouGBsYEbolzxxbACaatNRpYoOAFXf8WfoZjFD03O1O0
vGw8NJyPmVKR2oyiUHm458Icuh3I6C6dqutiluncj4c47PwXNQpEB0m/31ugzTfr
ZpYkwPp8MX6mmm+lt5omTUBcQ99Fe1+x8BzM+K8RO/oW17iEshRR0uz7rOaaRcVt
dj7snqiX+HXnvAuzXwBHnq3GgPxRo1l8wXyV3TpHdQLyzSOBTOAMQvBNnY1Ip6N7
NbrKFXo5LlY32SzfxZZg1ho5FNhFhqxF1Z2bSR5iuuxmm58jNKC7qJ36EaEVbGkP
YahEtMdwflyN7MAZM6QMBwhqMN3SSzGhgW5ER9QpwlImDwdIsH0JJClsSJ0pb32v
dRsM2M+yduX81w88jyW8sVuxKwEzVA7rNG/2Y8UjdQHeYvSBtrX4XxnWCUwz2ByB
U0YGOuM/fDjNSqavx6rZaF4agSlfRfLMl/suYe0/BWhPFOb9pGFyAQ2bYhOL5rhS
CGcPIZka44zgbkVUQxrheKZ3ML959egEjcbinAtpFO2qjwNGJvj7k9QFpTfJ6mrJ
tmzneky6qp9OLIUe6mH1tVVaNnLhD4oCgB+HBgnnwGeUP3YMDGVEbbrROI8ycUri
HzxWO31Sv93fFbjcNuBm5NDv04wPZ/dQaFNVZeWRHtC5TVVmNguV452Pz5+Mb8UQ
aX56h5oCDlACGJacqvj8Kzj5PhyVkAITCFP6ScOhtWOq+nTgqItpDf7v8tOxp5DL
cJ26EYmvZCSu0UJG2rZgMB9kjcdVT3NgN60mpc6MwtKN9aCAM3iJN5quZhiXQdEG
aOIHbu42OKD30Mw7nqRtib5lb3+NtquT0YvYOWzIaVReRM+sRQKrDZipZBh94aV8
vRPsyG8zWS6NQJZCr5tMjDLcJRGPH/tNSv/k0Lk38/pLIrKPYV1cfbZyh1zCL6aw
p+6OQwVbaKhf928JNClJsFrx35itqSfsNbgo8iXOSRR+FXsU8Xfo6ol9M54gztoU
jttGmirlW8MuAhNHh9ymQUt1aEMIk6i0oNQCj8WubaAjhZC1VdsPZEtNumBhBK8I
+fHLnjhh6Rnyjt/ykursZD444Ym4CtBXbFfI7VKekCHtvUbQ25FU+OCsAByUnzfv
MLuzzkIkOepe1ZpmCeMIHjHiq/tNZy95J4lmjCDVK8D1ZY8dJOzs5oad9YJTqUoH
TcOeO4UGEjpiyNwxVvCADCRQAbNW8pjWJX2XcHnkjquLQRHcrLot5x0zx6v4J5cw
YHFDq/pWUNmwKtD3LcMdqAhcmSpyhIzP5Hw+EI36Wu7ggdJQNnvwmsAsyvjj2mT0
Ivxb8ofxvJ6ieDLe5rlMUruepsv1jueEvYb2VGxjvMUqxHqry/hlPlJoxC/MDWba
z1fEdhHStsMXcOA5/NvY9kgbFxS1eGKEPMTemdDASDWBWNA73wwhSLPx7qPydEPg
7FrAm+Q0fZP15XZ6YMJhxRzpp9yxUkKvR8k2rDvj/dJFY3N5JNWfaJ0hynhwZJCH
OaMENAfdofmRIdFOnEFIPyOGTu7AylfWicYUVv4EbcHucUjZxVJTzyfC2DO1uZMr
Xqhn6bwC95pcnhwGZRKQtlbPSatHdMzzopqJjtCEevBnWedFZwJpX9XlYTziGZ2d
dc+DUOlAXW7pC+0kUDk+L/VGurhNZc9eMJdkYHUfpp+Whcn7g6xyHe6FCRy17cj7
CTd68dxa+Kmt7emu5559a/YowZF2FXj6Zj8Y+ugZLEPHSjTsjYBiy3kW4EktRxPJ
AXCIX7Htq5ooe3FWkK7OSiRlOk85sdPwsBuT3gbkkX+4O4gtK2DKD5cbvLtFXeXG
rwU5mbVICz0TRcMmlxCgq2lS0YIldKZdTV5nBu/SOkwoo3QHLGsVOq/MT45Ld9QV
MgMsBI5a3cOcC2ZVAFpQ5qhcUjyzrZhgdFGFYn6+y4xQmSY8+ouUhmtThJVFDE7c
qbOfl3K6QV/KzMBPPjaqwHEhJkWxXS5TwK7qWHpB7LD5SruZnclBBbEfhenvQFkQ
IS55BleRYNlJuhIPfvTGvrbDJuTNkTQ8fZB+McnsHmhBYlP+0hTlG0GvNHqZjMQI
79J3juYmSsGX6KcV91wkpeH3sXkBB+yGO3ifZzTKjnjvXUUkplJcdQGs6rYJc/eS
l81cOPuocbsHYQceYXkB+gep+varOlS3CXwljN7EXlvFVPUEEmG0xVUpt6c0fYGx
Z/areF3NkL0hBpqs0qKOOHD3NWURrdiaOOe9In9E3gSxWjw15n0yC0Vy5xQE4BQF
5kqA7fq0Iz3gy+49c/fOiejHrtIfGTq8MaAYEA8Gq+cc5G71ZlEaJv/rW3Ipnihl
ry3LD+qFFePJ34qEB+QbQS8ORPamnHGbN1w9st0td6NbUMtKcU08HyMShIaYwnV+
0olow0Q5ewKrMGwCBVv00HGmh4Xbt9fJiNvXs/7sicmepr4n2grWfRGe/k4aHc/P
VEGxuEo0hy0jK6HlBJuaV02a7yuHolM+2UMO4TSpZoO7P5fHF1sEPBNIReFEJqCM
cSq5XGIanXUJ9+vFosJ3hkKvN9Dv9FOIKw6HgxuCFOLGgZzDZOgSt5PGDKjwWAO7
cPHuvBThXFjRObCG1EPk/zU1Xg4g+8zsTJkBUtKKJpgWFJjRiKurl3BgHJRih3GU
+N3kERzii2eW8Q3xEjJVwg64XzjeqChe4KJYNrIKbSYnHMGeei624yHX4eFd66wt
tF4PCphXx1qxkLXyH88W29a4hQ4f7Ay4sNqe/vuJjTXVIXK1omsckD72V/O6X2Ol
zQ/EFlENNMITFjc3AiHyYDBM9I0bdU+V1O9RnEBrH7ss8LjM29Vu/DkDpkIubFqx
og65I97HK1XQc8C+mAJ66Gp2owLLgZylWHNUz2rUoG3axm3/Jfcd77/p8LLUXN8B
iTPKOxY5kdNQCyaC6qBwTVKJX07gOT39l4lgQUy7pIY2LR2h5aIURuz8Fkiq4B+V
eGVrkw7rCowDB2PGZ+I8MVF36E6b+vLtsGOoyWPA857Vd+y5z0Jf76Vaof56f10u
INVYrrEcx6+LlxpHTqY2g2445VCyQ8tIHKy8CmcgnJeRjZfzJ23BtF9iHcEVNAvp
ZbtxtjG2M1X5F6i3JhtPDoryxYYXCjsfW4pda4xLgNwDB3ylOqf2GbWUtDkT63Qc
b/hTdjBz1dY4o2kkj+H1oHyqsFcPaKf806zOVEPU8L94Vx30ss6J47iqjt9Rg487
bR/z5dvoGw5DJbjENQSrkYlPm3TH5xDQ0w8SCNqtmHE=
`protect END_PROTECTED
