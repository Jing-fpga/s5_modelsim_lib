`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zw4EDJxCZJEgM7s8KBDo+LWRY7oUSCMVuYFWf5JzT3XABRXPXrCH3ZsY4yoVyczx
Ln4x/XEigv68uZKgiTXzeSidD2X22jqx94WeZ8dOg+wSBA/CKLIrzGLioBLSYoGE
9Y/VDrFYZTkPWmptr395o0e2gr+Cm/ejZIFY/aBodCPGxF8lOGDtyWamZIIcQ2CD
xufnpYJEo9u2toAKSCABDyYgqM/SOUaWqaiZRtULYuckjvJ6MPGDlUGWhKQwDwiC
BC5TlvzRA07Vz5qohztNGhJEL4MTqMecnCMiAzUDVvjmbG2eBWSty2CLW3QS3RI+
RChYV+RicGlHe4dub/Bcd+cUQSEVJewJO4nq2/OOvmdCtRxzl++8uri+5JRc4GCC
CKdIX9sE1sM/E2dRYlsK3hAuabPBgectyVS7fWyvPsGF7+nfS404VihFogUCSVKQ
jugdZBkC3mu6N6SOjZEfcjK2pD2ZHI+CwS5j8KgKmdroXPLGSdNUzqNBWbdTGG8u
FVw7y0E372rvXzx+H+g/vovVLy61hpfYi3XIzQSdAaXCbEbADINTOWmJo3RBgCRy
2QcSeVl1HwJrWW+GyhjMsrGGtEc5AA5Xmr6VLbT69fdRFm04+kVHkrkoqSwydz6I
t9/HGSYz8+jo1FvR2zaq5CqQnk97GNUHmiQGk7BElxpOhkoZEgAdTJ/XevTp51xA
DIGGRR3N0yui7a1I23akAv95jyhJ/+6/ZZjpBWFdVo7bpstXR7GirU9ZAfexHGTR
Bwpo1gNeGgW1YOMeBqxbGizkPVLgsDvKwPQtZU8VZBIAvtmYM7N8QCF8+bNDb9pm
QxvlQnxFubtZNPXkqQSCTOWzkoqZZy8tIqSDDkNM0d/RTDyse7QRsj2U/4KdZrTP
IQx2RuKPZqVw8k4e6BVoDlXj1IoFzzdPzEEqmA3CZGDJsVAaUBmHoLDiULC2PqvT
usjjuzkCpNp9CcHPgrf+fQo9zVR05NrY4QUsoTbf2pBWGOMSv7ctLXCXcWpcfXio
2Wg0aaQhkHxFcR/1NxD7ChnKXlbi5P9xPqukDfiQs347GUZemMIKMIy/ffOTtZG+
5Xowf3eRKv1QQa5k27LH4v8DCdmts+1LDexD2AFAJ54iTTYMAfG06+lR68F7nJu3
EZrQF+jU5xnYf5YAQ9M2FOhlP7pQyXI3s1t5lj8ZWTEwxJcXcT/Ka2pECqAQEf25
mgpYq1kGg7zNstK6WbF+Kv3zCDhDnz1AcXXrietDyjBoJBa8iIFrwotATpcJ4pcW
VWa59TVdcSMctt4MwIrAhs4GD8ZdFK0ZqwDKiV35s1u7OikHHpUeNavKu8wn8GkV
oQg5oz9M2jkXWhIp/7tiMaHShk+DRybAfhHrkltdwhNiyiptJIUG4JyVFSXiCm5I
0CIowRnHzf8pLuwCOEgAGjnnxuKMLAz7LQ77vtvjJqfflPLqx9RgpFxh2E7hoSTZ
FgupSE+3bgLyXtCM4mYu3uJbPOTjz8S41Z13zEsBw03igY2VGB+FaCWLhnw7aIA3
7GbLMeXvkGzDoWZetZuHhLe1JssFi4W1T7vbxX43mJ0Oidf12QEwuZBT6W1f66bU
UFf4cMh2GLADdNgyOQJFq5j8vcpXIk4eIZf6ablC+DveYRkag2s326GPUjci0d+Z
1yGiyAfyc3KmdAVkn8nibieYcbiW/agJ1xc+MMWeYrRIIFKIu1Nq0hbiQuhukIu+
YzG9yze9uU9lhGy+5Pzr6Znbixz+wzCLd0mN8Oa8rCUVsHi0K0IcMU7bG3TnwuE7
qJQfrYnD6I7lWhwSVF+JG8OFYvw69UDIe7sd/3JSgTdJg305eQ52ny5DGn3gQdhU
alJwvjHqBnQ2DvdI7CQevB9nzz+eURocS1YyBT19H97riZCfE1Ft0zFRpfLJX30b
A5EcWdcMuviPfki72EjHiXcxEWJAvN/itBqIYOvnYdMut58A46zoeBpAup43eNCi
lM2Uyc0MKomz39+y/8RWE3dHO8irJESOd4PV2YIkLDmxm1Tl/10Nlhpukq0LD1vS
RJxoM6cOCbI0jeKozG08+jCoeJkmTYM++lDJ0xCNZMHugVKq18MYObo9aYD0Pula
R4Vb1llGRKQNIfBWLBrduOJVSCLdqjJ5brM+VNrCLZU6wK6FhGqpjeRQb7aLR+On
lcP0UfUhjnRsSdOdxnBggFX/QMB48kFh1snBzKNgduvTIGQrkxGiRHc7NHQd+b2m
69kCVaEbYMU36iQ6HNUv8zzVa9oTyU1Q5tLVu9XjzlCGVvzf9PO4RRXsap0f70qe
qbIfQMFqyEjQrWJ+LYemuybbNkNn7T3Uvyg5GAB8vj0UOlhAZqfuG8/Q2TLp7yJr
59/+Y+LCGQrPwuTeTzIobv9Er9Pb6msMbrRhQ2S4mbRDnUSvQOsy5oFHILpgz09+
lNBwv45j5UVKqn1yfQlelbcConaCd+cN+WGu1oLqNS8jUh4oanwjR/lbXDbW8S4c
Jest7iHSB22zyxqWgpn0WLQP++/os7U2uuwZVYmrA35PF3uFH3Qf1Coe9v3Ti6sW
iTg7AGe2jPWgPuwh/CFwHdSQnbhg3HKpQeoNnGqR/+6GVZOV9wjRZUS0VaVPA/2t
FkzaLMBF7tU0t0DFP63ocuOTxpFKOGmgS/tJwgbnT77LAWaYs8OBlAdkF7AQ5oY1
44XoX42eElQ3gs4kQ03rr4tSyIuif1V3NJJpTNG+Aubpb/caFv0EgdyS2fZb2wq5
0GDlZ2wk/zQLKgWQgdMurm3xMmIH3rUsNJ6geWhwhkXb4VM8WaNBjiB4EEUSMpmn
RMYwaBGy5/Q/STPVhQFSsLvQqB0IGyVjzsU9r/0feOC6UuXsMI2Ybp/1fi/oFURM
RL6vG5VX2+iQcG5Vx1bfCUwFGr7pb9MDZzUalMWcjcHu0x4RbH0DA0l3twJCpK/s
CPK3+mkTN6/cIPsuoZJJ1VYK9dcqektqCV0pUX0kIalMWXCqjkl9j3VIydXJrj3j
5f9j509RQCp+d4zQdlrs2Q7RPlESDLJMKkUtc4u3rPEZPkwohDvxXUZ0Ul49uzQ3
y+N5XwHPHEdAEmZEEqS7biSKH0NN25UgeOyqmZZmIGPctuRWmcj5dZlHamohWQ0r
cPrqqUuEYfVKCZDsOd+40mhaAikQeqAHH2gXNJoN3bLep8Hjp4ONFZEqUIP/VW0Q
BCxsJX8r0Vl58qnKh0mWpawr+Intivr0SOM6GeZbgEQtQY90z7cjbf+6FYFgFZm3
E0aiO0Q+9+tvpfHr+XHY1+k3y+kPil0dMBoodnw3sIH3xR6GdJVcfSourRZugyr1
`protect END_PROTECTED
