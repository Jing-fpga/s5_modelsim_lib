`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h1mieRJmTd/PjjX5Ggitkh4TZYPXipzeUIYLZ75946kQIM7Py1uIdPZVSSSSj1Le
gCWr9Yqyo6DHFb4OcTTGXjSy1VCgSiBt2cQWcuVhjIkfpUD8rB7XcPv5FnCrR5EI
49KxTQFflxbM3BV4EogklVs8qiFCqeDDP0EcBzwwBn9dzYKRYIjZGeVnE1XgD6it
n3OPx6jPXEgsMGUyBX4oPeXLNHWTgGKKNuyqLkHrdyj9ITq3GELnEtXFaYjikfZe
aOkdeiV0UfjMYsoJUgT6A8ZryebB7ULscbfJwm5WsI5tL4BAShSE/7RTtli+Xdob
HVY7toOLK0/CLksd7QVgFikqTzY+iqcRBLZWxn26vJlf6pySQ51db6RBkgfXHOkG
I/wmJOkdnHaaHBL2xYvRlLQiqLIJ4jkThg+qh4g6VY/eCi8agTZVIxn7ZGkUhuJK
fGoy+p9ReNAuN2JhOYsCT9vWEldpFVSbH9kajgGGnrgVOlYjxBK2kdhXpEs2qWLx
ZGGXpFQYZv0YEAZcZA7m5RHTpiy/Of4XdNSWrMzkWKQFItu8jBDgOqGaaoK+s4PD
YJjT9eA8v8/TmPtLLp/LbGnmogp1zWD93pam7aoRC/Bo+E+nne2Nw5UPVLt/hbXT
WCOx/1yMn5NPhkrplDZyhRvny2hzUzsXocaJiT2/D2g=
`protect END_PROTECTED
