`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
flFTQpgVN6zn5YzJKYONV6GJMJCx//8DErdZVoMn8zcgOVrp9KPTJ1l0i1qzSBYK
tE9BEYyobYRZjf+2BmbiDOFLKeooBCNpzd96JXor1TxBc+Q/Ps3fQDKZV1t3i4EV
nqQDsdK36IMfI3kdpluQ7yR9VFi9/rQteXSrfOgawwHWvFlBJyExEXFSJAOKPkEI
XVv5QIpuKzVifE/otisFvxbESjCDdd5cyomnNsV2BBFgeo3l4vsD2Eh60NcAMK39
xqH5kN0KWbrifWo6N3GzwtmieoBUJ+rOpRbAwsdYVC1VGXPPBySteYCVXqjV058a
bKtSOr8r/PIRJm2+TVcoPog4uSGS18toqlepcbwq58zwbrW7MaGL41PXq2Y1TMt1
s08q13iylSWEweJUfNLeygEwn5NhxCv8KTYp8KsoGW+CkM4vAh8fZdffvQkMh8Kd
wz4cj//iZFHsNugtwYi2GYBaDPzTSwAASVOTa89oKk+QbdSOG4dtHl8bTh3OySuu
g6E4GkB1/Gx4VevObOLppOOxwo/7VVuzQYqslsmrUbDBgQjzxoJyzfEGfmwEOiRq
+YerNqUMk0v0jL7kZUM87E8yxt6mOZgrrVIXHg7ELv+XJEJR67hIGsPZvtmXBKW2
KCdZAtL6QuYtfFI+PQ8k6NViUVTe3C96LbZ00FqvT/z4+iB/460/VcrqKnQdBTHm
vZIbcttAeFsIri7vFZWdqppiqmOAL+jo72xZjepvZmeVZDACQYnE2bCxBCr/MSrR
vQvYq3Oga2vuOGrnBr6t5XyxEAXtEKqiNGcFgpWRdsFyLlSCqc3b9Syql6kDV6kg
cOw/uGikchqWq7harZochyqt0HZ1+bFrhL7Mh1GBP9zFwJVZ6myscO1Vf2VDcCm9
GGDlty2/GGD6NCmH4bf6gZ/lkBkrSUiO5GsY3WZZYYOeok4UE7pckk+y4gk3nKNr
zk1IWQrQYENLvACDZHiRqaHE0ogvnXH8TXHG939SH/B8YZALcHcZZYde+aXr7yYx
8LS5MSOCsK1H/j7XxtgJK4HQZ6g5j7cvK3X1xNYxtV/CiS+TczRwbMoXkgTwxGiB
F9qA8HxnhpEK6mqT3KKqBpTI3/cO1E2QQ/UUbL6lEIDubxJTSIc9vbzX0oQxhaq3
GMK0YF+wnj8anqTjUAI5JHM+BMgakGuXhCWLTeI8Bn1Y7OjS7wvtMzj+D9r5y+pT
28UqA+GH4B9Zo4q+q93Gh9Ao80hVuVZbw3eQJXuDfSoP/1lUhePyDnOm1S3wFzna
0xS37SRnq60iyr/712jiMCu189BgMnB09b/VZZHTaq4UnZ5S3J69/Eb5zGSQcTkU
4b8yHB5R1ImGO7pL+Da64P7jRRO5zQH0u+njYRS5G9k2vkIp+Nj6ez70Mkp1rglA
Cr1hxggOdfWZN1VX48ksJvh5r6cdrEfhyc/lHWFHMqhAi7n32qRFXaL1dwOCicAT
V9aA9uhwy0KMeCkKqK0Q6s6NUVqCVTApF58ExU1LWSOuIC1X2PTvDtJ7TLjkszbZ
qqAYONdY6+Cu404EAuKvbetSMcp4hxf8Hf7pK19MAu4D94SoylwwDmYqldvYjCaf
LVnFUFWQRThTwG8kmJqnwq8NA8+giW7qfXQtwKjKSBBFLNmE5nu4x1RqU5Ij/tK9
k1atnZlk027P1r5fd0F/1R/H7PX5wuVq+0LYbKLw/fdq43DMnbEa91pbByW7rvFo
nJ6ivhi8txEpeqMLPB3vGLIfIFue8US7dM2DZMijiWWFt0hBo0E8fa+YOi+3Y+Gm
iCf8Q5aupQilz5Im4ambMima02lwhFDmpyLBG6BN7JHZDKMciXIynVMLLuLxUD/w
BMFld1F3YvvT7k/kHobUnyVna74pxktuBjBimsoiwts08bcVpOX8B7yDj+pe/9Bt
gpioF49FfMjOaDv8ZzZC7jcpRwacMqp0zImEw16vA0cpEWtOuJo05gw+JihwRypL
AQFMbz6VayNn1LtHCI51ZohJf27k25VoPuEYjo1ehnyDmKflUs0L8O0ntz/EA2Xa
7Bp3Ji73vzuz0pFHgoEWoEXp/qBI5VWMTzbGsOVkFkowdzJp9HgYrn+EhPJX6018
/2GM0D8JQoysGRTNTuNUBPcvzBcGlex01a94McswA6uocYpXdaM3g5XaIrbyY2w3
MfZtyGl88gfCVtKadKI0ySGImE9C54J/ciP/fhN7NhRI48chJ80Bsmmy0+pVh6I+
zz/Si6KsFaE6Fq36O+8+aJog+YwlWeYzWFdHndS6mqWsBy5y84kDAx5kKhYomCNy
OuSLndAsTq586y6c/GAMIdMrkwrA7+n/Hoc2foQYUbHA8fo/a/8+Ml7s+A/JqCAf
8z7WnYp2oITqZT2n/0b91UO8UC4cDANZ303Q0YvKoJzlg9M/OM618c4iJrBZEDrU
XZAgM+dDdxFuKxP1Nwya5pNeunds5yxFA9HHOXYluZtuYxNpsrATAgEupa8Lp/v6
Vs/TzMe3aqONPCxJBD/AmW9s8MhGtHjVLaLkVrrKjX5NedUy1uOD4HmZlwMGebSu
TsNtBTtUJwT/770XzsRFSpSnq4wvPnFS/bHg5SI3qHpNB9mGcV+/sg00sYggSlUB
w/Ytd2US/7BwU5N+LNEZNpgd1Jn0X85cq0SXgTQWO0wtjE88cgPHHxqDDHeHD7rl
VC4ptzOxKBcHqK/XIOTJ9T0n78DzRdoGCJRAVK9yA+y6hgHnnEe9ldqXuLWpIfco
DlQVEXvnqE6EMtDXqPfvaNWCaJmqKt1A6tj1KnCwfG8ZkCDfjtxXbJfNmrCZk0Kj
4LjOZeWvY6osUIe//HZ26P6U2uc/FGE90CjzYIczzMnW8rFw6jkMRKUH2XRxW0M/
tM8REuCpvOJxIyvWazAB16qzkbKNPkxTtfMi3yg6PSFtymc7DR71r3QpiCeTxfEK
Rie8dx+ScDpB/CK8u+7Qx2Koo05HJv3Lhc9iMaYjA3fRzmjJ7obsJ4aneUMadmA3
nOlPJtcJbWF01Qwa6Rob31fT6c/BO/LxHGaqCkhxWh+g6CNSo3fwZ5X9iJLnfM/G
H3lm2D/EbXQ4sDgzfp1wSjh0wyZpRWRi3F+CUNzMxt8evBpnxsC+hsv98wWEyYMJ
a6XYNwKpAm0frUp41g5UJSl5jt7dE/J4ZvETtYZFGlS7M+2PBJw0kzO1PA3clxsi
bfk9pj6EW6mzScp3CZfJXKkm0QPXXc7bPlEa9zgbWrCm7Y6luR8Z+5I+RbGlUoby
DvvmT3mYOuOk71dzcmAFvMmk1YxpqmWF8IH6tEG0F3Q6vl572uk3PL4PoFPHjTsW
9GNnM+cQl7J5GPUyoHFDNw7fiJCpK5csZpw+mqtbSgBCPygJ86s4RMmtnPQz6IZW
m+bXn1Q6ZVplhU37ePJ+jpxs9+C5F890y2PUzGCdNY8lvM+3qQ6XpojwFjw8RT1V
+BNwoIMVXZcNudcg9Ljh0Fqsl/YG0ggOm73QIwlItyXE6UOuDpNpNKpVOBy+d+TR
mYODQZ1zebm/WHHUmVCtXXBr+hEeffosYSyM2GR+1WOjQErKSxIESgCO/fFAqpw3
8nxmJyFwns85BMqc6VuGTyMQ41b4nL6KBlwmM2Xn/iZFO49vVxLcBExM7ufw4JRd
Rcl/5Ref1Lb0CVpPegWH67hm8dpUOsqXCKl01HDAWC4ePD9EsRhzyHEEIt4Uh4pC
CHf8ZX+TMWGEavcWAk52C3Ucp6ooKHXRwKundr0EzBaS1KxctrjPSij11aTESlxg
uw9NITdpGh2OOx7ugB6ga5Xnc72XrD87OLcq9Nvtm7viFDva3dv6+fcJ2adfwIOl
vGkiaKVfTTQSmNyTjC5t3kkxF357uTtjYzzvQbnRCPk424Yovmx9O8cwZ/Yi2tg3
vPHtRcz/pt2VaiACFV08bHU+t5jLh5TbhoWwCBVUW7tTP9ExMO0PsQSmKYCSu/kM
dfeVb62ypo6UHIak+eD2LU114uXyqp6GtoJbGLDbwhrbqJxAE7W4Xts4x6wllMEy
klFTNIx5SWTcW22iO7ZSKiL+NlJC1X7WVN/j2WwhVqDmuJwcOEQfiiLWqzfsQ8y8
UMynDop8YjvFsjaNGFfTZlurcb1TSSP5lsaGdG+uf/HR8CqwFgDmzjZqKV/yoDjM
fUhrU3PNe2JBHWE3/Dxf4DmTWNoyNztiMYabBlQHK1NU3gMf59Ubse9OUatGQP+P
+e2PakojvMY60T/oaJmFGe0e1atViJ/g2Spk0CfFGzwq1bMAfi+tzkgDn8865SqD
4ksDcX4AYzif/jLoshE9Yh2d7Nd25ufHQtvE7ntLxYQaMkylRBowNvaAV1lxT16Z
66Nxkx9ehk+yMiMhHOKYQdjSWhcdAAGCkOY5AEqlMPGHX7aih3GX+Hie2ds27pKg
JGpUxyfu28moju2MdvyFlYphXUMCvsfMzpMmINt02JGz76GWzd9sSwAS174cTtLR
XG+1u/qW/ZblIrOCmi7fbyBZ0Xs54/+m9Y7N4jEx+3Sz9JAVkQhypazEaSyyIo9b
EBQmqRLWcmFDCwNS+1Nf25M8V0mvPQQ/XGNPLr+6yY9ZWGN97a6G+qskLIE9NJfz
/jWzo7mnUCrprq3WP07/uW0PZf1sVN6fh2HAulk1FKyIapGXATrl/2Akga39oBXR
GksCqoIkycJCBf41Z2EOJImldNxOPLgIeZkKy8K0i1JWM4sGieT5jzVTWWjlbPs4
N7qjodJ7RtTzIdbsu59LohMO8pPTlitxKbPih7b64fhkSxwH1xTfNqqVXcLPJQYP
qk4f0TU1QO2dzgiFJTDUKxx2VGHj3YORJRt1678JdTZwzmVUBSie45NQ3WMIQt89
+/8MMFrnPLZyaNKWRK1PDO3NJxPtNTaqUOD02r5FwN+Ut70csnY+lXga7xMTev3v
jwyH5yQpiDcGVlxUBQNENzYHzZiOy5VkbnxZD/HcG+qVAPM6nLNdnpsY8CXbBnIg
ZOQoEt5dS9wF4ZpywXHTLY4PDJhSOzk/0g/Lfc7NgGQZpw2R39ePAjzLlU7XhHgP
R3pRlUE/0RwtJvn0B8Fzum1ONFSCmeZ24lqGnZ/QLEAK6CdmzbhqPapTQ7OufSMY
ve8quOc2OkS85IqDNeZcAlPEfXGQccSLX2I0glcc9pGHJkMw/xgCnKQdx5P+3TJ5
71u0X3HyLJLi3T49mMuB6Dqir0smMkIl8cKpakfC/w6Fz85TOU5NrbBByF8MsRZ6
x+k7g9OvjBdLaTDciZCR2aEoMGlRaAvx61Rn4U90oQ/dDl7ymaMelo3kUJy5OUgi
jp6HfkHBs7+ZnYGQiUDMphH/kviZTXcn1FEBfk+81x7jyKi+2vOxchan0L1AsR4j
kR1Tnq/t754NxFM6S4zxDaSDIH07qKDWAZDxdVI18+oyHXYjPEGpyNaqXOmz31QE
t9/Y608Odwwmi+pw9Za6R/yc5OICqvJLBOf58OU43JYr23IOxqNH3/b4dpoU7ho2
BeJTOklM2I2rkZlUnPZjV4XD1jNJucYX9NcfTNt8PC3b7QZC/c9Qw5jHMYMt34pv
X3wIjVJpN0gW3iOQnakZm1n/Kua67tJfg2UB4kiCY45pQ+mgpEkzJZDzHaQ6xav4
1VehCw8RSIpB//K0qhUVmR7SQYAPi0zFFrQnrf9yfVDL4aoVOtqhomPfCTp4yZh1
n+NejS5ks7mHoEPWiWWBxZchZCPDY/w2Wf+zKwAY0BH1h+fKipbGCfabAiKmMsQn
UaBYwlvow+MKwcG7C8RJl65z2iAW5vecW5i9AOn+f8MMVJM80AJnhyBLxIfdsBkG
ms0BeLQIqtc6zrK1BfYMaC55I3bzPnqnkCVXqBxNVF0vjcFulSDnW/veRx42Awr6
wAogqYSdN9Orp2jEMsC0sMZJKqLpxm8oKslDZ6DHollMZSybriRamlQdHz7pBgJp
Io6PP+eT1KeBU5Y5GcDV3Lfy3XTsrSBjja6Xh0Uu4OcCSFLFgbOKsiLZMgd/rjKz
TFiSEVm7y6Pe2q0Fp8GYk4Kb3fE7rc8jypJqrNA98a4GiDt3+uGgxj3HkXyLNEWx
V2ogRPB+TOeeJ+c4C5kbhQxZ2ffALqHKZ9QMhZoxAzO7tkNuU+SwJoqwErUloQ2h
e8OT1rve+KJB6dK4eEhzdxeAjrTFrx89JWSW1X8wcLTMd5dMN5K7HyKcn0XWps6r
JYccz/z2LL5jZbQv8gY3Uwqjil7fIoeMSQrRnKdICMThqHEoQiWvRxfa5UcfxL/D
iZWyLSm+c7VeXRaxEX3X1ImxXztS8wtxg8FEPHciqLfCKLGve0ECtxrJmrhK909H
AUW1/K0Mp/65SIjSt5UmFkcqCTTCF2i1rsXn/52hYyrpFGp0QG83EHz7mGlOFYaY
IyL/3Fx0IfYeMhdhhxKyCKp9FWU3LAB3rXpiu0olYKZu349MS5xLQ3tBGCC519q2
Pyy+5ISktQ2OytZ9ncNhmb9SyWjax0zi0W3irXIPAghQN3330NDc/3SNMBAIjPor
CaAkSogp5fZPPt8CopVo5WTcFJyMjUkkdJM1/ynJH8nnWPTPcSiM1LSO+qBXnPgZ
dA9DypMkU8roziDuK6pExNB6Y1M1tHejYIbL9zTzYIlM52yBkWAWdbSOUk/5vR2H
zdzZgDFScjgz+JzYZmypgpxEsqQ7m0AR6W6rDBQ56Jwethrsam7JZfassBqjyVra
fq4Gf2M9orTYpUrXt6v9Q/GA4KcXKdBBUQPox3n8EOQ4dGc/2k70V2aCPDFS3CYg
YXnPmySaan/Ob7Hl6SBkPtT2MdfeVB0w7BrCBbX9TZoA05CKfEHDybRscKShKmpC
s50mI0BLcZM9bIm4aSscJ+Qr2Hx7XVWKL/4EULoyM9XQOVRq8sok5HTdKkXIUFdD
UKJCQZNDFSCWGQ4HPnKiNmm5IiiT/qqobhNvj8HNQERPN4In2iiD6mZTDffCpL0c
Tx/GKZ2YJNR7AYod+oVgfUEPMyoiGnB7xdnSP73XZZ42feRWtfo8JJ2tpBEXoCGN
PvAluq34t6KEORTqv6sNvotv8sBkgLCANBoTp/qaGMA4SUEETJt3R20cQXeCcix8
cudZxqJdSeZPwcszoiPIaxf7L5mBjNaBvRdf1bEwR8OdiZOfrNwrgV7mkEmFs8rl
Hxoi4GuCdeVJI4jXkkHw/nYkX364ZYPm0XkgdyBhZu58QdFgEWCIgFWSk9wv/x9Y
QjkuIf+zxNeXTX1B3BE6Y5uZzBsQIyjZ5/IkHFBm8tOC4OzHqZQ9VTHJJTD5bYtq
Z5cNFhBGo8wyyeEruf1ILaYolwA85HEGMr6sZ9ACe3u2dMkadsYi8l591/4i4yg0
BtDAxVqOa5tmt+mnBlBEbjuVed0Wl+gKs0e0t0/x915GzIT1SKnxRPcukd9+6XnH
MmWWe9gDUgoQH8Boe2RrNG+3RMWQwcVt/LwdYNh2zffQlV74K3FFa2es+TczbcNX
`protect END_PROTECTED
