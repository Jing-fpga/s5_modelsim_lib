`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g18O57SwYhUSA7W8c1FYdh1AVviS2vzE3yPWzfkaTZsor0HO8IpTvuvvIrnrkNg8
+Tl9FYg3KJFip8sLu5mRBoIkoZAGuPPm+YLK1IQWzTSzHwmk41R2DHlpoCSeKsXV
C//MKpffHjOTK9AxiPmX6dr2PnVOkBPbpL60m9jiXlM7LE40Qzbj3a3d3aeEpcVu
5ufth5QwcYNg3HuviOrZ18s7SoZIceEhIB84uvYox6zsMBTMKpnqlhouNcYIgMD+
gV34j2AhETL9YhkaH6M3HRSI622UmaSeDfjGalYZb4QTWsK7mZHc2aTWIZm6Cmrp
YgDqCfqcAy09UmnrMhV9UEygDybVfEA12b+4eXTWADPuZ0Cn12P9QeZRTMaTbYP+
/mbqsB8aJ/oQsbzp6d8twmfZLgOtXwPDowjjyscmqcV7U5P5h/imKtkJ42YgUBuE
0EAHhypWKR1hAnyj3mUdOAIAV15PCa/esDPKwGcpXCfhctrEQB/vasswzJQT1h7t
FPL60V9IQCPTCAFIiEI5rqv4tBRfG+SYdeZSCZzMVjAw7r4rut9Az3eyDoqOPu91
MMq2vn5Z6aUz4sT+1l1MlNSjRh9WjCpa9lYJDnU8ILD+Bxf2NFPYZdFfsMtbf2f5
MCmJ/CpYqIKFJUc04Na3890l81DyAejm3ayqv8q06bHjz6DGERdZIRjKCB67mzJP
IaDjOdmRTRv9AVRgPjfbBjtjcxuyzl6hudJtbEfyaiaGK2wUxXS61lI1xiUU5Zia
AYdkh1o40YkCVvaVDoGx1yL9hc4lVLMftML5IDw4IlxfYi01Csgt5wkQMULYrw9g
rIzWlAzSlGwRj/7bnjc7xD1Ga6w3XvG6DM9yb8LEdQjuaeAaY4oW8pdlf6LfqHac
x3c3V6yOcr1aWf93YC5Vs8FDIRLQKF/UQsA7KgKs43iINbEG4Bhqg3Nz4g4BXN8l
vieoIY1WQ/QR5VOuzgqvCwPmeWEXaXk8ZQvWjb8P/gFEpueddBX5WHwORDUuOiBb
yXGPAQ3HYff1D0fR6yY1NJuL8rh5ZQGLPFZI79Px5FGsC23B8lBSQD3Vz8Y36Q9E
zXuO904g7Ex3qHoeGRw9lTTp7bGYJDmnQyuRAovAyhgVDkFqnNBQn+D2+QeaSw8z
Cv7+nN9rPMVsEeyNU3tYBASXHv0W+Z9BWgc3zXyigyDu70Fmm2kNhmSSE24f9uUm
o9G4qHnFpYP9FA4qxvnmsw4dhmlhmdzilPOHRmB4bgTPfa1eqDmctTDN+Yu6DYYh
4Jwh5/C8VqyrNsfL1CtTyU3YnkMbC9/DLZdMpq42zWHihQ/t3FLdvcQvzSA6Jk7u
/efFu8rDaWItBvFIantftG5VyO4IVwyRRcB4i4LOHJHL3SHM+qsSTs1l8VpCgqtC
mBBwjd8VISmKYWMlTQCP8Zf7g5Ot3Yyjyzv1VVm3P+nr0Dg9dILXCJw1mdp2IfFF
eY55c97coSb722WCgmn9h/yg5xFBPAPF/suChvEx9FT4AT7ybdYQ8KewHFGvsUSI
x/flODullV6833ue2JcKOArBFYNsZeN7w7ubFpHHrf6JyVYko5S0QD+iINP16TLW
igWQ1O+CkplrHVQwkI1pfUkX/JE+YFYk4dO/vXMza26A++Q86evKe16sxQgHGFKe
YtoI1W66A6Mh21ESNZ/gYn40AcbbUaItfo+9U/zy8LFQ28c1Spu3S2PdhYKwUkYS
HjAml89yJsuKiIlbmwK1ma9guxtNXazumjyI6jZgWllF5103JTGoVkwWn8e2h/tW
6mH02YApQfR8GvUN5i2XSIK/Bb46pDp+QD6UNfyHPmT5Ok6t4Ar249kPPnrjeJLu
euE+0ANjLaFMwF2TcjmknA4RZMCYs5ixE5I5K7M01U42Ju/EDzWvH4gVFC3Qis1A
diLe2wgJUmRTCE6ysJp2UFXovPlvD8yWWcIPnIvotSLErr3XVYcd6hXhrRr9OWqn
EUf/heQ7g0uV+ZpmtDiuIwqFZ3oJ+5GEBD4muddDK5un3gmMDYIC/XZkxyIBjRp9
xzhAEBNd+HtNUEvaPOCs6K5NxTa9nDD5pBvTWM58M4VKxx6NtBqU9mRXWv81wP5r
2hHPENRW2SJ4XKDOqZg7Vu8hFPBeL8oVkW+Imm+R1DNMAHpVbSJVW7SW5s5b6lOY
3utucSJge7xIX8esjvxGsELekxA//YTec6f6AIdtwv1nGI4j343eLIdZsqjbh/L4
mg05PiADiOcZ0H++24cIQ47Fwp7izdihR4ckO5yS5SoLLDpFICa2AunHfH4eUgSw
QIezg5IaUXAq6eVz5j2ELbXjR5GmavC8r/b9El5CpUQwOaky0M1XACebcfxy5w9z
WiShdBXh9spwnJWz4aOv7MAfMyXHMzEPpE9X1Xwvh4XI2SJ7lEfsf2PN7GGqMMLT
yUp9NgAMnsdUUAfRzTWmnJ8G7bM+QfqSIGZkEMz3YoBB9AbVgkMEFw+7tWREPVbg
sQclb1iX/ezQL74BBqW7xM5sKVWwe4STP4Ot9h9pNIhljLGystbIvxqnrJCEavxF
mDU3gIuF8gf6B4Cijj3AJ66+m05c0N85VdGgpqnRJXN1JvMcY803epEfXonU5lGL
Gw41U/WZOHs8Udzy8ezebmXJ/FXPofWvs7ImgurYiGUVbaGvQe6XDDBUMhQgt/Jb
g5iKKs090/gv38C+TDj8Cvt4v+CT80WqHLxRYgBSxks=
`protect END_PROTECTED
