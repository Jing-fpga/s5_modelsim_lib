`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vXAMcRlSqQ5YBvslO85bMuYqhst8WHsFYgDuNA4VXLEkgr/8WpVuaVlH0RdyQerT
lfEHQvqX/6Gy+aKAfWjew7vbeqMP9Eac3M7qkQJix2XN9G1BkSyuPOzsyMd6x2e6
rHYnsCUynVFNXmrdon3WTC7PqHX+kjLPWecZs0qhnVXRQv5DMeVUeldpscrgHgBw
o4GKgJqjU4K6HRNfczjE0Yyif40n6fUF9wT1BHirdPdpf2cItgoL+jbiw64XVt72
8Mvfr43FNvFrSGV726UTu3MUq2H29zX+7SM4+8zlpPVpLdB5KzZWpEYqXbXQtR3p
/CcxrNEUeLaZiyP5nN5JreMbHO928bfxRGs9AuO0D/M3UbfUUHDVtpNoRgwK84/3
Ck3JXeh82GXKa+GJIBl2RrxVcaFhEpoXh4a3y1U03mj582FSq2G+KBXNj0Lou0tw
ysj4UM5eepqdps7oAUDNlbvKykGQhgrU9adZgAkFGRbLN3spGacPOVXUFHV4e8S/
Ogjb1MeDeObWYr+S2ygK3QPULdDCzRnl6QCMwyhme+3nRdNSlO0jHy17x9kjwJQW
nZ3ON9lqtC7a0ic8jgRv1TNnQ10nhiPjLyn2wq7Ba9ycjrU+zHSM3+BmAOPtlSoV
unwejg2i4rpvEaCelwEvUCkEZ7bzEXzGCHJHSAjxZWx+rMQHSotVOmOyLuLz7d3r
/i46Hte3w9YOvFFOys0zxsXdwxlRrJjCBuv5e3MxDffkttIr+EzQWXzInFGnQX5e
QpZIsT/HBNLNiP3Q03V7cIGyawiEe4Y2sjJT8z3hd3TyZtp3MBxs4PILlHm/zMk/
65Fe29VuT+obiyBP1ndRalpvFA6QhDhd7MbMT4NbVKppaxA0uoV1GXRf+n+T+KVr
KwLIH3F6vlBGZMAhi/h3+62MXcfzAVeLCZvg3BBNMRl17TRb2FY2ULsc4G334FxB
JKRU7zQbpKUp2dRy+vxbxOsEpS44sJImsQrMzvA4EHxEuoe4rxD3JvHYsAHqww1K
wWrT2JDN2EwW29bklHlaSCWxtY26Na6Kq6ciiGT7LiLe5HkvV67J86IeZkuhSdFC
bg4svfhKS6DQ1rN5f+cK9Kz1+4mrrwrWf7sV8Pk2U818gFOobk5AHOLss09hwamZ
vn2cy/+WzbrGWk1jLaeKk+rWHDFbKJx58h5lSCONSpjKz7lpnBBPAW9I40reWaKZ
MHrOybvAH3LRLIDR7gXKaTwMMA6+yE1UBvSrOscUsMWFfXHy80qu7gtrnjlKhXAu
603Frj0x9v3ZEraoruwJ2eba/Rp9YLEHCa9INHMNom7/q4OjH5ZdHqzo77c5Pejl
xOgJgkv9UnZI2OtehxDhoCm40XNJrgV5nwqfuWxFmm/ne0StGYmrcRyz/W/GsUe3
A81cKQbIT09Xd1BXYO4m2lxBtaHnubCmOUK/EeGHXyY=
`protect END_PROTECTED
