`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HLtyQm9xhyGp20Ua4qIGf+sEJlhAFA6yW6oZmiYU13ZqPDLx/s710xEVO/J+Qn/j
Rn/Y4p2lZyZFyaksfyNKr/w98XZT9KkaWkCoUMkocmLCqzi3PS67wsnbYDRfwdsy
Od9yOz0lI4vhFAghDG8vruhGhGwuGKfmjeK7a5Vj7FdEOI6bUWC6E98X167WYipx
bBn8SxQy94vcl7wNNvFWIbeUwNwOqt4db05i6xIQNO9zyWFmbHdoVkAsSs0ay24L
RtdKCsiTwD+7ymtcrkad7guDLxfn/dj6nt/Iybw54m/7X2DvcuFRwRqgxnNbCriD
4YnL4Eh3D0pt58zr9V7JuAXyajBNj3yjc6bl7zOmOU/+jthtCNCNImX0CyVRGhW4
B1mV3KU+vyvcRxoljJCM2q4iS20Gslj3Ey3hkYrFmNNcoXfquQiTg1DkFNj9f+aH
6u42gOEGEdU7Jxa0jV66vSKVJ6hGbH7JIu1sCe0QBdNZDON3881omfJrhlUAU8Kd
SXfQEK5vLBNF4fTCNZ9DZHiCh0BT+vbePpAJE5ih1e6OWlnHZXZJP/q1zJFcEdDy
RVm0dO2c8MBX1f5m5VrOTP+eCid/9ANzVVIEo2Sjj9tJe1FdWo953rHXZPbzB7f1
R2vFlZLiWahaRuOMRraIMQJRlcgdid/2PpmEab6ZPkcP/E/aqug4srF4l9b9XazS
EANrA0NJMmBWDEactquT+bTlDOQ3PI3N6EdJrURX8EKX0Py+s8hx+d/L5RPWxu87
w82aIBlOLqQhBG649LUoQEOv9trWr62KTCz3tq6sE97XtSzx50Qst1dbOkebPSeA
AGVAUACvx3UZ86W+jma3atJzplcNC2fnDwhrNNFwifZ8oiPxxL7v6D8GIJOBfk9I
gABKe/3IW2sMCuCMfKegwq6qWcmogXtd3MFiEVLWKQ5/ubSXhHV1GFCmjAO2a6+t
dnnVhdFulaxQH/re8rC/fszW+3IcEiD4sIW68XVRpNf6rxS8Jg7dcBxgfrhNyUHt
fgnAjavkFXJ8f0ER3DXuraLjJhnpzBJGp+hnIFjndrerkV/6G2BzjuLG23n3hvbV
1VRG00q4VOOQ4QeT4Do1aCv3ZmmFtDTnN5bCVXsMuLUErrRRlultFjyUNbaihez1
PwBlvZldz4B0qYDV0FqYhXzIXPxslFw6IG5ZT4ddUsuI9Ds+NH3fbizi5yLnEBS+
5xQPPk+FrZUQj53u1GW5Hid483uw1rnB35BUCu06lR2/RNnNfmDTbkVAgS7bFbJR
CNyuCCx9+wQ/phnrNC8i9M9Nvbe25RoYAf1jdMfTTCLBe3QlUKjH6RzldD6LHiTP
mA+wzP3kzUGAtEYAOJdtoicc+odVQ6Ai5CvYZqsNaiB2pGRprMMvfnGSqtub5G8J
vQ//Ruqjf2YQTBjbHyCObqCWrXwBRwuTTlXa3h4hb2Yjji9xveMj135SEG4hiHNA
UEr7aFYZcjucgCYRCQKRLKcQEIzKTmFjFCvY2MtZ+9hrduobX3uv/5U2sQ3ZMI6c
Wa8rCr8z/wafspGlfZg/vm/H2WMG5SF2rFCA3bBW4Q0IySs3z0H5inEqdI7d05Jr
XJ3QWMPUW2LTbLRADYYWTEcUfzwFHgP4Cxeo/MZrl9ItwihcAfr+imcPpMxi/Fwm
oUDzyhG2H/qV6ssu23KGQJK/lEv8zgwji5f/G0rOspDjFaJuR6+VwgqwoxnPxilB
wtc2oc2aSULOY2/pa8wc3ygQ1vdIqzv6H++zT3oHv8TH3vNhgleunD5Lw6i66u6l
zuOjIpRZQifvZDles5SKiQ35U04NBScaeG4i75ny/DvLIn4npY+VUEja+EGCLewj
xz09pVy1gUPRwlL/NISmG4IzA/zL8WClIpAidoJznK94f18siCmgDkFTxVfmKKqC
guaYvygla4bpGPr+EREb1Uj/QtCtRJwJp/q6YOL8zRCdOwSHAPkQW6N4uhoORIMz
8SOLvu6yICpvsTJlNNvI/Wfgj65GQEWX4wPww2mE/kWxKcCXmWkmMx9BxjuRsqvt
s3kt+5A45RDihHX4l9fJPKT8OvfQ+KiP3VYh7xpaDNi+l0KrowEFy/poALCOJOSe
lzI6RgbTLvrrDC4ekABQKz9s5ib/rlCrDwKlI2P0o92CoUt70w7bpx5UknPYWNhf
u5ok16GP6ExKTBvLoNBmZD/lZNTXFVAfM4lCvl5eIVrCago/FmWnmC9KxzJJlLF8
OoM09UQYUhAmQQroFpIJ13Uhl+H/IJpT3iJoWi1LJ1MKZicM7RmAcih1quAcRzGH
VUhZn5oSqwDjiTHG7wDSfNgjOCVOFuiCikAFuE9NDCDL/pGPco3/2K3I2A3OrEpV
j/Eao6FYzu9XGpMr2Kl5LQ8b7X211pW+QzIHaEw8AEl/2ufksolE7f+iAZDTIoR2
GvG+TzdycDpjaSNzTx87rgYqOfWpOVwh1xyk+RqmOahxlUotrl00CI0Qp5S7OY/1
UOdEnRywu76ejhYmLHeU0DrumP4VIWsgZXTROj3DKcfjC+duMgRzqYgOp23pMzMt
rBMxwRhRasWGpQ3Jll9KkE4URDZgvdJ6N8ZILcFYglEA0EQTIue8fhjD+CQ6zR/P
Uoy5q+AonbEDrcuwIZPf34bcuYOzUp2PQ/QTs/FD1/Xo+xml3MTlcitD1JYKDqUl
M3snZjYSx6Ou5QYZWwNw9xCdsZkfiW00CZy5uWIPK5lOdf8iX5j3vhLmMVDAN8SZ
zLb/mahDAIqlIbcLm/HXUH1RLPtml5u5rkw9fkgEUPBrFAroltYvna14tgxkQ5Bc
6Ii/xxLYBJ+4uPlmBjF98CPdoYltRYy72jB9O6U6ue8RgZiJ6ZOVpZ8ZVzo5JaWB
K4oijUPq6gPf1CU9z171MT+9mHLuU4Zy9HfnRH26zqTKMDdvHGn1PzTaxGuW04vR
8e456uu/BkVB8OqYBd47AiqzrE0HnAWiQWqNtTEVVBLJsdhRI2HsRTqaJLY5dR0x
pZviXf/bXWnBJ9Afc82tOvH2tczKOFLKsCy/BVVyr34LMYFJUDmK/s3Ewya8Lk83
hPbsajCQuvmwa2aKsXaIOZ3DTfSsyvvyJMZzFY5RFEVOkA1SZDMWaI2qdppoO0OM
el048W7WtpvOOOBdEvLfVHbMJqJ9sksk8wRjU6m0H3Qfy9QmIEkMv2MTLCVNYMeC
RhpaCDhlDu2hF6MYlfvesArU0Xkzp4USLCTsa5PhvXaSpwURPuwtzEZo2xdLuGV/
5ENNWuPfWCc1xpA6ahKX/leubLbmzcemgyQe6PbEq0BF2qnw1Kwu/+Sm1USfB6ci
h2IvC+EmOC848suhT+CJW2Pr4347QsKbuDd4Ie5y5pZWNuyqN3viDGudXdW8LkSs
3q7zAjcba5JnfABwINuns3Ha9ja8g5yPPmWPS/XwaB7+CXF1n2aYcOILj9qlrXtK
UmQetC/bc+7jeZqm/mt9/+0TC0U8jtBSDzTUbqBskmMf/Td4hUtseUB9HkypuIgM
+DKQdpALzG0D3O/zkCTGrASWy50V0ozbNJYV3cIyAjhFVEaUEk97A7AWbz9d2QIV
6W3ApWQltft+IUff9I58Qa3XX7FCR8VUMNL010a0WJA9+rUb+CiDF3li+tk/1hpn
w9QDnboUw8ZBRCD0KzUvKxYQnGvFhrVN3FVDEHk7vsuamxcDBF6hcmbhJsdoIvFL
BxNZBHbEUOmvZhLqTpeJQNI/61Ckk/GU2nNzJGjgnm8A/D5RyLH4yzJ606X7unH5
56kfjhc8woJgPYEV/ZyI7uGHEw9zejlCtVRQPflwui/lntTQVIm9bQDsFhwm00YZ
6I7r15wBfrMuLuHJjKtUJ9KiEHnFUkXYKC6mqB8h+DXLoacQvju0sUX6I35nGV58
Wc53wJ3wvfJfln8iKegAXi0FFuoWZ8WL4ByZRiTVtzhyUhHKGM64ZIktU1xLfCa4
mD8vAEPOQuBiuLcl3ubAU1KewkeexISwFpZ0Qyvi3gwsEbRTC2r1v/KezQ12oStu
F8hUUaP8dsvHVRXEAJecEsx3AihGtsyrOYjYWZ3bU+DuUi/JbFVV4ykJwSXic13n
WZraxmn0zY3qnHl+gHzKtE0goi2zSGoRHBS14zJW1cTeicZ3O+A+fJQQ4Q322nsH
lkXquUQbRuNvJoq9afTwzoFCBpTQ1V0iR8jQYws2zGAbFCUmhoVd/qMFZ2wLBsef
j3lSdRbhxZciqqrMuBqvh8V6wKloqj93js8xjU8Ke/TGqCpbNCNEEoyFTxaaK1Fm
Xa5rgvy9xCoQ6phs+9N5K2G/ST36S7jD4HDQ+2q59uPaAaqwLBMPZLnl7OEJmHmd
pnbeuoTao5yrydD46e49VfIjqN3ESQNeO2iYCyCJKKFlsgSBXNgWEA7mMC7flZ//
kF3GxNbhFam6PbjufbEKXfMy5/KX985vEpv1AGi5IhmM3nyii9MXXQ0gSr/zXPLt
1d3J208eJMMCloic1k6lV+lEpkoAdLXXZTd42aSa/AoRNpzTcnHBnJpeg0n/GBAz
z8/lq8Rphz6DtoaLeHD5MoixKqSlv7INxnSZl/taNKbTIzHLyu2bTDf6C/0x4ZJ7
kglu8ICxtf8cGGsJ1YGmt1rC8/NBNw7bpHxrtUfOoWVI0cqETL3wTsY1AoA2RJV+
Ui9aGaBMz+hIQzJvhCKEAgM1wTs4BhW6RiEyic2h5YtptzbxnlAQ6ZwAQYeTkgwv
8r1UaqECX2yR9d4Dd5q72eoA38uwKjnsokE6r0iGtk+t1L0caZLcVyOztIUrCV+D
EZJq3ZKwUAKmZAoA3X8GxaCGExC1sKaxTmKg0esX//TV9J4BLdg6omnQqcPUHmeu
GYbQ0lQvhHqLk5d97iUpZBCCB0q3MIV5SclICsuZk6jSA7mRW+sr1moOR9KGcCTP
d37cxORTP3FO8f7O8tF5pxQ0Xd4jAuNwhRxDOHDokAxCt0MYgq3RooJczJI7coLM
o5K58GFR44rN9nFbkXuwGH0nqLho0gD5qKaTN4kv0eHbyHI+7fN/Cx5t9t4klOtj
o9GBFOyhCNYJYkagGDiDysMHn/efbpsO94S/4x4/7jg6bsmMZzn1KitA7ZPb5IZF
IQitmCn/oxklfhnNmIps+17xOeCsf9tGV656jNBzkSmUPZVhJYiipKNB1JK4EbG3
G6LIkGx4yilSJKvy/v4rOqvIk7fTY1CgAzFykl7y45lLsR390CfsZtVsDSl5AMN9
IjOnLt6c1Q9IFYuIy1MGcXA5a7crTOudYd8DAB1K3ydYG8fJh4AWtsAlas8cw3R9
U4i4acTNerO7DNOCe+M9+CXlm8//UR2yiV53jcJlt7l/urH3CTt5ADJMRVMkykoQ
/e3VYp6iKsd01aV1xRBEI57xpIeNq1wAuKP7WNg7WRoAl0pyHxT12/ndiTQH5gRS
2hV7CaR8tP0Ob4ahlS09WtV1NC7OvQMUTTVLBDHOn2GFBFyggnuOy+8tyWjoyP2g
K0OS5PzWcZqpmwHywKdqHDqGOOuR5dWhd6XYxkKlVIA6rGj94qFdySS+ZaLjtrzS
4l+BX5deYdjx12F9rHgeYidqZPUAXyLSKB+HuLSwHnjsEVJ4OaNXGgnGQfYKQCrG
FTuTfltbBcnMg6w15EAhdLrjPk376L5xBhLRdUNflHpZ9l2rtklYqxfGIqWbHvlW
HAAMpFHIzOdn4OXI79sTECsC/TfiKm9lsK/Mh54pAvHvFV4+xU7m+e16pIy9V3A1
wd07bozzaw0Fs96tGNn+PIXYxRScHJAb4jNbex5fm3bV1xW1mFsXI6rTEihCfEfk
NQk00bpZ3J51FqKXYBG9ru2DDAyxria+kS/jSN4FPRcFT9PfryyUxGBlpEKL1qTv
yVa7aBMf5Cc5JabVJXa+TFslMUfw6izlrTOP86g7g+crcWkdQ/G8SztsBzHD+ta/
1mjR4kTHCXK351567nx7IQIVM3ADN2PpjyAwxOy0Be6xbSL4RtH3kYwGassmEan+
NTMbna+emzPcVHXQ3Yy7MHHLJt8RLtVtRnrAQL9fPmDn3NzZdGJaPcAPy+xF/uu5
/35If7Go8g+5HYvPedCF0R2VRvfRaSX6kvIEO7JgTc3lB0q4TyVQJXu+Yqtf5STg
FOwSFJgYiN5FetwwQnvTkMxGr6tbwtol104Av0TMGz1NIVxd18TbDP/rzZTViq9/
8n8BUk1zKixTBFDHkYgmRTwpeVJtVCMU/wg9fmsduljuq829nOxAmcFLKj82vhfM
XaFEKkb9x+BW+UGqUNoaH+6IDLtyywkyjcnc6OvF8sP5vTTUfmsXWWFrx9pPf4NU
PDrLXS4lGYCDJ8WO1N+4ibLJlq3kMUYb+M0v+N4tw+TXBgMjgm2TsEXTjF5YNX4K
WsZf8bmWz6zZyHIezolf8F+3POyy1Rn1M7dE5Kw8VY9xGxCoBGwWa4yBqUaYqleS
eojR8wXzytAwBrGBDZw5UxjdE1AFM8yG0U7DKq3TkjPiQHDYXsw70HR6EnjAfUzQ
hMF4xtUWYiW8p8v7PZlyShUgQpeFksa5fku7NZEwTDfiyh+bqFeCwwNohYApuGn6
XqPXSNpCjUnX/W0PhYNi1s3xeVXYej5NMGO+5tEDtAL/Ui6QKfXjv415rz2mJ+ib
PcdzcmqAFE9TZWN5F3ddBeaibH4hI7GxOltd9xhnPkxxzKqNiNsGMUwm2Bk44wDw
MigEoWGv0+IA6igR4ByUzus4xhjb84dGJDDvEsUKqbX4kjBK1wYN7WQcIXPrMpNZ
YiFfzvhjoGSUhuQeS0B2IsXnlkr/yyor1Lsle668N3ewfkoFiusnmoftvuv2TKti
vXtqYs1J/RdHm/gaHmdXQ6pooPqgYy3wj5zNBnG0RvMb3ZcnMouv0BWDle6QI0Ga
dLlbWGB8DOfxUWvCpZlM2/nM/3bQDyOdZsz5KJdxkRUnpAXfocABTWiMjhIkaEF8
SK8H33JOUzwsnvNlqfRc/7fWKea9UprIB8JAH32/FrNUI9SRPy0ZNnzCLHxd9smR
buaovjx/1RhUaAAu5DKhSNsQpV0l3lIsxhIttPC6OwahA68LZsKORVsqXXP03A+l
zHrSaiMhC+tvd6j4bJ2t2j920fT6a9TGx5IUvJSG1401jh5XCosQqkuNlcD6KsZ9
nu5B5qSc9CELWBFiwwDF9UKld6MLcSwmHcNw+78Srom8QH63NMa43DR1kQI5Qezm
Swpcmn+ygZsHv8onVtadLJfvjCirq/noo0myXu2FTimQT3AYmHP1x14cZ8YCxf3z
x6B3I7HRNmwT43uzm0z4BOSaUAKS+BzIoR/O+trSdYaIYNSF2/03Gx12UcI5fwAZ
AdKSMVjH6S8yzrQ9a4izF6L9QPAFLwO2mrCbCjJR/qlhRjRJyKG73BvCeShQzvrL
vvCRMPd3+xPT5OrC4BZaUe7JWGKWT9MCaG1EJveede7lMr7G5IE5HouIqxfYZON1
E1i0I3abQIgSabEoQKVPb6cpT+p2riiKDtIHBOVfgsrvVHnjIb2uWfN2iFdawM9Z
yHCbJYPqkpELBl3VvR034INS5DE9vZfVdQ/O4WVqiwLvnUULdi+q5weceaodIiIy
qyoLt938fPw+8srK2+3GBAMhH8Sfkcg2teQrejwcRpc9V3RX6ZnBBBgCWdHHdh9G
PRIp1Ige6URaux+Y9nbqQBY3mGTp2cW3/IyF+7V4t0bVMkBzc5BzhiCDU2Pkj8J+
f2R2GffIKiXGp0NVfenoOPFwztZaA4d/kXNQnijbumhhb4nV5VH3UN3BBCqbhhSQ
7AtgWc0YqQj20IU0Sf0MsGvSECclqo569i2KMOhP/fY0RRtvf9+AUIjdB9DnORGD
6IG6UdhxHWR6R5SQ1f0rFEvmkxs2h1FF8x8tBzSl9+3JvmQrRKESblWjzIkILZsW
GLnBf48eEvjL4r1fmyxWzOQgeCgWkPmX878ndUT/iPFp2EzTBTMVUGBjj3Di35uc
UCVWI0I7RPNfhrjj83R7h+WSEvV4i877wDZjOuvUkDhoU+tUfLe7XaL+XrTmjK64
yIXv2tSBBNk2/7Mq9LtTQXoO9MmZkNyW+CvLr+SXEF/pE+6DOXZqopTJoLhk/sWW
Q5djZDBnHqrxvr/YFW3fzR+OSBwDpULct5//WObe463vrzCdLJs3klT/eCobYvD/
bF2vb6aE1HR8ekLxmZoG5Rp135suT8DERo4otXRAn2AobPPdPfMPp6kX/4P93q6T
fHuogCSGqqA6LixU8PJ2li3CHo1jScEwNj8BCqPRyFlN/9YHdAa6CTU3QJAJGjbC
6N5EOG6nuaJIfkMgSceHbYtnEcBplGp+T3OuvS7d0wiiDMVRlt/G1/Sg5Z0IuMRZ
6LYLtukkBSlMvdx2g7gYGFYEEqiCDgG1lXKkBtKdGmdvLHqlq/89aJC38Z44vGnn
Mi3vLhJLSTClJRfoz4no1+fpbtNu3nH7X3ZOEmSPVgLbJSNJUfwXuo/o0dFTwOsh
d8Qv73UHdeLKv4jvG5OFiYTLLGBU2kbJUpR/xX+nlZPiWVL2N5+viXdAni5hS/oO
NiUPjiDm+AqPF/7ISdAzZJFiXwqx9kwlqJJQrLtFlx6D14brokPhCaH9ii9KGuT/
7ss81CJK4UytCiIaBHjy1DdJKkXKRgQICa/697r1XNEmqp2I3daa1HK6b/2d50QK
J3Z9m1J8o1k9HBHtCUfZFEBNxV3mXqN3C7vl30N6WKQbfRVDlZhSwtEKzBhzgsQh
Mx9Ka23mNg5wONyG1Kd5KpsQtsbNCi5ATk8FT8lY7WorNja4oxhDk6Jl48lL9JbD
3/wTfaRkL9fkVJHG3eXJUxLXp1ltqxx+TFpdZYM0M1ZA9c4tvBJ0uRCkySPfeFO8
cnvJ5ydwjDUZLybCFb1P8OOWGA8rZvhpotzWWt08ETfOshEwqBA10Ff6C5NILRaM
EH2PLoJllBGp2K22HNMR3MSjiqHQoTCqMYa3mJQT/wttAwakc6Lo7R2slvNzOCOf
9vfXKHZMoq3KdFhbssc3WYc00yP3/4fBc+PljhDI6gV+ugqgQ4NqzUp8RILJ0Pv4
4hUhpcjHtnC+p9nSoeoDZDxDPyP00tQWbVrXptsZb//xkl0Q2m0AAxrhlNVPgvMB
QK/1KwnxSX4SoxAMGe4/ZrVBlUKuA4Z0Xim2YWJf3lmnX18mkiY/JFeHD7DUt6EJ
TJBhks2BltfAXCnCLwvq2TLHRv97YsyGR/FYVRMV/ssfSCSdOSi8Nrkrg5J+cDFY
bdEzZhKJO9YAtZRSgCvK/r4zJVl4odC++IxlYcFfp4218z5Cz2wQxkg0yUFnuwo0
ANFhVUS8LaM6CmPHMDQ2nnJLUoxd2tDlpftXcjD82lpbYnvh7SrQkMsAcH9ThYVG
qKXCTrzjponCLGEa/zTnd/YSlTHJIrScU1OApTV+I1bDuEoorzeivnNbL4re0kRj
SSSjVfsdugsDqMZDH71DIzYvZ1N4hxFnBTLIvDhnVQzS/CinuvXRseSmGGorYiaO
HgzWGo0vzoJhnKPusc5PFIRXTaQAM0n2MQTew964NiTczQ7jucymEpSSmg7RtpVc
OM2pIIbvMCa4oGgISTS51wGbJLcP4X3lEYr2Z3fzNVpR41I9djROWCZ2nt5/8sus
Up8dM49DVB/h+8sMKCRMfRGXZ3v+xy/Er7OyNA/kW5p7CSvKvFKtNwRxgEFryW5k
J6UL3dKQnqD73haAKY9QvNzyh5nLme6VnUg7ZyrfX+cGRovX5YI9k4OjkXxOByBw
RCIkK9wz2z8/fhtCVxnbV27rp6Qj2jNo/+wcPNV5aYfQS9/zz8LzVb6SaOqwLUt9
+dx45iVwkFXalf2oDTVVlVlU14czDWVBc0iacn4kQRKBpehOwOw4grv4GyVbEEjN
4IPmHvgkq6adHQhNu/z6SLAId3sSgEyF6pNPgOondFHG6/x5ujPzMWT/gKMK7izG
feIEOOdBhk4i20Qv7jBsIvmT25A9SLzets5h2FNgSEtNB7FfJ3gqjFFdAvzeJdFN
JvfaXk705sCMal0Vi/4fDhAZ/tapodxlriacicsdXPEXhNRJriCg1MdgKZ8TgTlT
L4tfay63wsGavt1gGxnp//kAu+67JWmVdRK12JcMUhh1mgkYJ0BiXTEKdxaDXElT
0SNVrpWRMEbFFdHJ3j7f/6FFw3TePRaIixAG+viQSdSG3Kk+p4eClR/X+YMr24uJ
+EFveB0Znm0ryWW1j2ApPFVX1DjBVVCEnz+QulmbIFlRMkTSvZmH0W9/AYoDArGt
pvB413nw+g+X3GUb7i8Y6vfkRNa9Did/9UUtKL88TLNoi/FCKgbJvey6J4+KtZ7p
+YRD3B7DOJ9bWQgeEAljraR07VUuZUVmnzyLIEAH5BassNdocDLNLLDYphoDk4FL
huJwdyO8icwy3Avy6jZh+cRGiBwIDxxC2ED7wybAIlzmls3MzFzMHYXHfO3EnW4T
CezYamPuwjOdpS/bMg2QSgXnahq6FAv9nbG8K8vNbJLFStc/tllMiyZ/J7PjXC+R
GCUxl8RmCthFELO5pFSaBzIS8xxnONRb5MVfAp72BBMxxwMx0ojFb/FzVHnTrnhm
5oT/I/x41IoUMlNpJlZBSbF4NE6Cl9zPkVu82AWKLKI8gWc9WsQFOXxnDjvCvAyJ
l+YK7ePBAjq4CmM/FrV5cO42t+GVYpqp4aNdqAEnufzhoYEYgK5GnOWvGzLIj1Ra
rE/Hw7+cx4/NcqWz0moaHio0WWcjGVetNPBe9If1DhrPwU3pLigPBVKEdRmgX5+d
XmZfpOY/JwrF0npu5QC/8n6IR3RqMWOfKuJNbs2O0lTIkX99i2KZT+xL8jIxNCZk
scHnqcbYfSwR/+oF+EIKXLHnG6/PMIIQu7erJC39phAUmYj66A3dm50pSoAFxjVI
MarHH0X9sCWIUafRQCWxTGpDq6o5Vo1EYDJmtFHSqSiYpQ7UNMksLaE/TglY6+56
5BEiAjFyh1E5c+LL9hWW5bJOdRe870yW7F0NdKpdI7kCqJD8w/cR2ma+M+tTZZsJ
o/iewGnzOTH9UPybchd4xwzcEN4tBzgYkpjsDdwqSyJk667bW23VLX3Nn1TLrC2H
O2zl5R/17Lg0BD+CTOXTMn4C9MXIyLVNNSRisL5Q/XjZTmJq2zduI99+KsJWyz5d
mb2uDBpCQ3zQ4GB0RMzOVPmX6FB+hb87Goxw5c9GrnMs5j3dQnTl5X6ROZU4N5/o
VMidml3KYGUjuZP9aI5Vp/2d2+A3crK6bSYvV2MnGCxq9FJG2CiAnn6VFp/FMBk0
flpyJHbVQMF5QMZQV0+z/Qe8gjC9Pvb5mCPKNDE3yfQzluvf6oj883BEhTEMOPPz
l85kTM0G3rl7/Uq4av4DYG8AaBDTO4HFMAp9rlTpgijR7rg40nMJn+wqGxLniKJ/
rBR4vrAeBaNv7KXxnwx4wEsKH34g+YOY0H29pDlVax9TDpnEpcggH6n3olsrO9m0
BjEnvshklttVEYPE/wpjFI0Z7xTAIl2yQMGLkZkR2DGMma2JnEfpWbQBPUI7ePmq
A3ppwhquQDm5e7XyVHA0k2irH6L+qtgfGNk2t8sFemVoJPQOYaYU5Ygfckht48qD
qEGzTDR6rOIUpcs5b68vWbsV4Zvhy6jwKLFm2moxDrjgM00CksX6nH8Ar2mF0JZ+
PLNCn8zb39o1UJk1KeWW/AM+80xGjWDzBDEoSGqJHaCE8DY6DZ72QUiEaXCdI16a
cuQZY1aQKamUvLc5HGnqP7MpHhkva7SfreUF2EcudUHSmhDCY77ZznCcpKUSruu/
UjYW5M/PEgUrJhfaBObGPcXSBBBwrCGYChdqP3otVfoMyW2qnsA4xgO/O6A54OmV
8CUUGiDJlDwF8uqAEWtngbQHtT8hRVofbhSNvEHEO/VIKEOB0q7Y/+y7+pH56WyV
2TJaJ3S3KCDB7SJFey7IZ5bIZSRrGb9GhtLIHkXyaS8qAi6B/PuDoJIeB/WmwN6X
aGdNqmfZQpqMbMmxVzBU4uYiQZoL9EFCP/2zac4kgxZBCH8EM6pt2dsQWfC5UcbJ
1ztWKh8w5tmmz/saA+r68/J0HfEJJT6uqpstyKr5CwPXQAv21TFR6dyxomlEYEfI
EroxRuBDfb76sddJqugDuSblSDE56kkQLF7wr+XpPVWlNSowjwEgb1q+id6ryd6c
A8VPt+Y1fenA3hu6ytl1/Kk1BJW6PxRT7+Bf23XiCwRbHN11wuDgKTKFUQD+k4sD
euE1s0xQvWUIf0DIt8ZgkAlbYXTH9U0b0EpV15ZtqN5D8yxF9ZulUn2wMKwImjYv
b684kFf9l1Bo6H1IFqo7dKx1+g35oCVaNIUE3ZSBilbiUUy3TWR7/tU05/iK/OxP
8d8fw4FoWYmMy++e1HwuGg3xKgjj2IdyBGvo45glnkHL3pbo6djEoAGLzafX6Wu1
C2AkSiSUcRYmg9GAWe0ILewWMlZvkz+uE41/cD0kYKjnZBKa+dxOndo0evrQhAZ8
AtIDcNfPFhPuqWXKP3GFRRpcHyMv4fcAWwJoSxLCVrKds65ed4z3kUrlXFXd6obL
BJww4Be1iMOEfNFaaO2q35WyV7TaCfy2Su1quzEuvWitVaPxOz3dFBpf/xEdUJDI
zObrhOijQ8nWlUbW42wSya+hwPvODIZweSIgFVANpPTFAVtRGVY+QH+mktmecL9A
1H++4TLvO0ELokSkCQnAAlFS/rNJAxfw8qx5lU0a7AE1VGQbJ4ZatcEwqgS32SWx
SJ5wOvHACpAwOY9MX5xIZwWvT+E7J3D6VbbiPuzBZCFDFxoorbPaxpasvTlgvTtg
FnOqSms5rJITWD6YKTKKeM++9IQpsBvW54ma5w1YZTl/OflLt4zP7ABGbey/CUcc
rh0jwvJVmLnc2Xt2nP9lMO2/SdamOlj7mzLA7g87wwr6AIo7DHkQw3QzPFhQ8uyh
cuvguEMe6DwkMCITsdtDeD/GDGFaaRUqwCZvizUZYBJPYHGMCFuTJgzVpHAg/0JU
b2dwUjsFqq36WCCiMJ7ROyTyLZDdJMc3terIy51g7oMJHlCVOZK7DAoPwdvjFCil
MYS1hf9BbpNjQIKnKCvdvgC4uT/NrxscuX1jMAKQYB14TxsvmHUwgcfRSgY27wEb
69P+VcqDsa+TUJOAVY3QhgsifsHAqCRRf9naADfG6IFGpwsIbCdJu2FIv5fiSG86
YR6yI1OyvOuqeaoX5du/5ymXCEFepQJQnPHkplJJPca991mhlH5GpyVd3Qr7rc/v
y4pjpvmvzjzKgNPMV9x/tJBU+9HWXmpHpMGXLmvTkrLpib5gQ58j9a44Sv+vc/5L
WWlbs1CInVaXQoExSahpwmBQMRqsLBO7KTaaD4g5KcWEiUQe4gRFI/Mi3cimhTrv
i+J1MtyrrTdWS0YSxv5tROvCq9hItkYoowREUI7BT8ylfbpXw089VDJKSHyfDea0
Znd1ioaW6AL7Mpq63ei/KJ7JtiBxl/jG8xCET5RuY3u3/rlBjSy9B2ZGqC9Ii5Ol
sr86VXb66pzqIuYXtVeVW97jJGxP+4SPfUmKZfVWyfZz+nQkgqZffrVkBm8BeqjY
F+446OZBfQNZ6nGGT6MrkgB4rAo3YVy8O+Sl368JxImsK0PmpW2fAhXFl/TubsHr
KzKCFK+2xbzw8Y08BuxsvGNFbLk5u/AuB81DeuPIte+xGWThCV0mQ729MHQQxOPI
M7GxiSPEjeK3UPfXprGFB5w6qh2RDt/1gJTVJm6qvmh6XfWD+uOc8Tc4ywsR5rGB
4ZiNcE2w4dCozw+I4/glN0/zL8r2kmsn9phz7PIcdL79wOiRxhS8EUn9s+mQWfBr
8TartavyeqVErkLz0+A72Ph3ajiM2hOUw0C//P1RfBh+58B4sSTAT+7S9HaVMPWs
eUQbimLUHTs4xHrhgFpf8hikMtzc190kuX9BvJX2fOea5dQYXgzvednb55pzeDeF
T+UQdEx72s2RnP3LhzvXnxzNd9L6WF+LJNW4BjwEbTh29kLHeGWto8Oua4M56sus
B06cY4305C6pj2zXMo1+FGS7qOL+gMi0cp+07Gv4W+sNqyejeq2rH14uboOCCAIv
3WhX2c/n3yKbHsbpGOtvBk4AVj9eCWWk6lcf4BmBIVOCSaqIHsrMy3MDtA46qBPR
ZHHa3EsWeIGwxoQEiyDVzeIsgzF//02ali20W8R0dPZj4K/qqzYftohk8ZzN77Sw
LZXjtde4HzoP1AEXYQ18O2dy4LWzxT8J9oheduKmvhTP5utGOj23QA+ye3+qQyEH
4TCVIC6eLRHyC+Bsj8RFdrb4KgHpqnReBKjTsqyGt93bCbrUSH7EuD0JBB+lhBVG
wWgE5jWgedVfG9FuvqglIar30pZEwvx2+V9S0T8Qhk4ZQcDlrpmyziiUC4j7qxd6
mwetG6km8IAjr2Igi9JLAZeAJv1XwGbmeGSZ6wZI9JM3jCjbqIuk0UVfwgPvEPbA
mD3itVnLmJBqVlbSji5QPZCiXvICnUzAZtyFnNqpLz7Xngae1nS2P2FGVBkRn/Ou
K9DkkwT7I3ws+IOjs7xNT0ZwciEBDXYoO4kpNcR90eMZ11vNP6odsaprMvfZv71C
CP6MYqZfWwEPfv2rj8eWHshEdh1wR1F2adt1lR/+Co7zmmrPlWhw0PZZKBnZK7qj
4eDPPI0CkEFb2elNbgq/mxS1yZbsb+1T5IOpEzlAKCsX2glt/UKgvU1Qr0VMOfWy
uZy4TOOPM6YjzCklh5zjhxzkEW8QbnTVVAcy5NH4yaybPZALDpFDNEkNRvziR+e8
u8OzR/fKP2I/d4Eh+0uadBG6rOzNQZokr/oxxdG4gWRLGDu5kEDmqEgXbSS/oqMZ
yK3eTjgJFC3egCKfCHJYZgLjV+CYFX0DemETen+iq6gtVqpsh6FQblzkajLW678e
bzn61JFIJtOROSZB9fzAhNsRU29jBhkjyNdJa6EHa7YbTVdMZSkvamQAgMCIuPSA
BIQCuRmFMFqS9sSfULA6YTOFrSiHVf+NB+aMvibkhS6KZb798dfYPs7WFtKDiaHf
rjFa+57+iuUQ7gsfQgoEyAjHvUs947S06Zmy/90JwAlfeOUjcKBjBE8XfhNufvlz
+9R9HaUo6yHCtbSouZqgvQgoZ+6xSwThvbjFkv+up4JQcdYoLGxE0ROZWTAmZmtd
2NmpgSO5/SOzioQANaGbkVR3Z3bQiIC1eHgq4NPSUKaakFdSIIpVtJz5Km9r+EBq
T5UT5dGcnSQ+Zkvus7R2JRwiFavueOYvJiHhgXltilRS2D783qMSbxgyl5RJhkB5
M9oXmwydJZeNdw65tvglQqsN43klDHnx76w+KlDtKeYQd5iQxwSnoyfEOTKJfxbB
3iFs9w/5Mq1iosyqBwrveGgJIDhCQ6a08j7igK54JPsH9T0zi7eaz/GsD2tQdOLi
YIhn2Jubk0hXoj2aqD0JboLCmusboP2yKREMV923UiBqP/r2rYc8IB6R2BZ6LNAI
SZxTj/zWgy+lGmrD8GInw+w5gamtkA0jynsXyHrI1DPHIlIcOubwuZv8duhfg3Mt
CGfyIiuhE8Yo9+aihNcpMICnHxQ0KgHecxB4lr/gK1/eAwD3VtgjkTuQ5PWC/Zw3
JF0lklkfADnFN9Tq9af1j35pCr42zTA6eiHfvdnxaQ8J5kzh9t7GI3HsFWUHIZkX
cjDDnv4Wx9FqzwJDHPaR7PXUY42XyNZHdc6AJtomhptAsQ208y89ct0rmTGZ4Nsi
71EFcRXd9VscizWqFfq3CnZ38sVIPdl2D5NDmyh/7wr5JXeWvrcirlTMCYrYnoLb
maiB74Ew9Kob3Joq6D7uPp9wHpTuCFPKpl9q5NSKsDPe7FDC61PH75yJqGiZ/imh
UJ64iNCFPQnK52MR+VQA66LulgCRrJKuEJHMxbQW42pX0kw6HSCjkeG7SoNfRj+W
MlIujumTQPsTR1/Z8uGqw/AjYpHDEEndDmh5Dvf7oddkh0FNcIiSodKQQctLYRBQ
FSMTBS+P5uYdof06W9gFqoZMKxObpZG8TH1Ec3YJkxs6UAfSgocWCnjgpXVxXIiD
tINS+ySH4jaXktpiZ147chqmlVbH9pi4g41WCROxCfGokBtHUz+R/+K9m6IdxFXA
TOKm7v/Q5OrZssDA9V7eMMG6KCcmfZpq5vQzKuaQdbAsBWbbZfO1cNRArC0EsSI2
+Q6cUQ1teFmWgCM4hNjapxeBJxUQzVrD4TjEp/qJshzOB82DHiFPDzZRaWIZ9soW
JUvgvwHdeIxTYjrvtl3LAXkijvDQyiLBAYe2QmJil7khdtE1Z3jgCYFXOkFQXdaH
i5mY/iSsLv6e1XBRQ+hcbB7F2GmvdGsTSf4JAlDXA6bp0WwVByKRtLSXj9K3kWq+
Mwp0OesvxCNVOlVUsBXTHTBBhjUYhFHwn4JX7/4s6Sv3skHycMuQXZj4XgyFks7j
+VGqs0aigiFux0KBi0LuEHOONpB7jx5p5FhlGWq8Oj7OPIBCCetmOK1cD7modlcu
Zt9TNZ+e7Qmp7ssDfs3rH0saDT/HqHyDsitpKiRvVrnPRJ+c6AZn/rG7Ri+gkFOH
YXTZkpFXR4k9smdkRsHU8Q4xhXC6G2UcxeYgnAtDJo4ow+caxlb74VEt1GEOiSn6
tk4vgJIR76gKg7KQceKAD+8ufoF39gAopjq0b4lssKG1IuzrD8A1TFzee+/zopHz
0PVSUE2z2SiXc3+V/J1J9ISk/saFPcNWSfiSEaZsxIro3ZMUyZykOhjN7g0x0wa1
U/SUCNgcgya30+OEdW32J8NZUHFmoIGlaZXVunlFRwm5jP6t3TUHyQRUV0EqPYeb
QVSK5IfCVKxoSO+hwtLhlXpZhLFKs6lNARpE3lzKN+RyYTS1wqRISIZB4bI50vwa
0xPruO2BFUujNcygSJ4i3fEckTWTEU7KHRUJbaRcVZu9nxZ2V6InHzyrhbXWlpL+
uENrHLCuXOG46PG5SLHTvnYoL1El2FzSKappb18YmSUXvzK9TY/9WjX8N9ltvbt9
bDMMXVHfPR1PeHd720rr//ybyBet4qqg8Ihcs4Ok3yy6Zbrz3FpPGB37ZA5Ba59M
Benk0Aj95p8S8h9mQVbsL5Mrn5GgOCIVOBIgfLQ+s5IsayPxsTYpYsmpml3UkqUh
P04HBu8mPrYH25eK5ATNTSyV3+niKEogirl+bcdtT6hFmz8e1n8iGAsBj4WsQme7
lYroMZ+vToFXFly+NzWniEcd+v2PDrHTSCAkiIe2u/UjAaJe4gpmNynGUIBHpeVs
RjYWyb0WGW4mNDKnctD4fFt2wFgPiM1hj+W5p5/O6PRHC8uZ0rgo06LKCfK1oBBB
fGayrwHK+KltbgyaS/rkj93TLYO0NpqcoJij3WTDYyc9bBSq0VxbAE3+v75uWf2H
ZL3wjETEB5ejw8pujLRqy/8VrLKVgrFW2adocNwqWL3ECYXktwgPZwHml7/f2pBR
oBA/c3zqK35Hw2sPENiLaofdb1ZImOKO/Lbg2txJPJqPN8/tnId7VFftU8zh+IVI
aH4+mMqOVwecNwgvhma/z7hgCQx7hyIrcXcL+5cEvkL8Af8kst34YQrq2Pehdx/6
c/uDoR8Uf75KEj/8oncyjIyalw3t+W9q3NsDsD4cdFE+l5JMQQWG7Vp1ZqEh5lDd
DqTEH+SQ3yLbbJWZIO0URUkfs8bHGlZm+u3lziua/z7jX8Gv/BUTXRCqR1Cy1PPc
row6m67iebGMTrqKIvgSVpfZJV2YPvltPkkneESL2NNDBUQKvxOUhK9kTUtV/uHp
/r2Ucv+F7VDeDppQtlHHK64+VjJGG1D8UrN2/32uvq1pmEpSryAjchYMxgaDJJfL
0O0ZiJSQJ11ehpMbVIrJ+4c1WLEirsE5aTkNLXz75BnAkU3HeD918rMQaoYdnpaW
qDGXTFgXWfs2xyvxfiO/wTuFmMGoJBeTXF22wiq8YlxvvTOaYudQA6+VLuNC/Oad
A4kKxeAF+80uoe1T8YVQw8TTj9jThddGMCZW0m8+qxk4Y+d2Ux9bzXwAUtMMy1kz
aLDXFsb0xyXf1q+8/Zo6YeYunMuhqqUqTTteBZy8KqV8z0EO5VRFXDcSXl/hBkrl
n9wZjtxEgCfWlm7zVSh2doBq2+kpYkReZX9CQo+3aA6vef3iQmHmuTlWDopzOiXK
/Pwd5tkBpb1158GS8ZMr2+17GnECpfQ52W4WGJWmB2zgzCviI0c9rCHbE3IOGBJh
n/9ZyENJZdL14X/SzfdqL6r8HKweBttlDi+UNAPyyIS0IqOvGJahsy95Hx6ZABdb
KtEzy2hoHyYIS3NjVEen/mod/HeYTI5ksIziskl4znICNxHThQNXjNjk+aswLTRI
j1FyoDoErT9Fc1A8EAzhWMZFNm2dWQrZvP+cPZWAj8p/hqlISYx48qvdYpEiSy26
37mBbHw33XZ/hBDss9mmECvnIMLm2zL9+WMoliG3HbLimDCnERNEjSNJmarMunfc
O0W6vkVDB9pyXUh1LzE/MsQfTGITFYQEGPuDE7QIkS4fQ9waf77LDHsyqI/MqEE1
RycpLkoHUA3DGS/S4B1SJQ2Gu8IX/vHHQHAxecwgTIk//NG2KIHZLHhgHxZr0XYA
vLst7JGOU8xlbLBqMiRQ3ei8rJwSElQzaJylDyzf3gBqSEqq0pAbNmQ+skyGeykf
92z2+gWCH3Cg2D/1mwoKjEGyQ3FP8tbzEC+doToFXypNdvVUP5wtnt/rhBACDqCX
7mu748SPOASTg+zFBn1eWL/ql/TSkJn4IQidZ0tC/i6pKjcjOhoV2VCu897ovS7V
LfC/VAwi95hviLxt7p4ZKrgxHR7kppbtL/ndglCq9bJQbUgt7otGu9LVYsX61zZY
9qfJ/yAmbN9vF+/dxf8p/Xsur3FwzUm0mBQx7tmHaLgCbhlQZPfGWCLoJoiNhoCS
bm18LTsCKJtenC6yglxMRFRFeXxb19Lz/SAz4kw3zV6IyGG5VLKpNSco4RfMrHKf
8K/RWA5EphTr4EHFImEpamBYQqXZwyUE1yWFx13WpSXk03oEhOloiZJQrnxaiciP
GTuV41agXiNdsLoP/PVf8rFBO0+yLN9CXgU6+IxhayNoyGTKu531kpqRHnsrqujM
dl/rv+LnYcGB7MvxtRxVMFmOAwaQefBquS72BZKfsbof15XfUqeiaoyHyppqg7li
iJU0U40o4b7wDOCfHyNqFUXyGoY5VWQIVN81w0ccXDAZUm1Edn8ONIKSAOcr7xtJ
/sJUpUWa1S4y7Db5VSdIK9ZuaRQLEVgo64uvqISYke+93bZSS9p0K3jdPErUiwEI
c8aX4ETJ4kd16QJk6q/U1dpWdSyF34u9wyDPPCqXPNshjfh7qF1e8aq9hU5K80gd
fHBYKeJDQxm/lrjWrYLDtXp8ujcRX7xxXQYSY71sckgrSYh7LJYXmxnRSx/Woy5g
d0fkNiZkX4NT7/fF/jS38cf3pmpAW2aqs0ckSxs2bQg8Ti9PcQ37V9OMIdCxt0Lz
WNVpq1rfF7JVcK6twHV+Z/ZrhOiaztYOrcc7WWGxnElk6QoFY4fQCA2xKeBVowl+
ykq4rk7DKXnEAlDkcenQekUzM8FO60wrdtEPKAZkcqT0YqX2E3f8NxeA63QZa088
lmkHwP6Tuc5TD8v9+iy5oRpdtuPce1MjTkQPGcNTASRs4ShXUCCQoTxYfeFE0Ynm
UOl9V7rlQm40EDR8CKLPFg3FsL2mYvvdnqLx5cX+c3GYXwYdCiIKMa1pupCxxQBF
U0iK024bVPk/Q4v67xSQqcmm9nkCe3+OToSaWE9w9lgKEGtiafGUchLDmvvKX4GO
nCJ1vkGZXxpbLbk/T4WPKR5OlGEOYj0WzJIyHSJW2A3n9XkVHe65yCSnHAPKEMzS
UpRSUUlejWxuoGiL57AU/DgVqyA7/b+HSn5w6xgHurU6M1s06udb2nlJ2Z9bgysG
8UcEZuguAQa1zOYROjh83e+rY1t5nmVS6ZtlRQLyLL+FnHyl32/c92cm1k/HY87T
OzCDcwIxejHghtWCwtP+ykUoAxaeGY8alYV+l8LtBfY153G1QMRwlRWNKEWxF8Pj
++Z6dBmI8Acfgsd8sCVmaU6c7Vf6g/nRuc0mMq4nAx3xKm9gWIV8MmSgaJMERJI7
ldunupB59xkga7/qDDtwUDIHOIcJUxLOHcn5gko6ixZTwDIXd6MNpsfpX8wkwFwr
7inH7RF/zc3e4zDlExfN58ugFuXOpuHpt9oKXU23NIOEjejx/CdARVqkwQSEBaXh
XFfpkQwFo/CFeleoMNYHs2rdRTEj9G4DhL2VBxK0L3EIvITcycaKEXtPGGPWABqS
LhRlZ5YhG0OuVDNCLzfQCHfOZhvdpUuuxZGekoq/LTRBtr5b2BtysD5VVo2BsqYJ
9fC2zHWSSAAlIZuOt4/SCQyOeXFrFzKrrD3LpGB6dPDo5TpRfv3b+Kj0Be/kk24g
0dFzPfuSFbB9OYeFiTygq8mb4fOgUpFjkH0ArsfeSPfc0daqdjSnrdxWar87Qkva
vim7DZzyoCPTRtuGEl9ukXVzDvprpWV1Rv34dYanPi2zkwEROQ1iksGb/hK3opRA
EdYSfcZG9jCdPusFugWn/mwMU6yeeQu9OE5t5OtHTSAwuVHz/lH2pSr3NvyT7Mpa
kS7IZHBqh09Apdf8VuJ2gbEAEx5R62RsNFV6NnOdvpfScuIeUeKxs2pic4F+UaRP
lceJsOxbFyY88w9rVKQFBzpZdC/e7QQe+SOI7viUxfygqVYrvx8JfKR9w6foBTPo
NDSdd53ZYP4JLtzDCilmlHaDBDHKZ+CAD9bh15qLb3gPRo+AJxoT1Oh8GSgFRkyt
P1W4j/9jeJ51sNNEyzqtzbpdcEbIsc/yA03i22Dsi8TlFmh1cxQ3NVa7vvE3PMHO
wPZIUwECPPveVH0lhW6AoX4hfFSuA7HQ59etU/OjoIDFxv51ERixNk9DpMcNp6GN
t/ld8saNsEw789AJjgoQTJTU35wM/qnV8cZy3y/ypKAoitO79oWVl88CmmFPAaWS
D+lHktmKZNBzlykIiOwDxJawj/4byA5OUd/2A51bi9e/p05/WoPX+lpa30ptKWCb
tNmCbdBjsT4Nlb39A7cy51UdwyUopwsH7hczVTnB/6KjcT+ZUDr3Txngrnb4msyX
0l+/M60qqu9NeLdVNjeUVB80AjlE5NVCINLwC1QrusyfELapmMuzBORoJYzN0Pri
SrsQ3o0Q0OcvhQSrVu1yIu8TDI2SECn+2VaL73j+ml2ElDql9FOINvA+sAuEMfrr
UijwVZ+eE99Nx/5wVMObBpepHiNys8Qse+NPUu8dYaF/EyHFUaO0Fy19Lxl9dxy1
gVbkr9Gq/++GyMk6fCKE4i9seN+sEcEFBTrojCEOxUtoMr7E4dd1kA6JDO5xWFNg
2JXZDZgfUkZXeejubqX0028w+gORA+fDachipXJ6hY/xg75lMHJtYKJSBVJ/tii6
gDY1djJVTf7fnbP1TJz0LjHl7GOqO39KeAwxSTNwJqT7Pkr4sJ+JEn08VSnExqXc
B6GNxZjf98YuwWpwyGJqtNUuPc+yRGiq6pYeblu4u3e6PtDGwMnEuB9OplirxF9Z
I6WAH83XDOIpTrFDDNhkG4bokQH6oBwnJduUThIoS569RpvsH3k4udr/W0vLZbT3
7AsVL7M8xw1xIjjfrP6yeI2Vz4W77MGWLQto70Ntn5QlDV58kHR34xJktwXleZKS
kZHR2jETHhM7jLhqCaYzKODdFbJqvmQlQIHPlaenTfk46xa3YLV6o5ayccIlBRfe
EPBjdw7hDJjCuhNR1JHoQccOa/SKSKvWZOJ4uX8T2VNeiAsDmSAxSB/HgM4LObry
WNTBsGm9YCDs92tue3gcve8moMJjqlKygrlkMd61kDoTWAaEopLjyD3hbVyV138h
emV6MWj5Rm2BZ6tyTCXoL/xNxESD/rLTKYOcYERa4gbyXlsmoz3IC9irFq1AKYnH
OLEDxthEuZgWw43BamK4GwQThhOLvceIB3y3/TKtaXnKZ7hamwMmcDZ6VD2DnitJ
J5shASdChvAfWUsUmxMC1L6pQsp13NNHz/8+yGamc/n6KTxvUnThgYGc3y28e5sV
iiRPEJvCM+CCVuwK3YphU5ATRjjEjnBKqNZj1TcwixuGILkSpbZoyDTKeSo17GJX
sFH0H7z4P3EmZA85XOH5GKDm/iNtEr6ANWEXLOnUmymB64WdwzGxoekKVc1Y9M6L
7jb1lJJl4l7PHE/4/xjx8haDWphGi1IuUhB6TfsUgzegFkTfK6Qu6rvM9R8RoHxl
UyPHIA5NjbHTB1F364tP9ICls1XDwMiWhS9v2weFHRRBAybRfZofUAVaz1WMw9kP
jJAj/Xbm1lQqLg5gkwJvcrJ8hKYiX7lia3i2R7xvRAYAheXKgUzZqfgmAhDCggSP
70OyuJ6wJtqofSXCjAbcj/SCiUh1qB/CyZOkX6eLB0jdLgeaqNd3zvpSFTuB2T7y
Yb8o960PUoN10PNC8lMMf/4aGL0VLhnaiNjjD6uYJ4224/Cu2aVfts1ArdT5ow2Z
1Rv+5ybL/Ar2DMxMcVJ3W/uYlCKT1B9A8Ms8F/MDVsWBmXL860bqS0lBMW1SBWxz
ef2lkQ61qqMPKn+2R4XQEfQ0rLYNzmtqm01p+NW7dSM1+qDBj+3FvpcqPSd2H5M/
Xx8ZVgsVZwg0yNDarpynilgqPAAK7/G9YIz6bFKPTM0WO21oBY6MkRTq0WoZjVm3
PjFQWeDK8cgE7Vhqwf5kqXSnXVk38/2k8/XoGXq0EIvTBoCrCf+S+8bW6g3yAWrn
zKCTDORlk+aD0zSkzJMccJf7YQxLTzk25YZ8DUaCixNCxmLaWHv5Mhk5DABAB2Ut
fdBgC+j5pE3rHiuUClkmMzCti5biJeKVGqPX6loHyetSIFdukNXglo5IyZ6CcOVf
qWk8z4ECHonw39RlD/7dDQkjPHJQ2F2VQIZ+FlcyDL4ivzHbkYkHNQtDSMENmNoi
nFAALfuSVZXVBe94zXPNPyRP15058I/HVyL+drrDdLpbZQHqlvJARral4nOIO7he
ZJAl8YrYkr1FAXQRaq11ZQYHW8XmJXhaGwmQGnkDZNJO2YsFB+BLvPKmSP0Qcvq8
idGlNKnhlEjuTlvOjTky3IKLPdEzgn2xDQDfJCjdGLnNP/ZmnRB0hOHniyUOSU90
kUbY05Fc4cyVNVBStRn8FmKBJmx0NlszlJlTfoeTKpSKYeLtFqy+XWQtJ031fP74
CWS+k3bf9RpafNVqmk286uOEPpFBkdvJEzF8X/Eg1RXJ127ljJ3nKahB9f/+DIVw
aMNLt7sdmrxoO6nMzEpHMxiB4kwfrbMHPiZUr68dfz5LEbhsvs/+POjIwXkL7Qun
zPo8VjLbAXszhGn1JMcaD/URSC6PWplyNHp+06UPuJlVzSsmjUXWLpGLtF7379pJ
b/PXe3/zTW2mW1gGw/VyXA3mZWBJFI2V6nBs0uLQeCYsWQiqq5pY+KeDtDhzc6ik
qH58LIk4pXu4AjthKaT3SkS2JGrZ4P8orWynv2/YjejzXEKHIryAD2iJL96T7+sb
FXrZd7Nj3RSPoES4+dXRIM/5u3mYEZ3ujbHvSv2InL+hmJNm6MjXYrZHchbkRiW+
psDwGPS/C5/cWN82nUEkP1hky8b2uZDXyh7DhWsH+DOGqA4laQXcCyMfQCW0JvEf
apdtPoKI/K03LZQHTEpsQRK6YBAhTGDAbigj/vS1YegmrOypcUOf0uYZZ3sqXpKB
iXem/GASnuRM7WMcLMk4I9xUQLQoVxXUpmdz8eZFgJiWrXNUuktS4Pg7GycT4HXS
LNJuWRYdXhTI8afjVZxQE8xYuNnMjSnw8PPbjpZELY2OEPsvNRP7BRUWb9iODXPY
bOTF+ng3t6iJIm0FWYdKGYhf0ytSiXQztdFRvklgDPC3evoS/dQQJ5DTQ1KkZ8jk
dhxvNJdq57OwdZfD59mFemlf+IHddxjmYrQnomAu4BiKC9hrfWImPYGHK0HhEExD
pJen7Q1aYuNLCleT8ys035U2qs2mag+/JeBNr9/Vp9KhqpYkWbTiRaxbBjyzuU7E
BlEgnaP06OrMQcGF6coK+nFCWG3Wh+s1NH0ApLt0q16Uip1poGDHPrmtYu0fKj5Q
Q/LyOMxzzDbwA94Ox3Pj5j8+f6Eqw2vWlDjHZx/XGpuSzugwDSqw48CTeOoAmZAT
M9s/UAjtoNNDJjIhEVdvgJpejzfmVib6wqismjk3wwwysOpNTgknN1EW+kcWURkf
jSnyyQUWlIMWN99smAkBxMH63J/b/rRy7B4NnHyWm5JtljyIg6kdY2CQqo4n+J3v
0moWxuZokD8vuZMhODUCQlLtt3vuE247NnWgEa0bW9ZZEKxfjROA0rJY/n3+gP2w
RUzwRVcpEX+V4x18qjmhcgzxuTt62GyKyL30azCbWrPZKj+hA2Dhu0xm3+MVM5fO
hXlTPHbtPUowRM0wLBAUh3msx4/O4ligJVMGIvJIwQyPkaUEB9pJ6nN+qPh2zAz0
HKCzPliGkU3r2mNBPMsT93mR4Ds4hVZTO1lSHQzsesv+KvV3jLJWvBz4nZua6x0l
k8EchsMHi9EgwHuUe1HefOcQorXVU7ubIcvtTXfohCY4xzL5b/TvQAEVmga/qQGy
bBqu5FRuOfetk+AcUSnFQQ0JT7hUOaqBwxOk3MPRCzVbdqMq0i77coOVJ2nYWXRo
5xwd8PN3opB5CgFyXlk5KtYVcmwEJ4rULTmqlZ+6FAk0TCyZogBxgbYrv+bnFrNg
dw2JUaudZ4g13qQaNuMjaso3UOywTzlXEbNMPX03/A391GDTo/G+D8zjNWa8Q0MR
ekK/3q3Qj+iIl5MK8bOzyyJZ9q0rFr0KYcu7meXqCwRAswlKUAfmYhtyFJLc2Ywy
le6CGUqrunBsxx1LVaDdwbOslNzYA0RdDh8wvybR29sAh2mdhTHFVA9ZC4AGhVaN
Jml22YkPuPrMPt9LHz0LDp3Pi3zbTZGUPWQIIP5v+lBnONqBAjY4J/EAY+m9J1b5
G7E1HoiNrsoujwnlAn4e6PE6fY7/TuJ0zO2T4cLgrIaF6SRfFYPAP2Oo4c77jtVI
linXAT0+SNN3N4nYNvYbpzMkU6xgUdschJ3wbl7byf03Y/9shTMAGsnuuISbLsya
IA8uG6C4dKBNsOzynJPRCYgJEoAVpWH4kTmU0PZo+uF5jzk+eFGjnzCFA8cagSa/
ARHH3k1WeHqbN73Imf7xY9U09i7WZYlkdP3tjevUic21yVTL+Q/EcBEsZhTMbIMb
xRlbGmd+DG9LZ1jq1au+WRelXi8rSLYhS2vdVTsgXK2Dn+opptTc5x6N9x+sx9mM
HnR/MEt/cRIjSEjGC86Acgn0/NdNTvC0kBzrvqfZmW2C6wIEOxMTTihnhIyaITTt
8vCsbKpVKGEgrd7R3wVZ429wIHQU2Qstg2vLALfS23TGKWHWfj/ABgV4HWhrWtUd
d+PmlSs9HFwaA6hWpzIYxYRzAgWtqUhnPQxqYGZfHO3tA+GLIYUox5KUMGwnJwWU
DIVFovNdmcQ7rXXA4QPbmhwcvlMvjDrUhF+RvFqx/dEvOncWi5YU25uqcIuIT3yJ
EAXhqj5bosxbAGPR/f6KJoL0sPye1/rZcFe74p8jTtFrXE4lHcwZAix7aQdhoaU0
dc2OHqwOEo4SrQsxmBI6kdY9K7cmSq3I4qIhufqD6pwl29Nv/R1LEhG1DKbRAj4u
R3e7Gp4XJGXDput+oOgKz/7kzaQtChS1kKCF7g7uGJzJOii0/d41bc0vyI1AVwjt
lXKwxGv4Z0v1PmhWiyH91pd73lzX1/4s9WJKzuGRjGQInMnY2puU/KrTtHKZD3Sr
6d/plO2L0r6qFvowZNlvEjHltu2PphmKfnErkg07RVUxOpN3IaFpgMNqN+IEuGpS
bji5iHG6f8U20wvXy09PdxQiyGt2iWeBVHtjnZ+W4kHgbH19td9OTE8Z7Yvr2WoE
XQM8oseId+7t4kmY2B9mcoZObFOlsDYZpbKlMTti6DHFAUZa8sN4ffr8t+iEKwpd
Qcj9xCkLUES4lYzi2kZaYXtemJ6pIXhsXGXoAc+syYuGaE9jKedV5q8Vo0ujGj2n
331/UQITID7Xm5vv+QGi5bYIqH7bmo1BDj/nqEjMb/pZDgMXCPdicwDG2GkkGcEM
u0G7K49wLjRkACDX6GIhecc6mzI+WeQyMXvw/8T1232HVUlmXKCQkZ72oQAKTw1r
g5CRGljabC7CyNCVzpw88mWvf04ZHEDwJIlbZD2GDSl41QMPVplMzm/U3yUhoLBD
nXt3+GSxxIYHiECpPfCurTFTzq1k7DWdW8Jt2VqELWHjefXfahxNLRHTeowCrrgm
S58ne1dE2Tl03kjdqHQCqM0pYKLbyD6SXA8i42yFcQ1bzsFNDGZ+2n6ctW3PvZv4
R5s3qT6Dqvl0RtbqKESGSaO6lmA1n9miMsnPvBjR0T127xHrZiBPsnGniAPWj81r
/nqOA1vsMCg3jUVKlPmgDcaiBi5R0xDop3myJ6YbioNUUJ9LHuTlvoavvC6P1Hlb
rtGRSlZgMy5eMziMWgFL2fonO/t9sgHB1np9mwpPqnjTFs/AcxXQK7pxrqYgsT/f
7eJop//ErK7LC+twfgH/wxk6k1Beh1CPKyt3t4yo2xIJRSswxkvirsEC0j0m8wo4
ykBv4XRmpsDgUQXPZXvuQtCy5oC2Bi+uFWbyZ1c1MapsFFA4dn9xHBdb9EqyltHR
2M7mVDaQBuaSfEMkJx86O/keDZZx22tFHefvYNAk/IzyAoI8UA6XWiA16NYnStrs
XsfR9pE9TwshePFADit4k88CgJgzXsyiB1kRWZc4Lh8+APQ5r2SnXJZj7MbU9Nom
2P87rsua/tPQ7RXHg6l/IcO9GpfmIDX1an+p0uMmnicbEUMIW2TgCIw5fEN5lcn6
5bncFNCz6Ch4SyMgmy+Xwpr1Qtd93wKYbuJzdwwicBnFOGDIJwXTB4rEF0C/basQ
N+kD/n30SgBCvFhrm6nGznA1MDAueKPuMdl2GAmoW82/+J/OCSCimp2WvcoGe53C
P2R9p25sL7E5a9yQCsadVPW8X0eu8KVEahOxj6TIfh6hzfwRM8XEpdyZd7B+OjmF
CezZRVa4vLv7Imin1myDV7W3nNlKQopYcsIG2Sf4T8mFFp4BOp/3CFoJKn19G8ox
Ygq9CGj4OMuq73OkvKhW3Sl2naKsmw5pV6lNhIDfgfCC6exdlXxRa626kksxMSEb
/5ZHcSEZ8rZjrqcFxLkB6fQn3tHwdGFsGE2tvVjcXBYnyIAIvwwz8eavYfD4dkSz
MC5egpITdAexu8KQblb+ajTURvVkI/BmQZvjZg9VSl3+sWa6jiqM9/Mkbxq77wne
3Ojo6hIr/ejeP1AaXLoquiu6vBFFPaMqDKKt1jSpalU7iDlgl71JN0uf6xHmsc2t
ESH1z9vDmYadJAl14mE5Ywfn3Mc2e7YhpBdPFpc5OwptJcufq/ntk7G1qTq4Mev/
CnYhuU2v09rAZUiSlzvSKUCzS9Is27pMKs8sPEy5HumdpHfQ0YELfhd2fU82/xO7
TSqW/6AgKFwvWvKxXYpftUUCvyZ+D9R/ku3OFyYFwe4TYDBEbu7Cf9N3SgFcZLrD
uaYfVJsEcMsMoYCxCIeAnQwmAtyJyFsNEVK6qGjyOUjy4x0F7gdv55qhuENK1g8T
EOnBJir7TpCRP7/oalEmu1wuqjZrWPU7dlI3n0JgwsfwBXM/iC9WGlUalrtMa6FW
Fef89t/8Gg63Gz4Y4c0Cb7+jYBrh/6K1nb5M/cZ6akI9HSSnNGfHMhpL9sqzsUyV
Kc6vpeeUx/h9qf0LA5nm3jp+pOz2xHVEHvF/UPhWBIXiB4MiGLwAiMLhHQMpUlOV
yrgby0hMAxk37LUUNnfpsUHLe3BHAI3dMdFVEzXtHK5Mu9wOvWd1GUW/arIBWrK6
+ZJGPRx2tJa8NK4dOIvGn670OX2ue/GqMYnRnzAS9ov7jdZTaOozw+knKjhRWjDc
zsjr4ADSQIYH3R1ZYPo3+sRkwzqcb+ZDCj2/wQVOI10RvYtF7kyppSBrRZ0skWuU
i5/a/P2NI88T3Gednaq2ukercZzlwRCKvIFcyyfE7At1i40YUuST76BHGoG84Lpt
1F5lFq4kNEc4hTf5JADwG0CKTEQdaKySEJAA9PAIkYixy0pbxN4cPjnlPsVS6IKA
iYqXvN7PF6ouFvQ8qGOAHdI1cNaPLE0N2icvnz/rD+uitFrxbSFNWu9JwrTtWtJx
tA+jPgH1Wa1opAg0TpMJzcHequoVQc32Y9t50l8i9j/DevdD2ikeFhII7IveApoO
tQhJSyMPejssKk2HuEkKFGVF1hKMtSfxP/Vn7lHkZth6bucNYGuCCGQPDMPM18Ex
qGXlYOP0a9+H6SIW0D/Ysr9SKr9wgEiTKj/+1j2lPLFSQvqZeqVsDR8jIcdgixbU
YG3e29sf0ie4jP6EuMrUHlcoLem0ieuvcT3oOV5DDoz7Qvhq3Qq+902pIKJnkU8h
91v3TF3tHBaJNN1LWFLm7OIS3INpGQxwKUCblN0d9nw2Cv4EocCkOslg59W7y5Eo
pUfhpfeflj4QZu7cKDN4l4LiCjGtJI7Y3W0gutQn6U1GVWt1xvuSRiV9mGjXdlHj
XYzh8ZT4FfmoZJU58dc+nyoFF7rrtvGMtGl+Ff+uKC8vm1Q4hVU7StXqcVKLFgPV
bkcP+fw6hGw5D2Fo1tFLuNWMWXZtdRkLDkXyRD3QaqBdkC5QZH/GJWQ424CNoDAe
/PMzbhIuDkapdbLxHCbYfG+Fn8shBl1w4w4LiLaJp35KbJ/3N5PfTXveQ99XPbHU
RnQX923pZc4sNTgXgidOm7IdgAD4BXo7p37meGEqirtVq+O87xO1gPhiw0dQT8/a
xIXx6lxGQhOIh577HJn3q+SuexDVg/mxwdcrUOMO2mMr71ClajAofq58ZAsEn5cD
1686JR/M5XlBvY8QkK8e6NTG/WVdysNkOHKXNQfCFNkjvmbdUDO5I7frnPZ3Y0Ip
m7Y5TMFB0q402nZxmMpTtZL+L8GcE4rYsrbRtD+NT6tQkxAx2eLdmIQmok3tUWRp
RV1mTY1l9P5DMkikXdypslDUNBJvHPT1GmIw7C26+G3A7Oq/Tkj3EMxKgcjuZQ+x
stsNvwOYeeNSrSlhSuD2H4XCE+sK8EWQAQoVxCSoc9Cqj8cdlJfTdasKUitAfar2
kHsISGOB4Fq1z0vEt7NzrqKbk3t7aQuWlRPOVADRUx7kf9vtbVWauhABy8sVpxNt
/ExtuSxAkRaoKqErJ4uOmSHK+nrLIQFdi1CYJFbOtnI+rW4PRK73qIQQ0GTg2K2u
izPKVJjkJ0BeS2WwdMJaOVuSJ8if1KXVhZIvDSx9QyWC99LKC08tfN5oT5tFetXl
GZCz4vrQjNOwVmymjD6027t/k2hMa9FVXP+sWRLFHm1tBWIm1lXL8USRFn81nuS3
Wx5IshBDU0Zi4IzTe8YoSsYBYp2vFuGPvVh5l2roN6WTGfWgm4RY1Jrlm97uoSRu
oWE5j2QoJSfJXyB0GHCp+OS96CuuN7lfyztakhzjZgoDUmi9WI7ZI6WLATQE2pDt
Vj59eMMjTFla6YTnCE8C1Tt3zlfOuJ+GgTaqjX+BNk4jGh3QYOY++aEbtVZ4ttA0
x+1cIzMqsAJ0R7z5whv5n55BsAY364cwERFUxaTeuXRMNPeo7o9nAWQWzMD4pY28
PwyzIeqGsYlotTpAv4DPfZURC+10J6xRAC0U9RpH2AzxW0weve3yeoCwhOYFuBwH
pfuBTHWSRrUUsbKdOLFYZ5CaPsnoABf5iFaxaeXcsVEOH6T6T1CAL/+ZTAZwm6JX
1DnXWMUl63FXkLA4Tp5giXTb1Jryce45iWGjke1ISNAStylCtpp8Oyo+xYpOmk0L
EjBoV1S/6baPUs30v4xhP2QyiK0x7aI3gk6DKavScOSYw7OA+5i51rUHHjf/W8+/
0JGTacOh85sIE/SxN55KvTZxQhEbvDHsYYtWGV2dnYD+OBKRGxXuiz6YABFfuQUL
6D87eMcEGRgbOGClUoSd5MrWnRliyRI26k//F8GYgKXB/3J+bLAR5+BbJJt/w7FW
YDCQ0CSvp6F58QAdxNLUQaDGeyooPFXAhdi+dnE5lXcqMyBThvrblWnaVHpeyP2o
Rf2SisbzRs+WSQVyv6UW1IZJyEBUywLnKYcuHIOMfdXV1w8eyc3OQzlREeSlAykM
JardZZf3rInhJQalqncttsR+4rtLxsHF85B7FWes/Tw0nLUkoa+1m0p88vBitvmA
8Hxmhno8rJbB0VjaI5l8mF8sxE8Qn+hkflfmlsHJHTCsAde1bmdrZL3IUl6cTMSx
Yg336KIqOjllXz3EHzva+q9OjErvor2W/9UkK/tNF6Zo27AzYFy3EqFOHrNxBS+M
GCVJCGShmBGdKAtbaNKA1ouR78zh30zm+5vrcOUIoCJUyj/BzG+wwxmVTVavtPGj
ECdRvoXixsgiNzeMis/lSiOHcRzG3jmobVG5FR14jpt05gTF4jMGyWci21jXHKeu
o8sU4gZ4h9l/Q2XDsRVdGItR3maa6wDdS7E26QPLhiGzrFyGC94f0EzKqjqfkc55
FtlxG1XlH3ShuA3aKMmMBew/cfAPBO6RkYPM821viLnmxStAdAuGBgwNTQPSxzen
2ClAvdDMvUJN6he5CK09Td+enb7aFosGIFzv4WpRVA2JyeNpSRXje+wY8LpVFTNN
4fcCIvC/Zd3DZ6iAlHeSQcpWXoZcYvGL89pMnC2ZHVBEjKelDXDf+LRHCHk2TnMa
XDGmc7C/U6NRL1jeFkiDedvf15nfT8pHEiDYBbvD245VaXQphv8DIpliubKdAb+L
9KDXcFqcwScwGMVrg6EurtBJpQoItaiw/DyuR14uU5BIh3pj7ijd9ADcQvDedTbt
Fev9VlmN9IIRRlHoz/PHvuP35ILQSPm4NfehxpJtenzdnOx2bk7m7m2xCMkv73ew
vwL76u/8zXnocTW0DSdyBTXv3pHKW4vJU3toOko7SeyhccGe4l3oUej7xOxYzci3
jCGhBqsmzzEudBFLBofDJjPOLZnHvhdvzW9oJZY3fFJmBHOd2G9x4NSw1R+HnWMJ
EwKbrd/OW3Mzdg0wlb7PZtnbqJLUL72GyVtxPfpCVr5sxgHZvdVdhR5Jq40S3YVq
ER69VgZqZGEENdA/lQ+1PUzCCseK42e9f+XSR98WXHbGtEC6IkVaiuPITXXQ7koX
kd63fkGiFPp9Vk4TTkxdcFkW7463qNKmxmHjPrIgyCBMXLsivZ2OtckJSFPDNwAJ
e0XjBsX0xsC0NbcbADWK/6phjHeLGxMVAl4aUPTqv5g+8ijfoI+nA1+1C1Y4Ne5I
B8Ei5cbdl0d7JJb0JBfDFqShteM4itvZB9gVYsJDTFuFC/LEQh93k2yPoDSZXymw
KyEsUVdFka38dh0Usn3vMlLb9/jqJffVS+LRxvgK65TnDvAXHT19mx2Dbw+E66DR
KkpPI0F4SBXFPkCX7osO5VfHt68q/TCOut3Qgt9ZoEjh675J4nlFG+qr9NNuxwl5
vt9NXAOwhW77zknYZf84cP7oNR0MIuQi8lQ6epvffqnKBfuqHp798RPHAuF5LZq3
2Z1XJo4Rwyq19kmk/Ch7VJRLif7NOW0cKEbnTm5C2L3UW9ajoVu2+nuAbCjsVDaR
kK9xVd3rk/jeTTtnjNuQLs4TKQgOMY2wVYmrc1XOnhyJT4xv4DAtQqyhVT/qKusN
nrHDoW/4FKf3l8O0QgeXZLehvy0NqC3EYiBU7p7tyGYLOPjNwnwaDg6T/g4WNY9f
VvWQJGyadaRl5x8hJZHiHnhP7c88Z+wzJ1VR4fkT8cPH2dDe5Pk5OC3yNX4QcPIh
3PJRCO/ObuNBRTsoCrTN8EyPK7AngpeHw3lD4Jbi8DTP22/fRp5qQ3BEFm/dFT4y
cHsXIXZq8PS9al4IokkGfov5+ZpUJlGecK5QO1rkGLBxg8Rj+ysukxns1wQVk2/C
ieLD5ynkv5TXHkfBaXW83x2V4ejViwXhDD/hP88KGn/oTmvUPYjDQ9hY0dVX0FRT
Ahqvn9kqRl+Xftpf10WQpugi6JJ0Z/TJOcep1ih59Q+zBePLzpoSuzZd1Mg4nrBe
8WSktzDfUF1ours3I2UbPKt7A43QdxD4M7W6ccrnSm91oBq2x2a+SvwE8VrSc5Qt
1duKOHTWiupb0iHEz0J8xUaiSsGjpoqRzzP8SqsS6ootHOgHF59cAYA+EgHWhNWZ
8dGFTuxBXqsVp/6hRGfIRaM3x7j5eN4EzZjZHOYYSfju2+4OUPPVn+NRQK73/v4M
bH0cqyxiZkEe0a6W4X6rMMBm6md6g+EEFKMLMosZeV67iaLabbrkaN6/1l29oZSI
7+5kI4afRI5u9LxzqTLZ9uoJ5RfYXfKHHXW+MjX3Rkq24wt808ouDYaC49+5BxEl
1UBIc0IYkjP/HyVAHXJe2qqJvS90p2iUwtYxmGpZti395BeBHkDwlphQQioyIDiD
UyH5FKocq2NrGS157Dx3X3uj9QZkXKDPGAQy7th+gRNYkRxzDEfrjRGCHWqLn76j
hqglraj+r04YMew8TMssetp+5WwkfqHzQAi9qNLqIjbcsnb5H8ajhNc07ibzRf9c
Pp20bpDyAPcmVn3sun2QfkZFmlnacWjC6RWrpxEr3VKsISNxrkOkIojVv9pMYQt0
cXOTDnMwN0Ttayp3x1101eTfViM9JbVJHYDEtjCuwy0BL4FA1vzOqozbwsx2dt8I
9ndfzFF4UpXhyX6dPpolJC96iBAODzWGLk+YB0GbrwBziqBnk8hyHZbcTZayvcKY
E+EKTQcj8WPeQJMf9Fc7uh4ZiFd8RGgAAYfBW3/7uYYCwWzQMcHO3rj4z15DDnzR
mU4H3+qnPWspFXhiVFzNxmSfqqsDAoMmYmqUZzRul6t3TAjrdNeGRZcVSMLiqWWF
z+WdCJ0aIEf/bbS+Ski0/f/NMPurpGycVvcR+QjRQQAERfoDjcGMyyXpt/OE0ZxS
R0PVJOPrp/CwMoVQmwvwNl8IXVSCqppcflW9M5bUe0kdLihbY1ch6im4kxpD+inI
iG6Hf8xF2veLeiHxoVbtGWOOVhjYOS7G9MsTtNP7jNlIdHKi1CFmtPbPqpMugK9m
Rhol35tp01DX1GrOkuGuWZOdPd0rTnRFnvxx5+1WK9ZLk12eP+nrUAZqiZd3DnEn
DFETmJ65GrS1nIuaa71cPaTFKXAPoTMrS949dSGMDSsqsgtLVMgxVr/IYs3gfU7q
V1GbEXs+dqgPQDrsIdfApGX3vDAFUq4Y2jD1ftV7922SNYPqWfM6v4Dc9ih2r9Kn
OpINueLPbvc9xYeOmuwocJkOpCwkJXBeemaofURlN12QqS6wV46IQWpfblkwLcTp
xVLHPevWtfvhCt78GSARPGDQWcsWHXZVX2A6Vb9IhEPMovTXk9Bi09bDzR4uKe5A
jjSQ/Z6BcvsGFUJIvKTnRfcnu7T4VDoDEQN3noSODWEx/+04YGxZv4UyC2KTwJ0C
u7UEdZcXYMV3R2WDeYCzqCY4q5I4m3/eke7B3PiaqDFZsFTe8Mp/EwhSj/OPCyWi
mc2eV6CZs7TCDtUP4dHTWiYcsQO8Op0/HIUHJAtEk77qOqa1DEvEQtLyTCItg69g
Q4Pvw0AeDzj8O0bqWng+VmubYkw9LKVSw6jeg2Pn1zNqJConxG6Y6dLQtzFgcP+F
wIVeZPqprh73bbvmRD0XKEnr2vc3ManSmAJoZk45LQpKO6d5kfyHaP+1Znp2sNQ2
Es01ySfIqkOVyMffQ5dR1ai1UK7dzvOBsDuO8yRkb4X2hFkfGOqdV/sXPPCMVo8I
/2vXFqmQRLWp/8kycNctvlayMfXhOGOQf7+vniMoQvF7/hOdA3p90UUrtT4S+SQC
OZH+yfi5XQIvx1T8z5NXVwi6Z2+siUjQJuHJ7THOPFlxS+q6+vv0UAXpBJaodIPI
Nbof3TOlYdEfBAbL0u+C6WFvIgPtZRtFUxQstqfe8PRmTNPJTXnO5XzzNyG4SvOw
L9a0nZZ1S54c1aeVWt5VUMjfPO2yoD4959fp1bvjptaWwvHK3LyGWKo6D9vqIp36
iLRXfLJcY7QfvuFGAw+QOPvM0SgztqIwb8XoeRNTZyB7AFoQpXKg1VGFct9Sltry
e0x9E0RwyHOAHwG4yFruHCCEhsYBMBp/9VglWlWkbNyFbay5Ah7Je3Jbf1tq6ltd
V0eZksa1/Gp+0vcUPG/NMrxki/3AUmYEjbiwGDDStOM6J4z+AHuWdPSCtT3KJh+d
bSSphE76+YLXyLxe4AGWDXu/ugECydDbOLSyuGC3N8qXG+8jEJIkOmcltgKUWamg
Kh1TW6HhGZj3i7POfp1qaFJTNe+i5DozbHIMFRBIwJN3n0exWBGkIhbfhdrrffru
Kudx3s5e59ZG5/DmLMZYnTRNGk/qUnlNtaAvVvntVdMmgzfmG2jjVIkDNuIUeCiL
jyH9wmpnNFVeVghv0URQqXPaagyw7zng4veAFLv6PCIAX+decjyfxT+xVkrwCnGP
2K9YGBQtXhFMMediju3hXvHUnhSFrVhfQl8auINpbgBn8jJnKCiSaWF5zlOC+WML
cLJHMyPvM0AATpMNtCI6GQPojlULfNWyUdjc1sLuHnrGl3iQuT1+cUPCpS6p6yzy
XLqTZL3Yk20EhLK5WYcXEZCkAqiXHtqNw2rDudazkGuGJPX4RA9aO6ACZ5vidcGF
Rs1YaQGoBXh0ZpHYVPtiQ926sCz1qKPi8z7luoRKy+kQZydCblPWtDNtaytmJf1E
E2dMmQlhz8qQ+wkgkVyHDRpZZs/RXVhx9t9V/qNAPtmVVtsBqYeiNH/LfwMcLaCD
FDl3upkD24aRZ5zfpemxqxm2r2MFVdvYcnuAmoV+E/n6PyQq7bkebOyKNOYJt+1q
a3V6NeM7cCzuzH0a/ntOO6PGjMyT8LwRLn49k4fayv3zRkYSknxciNYwX3DoqUxy
tBRWerBiTZ1kJ1xkhvMuLJkQwzYGjB752OwCV+hDPgI3v30O4FPoE1psNjtPKTmE
W2k+eBrGA/JmGIn23TG012PNPz7pZ1/pOsLkOE0QFWuU2PfWBtsvV1Jp3JiecPhw
WCoHB4KRwxHFFft/cXcR0uyzBgkSSpAHPFOqrq1Ibx9mJswKH1U8+ADDHr42m323
QuZdKCn0xZ/wJT9nPUyS9Q53fOuWp2eXXDJnlBkKufyJktjktwU9kmOh3xht8yTj
I8JfTNqFUW5hq3PVOEBEsN+N7QnSJQHVL6w+6ZBpkakZvGyd3r6s8JFb3QuSuZrO
b/2aM+ZY7utxXCUc6ZUA6EFWWD7Hu/7XINA8u7nrQpW9Xpm2Tzlxwg8l2WA7/Ona
a/Yj2auAoqbcGTZySPyoz7ALeL7UwfgoIomnEfVZd2FPJrWq3VAAKBMK3V2lA3j+
3skdyxA+s/Dym7Rs9ba1f8qg6qwGNr1w0GPitgQ2r2cYrhGRBMmYlOqjA3ORMB9l
mPHlOguxY4IAybrYrdmqHqYnNQbj4IK4Opl5cMN5/B+D3wXTpV9J9nShvtU+xhnN
fYog6kJwoA1Ug7B9qoqZTSkhxzXkgcCglg/mZuLPmItbM8Tls3A/8SJkK4LACa69
cQFARrs8qE/BqinNKl86THiAUUQIMKbvNosz0JBIyVs767w3+WLZ0K7qlRkEVGcu
rDRuP58d3xZsNqOH0ehh/MT1oc8xZJfXzm2wSQwdn/BysMa1ld8LZl7NMTOlNX5I
dNkV+GLvapIpivw+Bq9fNEkfLLv3lT6xIINvGJfbW0++cdRzKftR0zowHBIWF435
SHx+WUN6uaNdrC+9LTwDki3fqNRIcGnzfjn0/TRWGCe2TvDkx41xY/BoutLwywo1
F2JX4VJ5h0S5NjAZ4dywtIaIALzS286LQ1TpaMwf+whWpqgYOE5B+4/sho3plvRj
pJlwXpYJFZX7ZQ7aAJobXsVejtzxKJgoZhuVP5JTyvn1RQT6jJlz0hoKMaG1rMS5
AB3WzLSnFLst07RdWmXYAZDGzPnbv1phADtIaJux+ipHhc47scrNQNI3LtWKWcsd
sUoBREevNuSWOl+vefUiur8Yb+hZ0hAGIVUk9KL77cNLHfVHirDHYNdDberJ9WtR
VRmVxH6TDHXpppWTXGqQnDPLuPAbjW1ui3zZw2jp+nvgIpLoz2W5m6wTak/gjmu5
g/pcXDepu92kD6WxNCTz+l9mjSq1fbAcz/gPfwF/UTfx3p7Udwpt8YcbXcFK3S/d
4SA8IqrCjthtrAFrCBL47Ce6GQXo7M3QxbZELmX/PugGeSAkN6PG5evH3izlfZZW
sjm49M0OeigkpjJRg1wV7o43rPiundKVEOJZYg0AleYHTAcnJE3faiDp6Upc6B9w
ic7EW3kAeB2wIaOqKi7kU8vHd3S9IWoFLMLw68/Ha2oMbSEMmTlEXFH6G8lPWC0y
1NJsOUhlmm0QlWQMQXoawgGjgYE7bCViQk3lS0KRxiLh2JHlxvY3SDB38kG2DN3z
aD2kpFBVfkmk6S/D8rI6FshzXLJHnDbee/N0r01FI0AIwN+kwA4Yhe4BVuJJVgqu
nncZvN3QINubdNSwmOBaq5p6zaaWKUuP5t6PeUGXg1rl2o75HnB3dWzhRc6RJQ5B
PdEBL5p8HiYgATNl1PjNfT2vvTMxILJNW8FanN0yqVJSZKFM3EdLCYwCrK090xNE
GadOSV0wFSV4weCHvWCQ3Nmv4m00pW2bfzeEqgxdCiJr+ErOqECzg5FjC1dksHa0
zcTr18Y5gc7PVIUSF3kfIoUAvko64LCNpRvX/hMlV+zVEjbG0KvSikjjiWL10g6O
9MjCnp8xFjpADieod3uN3o/DsuassqxNAugR2uJJFsTDFGwqVtJqFrNImjuOXnnW
2zy1R/ue9ZOsznA1RNW9/JSkK541PRp1OaUIjgPzOjBMCLCo1JKWVZzaq96BjlBz
oIaQKEDa3mIFt96LONlPg6vaKjt+Aqk6saqjxXLhOFlGlUwFNb1sdLn/UyUy9jdm
Wqtlsrc/fZkiY0SityCzvXX2ztYJMCl9zBZUmXQmaSSQ95GlGadjZngD65zdmNCT
lJIvJMsfTiQyyabQWoUR+dFQeNQOxGlxLb5mXO6u+on4gfG0DcvCaJ4jK+nc2OAE
ZEm5/Ax4+UJSWTHz/xL/yI3dNLG6t0pOy9+nkh08rfaFSiwPpEfGHbxQbxkNG3k/
nTc85xRGII5bXbDmHSPoOwaClMZDihzF2Tb0UPzQlaBaObz3a1NCX7p1XZAigqnD
hiXWzhp0+8Pen86HzWCFh/yC2aoDAMHABzVSw4vqJvk8O3vM8kN0ZTi+I0OBpuGu
4/TuS8fLzue+ho5jNiiF66IFPXrgY6vS2bqW9mDhTUwfDSnQGrO4591Nw/kdrV5L
sZ8ONdiP2m5Obw6tnrKvAUgZvNVRDyj4kRy8YeNuWfcMMDmHnn19wIbwPRnGE4hr
7lbiz81XzVAzaBrzz1xpbbIe9RJ0atQK8L3Bm6WMGa4wNYMh95eqA8GC1RU6e4MF
sHbNsjOEa2i/Pi9EKuvyc+EJuqBh1IB5KGRtemdfkmGyi8v/FQBrqDPgpUeCJEb7
K/P/wNsL0o/qJOCnyxSUqt6S+JV3rHsrnQjMoSsx7gmmBXCeOEHSaJfuQNILpJ5m
9ejcShT9XNRgRs6uLJ1UL8E/G4XkZ0fyLrqcaKiw80xnoUlq7uzBv3EKbMju7yyq
Xl2UmJQMZQeIlaCe2jXCmJBrpA1RHw3tXHc52r49afyV54yptFtVyv05xxdGihkT
pwIFwc1v6lJGtNy37XKnnbyxaquRG6sp2ood3qy3yMOpdroZcnXrHHi5rqh9zh/8
xQrT9ggy3mRCwfoNTsglaKAwC+g/rOGRhk3DYkK9XQwvRpdxti+yoNsI10veInVh
squP2sSS3c2726Y4YUbEaSqhq5qvmQoU+TLotuP/i0Sy6uNAXsQCLMskwYZi+I5f
seTlIFz3TitESd7ogOplT+z2aa3miitlHQB9Q/twhz5YTLHgfdBNXQ5yZB8osQwX
kxTKoN7FpJ2zP7qgfqlF7krrwpE/fLmUKRlHZGHhnI1dR60B1iY8f/cVa0IQ4FBE
27KruwGT8OmsapYU2CUQ0Gyzn3deECwjUpKqW9A7MgdWt2t2pyB68fgNBe1wx1PR
HAsIIEpWgwD6vNAPjdbuvX3kDV1Ccqicmh7zEjEH90GoX+Ix5IxawTjDpGe3cp0T
CV7PpkV7mKvVbn+RblQ24NEyDcqyPyxdPv08nSIWcSr5CMUO95Gw6cst/c77eJhu
vAAAgbDK2ciLolXT91cXM0MhFdkuInnvDXEgqS/KzKQCXA8ycRMdbMBpwgobQjOs
2yyFbjn3glOnVr/ohR22x5uSFx+H4KILywLdCfXiTFiEsi8P+XuFuZnnD7Ns4Vy2
Yi7jVDzSq320JV88aNXS1xWjLrdseUQzUZUc010hoTFy9Fq5zGLTWD/w4fubboXU
EafSkr1ZktsoXbZON9XRNvndCfXQUbIw4VN0TmApurC2PzsiT/nwOv5lMOqgD/42
DuNCgVJC1Cno5pR0EcWeL6AW3aX8ZOPZeyFLdt6rVE4ImUmAD0oU4i8UhJ729xR/
1AAjfjj/CC1qIAzdbXNo3U8QjDiLGEwwmqzS/kq5InJ1lGt30WJEoucqkZ1i7fYr
L3o5Hh+Xgy7EnR8Q56V5fAnOTyJzakWZ4WOER2p7uEaIJ3c/dDNe45Qqy6S66IRg
Vcajq6HwXmHB5HKUgi6rG7eBi2iHnJ3ojISKnkDKgbOiEwauiZ921R0/TtzdEWGg
fv8KXq+U1zxdFJriAs7xuyjetqjgmI6tA7YbRkZTr89hZpRBYjHxpa4X8E0HbmzY
sEhdqi4qhnCcbOkuzjBw5ZijjL6JaM6T/ahKdeZB9iilNjreBpPCqSJVeis+ef6L
j0p8fP9dUAPESdJF4w3Bgb2pFpCe9twypO5WFLc3wpnAO96bataI3v2dCBDCwkkZ
bfV2Ebg/JFA7UJ4f7V49R5rccezdIO7Q/lIuWP/WGMEBsxXXtaitHbxy91RInrRf
ZC8KNV7KkYHG4CD8oy0m70GvlIXXxSeOx7Q25o3ymuJJ5tfKAZv2qagSNCKAfl3Q
UHdCokt782tcVfwgAWS7+e60tkqLApLMBHRwKbYf5GYXpEpc34irqYaLkkKYg173
QVhAaN9BSnOSHkRARcSD51qTKZam4wnyYKAekII2gpLC/A9azopn+dv873FKeWnO
TunI+76Vev8ilv98J3eDyhX5h0rsh2i0PB5Kr2JYc6Re4te4u2xWHBTICndMLhNn
Q7WJH9ww5o1Ja4u62RpVmHQzFhscQpZpwjqLeXN1LMbHQ0WN6oeCqZIn7kIA9JOk
gjX7L8sfKgHyNg1rnuiYPFlRbCkNbkFGpmBtDxOWoe4WQC86tcmrVhnTmpbyMO6e
lG3bjnAH7vcsfttZ4ltNUDGSkvQz0LpGa044tg1rmWkY5COxbGduvRoeoGh58QGe
DJTaS9MrG7PzKQDQXD1NHUamNs2FtR4QCwNkKLx0Oi5/mBJC2MbSFVTBvCeMeVgY
zN8176LBld937a3DHklxFC3uBMUy3pAZEzxgRBuEPDlqftjo+rzoFZUjWNckwndf
20bTDQC4Frmj+LNFYB4ra0dLa9WY3pZ/QMUi7dRTtn92q3dgLSeTGiXsu6matXA9
CGSesOSGe1g8eyIRItAU9sSsTrAGEhNRkD+Oy8x/bfW84nXafUU9T+OJkGmZjESV
4NqcJXEuI0uAESefeBAjSBMURz1uoumjYiXdRCBqDaavfJItgWuBndUgHoauWZI9
PYF+ZdNPLkbiMCzCtprGMn1lh4f29us9XjGrMmapgUZKrpNFm3wyHq6KajiP3H1M
tVo1ay/9Bji2yj2bEqp+JejmNsdu86tyQAaf/RlZCV2KP/v49Ayn/PaPQ7BdJFFf
WXa467nz3xYxoatM7a1752kAqPXRTPSusAgFHEP5yjZF0An9OLCDL12mmr5ZcwrW
pku/YaYEbdYQczP1UWsEj5sSocVKkDOi2qzK4MMm32Hp6iARK0TzRgqJk5NbnXZQ
6PttHouVdXEK5X0Zm5W4QkgA9lWF5Wpi9P4u1TdDF+t7AxbrmmAYfZlSnkEzcbIt
kdlR8MsCUVA3B7edwD8TUvVaPDdVui0HvGypvNV1Wk+rX/InQ4txdCDCdEdrrXG2
VNvX49IIWqG2yFp0Pvb9h3fzBOJrPMY1XW07u5Nn8uRLTX3mm+6dowPc7c+StzWk
oIb0ePvW6FJlG6D0KXJ5HsnzUmNh0vDPHiHeDCriYB254LlDY6wqdm+7L/25CNt6
dHD+wdMhfzU+c0D16g2fRpyw1573akkWZZW+y66Czvf4h4cSX8/EvgMmpNGRfeHM
lx1GCYJo1LORR6xj0HHkAuluUXYyosA29VlT9XoTwlaRgSOLYzC/+gS9faLSOUor
euN9SsIRFUSAu0eqIkDGXPboQAToD8ulynCV6RewUgUChpVMkK/B4/kgn5aEBaGe
1onImxZzUExbLs92wyN6nYA0nlx5yO2y+ipGAsJY0zzVU2g2z2m54BXszs4I9iBj
YOWH3qd5MC+RS+H5OsjBl7GDHHDlMoVZTzg/Hi1npwVM710Ut8FZ2X3cnCMYMeQ7
uvzNKXYZG1N6ZtZk+yej9XT1UYr5BbfyZDwsM8yQ0poErKGPUgzIDPITNa14RHOM
YrAGHYddHc/uXbLOjw6zf4/MkwOMasTukwm26AsngGeMJiwy9NLKT5VtaH+BVi2M
3QXfXxtrM2QFfmebuEwL48EXw8yzmTt0MeJab57GPBMLJPamOCdzpT3uCrhcKkxa
Mm614loETqjHYD/rLAPSHQZ3ccr+e9qJmDw+Nq9eYJGYj4qq6XNKVXZxOGgCyk7o
Bw9sqO5fH/A2DWHR52z/kNszT7PlR5nM6DPbfjlW2UOcCKQH2pTDVx5jRkLaY2t5
a8CwRl+O11X9rg4ZDm42BE9cYSjv8udLilRkmWaX7cCwXBgnJM9rgjujhELt6CKf
z2BUNZ7yDh+WPKgueXBY7D1Dys660zj7qHpM6cmmvhV0QGh2xqyQrsdutZoQWzCr
yXZVMtJUUIBigVFqJXLN0b4/5mB0osGFWKBEVzLeAyXGWI2wcmuf0mZw84ihqS5A
hoAPl1UTU1o2YhtKYMe9On38ucZavSLEwHlTY5UUktboBw7fv/3Evl1fMXbuAqpV
MKYcsACHPydRf/oyXLyrzxKgblofU1kf8dPDsIBB6wAlKrpB39eae4QOkvGtGZ3q
FYdnG8CUEeGUQpV90ncxDFIBJaTWj4pm7/5rNhIrkQwOG0zdhb4imXO7UAtiU9r3
eCMGSpjJ7amdJy1goQQkLlbwHJGY4o0fEkxiIzEPBXo62zsHnTEPNgaveSCN9q15
1hzELZ7ddU79cNLgTkT/BWdpQSE3Q/DiLn2Thf/BAJxGgXuA4xSG5DTlAUxoi9Bk
dwVVV91sRg/0GQa05yStwk6e3O0X7z5OQBARv6vEsZPmLvZWD4H7Hy7GHEVU34Cn
JFrMUvRPAiplfz7EZx9D67zyj1QeOGtGLnqLTqTyT5c1qB9IpodUh+j+rrnTFZnd
zbyab/Xp5idClj5AOUzvatncUKZjC4kfyv9YW3bOUeOuLsMRs/TIhWbuLf8cVXC8
LtxpORphkeTQVn3z2weZfNM90ugHmXIMMLfd4IyKi7VGtDmCqhgB61lnl027kqW6
fME40FV7EuYbkBRKlW1CpjbhU/ojX6NBNOxBNfh9E4J2Veh+kU1ZY3WR3aMHZ2IO
lOjw0j/9dspkvBW3s38cUnDCKOYSIHVlL9WW+0QDrf+jlYYLczkBwbj4VUiUZETU
MhpujEgnp9p5kxh0+fVbF0VfzhZvscoFcYM3C594+z/me7lsZgYFu7/M4Y3Xbcvd
iuXxDmTcpKPjyK+I/rpflA8nUqydJzoQL3CSy9lWfa3bUvN4M53lwwa/I24AlkTp
cl9/5NQr+/Zvyrolnl8ruTMrfRagOXm7jWsu/L391J5MOTMrD3O2DkCDqsf2iHKp
2A20AOKpWDXpALDOB2ASXO62v1/SoS6gyrBq9ctQoB+a2EiAg9cLT9YCszg/46Gg
TD+hL8hgeNu0hAEwphOy/Ej7E4XwfuS3zQyW5Gxf4YcScW1/QiB88w2eJU/g8Iiw
QOrEsBqK4VITPYdcCdiEw7xI4egj9vsVPg6coEvCSaYj6ymhZcAWGKJWWzWRjP2h
I/tog+vkG/u9NL4QFBfdIjc4/OBObmTdM0XQvYcfQVOUrVyMgI4Esasx14Ky+oiq
GuZ/THTvT4tFstCuSFTWTsk0DcyNjImkoRWnMvlfldEsAPbmYolIRZNaadwdTylq
gLTOMOYAQqnpn08QjWWLD8J94qiU7wh0484pZYpB5rqakyemtodAgZMimRTmh5GW
0Rsmm65vfSTn6dJ9OEtYVqXMnFMT3jom6Qfwx/j/3nZ1iEbViIi9uu0xJ2hIPaaW
ZHFTfu8Lhz1ipePugknN7IP8qsd7O++F7i/r/NigBkPUp0tfsyU8z/IZfdqVdc+S
fBkjhaGqybyKE1U/pgR9KtDzZQGLSKyPoWZset8aME+BWUYz8aWjKJLbi2RSS27k
9AC+uP1YEd7nCLpy8Xmd8ymJdeVmlJV8J90Kx+kiwEgToOIG7G7rv3+uxExaFTAa
OMy0OVgIxoMcXPCxwcOXPWmlScN9KZ6dWfEiOxAkVdB+vaV4kL9ea/Rx5WwjQbHZ
/0cWyOAGcStSPS/OnuD6SJTtskvpNRmHPA7pfazRjCcu/N0HWkx78rOjkPGb5jfi
JI6kr4mCrayKSCnsy3Q9UAfzsrzKh+42CDt3vJOGIkFilkLGz7ZKgFrrN+bhQMZ/
GYLYCOZMf0x1Tj5AAAeqvZcJpHQ25uanxKit8B6is/qgDgN0GnBErVlVOSAXFy03
rIkzDfX7MUuFSnp5HelH+PAoK2E/248w4Y3TnZ1Q99am34x81deMuU+Z+aqupxrg
OwjviGIH1c8LKSTpbbaH2GFUvhTg+AJofl21TjF0wwekbmNwaPJM3UMcOeNOkDzI
esgTiwwHsnhCbZ99XwjaEKT+zz/uVjBJ+Jg4kPeNXu9/OcQWBVD9aVNIBmGqEZcg
Sj9NwMOu/vVXPy1qeaoy2fNOLcl16c2C315enCGeupRLvzyT9eVvhIus4qD5x+wR
1oJ+ReMN88ysrSKlgODkd/QCfNHe6ItOBFgxeFl5Cxztz3TCAbqnvlX96qnvZOHd
zf6n6AV092ciIM+r3U9xChY3wAChSr+fxTmPYHs1Iy4lF/1ZvvL9MHtCD6dSiJq+
/PoOUuN2kumifMjer6tKEopxrTZJxSsfY4CeLqxQ+3T0fUgZ3JTkWU/SEh1UDdrS
/X0Wi9wLn7yq/awz2hrAzddCL4ashhr3QRtz5KQpqiOf5GmAn/1mtG/z4RVW+ueW
ySY/8rSXIgp3Cszn+np+L56OQqo6bajbJXsL0gtS1S2F6DKdXnv9tZqsQ9AIyLNy
ze+rk8J76WVYKIsm8ySVt0xY0SWn56nckH923rfKNk9ToslCf7WzAJuIGFn9D5mp
6iNx5/tb8nrPPfi/aVkKUoefRciMgzU/TFgHslAWkQKLHftr2jeK0fHaKY2FVRGR
57ad2VykmiJu6uWJp1X2JZpcnjgWYHV3eQJkUTOJIJmLFxLfEcxeskRQeCLEzior
nq00sX3q16OdFeCkcPYWt7mlSJpTfH5+QLXfc9bkMoNVKj4nTG3vU3m/GJ3vBuq8
PdXzicoZce5GcmsXHmbr+kxTKPVKLvTXgTTfkHYy+kR/e+ZghGRbzEGEJ75K10Ah
2ZlJEVomIhvlYK8nsfk/SV/BXqxD/qtYouNWjVLTvgG6Tab5NKLkfGEHCrtE+amX
VpEtjxnk4LrVQ9TD+87I9JemFFbvzTqLzB0QmRlZa8StPc67mkL+8RqzbPD7YXom
nfmZ2DYTah1IbZRC2GNxFojDv3/HwNeKS24aElZ0aX5g/P7oEszh+HLaj9m82EV5
Wi2xHImCVHsIVMOxUbeJCapPcioRyBQMQt52RxBwcsGPnc8tmpervYGtq7B9x1iJ
YIRZZFmFoSx6ghCP1VkQWqC2cUOW5iPxJtK5cSlTrwJVZ7TadamW7JkZ8ObTnJCD
/M6xAaI0ozwKOEA016GPb7RndrBQ8daqBvWY9WsrskC2iXTsuMtmNP13a1v5/gW/
+xHwGVDiK3jdk2sopLasHmab6UL22hvb/UAq2WRr0ZnDpjiuwKZxPzizuVK+4+63
MFX51jw7hjK+HY5yovgHIvltNsnh3iowLyn5fE6YU8TH2t1G38E8BK7wg1FmYOIi
W5oyQ/ldJEUTZ3Uo7yMoL6qS7AQaMavD5mgZ4uet67Eb5l7GE4xsIp5/6/7xvE80
bztGEFrmTeGMya7dWM3/KgYaNoVnhV2YiVIOBRviFKoWgLEShr9LLEcQTmWWhRad
5qnhM2CHiQAdfsfjY/qKbt/nzrWuYGz38ia5uexg/oU/P/5nMxa8jJqwUAgphllW
xFN28BrVOopaYczJ0QJSEgaIqnf/wC8V3beudetYPv/wXC4mQgJpjK7WKjRhelTd
frE5cHw4vMakYEYd0ytuS0dfdTFJOZRVh8tGQGpTlFjHosgaizEMahO7PYysrxNn
KK1EpLF6fFw0rD3YrY2MjL90na/J2Ag+YfOLWEkOBGqhuZ1JpOZYHN0A7m9O3uzA
CB2AVhM6bXy2RYR2ue9qATVyOAOn7/2DZOoUPLH0Vyajiwy2kKm/0ib7s9A+R4RS
r54HG/coD+/rVt/613UAajkBBsWH8GS0rhVkwXMl2ilxz38pc4qKdPDBlvHaunEa
5T6s0vlXE3jZT8bqbrj5L4Lx9A1uV76aaNH3sR/1MIOZ4TI9t4dz/fS9NxtvLiN6
cnXcttu814F9rlNned6cE607kP++Tv2pLBBx6HihBq25KVWzH/1SluNr4o4Q+D6e
2LsjMFkfTIpyYO4iK0clVpE0W8FrIJP40RoJPn6VllOkFDTbB0mAmT3QMYE0n90A
CeY9BtcQgK2hFEAD2mzJGCqY45ycN3hBIjVYzpObf6dlpNNkAiC+OgF8gLwE98t1
u6d4BrKkndiI3zs6cpiVf0vV6Jf/5MmXmdLtFjFQp6dUQbho/5SX0XSaHaPFu3q5
/RiOIEVy9mN/7aA2E1Cms0EwLoFLtXeo57Oi4d7iarjkk/t2gLWXy4M9DF1pFUUm
+X+/oScxRVnvZxODfkTzaKKIwebqn1YcdxN4j2CRETQAUicsaEcqapfnKy5SOA8t
nBvXvk3yEX1tKJAVSgCAybd0NglFr8FcNb3PHsiVwX546lkaDf+m5Mq81ieJRhRu
uv0QNrmPjtiOlbnEv1bXWJGEbYjTi3RFaeHxd5LcBD0/CPjtCMeJiEj73H6CnOqd
Af/LK65e3Ne09+KNtFSR13d8eFHjn1e/PCRuG7wQ+u8rPy/3BI7U5oC9FU77kTOx
DaE93ikz1ZZ/eWFaF7wRQye+M1M0trzz4ShSBUR1LJUzSzmqyOvi3voAeq/gWXjm
ngd1ZLLPK9krpbK+6b4esftcyKFRTHOcIgyb4lKWxIAwCPFBEz6RvmEiUQ77ds45
CMAjY/3Ra9h6MHgtky6bOoZILnkI2MDghZNj7/l00lZfKx7WROH1IBfkvJZhOaCE
sXx05v5RPnw5mVthnG38tRR60km8TDQQ2ZcAHNdPoSXesIi1amQhGD3TMEEMVFdP
hGPgiHE4PBj46Z1bF0gO+rN0OLUjkY29y7sJLUaw+Jbo7ViybLcE+p9YocExwnoc
zy5zBM60MZDv77G9e59JkWazVm1FQkWVJYuDtsw84wVFN16ERpqkuBoux6DSE94z
c8ZrTdNbZdF2EIvD3pkXDiflyg2TkRYE+TmGG5rhYbWegBu6mC8c+DIUp8oER3zs
uNi949UP6pni2GyOYHqBE/z9GiZW+ajM8YAVSd1vy/ecmz2DG0+c2RRz/XxYrlp2
R5xnFPw2uDq2kflPvPZlX50tJF48q+Yk4rsAtSaJ2URcdVmIOao2M55JBQtVskyR
KJeJDQnoX/mlGwuLn4x9bdG+TKGRPUP/Dz3X2X7aCok9amPVol5HWNBLq2y7rtWv
ixQ6eXjXUlqPuCpkIn/6w0q597xMtnT76LGjXuJ4R20jNYt1cPctaNjdXlFJXMq/
503JXaCLgrfNcwSg0G9fO6QYYQr4ywtiQjjIGJ/RN1B3p72WDT/FaraPz9atBgr1
4SMEU4tEn9ZORXMB6Vai2dAEXscK2j4LqWP3saOFCK8QooZG7YRRm20Wnp9iv5Mu
OHAGmyg3PXcBnIUx+E4+P03vjZJ5FzIn4+ouuTIR50IEfFWDdx7XHniagkpxZjlS
x/kI+rHJoIkf2qQk7qCb4bvNj++GYsFLs/kHq1mmLUVsmsEFY79ZmsyWlHM6RQ7k
pUSrxCH+/s9wgupdT8XXTcR25wXHd/HwAu+hMdzB0VkeYGl+uzbs0nwMtNV8GNSn
e7sl2L4L/0prKY4/FJXdTAELk9wBDsXxes3DeaeQpjocdX6AOpvhJag0aEsxIlar
F9yutK7jXbEX69PXSwLE4qvyTn2+DIAeCoU6+q/o5SEhNbHexbWdvj7sj5o0cZJS
2kU2RpHDIn9p4ReO9BCKJ1T2f0deNqVHdQwEoLvhkDFNwIyyIY4NNo7/U/2cPfPk
kH7aNpcY6FeUNOsfzp3V/XipHGhiS1zr0uDUQlHR0Mohk2b+WmAjxRzkpBiE/giw
toKz2UzmICfka2cuy6IZlTHlWvmA5AZb5Bg23I2GM0TFbEVxno5ZokN+Gvwtc6Rw
kwHjT/sIAuLBwhwJyKSGTH0q0sPJTjLGdPCE8ZHLw3CEL9fJD9Wsdbo8rj36iiZF
JaeQKB4V21xXp3QQ1mzvg1Bcq8v8evBV6dWAKAu4Z0vvix5LNap4/3zeqksqPr0T
XKgxx0aeXbqo3tGFbNn30BoS11HQdNMDrCqA5Rhs9sb84UE+D0QXnOo8N2uT043R
MA9AiVr8L8bKm3zdXJttsnZx/W5DEv3Rrj0B9gTcuBDUt6WhxpMQaULrpqMSVgvR
tus9U541zUZEdd1pXX2+XAvPDY/3L9lRPMvizNTs6Kzxyom28Fftvb1Qrik5j8Yl
pAVQgkf5gSecA5t7fo0knmLxCB4cZgIgGbzjPArHAlPB42SPRuudg9LDqmMFxMmg
MqfxjDkwaTLUkBr6lQ2BLtTluUH/USBkxJOEZCb2dfQdPS5UsG3acnSyZHY0O0Lb
A4MEyDcjj7VmlX0DyixC30/t8qWaaqgGAB0v25B43c/auLITa5HsKO4vtQd1Ec2d
FAQu30mXb5H+17mW3BqNJ25Hst5nTnsPnM9hLMBZK4152ar3aEwARh5i33QQMHTQ
5OBl90w172FZ/4KgdOk5TyoQl8vh1FzwJEBjrNPCZr1+vd7Sd5DxoBsipFwyYjRQ
mSguQH4sSzWIdG8pb5zwLIvMHZ3rdC39NBR3XIvhMcQGKXJlbTQvoAqdoDWGPsK6
kx17W7QUQwj0MAqjBFZA1Zd9Xa1cHil74caMkB4kvnzDtOUAD8CI+O11pEnfIxEz
Qiy/Me+WcsEVHJi/Ue6OECHazIopOxQEx98kLec78daCWjPAVitaDoXKYp4GtX1V
PbioIF/jMmXRj5TUTOV63j0Ijs/Cv2WmcHCJ8L/+IzHjK4vBz3Y4oPLSK9bNerRF
pLQ/q3MejliV9nnQMylODkeFVeElfYajm9TdTfBxOiaaDosI7oBXyXLLjDCAB4nd
FXUsYAt2UTBlsdb4GVKCkvA66QT2iWIfculcw9/EtanEVAeQPgIEsmz45Si7D51r
QvLgmh9Y/njdQ0YhHHEuSIoFAZUT761jASqp58gXd7fGrX6H1oceznKRNP/ISrPi
i6tRyR13KQMc91gv1pD+CsdHQrzOcoJ+m8zN+FQmefhgpqaaXAoAgKm7hLoR6uPY
HMJdj81n4uZT5C+5n9JY6r+tC4uG6l3Cc8aKiudu0Y5kspaT6HSAf8A2xhfpRIMK
BGt6Khdx5Dub7ryiIJNPQVsuKA90PM2n9wwlQMhTik60D/L9+dBbJFJW8/RrHNFB
rV83LUTUwL9Sz5Cf801OrTH0wFtzQCkc8RsE6fSE+iALJuCJV1uBh/K1iGogLeV0
JyoJPcPGgB6epuIss/Su/qENxHUrMUAIoD0MrZPatD/HV1zA+Wt0SzHu3dsK1qKu
Z4hQ5M3cL0zJWcukPRJD1uFQMhG7lt9QAfYXYHEoqnPk0jEEwn0KUa0nZO0Lf3Uc
h8p9jWCQkkz7O/Xg2+eO/HQ/2YdIaQ13KZnLZ3j4YrYCjypSF1W/xBQUjCJgfAbj
m+w0p/c0MFc/gjhi1B+44/XJuZgXbxQ0lcu5Rhh4ZE36fZV2uFYKUtH1BZ+fSlQu
44UotvaNqT6Lqnkz6e/onjd4q3hvBC5y6CRBbCJ4WQdRujYsUdf4ixeT6V5KEPpF
0AzXbB5jzaq0dZK/MlrNy4an6YljTMikXz3UNr28JvE6PJzp/RW+braGuQgLeGwp
b0GgvKeLzopKIEGdbQPSB1AfWyuDHcWlS1RKIguMXRvHLMuz30ia8NqrrVXP95YF
dpcGzGGiK0+TB3DCDITDiodrjxyFjcH64RHCubdWQpkvuhw4e42ILmK9J9wyIeyR
IV8WxsoGWKmcH54biPfBjPwQQlEy8rxFokxTp0KEbF6KzFLVcMPZsy1damH+O5VE
Np1oQYrUeaSkwcupvJLUf8F9Cw9mGW1MkaYVk8nnWr4sZ1OWifSqyxYrg7Nh4Mw+
T97Beoiiutm8wLOPd84y7F5ooFVY/oLdFFZWWe6clppR1MZysowaxB2s1Evb/Eyy
O4YbpnpjjzmYjN1b9uY4IZbNflf2sJvfaJOsqt7VtqyZsbOCL4AhT2LRxUMp5teS
d9W6/wR2doF6wNpf4711zyDiGkh0JFJFcOL460ORlFF+jIjVR6BFweSUwNCN5LhM
dMXvK1Y7tI3BYwZhrWHLPi5JC1Q8QBfuikwZiN/th2xzVReAiAe+ORSizlBZYKB/
3ZrEM3362MMhWj9npJtggqJw1y4Y0/jDQJPKAAVCA1R4XcpC/xJmS92pYiX9g0Wv
+UX9DGDiwapYHAcFWAy+46deobmbTrYR8zzpJmFUIbGpPkpZq9TrhKkZgqDbcvyo
zvpMxMx7uHYSdwoems66hpzOCJUpmxYIbb7sdNg8YiC8eDWzW225fOibqPU/XjLN
sNetjICu9vNLEtC/6lKfMENzVEDgzQGn0FJjinZLVxHtQCCGaQ7WHenxtl3GCw+m
sCPi/qMFdn/aV+Fh22gg1LWDlvLqFUaHiFPbUyfwkjERdFA/fObfDVdjrWxHYJ25
a9UL+14bN9yCDXCbvuktjfLm7oiiOq0ckKIChrdgG2T4AuWR7xpM7QtvoeQdkBz/
yUx/krsQHm5bnEoWvJMDow7xZWk+IvIT3zyqnvib6rRhG+8uh8cM0R3dJQPjdDKL
1EQ3MEkJLLq6U6u6td1xxbWK+ReWObamtnO9p0qyQiCeUxV3sT5KUhnZoT7UZFsJ
lVmYoAl4fhlTO6qRhDWdONr3HW1UAHm98EvHCDaHLczOp115H7Mwt2rsUXL8anBM
Q4MINcNx9nugl56Hlyz1EFlheJO3zbDd1TBhFLLcrR9R92aoUTnIps6z+Ct8p/y/
y4nlYDLEVjuSFrDzOIOcoEU4Op6hnoa1CEV8ZkmzHMgXrMDzzytjAOY8f4+Si7ia
7GnTrm1FodpjKasymLtBpkhIK9yg59kbkwUNoy2tV4hhsKO4frWWBHl32vyCrUKw
IzkpLBvkSJguECIRgqErwl4pP56MBMWaNy6ZBpFYGjv0yAkMC8dLAjlw3CRbKcRq
9PTY+6F8CWdN0fH/D3Vp3llapZLARlI9GCO/3pOhpQ+ifSSt8UA2GZbwQwcitYTO
kz87DINANt/TyO8pI91Zr7xD9S7qpjMdxgzi/eYtDHz4+OeXNnhZNyk+cqZ+KU2k
7uzAmYJVnedVONUNcTsjPTgYy31HlBKjBgxuvdUXNnmTW7UacmOtPYwFODy4LtAd
ZTMFpZhflsl0skbZtfdSDiZEwCjVUXA5srOMmrjSei8KUVUVL0zHryNQfhtHXhTS
ZCdHhgSKm9MOv5WK/EO7zNod30k6F1diDXWlrwQedDRotHfEEKdo/XwQ7BU0B9K6
VJiidBmvMNbs+cRJVXi0j3YDFbQFyu3eqybUa+YW5RG8CwHl//gqIxLtAMsL7s7f
hNa+iPKrFbimlWWmMDaNHas2YxQRnBKgbYbq6RhWn5/WCih1d1l3G8RQuMSJg3L9
c23kBx0TxdipNPtNuQv7F0D8iUE2QIK3u03AYqJ5/xvZLQm8WeQi99+2XQ0otxRj
zSt8xdssumYfTnfd1euygvLZ5gEc/Uj/FAvOIYEVKITiDKk9RqzQCw1Z7e6umt+a
ZjJp+zgPHm2/V8yIEK9mVjKfiTgH0wnqdZV5FhxN+q+LxUeHJoEkPBcJm7tgMzGi
wT7WWhA7WXCZTTSm1rMSBXkXATMzY+PAtB9CTzshYc7C+Czcn5h4Ba9j4UrjyA4f
RdwCJhms7Sw8tPXnovMPs1Lq30pS5tDI55u99ClV3mGiUF5dvwl2rI50FPj11fy+
jg8F02dLrXvu5U0ElUdVq5ND6Q+W/cEgek7E7bOg6xGt61F/n/+iq4Qpf9dAakGX
+cRbBTC/3b5LZfzqrLpJ7SJkib3M1qDngAAWAmuYpdPk0H2NlQc3XP/55X724rLS
Tez1ox8M3SfXon/pa20D4M2F6m0FCrn5p0u4sQ+wW6/A2cPT3okFV5EKS4yAgIZt
40zfwlOueBt+8PPwqiw4gGiWuEc6KlK65WPimLpbNa/5t11vJ47/iJVyiZSLiYDM
9CgYLsxmfplKvhth6O6UxBc/LFEekfrwz1KgCHtJf+MEAkaHjkmNQzMkD6GX3ek4
FvGAfWqKrfUPfUPWQZvdMg5pXDTlHB/r6gC97RnqGJ7ZIt9kHGf3VzE7Ip/aHv5Y
iqquUD6ybG6QxYN8sJEogRgAC3lmddb+zU5S0IJzBfQTq2I50HgAtYTFzZ4AZpA0
WP3tpeBGN8L3hJuup7rcOOUTFGycynnabOIucPLOHngBlgB7JXCKQ+LFp05EX5qr
uyxoyLXrf6nXr5r5okQge1nHaWFMlqn4TChCba/gDD020yIP1bune1tOY4uXdBe4
740T3ugsW1WG5LLs+9FaEwkgfAAgJ95PC2mENQ6h66zWmiGpWsb37RZQQRfPM1qU
/gTDf573nrYDvddQSpeyuFvq/56wJbdfoGIbBAxmvGDXDdJOJOt2jo3nsLQqccP1
P59hWfFEcTzb0WlPvLCwDALfWySxCjiNCGka9V7pIXdDlO5B5HkK1O2RFddGZ/IC
YlYmQ6JGKLRJq1EdsGo66L54t7aujjZvTHw8gWh0drnhayb592wcvkToa6olx3RA
fz6N/wJZdwuAZCrekPMfEo+gvGo++p9Zq+o7Egemjiv5C4Fbikk0/2s6pUQyryXC
xVU9SmOjekjjsuNR6+g2DSvXgkRwvVWmULLNqulwUT3MZrckGiWrRPsq9oh0lGlk
buIBOXtG3xgaSlAg+lHlhOdtixpaSqgOex7dOgQ6yqbDGup8hgt5+Grz8vrH8FgT
o7okBY1FciSj6m2PibtRgaHjqPAscO5PeAPSWnecSyC63ntMK5kDuCOCFaRRR1ID
FnkJgH8fF14jashk5z4wGYNQW/ND1RlgylfUHBX4eF53/22mpWvuM5yzB83lYQ+y
51J0K31JDqk6m13SslzPpTqlWEjcwkjCBYe07rh9Gu9N8qYETrCR7VSvY2Xf4Vvl
NX83wdQbGarz7n3le7jn6XPNK9CrVCK7nS1L7NSg4TB348vKPQAXj9zFCfLjOQUU
gBkhWjMiqThis8NCwSdrYCFRHm5MJWzZwtsUPxJzKx7jch0vVnfyloMxATF+RcXh
xX89Sx58x2jbGFl2TxB/eMbM2szBhTiFT8OQXEOKQOWMi04Ww0o/0C65wYm13oRY
dA4a5QHyx53jmf/vpYqlcTnNrFHbZN9bfenKoZB+xjtlBT02N/25eQ8sNvcj8aQv
RH4lwNz8vfWcN9SbqMpx2FeOL0RqW5NeNBauBVB5svxPg6ATLla4qxJSy2NTnrhN
PGI9EDOuuJPz3JvZtSglVOoAdT4t2oR/dhb3Q1SRmRpTV8A5pmvFKEt2/7z5r84r
yyu77jVDGiIfVaeJWouJkPmp0ake08+Drya93ljt8tOnkMWWqgxGEQ2EIDZRjhyr
7P+pShJVbiAEiN6Ov7A/Xv/NIxR317a/CxFy+UzCHqs6BM1OFyNvKKNE8O+M13AS
bVkcRHvGieb6NSjqilCFwipN2512lmI03/CJVT5CS1O4XqIlemRK/wYA+Y1WWu5M
HiiSzM30NzxrqZlXJX3k9+pomoWFwy8pbqOExg2vu+Tnz0n5nuz8mhO5A8Ba3dz7
v1eYS5jD1rq1dDsgbCKBTofh/Fpxi7zjwLwHOzmkyYcWAkaZF1EhndNScu50dnFt
N5ORu4zCykRQm7Kgf9CSfXAUPFt5HOnbxzyoiv/2b9A7BwHJiwVcAX2FOHx0DlGd
F5w7cmauculHWOOl88qDsObiiUIEDmNfzmxZSdzsIIEBhYaCCDUHutD8FkaXcFi3
fLE059ViVHPLuF0AX6CgmbKv7WFf3IVFd/OZNZmPdKWo7HPPcGzCnpj/4QvUYPH3
0vbTZ96ggnj4jve+L5ATRdiFjqnfh/fN1UjDrZOmgxHIQVk2RErwEqiKwbkKq+yp
d/nDjMvlon6Z2klQnuPvb1bI3uSvcfqf3FXluV0CSDcO6+QRu1cyXKVkWl03vNNu
B+T3XWk2fUi3sULlZXH04uoasSNeDH+UO05aJlZq5kmpaflJXyH45qQPpQl/bc83
Z7Hnd/9qQx/QKYovxN1ZstGSM6DiIymUiPMezDlBe5NeaTr04Wo+QR8oHbqxMppY
G+yQWv0uyDlYsmhPEt5yn+lUb0K3UD1eHBm+xY1Z+1UbTvmgcmo+MpONEExFnfMf
KJxe7H1oWpoOnx5ACv7NNYE5kfwLf0RRPgYzJVCRtlj5e24A05k5OOtSJteHjmL8
Y9QvYBGCbfRzOKhq8mVgSjmERKBDCK/SxE8+u/hdn4CmSmoAzI/5du8iEOrdxv1C
roijSRG5uEofC86+QryW1FRu8Kxzg0a3Dt+ITZ2fnRmlkS7PbSeCecYfz+W30PRe
BlkncrWq/3g/KPWmA3iU+CjnyD1LBBS7JzNIcwK1JGsIsXwM8u3oFcsNBXt6O1ye
+q8jW5umXvjOPsaF+0kJDTdv2bXmQKLsjTNxN1pLGbZM5NH9/fO+mq7zEW+drJ2v
OtYUYeQCY2Pv/Hev21/VovdWmLaCgRf1jXu/LxfyylvTjbswSWo54Z5MFbI+rDev
VaTOMcUgwnq1MF3UoBaF3BwC4865b3mHPx7lK4Wm7H6mJFRJTmyLnmMOxtb7cTQx
6Eccks4bkQgnzOBNzDoENMZqpfb39UBx/nTdlt76lC8twwsNckDSLU39Fnp6ZG7o
6aOR2r2eVBXallaYFqr9ttBVcIA8FRVn1NqK98dbTjIXctLR7kA4yR3j0nyty4vv
+B6PS+2ixooSqw+5MCtV2mPIt4QjgQTpyxMPP//1t0dGCsDGWWsFoyXpTargJ12v
zxIpNxOcbIxg+72ZB/B5Ve12nu9QcsuZFc5Pkv6xrz63Q0uH+UHa3AUic9FqaiLP
L8YavvqfMxMPlzYISPf0fPCL8I0xGo5XcsK/mEb1WA4OxFqDX/rGPCFB7einJzKI
nc3kEn5R9tVFJeoQQIzMXai6+pcN6nNQ78iSZgEyXJhaiDzBZBnb038QEWqKjhwT
V1I2Aoo/jwMX4gMQ2p11E/9Rg13cUd6LYGHn60HLayBmMGCqwClAzSEpu4AS1Pqw
o+HeuobYmpS7DjMfX7AgJX/BxlNzc6nCbGkRIO/B2iXtvGyV4KyzYOcTApw1OJNY
jqly51sNzvEqAPZxeVvKb7JA892Q8YlONIIgcMTnF5CmzNd6wKNXfDV2hhog15gc
7ac+2ANK5IP7QVSucwMDnr0tFpALcJ1HlxlRsfhUD/8Q4pgMpkAW/1bpXUQHpui8
g6/X/+u8nRXNT0SwcfQ751MjUDMkQiP5oG/FFaTOOqkeWvDsXgOdQh/riYQKyoJc
xKPogTVsMO6D8xir8f2QUS4hxFlbdACheK0CxXkqb68afDdnZYz+jxBjxmAbD8ZZ
L+XfprNBzTbkNOv8BYLP9vYlu7GRWn617TjuKMV7UQUbaWIYj9F74+h98A1xENUS
zW0tydVoZa7Q7RJIukoryM9jxaGZX/8Rti1MVeA9OrIUjslgv7rkvHFjjUc3EYsd
eW2T7emn6Uh5eocGuKGrHdV3+2DISrvTNtrT+7YveLnznEUKmD2X+vN3fGmbJrqv
PWB+U3U++cCfo/TJH8SpMKzUWWdtaBvWg/D9KghsGXB9DOPIA0rdrnXLjZlyub3D
yqVdOstGzxK+h01pDhhh5vj/J+ZDnJr4MyBQ2NVu0t2LY8ngSE0a4873A4bQRf/D
2+bkTkzJCSfCRzPWsOYy0sMfVdW058dLppY/QVSvfe2FcGVxanpIwgxCWDUDFxVl
+EXJPl/Hrfjcd4lOeK6qzJ7R2AGYhrJ7u4igBSR4gVVIj6j0/ZZoQ7pkPww6kh2i
CRHozISt8Om4K9jQLBoPRAuNkHQL2/+hkl04ej80zY7c+Km26hOq9BL0sVW00mKg
5SVeub51M6GALbdlD4aQjR1fUMauwmIroZPCPmnGJmrVziwb/Q3DRZ+OecEqDx7W
YvIst5N8RoBFCwXrYSpWJXczU3dpogDeTtw33zVwqFoSxOkak+zwqZ3LX3Yo7r6V
3Gjakw4lcNo+SPZ+xGf2RccGwNZZIQ5HyKcOXzUEYM1ON+FTLqEi0dcqnroEqNU7
d7iSoj2ixBpij9L+wd98kRajC8Ts5Yn+kuN4QsQZd/yoGLqiLQ0jVQebEbktF/zZ
atAg5WwC9T+iZ7paT7v20U6+e2kyu3LQ0dwHUHlXut+pyOwVU5Nlo87BUVbZtRdA
Ree7RBWYz/OglPpUpohFFXm1B3gNnSeVrYUm8wL1fvZpl+xERERpjWH3p3MR+Nw1
AfTyOs0BOZ09SVFnSYScSidoqaZhZEL92UNgKU8/n0RmHymXJkyLoEkMHs9WS0q+
Z/eoXI+eK51irzM39mEjJ7KD5ue/F1r1CAoVWMHzJ3QhYmxw9yiaiOEqWu+tlCN6
+EPJX02L5LeZuOjhcRbmr4RXRuLcw0WwCmsnumoNzKVNZy//9uqbza34FX+6xeri
n/WyEqy5wLZosNk18JDsAreWY16PfEqnwXV5jq5riOTlFTkNxWYcXxFvBLRBYnVu
1wmaIiQtR2Lceur7GYxsEJaVRkC6VhZeEj6HhkMimeRLfV+9dj7qM07cbA1ShXpF
dKkaGBB9S6bjhUXEZkppZlXgXv0CIVPa5dD1JSUE9IuoZhRIcIbAxlUa/kU1wXmt
jeEg8muKM9avCD2bkAL3Cu8tMSvVKop0CfyJFw9zOwJavVZjyI2pMxy7GBJ+2nKt
3u2NRX2qtSFn2k8aDHvm7OQ4im0K6m7j7shb/Mx90QA3s936xXQJu8FdW6UncZs7
aAYuGEXyStuDXIAVTEIe3hKqqvn5C6E4O9qkwBPAHU3ff7sehlSpYLb7fIw9fvkY
FZAw36VylaoyMBTheaOo/dbTFxidem27XhVNH0q4Cw25OqAYYZaPOTs3eJkKs5kf
64jDIbWBcztrFA/Db8vcYWxTK/DeUIDQCPLVY/yL1M6Dl4f+7GgErpsSK0H7cOOK
nCzo6E7yjLg96p44JnsGQV50DDULH0PtV38auMJwr09UG8BgsFZMoMrhgUkp8UvL
1Zqr3PrBXNshSeaZL7LaVspHJVvZyB6lxhtzxcv07efAEUXXxjVQxI8uWMXkcfEg
G2rwuJYtlFQ1BhbQb+XL1A3zZrheSeqi7phAq9xSdHWM/8/oQDF0BDkqR9bVW4/i
Xkh1Hwho1KMA8FH3Haef+Q6t8wcAySiuLoH6aRMs18l6wIEemFgnzrhnb4Zvppav
rc3f4ik4mMGbDQ26L31sc1bbWtjrXvZZ4qPgAU0M5hSshbjTTR6e9Qcs2x8PxjFb
8mIw3pNyW6RQNaJ5k7fo9sfCd4AyYhpHugulyC0I5Qjf+ln6Q0swylm+SfqxraFE
rusSzo7xRRAXYrjkrcc6jcXUXVjkDkpLzANifoslofUm7Sz3ecltr3RLizbcBHqc
5cudbDzYpFKTOZ5BMBX9ohii7TniksVUOkPibPRcB6659h72CvVQRkYJRoKoRuUe
VrsjVeCzbmZuVgC9UwlPKYIoMvXs5qcFNDeGnsa2ggvzBxJFudwuBpFFI+7jVHGG
SEh+aarqLiQR+Li3rMhUpL/J6FCnqZW2XetdzEPPTWU6w1mTUQF9p2Bio+yBkQiv
agMwgZ8kmX4G9/3KTp+Tx7jA+LkLfVACUUZHyeoJq9TVJgX+RakU2H9oSJuI1JS+
I1GfeEwgvJbEvP9UDA/sqZNOWm4cexygUSMK52OP2Ou5nSx1H0j90cSQtvHmxCnj
Qum7ri2JA6nwZ4pqRSY6qeoqqobwpXaDM/f3gVZ+PSVTnITbqTXXH1UpC/Isb773
xiKU+zbRiHd3s/FUegELN2toe6K80nNMtuPZoWuYx+ydVANxcrY0qnkMOZuXTZmr
U9z9Ez7/pq7s8+hBqbxGJ2Isw1sCVK9iTJU5jPVyRt9yqRntJG50mkcici7ALX55
i2ct2JFS5uUOob7wjSGpig+thNnAhFfrsCQ6+8Sw4UdxmJIBCDEKE6whMEOWWrYT
xC8ttXV1kUnYBNy1+Vx+OMwDlTnZsDL8VkCW8HKwbOLrVUB1tEjc4VcxOhLxeYK6
A00fbcTKx3wMSdLuNI3hfvZatz42tQE2pq1SNXneDqh5rrHEGvFBWKwILBG+uRFx
MRh0OxUE2wfcnfgUPQTkJtX7xB/6BZUuUEOCJDV5i4X93/a0AeQapy9rOb8LYhTv
1t+zWBlARvrXdaDYCFbvaq/Xb1MWInSYhzrSBxD9I4zh95jpDBTHLwTdASEDxrLt
/SMzpt5qHR+QNIqQIXJW4jCjSnq3QW+XdwD7QCIPtrIrmiaV6zcAPfVsM9HM5qiT
C8jMbtZzadYCUIRTvstHiDojeu6+m4SD4VmirAlss4yc3H9Qec2IJ5wB6b1lWK1J
a6UU7Qu5yhgbMXdHAMg0bXV3IayZlmPqnGSjg4QBPiWyjxL33Gu6aclUcniU8l17
f9qeBThH/3tWoeEJFNtp37Mb2ddCXkz2XjO4X3KI2ZH84+QBXBYwWAyA51OVmC2J
ELTw9K/WbtuzOxkzTz9eCwgv53T0HE0WBUgxhTFoOp/WL37DtWn1IW818TD4ZbAf
P0WtkjIEnkF1GoB00+NhgAFDSfWU5YDv8LXT60NeXyjmK60N5dkolj34PleT/s1W
T9oxZj5zcg45nF3gsZKuYwXywBJ2ua8J20vo7ylBkKUmZ+4PcSVRBNI8sr6d5Bff
uKgz7SOLkgr/c5ns+eVEnQhOWH78cMeokTI6SPDy8+c1s1Ho+EGviX8aBLDfHB+Q
/IU91QKVnDRJOwXCx3Yu592AJK0YWx1HFKR+pGsWsJLn8bg5NsB/UAQbWo2oQzU9
EYI9L5eohYt1tGC+Rc1AKjQ9ZHR2TXM0F5yaKiMn+JfwXe5KiAgWHmg1nC/tCXrz
4hOK+srOn8NnZyLMQIZTNFEWFQ64BseeSHynxa6CesIBRHVAd9drYXdT70osYFLP
/HKS7lp79L0utMAQrfPoD8WvKwezrKbvzJMnosX7JY3kJ+RWh4ecjQ7CoL5teLny
11vOvqhAFpexIXcMeTHbrofZ/Pfb2LFK4QyilehPc74YmQEyp5jEOOhMYhYCYTsp
NO82A8CTq7uFKIw34vtgKXYh8p2GylgQMd0GYOC9e9FYOsnqF9UsdoadZIDJ3yuW
kDEp1lic7mtv7vwhIjBL3CzkliBuEF2mw3UZNMbGQNQ7ZQExeR2Fb8Zaeva7zSyd
LAHgafqlzhIIQsRmmwSFmNnacZSRhkWW6JBoywcNw0Jq2V6Nzp7V95kOkFDAJ+IQ
NDNXYq0jDRvHGZ2EfXoGTXz3rLPY0RAdpTA4HNE1gJZOFjEo1Z15FM4hikx2DKNE
u1vKZzdq4WjmixTTuutNIlY1o1sre5kItBVl/i9RS9a8KUrO5vwCICwckGz2TPQg
jqjGMLf61QYbv+Rr7+tRoA8Zqg9CEF+SWvAu6af1P2AS8A4sWeTvrXZdlGJrJsXM
p60XaCqiL14r8BgYCD6AtdfBlcn8uyvfuj7BbW+AwCiG5/ppjw2hH+xSi26MBxMW
B6Sm2jb1RDLLZExxoS9bo0DsQ/LqmJ069pRO4o5Dqchv01yYOyiP0m+cZMUYZQ+X
5L8USKoA5EnReMFIvvPAmZXnmz5RrlKsttG7kNqelfqJljk6TvA6egq7VsU/+s2U
a4/ywnIIsFRbS+4SyOiByxWUf9jetA7/qynVY4pGCqNw5lZ0yP/rgvKq7cCBi5fx
u7cwfV0joNW3tMu+rWOm3Sohhjw7VejnYGq15gOoVrCYJsUqvl7W+O1yvXhv6ij1
GhILXzMd2IfKDP0NJO0/2j+2zWbnX9EYJvyj9KIdvrmubkvM4UN2WObtvyoL8kdo
IvbcRSL8lZi9rE6Jf/KO+zwietvemykrQWkAkXiJpp6O/yfPeF8Qgrz6WQZ3Uxak
bTxhkaPinvRcFMgw17svhEy+TXyTj1FOEEsaXWtFDWM9MlJ+e2vu4ZiPrAwmKZW6
oxOy+E7jrzmbCr3YvRy5L2Ap5eMxALe1VZ/KGqkNBT1O3/SWOnnfd3bDCRevfGcK
2R0CR6WX6t/d+QKyrC80uIbVOV8Noxryr2xd0aT9F+or2FptlkiqTJ9uKaYl6k60
lWJShImEm0hymZZ1JMdCYJ7ia2IexmgFF5CV+uhr5NlodwSZVCpZ6nHPy94mLNXP
Q5cUPif9iiMr/0CUCgnIDfVJEALGLMMmSxP4VeHuFHaiz5fm6UzTjerDxIwEDZ/Y
uZdqKswd36An0AvMS21Jlw66hZxXpM+yHy/N90CqfML/OlCbIEQwcIGcyz8kwpQz
dD9wh9SPvYaptWl0q0pJH32TmzWvrHxyrED5SVJDxye8l6Eh1Vw+qP8KMMX0BCjV
JM23RMphoygIgeHkVz7JJksU0GvCxROfn63MS0qJFtOgEW/09TzKXheNgLgFajoy
x7969B6AEqCldyszc/kfG6oYWByrsXMIP08n2N2hQqfiTtxCiLnwnR6GU8ftmhPU
Vx2A1p2NBxgV5C4nWmZRr0KWnLSKR5EbM48bZKy3jRakKpk/8Pgxhb8wBUVjmf1w
KZk4cXC6C4ELuInvt56RGDnQl7oITIHlBl0fz8So2AAsdjYT2ZFUbjVQw3OgF+9P
FOZRxfrCp/5FaB8Bw48ieKAhe7Gg09NDcZwyQp7r2KXnXtUZG4K+WF9v49cqGJA2
xlpuT3ZxEB/yL/FrQy3L7YU9Bc7f8JQeNLegskxDpUWxSWuNMi7eCifu8rBQ3T/k
uaSgtnNR3e2hAhsREgWoQ5JLvKv2FASOuAX+qP+tAKZ6H4h/He+K2dC9qiY2T54e
D6bWl8dOR+fxFaD600veevZZx4f9kdw1kIxrlVpkNRGAaMXysan1V3gjlKenEpsL
WJ85mLbHeqGT1n3FUoVP4eai5scbO3ZL4VAM2YYVtvvERR4UOoin8Tn+C5zQIFIi
nO0nGnR8XPkrTzIhRnjSSljRpzLXdfDxcjusahLamaYoibkMskprO46jfcaaZN8Q
FmnjFoKFEye6tqAHZPKVor7tA19gCF43hwn/tWEFsZjvwDgXKH0H1n+fnjJsJ7+/
hykXD3VWNay3npZa3/lL3lUZklSUUXr/A0vcAHW3oQY5kzgOO9/Npj69fwQJlmvA
8GsQFDt+0W43eojONfvLNMRSNOwFi28AN26rTgDk+6dcxJYAY+vG8yQVJ5kFaCuH
R+RQ1h+FpiyRcLNFAio6lxLv/DSkdPQ/JbyXVRwUXJJRjyZL7xyg18OhjfC8d8dE
Uedv/g6Y2if81vbUNomRZxsgJGA42PRyMJVJFvmVaP6srfN5yjAvjD/qjwa6yxGr
d3OBkPVv4bWqevSPEfHJln/DcDso1oB3Cd6pb1nATv2z+70mroZuR6Yb5HpzXEo7
+sq8jckrzK7kXKosOtyg8lNm7Vs5iEydJLO1yFSvkKOep2+aAysKHmAulQMu8/zq
+ST75xG8Tm/wObUl2I2O5nXTRlZPVO5J0Y8b+cZffPx8FhLeT4axGKtu0fntUI4/
b2fBTT/N2o0EBMfVEzKIvUFrqF7u6F7Wo9upmKC78lUUcfKF39Ss6aGdyG26e/1X
vO+78AGBiVL8jFfOKjkmkDKC4zx0aDVQYDYcr1hwMjBJZ/2zVIMDfM15qiL/J5qG
mckKJqB9P5QILT2ZcO1LYEz8WzcYZWOMV8RfNDfn+Rr7hrck6CvO1/3Y4flQwSai
93+leesnjnVupBszLlLM9z1znRz30HVxNmuNnFh/7qB9yVT6gBYv3Y5S6EraZFKA
b3/cAy74rERNY6pYIrqF/6a3sbaheBaUtV9TeLz/GN9TJ7o2l8lRiMGuOOVDh5KD
si/+H7Qev/JGYMn7dow3YDWWgw1f2WgFrrjF6AEaKchYZQw9s/kqNPKy8AnbPcXS
4uZE2AzMB60NDT+oIRZ533CWrxgN8qxyl6n9D/0nj26jPOQKFhVjLZv6E2E/OjjS
riPMKtrjqR+PEZ23MDb1C3LdXQ7iSTIZNo/Wccu25V8kf1RkkEvF8QcP/XbE+zW0
A9QtQW/IblApozWETF2JPC+Q6f/kqpBhmnRIOSbNM/UY3kCTq0vWk7NF8UXw11eH
rHuLWV0BV1++/hsVTQBehMUmOF68tdU8VuqynyaZtaNTpTSg+D0vXrA7/CVNc4UP
w9VAiXlyikR2QygUR2RkhflUCaZfDb4zDAvLR/yPYJlWOgPtbDfIgPV3OI5Xi/bi
jw/sTug5fXMrHFLfjv9oVqcJi1xv8UIgG0eLYyLdqABTjvWusK910OF51PI8CK6W
pwaOeAgyVueXCUI+nx9jb2MlfYYgE/A6+H8jWneF+KCO/1/BqvTQ0NCFUVkJF9Ie
OcbXtUOXrzgTJGs2t7CdViXlsgsap0VRU/v1iIEjyDTuq+5bE9TCTr3+nKr8Yr0D
QSc4UWEZAU7P/ZUW3S4JyKjo42andKBQMvNVCBJ86trUsWwLfEcKRWhp5JnDCmtb
Jza6O05/UWkLZtpIS5Wa8Kd6Wt2GGXzThr0yiAaEwzj7SH6+UuZHQYbD4Mb/05iy
y+elIdvKk5iZCHNCWOJBbP745RXABP60jp7mgXHNu0wCouQJDHowGB5Tly1bfu7i
JvZqsbkUotIcqAF1jc112SXv8bu7FeT2Vs4eN1BIy0y56eeYh2aYZc8lSvMzlOsc
/jBWnG9oB70GOX5TNR1XKanuTZ/xmlyYwlum6XV/pxM9FzlqxbP4PRCNeXi3HM3/
g4ADZJ+GIRBRkrVutqURKQtqN9E3gQr8TQzynJGU1uVSkPihm+7ehIxr7UWWRlWn
VYaGQoKNlogXBXfF94YR7perVUSG4oXz3B+YEy+10gW6PmtvXYCl41JU0tX+pPVl
20YmV57tbNr+EYiqm6b31dylQ2c3t6C9lyJEsgLyukFhwE5mWp1hrasnjpcXrf3+
q6hiJd53dmXeADvu3kNsAkc042oLABuPq306ImPAnBGhpkC9ePlBi5Bi87Jrwtyw
SoxgglgKZgV4+TLdoit78YoyJuxsaFrYt5WVsuYRgL86C36XrnrhiRJqEX4DyY9K
9wPmKfRLhMWQtbIT1M6IQIWeKAAC4sU0gLQW7sBqL1BFKifypxhgSKIm6fhOJoru
e44QjdxxmsX05SGus5YvU07FlAwoBFvFDf/Xeh8P8RL2GOW/xA17VoeS/7cBtkmN
Fd6IlatJAVFfHMixHzs6LIZQFEwPnKc2c04RvxN1JPtHtPosbShpPJ7fvRYAMHed
zt53GmcSHtLsH8QxXCYxxLqlen9YuDwPW2XWQf/JJnu8npD5GtnqIM7G4Kuf100N
zuYNUO6qmTj6WrXgMH+oi3MwvJIVDW6gIQHhIBKp7OtChPs+zvw1nX0Id5bOjyK9
v40416RbsYN2hILSvNUCzHpZD6Dz0vI6LkBcCQSB0lHPQXukG8bbe1tWRs0A5g8v
549zF5iMK1aFfOcxH1iht2ytbFM/a9px2CNAjk32m/wBrhontoZWIY+PUTol74Qu
uScMWMIHx/CphTVDZVvZvZJwXZ86+EDNVrOvtigjODIs2iQUP9depiwor+5F6jzE
ghAAw+PtSIcaTBJUq+CLvX8DJNJIrpgoTQJAwTwDbJxnz7yWBgQtTwR/pLbS644r
U/LFDAIpZFpnUkbA5sFVj1ktIlPV0nn6qF6ZNcEedLprMRGgtYpt5n10jHA7bDcB
g8g5wmBki4IwtTfGr/GbxlzHJLeRe6edfVE4ZQYNyGyyBE9i8e3Ps7gMmXEkSdCY
SzBMUh3bH/YamkyWFFk4xjrr/hqCkeV79Ide9l5kzZAUAkVXOevoV5b9QtpuW0cz
CoXTAPQgyDQHm6PNMy9jwoEN1IyIFpTF1T0BeMh0wRI1OVnrUAz2cFEFgCMvwBcS
AUoTZTrYUnGhTzoZHpVSCDrKtHA4T9zGbDjfy39uX4CbFZP1EsR9mpVE+0kpKENc
ZKFPVZR9IE7CmQoY0HUkSRFJt5qTXiw8ONLpqFQjvLbrHei7/hdy4K0+5B5vPThk
rT5tJJscGbwiJbBtQpKpcPdBwPF27yuNaMssK+JDwA4aXHjg+mHZMcGHK3GeJEgt
fiYJYxutpxSMUDCG/dp7YuETOUpSLZhnDzK1wf5kLxWjKlnEE2tnjQ8PuC0uUZ0K
kwFT3/JVAeOEdJQutftk9fczLJtc4+IKE27alND1yFBPKjuO9Nf2SzU5vfjdwwLm
xr1r37k0hgCWrIJ2OrbjqrFoz8GJXVZIWihVDlh7hBB7lJlJ4NJMMhz99vn5zVUd
j/AvQUTeraedpXJJEPTq+SRxke+3GHADNyzm56t84OLnvn4wD6Wo8SNXbHVlN+QQ
T255LM61KNOwZzc5YVHidigLa04MXwt+tbftmpguNRF2HABKAvapyE50Vazf+q+X
rt7b+k6c/8+Li5p8W95HCg5GfVwJoVjDJ/hyIgBils3vqO84RxFaF7ubtDyX9dqW
Rm/PDHqadLLyA87Pk4FeJlSqn+e5PND8+oYXQdOTty4vTKfES+VT+cmRnjSXWo/V
iqwAI8BjSn+gIggP2lNYTm8xjS3iwHQFlT7ROVLG6ugFvmb+odbkImcnU+2agCiI
7M2w9rrQ/zsmfzuSD8kNixr+MJVZE0h+e55SGnof+utQhAYeABgDbRANoVoq3pF4
C+8TP5EWIfpHf3OMCLlwuRafAea6eHcxAo4gdyPNf8DI8t5XHoom66hQhp68K0zI
B4R/l6LmcUqrppkRX8MhxnRVMM0GlpfX5eU2M/2igwrEU9Hf0ATFOPfVfO7B3fUy
trhMB9oVP6ccZFYepaNwBLhpVUxBeIhbk1YpJplXEd71hC2za1r8Y0N6pEi4rBAt
LFkcGbvYDffFO8ABH1FtSVnJlGZQxzVYM29HLBhmJbsGKaxjaryy2yYEbOOujhRF
BFcfu+dnQQVL8VamOX4gBNAx384piBCTb9HR+tsAgx4qYMQMIbiMXtJxjvYKmeJi
YZu6qyTLkMFYqwTSjcMrHavKo1X/Lf4P2DmfO1VeRPWAuD6FhwtT1G2ygiNMv/iy
lPQjZgEV8G7VSrFm0Ugd4N+MAyCTsoxrsl0w7Ow2FDPBufCVYXV16J27N8cLKYYB
rMy6HGnWaUt0CBx52LwXYyw+NFFy+WPw7NQgkcgW7lvq6WLNkuSomSBxS1OauMi3
kQhV2AFtt09KVnBnWVUtZB1VYhHq4kZJUIccsQjbYgnhSkl08YzxMZDdVu6itetP
AsbbBxRm26QpXZVyu8aXFINCzQQDCJ+jtE5I2afLkRq/cp66Jzx/GuB7NWlKIVj2
kktd8nSZcY71ff66lURteyB0GP0udFtB16rGaB9I4UOgLUNARbfiFajl+BFX9qF+
kAI/6senhYA6CiNsX0p6WXiitVV2a4ZJmeMKrDClw0VgXw/anj3b5Ixxdlg6BsGa
mYPTlT9juYuuwG76+cOrdXaGnIopQLZm3jCek/jqOiAXVj4wWqHtf7qs+RzuXBq6
aYB7t7LBAJ30Nqli9OO4My00zN7IkuGbIByLaIGzkyEBkMyo/BneJHUUF9cY173W
clSgdAcJfOmJddFbkpy+/3pfKsoIuzHBIKf8S0ZA9kMbJY9XOEW+i1B3p2kmh0Fo
f9whU3kyeBvrNht2dfu5MqYfmqSoqU/b6Up6DJjaNdfzv6P8woa0zmPlikO3sDDx
ZFoH0qsKWyCmsak421WEkCTtPEvc+9Bdg1gY8e9xJKl6TdIqYXCZF0wC3MhnZBtk
KnA3IvWv/K0wF009HnxUenCBPWk4hSKkbFNhDS2gsfouVkQcxp8AS6b74f+9rMiD
KJhhtv0D4eRdPBaHHCluzzluWl8ny10c7QdTF2BrEjqrMnocYAdo3ilnNTyrSP0w
9O7TlLON6KJ9eCoB2I9ht4qK0k26i62qCCX9CbakHWfECQDtV6zLR7SqxlndnMyu
nCRWefkvxk6ne/RS8mAlVqKOExEMASe2BV+29mpZRNUIiBeEN4xw8w4Q1VYqwpuS
gzvpcT9C5c4qD2jm0y4fx/KXOMyzqpfnHsk9S4inqmdfNupPo8YDQfEPiKwWUzT0
5fCAPx4XA0ESnxGfDNyoSxHaMajCjZJ3mCXQvGYLq+H06/EeCHHK7wKWD7RPWqOK
Fs93gmANNjfTO1+fg2GXtr5NTlwox9YP1Gnj+fnIjRCR2X/ONWYzuIhkBrnOnNmX
3Mp/WMEEJ9+ZkWc9WFaR7wyYJQcWKPq0kWcoKEjYv53VtHGOUUmXZeYHVD28/4U6
6ktxhLzKOyzkyB0UiRkvQhOJPv9saIpwPC+hoEQqeB+o+RlNNchG9+Zm9X8UKpsB
pjU4JvdAm4KgQc+SurM1JtqlqnoRXXuSVxirc24V1HJT7ynRpdYF4lFrM3Tvcujo
6FssJtNPThvUx6Pxf/XL2RTi3ZNtfLegQ1ClKRTCVswsRKIlARdoPXmbmeetcrlX
1v4O/WlOaNcNNPDCPkPTVHn3ZrlKMDlHnW1kg6dFoNhYvW1dVsf4i408LB3h8mAs
KvfSlQtcEZmP0OuiSod9rwh7zzRHT2iAOSlqLlWGT7Mxyir1Uq99JKSPC5ZkPk4O
v+Ai2l07krT3HPe7B+LojOmtshJzuveWOpmghJrjUC3HkSSqQWrUqdX8MMMO+fGQ
rpknAgWIGdBMc6zBWo+QUCZ5V2b1lXL8LgplnYQB7tmiggzaNjiltHMFE4wM4pOo
9X2nxFsh4/QA9PyAmndedQxzV3N7JC9B7xFbwUDN2iOjeW44Vby8KyFxcbDx+T0j
2EfMQEm3EIB3y67lYdZAUHSSGCLmK4n2nz+WLD5cj5GFZWHyMLypFtdDTqxxV7aU
8VxjOjtc7KSK1BHDWK2hMd3w+Jzz1RKry+ZvvMGzhijok8PELoFYTJ15/znX0q2Z
YahlAk7QOcutkQpETQFGgFCDjgSf5du/nccmjCeEk5EWRLUBmTZ5rmDf9WFe2IbU
SZOwXy1mIMrULDGlQ7FvAcdWQRmJT1rN88QztG/QDSDm7dFeYv+HnenSfIta/uit
wOHA8zOccpW5VGw7WvFafUQz36E0AX/CYYh0aVbl6U9Jy7ngW9d9O4gUGf8lwzLB
38nD2Qq93iFOuAawZe4MYRYgPdRPGva69xf6uwAwuxIaaAjvLyI/bWsgOeMrecO3
hAtd9gonYCH6A+8DLa6PfQI46bQA2hK1jJlCfuYRXJ1RZEIi3f/rbdGVx1TaNybB
7215Lt6TSyh9nah5zc4kkN5+NogUeFsG1k6P0+XQckVltniflVH7Pg/fQvm0vFd6
ARPNdZDsqF1QylXpxM4qsHXfc31BQBcAc8tbQ3jld1MXTcvkpKfO+bCpd9YyvZeS
RpB/O6Zkr6uWI0V0IG16SqDNTiDO9ktnbEoIWuPc0hzvebiK2btj7TpxTXggubcD
8fISSSq9Di6267g3hk313LkHTFTcS6v0DLHZC4DYBRQjw31e8j3yHxIWHe6CHqjN
kyIkAUBke34JVyvZXVEXIhdW+P39YzRwtyNoMyo4NTR1hn5NdA77IB5bkuNAyUzA
8lGj6SUIB9FcSe/jfMt8voFvo9436N9u2aOvx2iPIkhGnVjxme7HMUtXX4sAmfmF
7/ZQtWIP3rSlNQhQ4T1Uzc1lzh+tD+BagXXm1K26FoL6TqqN/w7zDzYPf/MgqVPd
u0B73tO07Ta+KNadOO31GkV2sGhCRAHqa8bZhVKujd/6anR51XpvlNUCdClNirE/
uA8UmwbU9YTpD55Q5JBK4RNDKdssJyQ0W8faXtqdqPu1HYe5Ligh2Oiwc7odeUBP
BQm68yvu8P1Z0WC/+xOm7JElx87UvxMwLqqVvoyqLYEbS+WKp6yKDCLqAeOuSdKt
/BXS6oheNuVTbSS4y1afGhs+23ohH9mUaNpM0ZaFA3OS4BEj5h+cCAktlcim9BkG
VixZmQc0r2KZRdHimpyN0VppRtas2GMDM30qEUGJ2q9VodzU3g5BFTwgeKWDvIoS
eXDjGPPtouV9m1OLhWfaPN+oIZfOJKS1UsgWZgaH8AEkEBKpKnxDLTAwNKUX3kOh
eyzczWKtXOtfIltDV3z7dQkoZjD60JiN/QN70lJwjHqDcS6mxV6XdKD6/4bXKvTe
eXnYTuLvXJ5BgmC/pyE5cQhGW+Mn7sCxprJ2rd/Ouf0zixHS+tsB3Pi51B2lTiRf
7bNhxP6GA0XNYfnhHefC4RywbeXYt/cMKk4I9GD2l0RuzrOX9j28z4Za3ptr8nb4
ImmCOHUPEi2140zRH+DCvdxwSwdzYGVzgzFLCLXgvZIPvB9s1M3BkHDkqymgE+ex
HK8iBAZdWx61xHaacs8R+WTA4DVCOKQFIYz/SPKhc5MUeRI/lZyxqpqwsxdUHIRA
w7ISVh2yL1d650x9RJlylK3dLKKFkKOAAE3sQRwCdEEPOfneGLRXOCqrxmShBujc
ctv4QTyFmpHwTqfLfBeh9cF0o35yBUOFxNY5tGojkTAOjpJSibusFXwJIBieps2c
sfzXK3RDD4lP+0RCYgV9rB1gIOgCBHAp3nevJBHc1fdzuv8s1QpqC7JnzQ5GQsql
sdkBFQI3FEKYPRIB74RbmDX2e03iRUGfXVPCoiRSZ7opxyh0EN0rHkwEba40ZbaA
2JyIT7DxcTyijT+8fA8dsL2ncV1so6IuDGNwiNgJ6BR7ZB4zWFxk/jrfAXtT0q5k
snhCVbbG0T7CwYVH8zQWmYxZ/XiPOcQGdM7IuDDV4LpWG4Z7Ev9odDBWvJ4k45QG
lCLKj7INVDryCe0huUCVPKaxFSCfjlQwNO2WtxyF4L3iO/4TcW8cqihRrrA1HSLA
POoCzLjCG7Jts8et51v86uxZY+W43j/mDMMwI/Nb4ZsH0qPw4+VX7182mCwWaUzt
nQ9C0fGcEaohRsQw/rsPORDk9uFiaDXSJdxtljgZyQU/uS0rVU6cQoYcyuzBILGr
aE9oGkoyLeDUhH/ERMXzcBAXWvh+Pv+Vu6T8d3J7ynQoooVP5Jmkgo4nOtwoji+n
11RDwZv807aTArzc3Dw/uapd+iwTGUC7sAgxnLXgtqsTzzsuYdLPeI2AfYgo3ad+
zS8N12h3mrX+JKaW5wlt6f3j44zcDCMP9FXpXUTazBRiCKH8KJwUsGWvKLW4WzM0
8OS2YsLkzGKgmE48HJkWyAEhBOuhNQjuNBJ6f5oGbOoIrx5PPR/QfOgnpDRLbJPE
5YlbqaxgoDMn6SY3h4BklEVg70EgNUR69GcuFi9lEv5N/j2NGx88RTPvkikGvap6
OEjFwXXr7uCC96oJ8ghR+Gur5zf7RZ+B+JNwURhI7Wlxg3smEy2jJRdjW6HVDJ8Z
Ai8JLM0mPmVEY/50z9itWXeOKnfb/PXxhrp94TGt2KgCdqgVeilSzSOQyv0TPpAG
Tv/9YT+8YCSN2TqOGXbf5jutxVRYceScmEUhyaUR3iQvM8mPsWCYsLjLpS62T2bk
Xj5l0to7mxo5SMrVvr2r/kctwZLnKQkvxLDiIfVWvmRCbf9hl5hPfcJda+kOH+Mw
yzFQ6Mrtgt7eqVUFhjpyZMnSiI3ywUpfl+Qws2xo91DLAkxapxXwvLytrkgOj94Y
LPAdXxnwU8GzopH92qFYdQj2jOX6PzdQZBp6r+tx1ql3BPDKD0+BEWkiL5LxmjwQ
yQEnqE7gOSMWk3Z4tIgHd5VCj+EDtBIBk+u6jFGpHb/bvD86Hnd6GYaAlPSu4pDR
Ya8sPSVNLYvf9xXK5z1ORv/W9Iwm4XuYqmpm3YL/jvX0VChugCxZre/YylN2TpKn
m5zcCfPBSV/5CG7KfvAbW1uHdcNXH8wblyFXrLDcDTR69nVNWZVpAp2K0YAV5QtR
BmzpdFREAskEYcNESqJETz/yG2uCmlPdfwI2nserFiAyUBsG6ZhRK5+77oxoYCbo
cqMzZbwlYUw6uMjPMKl6OpnnBRlC1/8+9xZIRLTNzDMRl4kvbUZDtZTnyI8jpVhk
WT81aGiFLx10BJXiuHF842muEe2v0x0XkIvpYIwi12FkbU/gg++CUw+MaBjJPnqH
ONVzQerdwOC/yZeYdvIBgwFS6A20tG+a9XNwZpBMXK/NiKRYdgR8/Eiak71NtbT/
8gt/sSnxOpsn5N/x2tWDbY3GTVlN7dNskuOV4apxAzPqC0RtkFokzKuq7mDv9Rgk
WcilVLFlnHvjDJrH17SZ/Cby+fs53erGA9/iy+eo351J52w6pEekx3b1yO0LKHIi
aptdvmcoobqM/t71fzjbtgOqmrk7FtnOlqB6PK8FN3tuNT3DwjWKM53FOIpbIAIu
XUdzp6RlxfHBXwoKnwE5BoBXwZdOmeX+jCRK4m6djgAT/zZ58mDomaX4DzhkMPf1
FZIUjBqJxCySWar9NaFD/lmAWJiyKIjRlSxf1wiS6ASRyJv/ZJdLYFmem2TZeJcp
Q5V3EvqoeICZwnD/S/XXB+kTJGfIS6U7EL0WTn4PUpQ1tjIi1AH/fprJOybPu6jC
JvxhBQUq6TcMhVnrCq4BLBHVveG1/CW/7k5lSSokIsxB02Y03e/wGqpoIDj7xNkF
aKJWeerq7p9RTrmDLwMBCj8st6vNYpIaEM2FiByQQaFj/V6GdFiHoAypNZT7poAq
uLO/PmvQaVpyV78jEVkAuabpxkw0NvNyV1uZNflRhLhnaeOyX0eZvxVErJCI4tUJ
yxmD2t/tBrQ/DSSFjbgANkkFrEpPAVOFU/G5saZQaWWsYyGoaejEZvTYB0r/jGuF
+3zTiLd2I0LZd1Bxm9LkeG4G4cYaZK7bJvJQnvMTM5zV7u9AG8jZDk+T8UkR0PxI
IBDSaR3g1cbnDYsrYhtlUYR4CPYvXtcoTKgmeankzfZG4LeAtf0U3/b/Hng4yEaq
ZVPOPYQdIkoiGjZPyhaQDFBEEM717fkFiP4smymZQAxEPBwKpIXYeVNOFFIbLwy3
B39VToUk9ekEjnUyUI9NTDADHeU8NwEOlgRctZDR0jcDnYT3TpAIHGwQQWRRkbox
zddt2SLpTWsy9voLdmxxCTuY0BPnHOOLYQKWiZOkBlVhagtMft59+NNpOLM5xZow
Q9uAVha+VBy7puP6fdlcrp38M/S7GEmTFwJULswmyHw/uYX7KJDgsFyQJBjIU1qf
/aD/M/cZCXdo+l2QeRlmjvPhFnNgFIabhYoBBZQ64GjT4zCCj60ajpUtVcExz5Ak
ThWsRVb3CZrLNZf5yRNid3nJ8i+qlhSv6vPG8JMZssO3zJK2PWTy/8QiAwzHAzc0
FKZyJ+agC3s6KW5TWKDDFyZARBYa5OQH2C60d5pacbh1PIHPNkozEY5JP3Vi5DTs
i5kXfAZ0uB1gE1UvQldIce6+1jbc1FPH+ui6g9J1fZ3t2/2BvmgzgSFI6tcXXnHx
Qp6aZOtYQVwx7hB2MpSSX4yqjJm5qBFeaW5mY52Qj24S+LwobMYL9Yiz2nIREeET
/FTL7M7OwyXgJFqhDCLR80xmUSn2C4gABnoMyqlhFW3KYYSFzcrf3vY9sDRJFNyr
mFOFwe/2dEJEBIZZ4/RupX1kJop+PLzgxImR14P/3QtFMzUmUpw5t4/cWYl7N2X6
eoYSbtKmI8lUMvUU07/w70eWKqGfBV0e3m1MuzaVC7hDCI1EG7A5RBZV4kXRV7CC
bl/ibLuzw4W7yBeNVdgP9OHV1yczLDpvAjvDGatBxJNF3qqe0ycd/gFz1L50hbKn
Qmrg861ozyFm6ZYUMtSbBZ5ZGhPQSt8m1swjubKztFtemQI85q7oGxPEuZhThs2Q
JQZa7NS+BY5dalTk0a9oytYY+7CMXhfN/04igXXT69afO7Zc4hc8je/MGhoUjT+k
xA+i0kMN/Ln9KgQF3c6WlRD0LaqPLI6uAztM34qsaexpZE4UUemIwGey/mEh43zl
pAtUn7NbyvQHxiGDo6XdSgHkkvKgt3OGXf8ezyjc5Aoa9TF8HHEKmwuVprIBl5GC
JukVNfvueAnYExMCjxHw7XIwS19vLiwZt/SW/5nmOthBuw76PB/7nc2/ZojXysM7
c5fDSUuj/0T2FQ8Z6MRPF/euVjI2gJu6YRN4h+IzTFXfEYpzDQNED26vzEIQ+arZ
bpzdEgr6QTJQk5+RE9yxmg4S+UPVgdY7HZUm6rnxzCOAr0ax+L/ihaL0v0JPne6M
MebhVDzWlNDOblQirCMiM70NTSP0Rl4xR96H2ccF7ydJFYIKrxemOb2OMskjoDa4
VF4kHRxaXSGIbZfCCufBjJpcil8BpG2l4MHlIUI96iCmvwUJ4wJLkQVLH+HstZMV
DrQxK+saAFGiuMX1aDskB7+Se0PcKDymdzkR4ZP/mEOqnqRlpf2pbzbLya0chOuV
ChGdVRuHqq8jZsNmYSBNUWwwPXr24GoLGAXcm1B27A0okH6hD9wcm0vu6TFwZTXT
0ibk4sutTVi5NxmsAzZZ6BjpwAzdi4x8JTh2gQwpxdJFsbDN6LTfXxwJMMr4Cz77
G/cE7L+VWUrz/G+Nn785BmVdWw6vl8jCCO/lLgE+DXpJXqcxDlqC0UmkwZI8sF0C
mVO3L0LmvzfomQE5nzki0bi3SP2eRI/mFxmgVYHBwgeb0si4YNNgtrgVpxtWw8Zf
FN4iIGWRspBYQe6qkOF6tO7L9nzXTJjWPdHExWshlCRvZzxVQNuVV8qn4pz83+F8
wxt/8hyyqd0H444qmaJiWWyGbzd7ubm1AKUoHmlQoTFTKlY6kzHkWH/a0YKPPRAA
KuT3UKRvH9HFewcyxNgGuhCyVs9vm2sPkbVF70gYcZje+e9Ccjc3Z3tE2TDIrSFZ
toffGqXS0FC19xzuQqW50snP4ZJXV+G9gYQB+S8ceAyBGPKXidTeNu10s813q0mx
ZHiLj2Fei5YxgR4WTnQVKh0bhqYfa+2rYJ7fps0ZNTh/lsAdV/MItgMzGZWUl5jS
ut6oOi5Y9ZJfiDq88V1ZWZwHb5EAQPGK29oeT+roNeBHTL8ws1QaPEUICXwCir5W
PRy73effmc6tZbPWhX6h44oapYHadKx7ZzyyvtTWlg0TcVDgwucKsT3F2zhhQO+d
Fxa+wMWp8kG3mckPaWHJAK+skG15pBbJCCc+D19mgJcylPkmaOuuVkuQ2fxE7bPr
Kx1CwL3ZXsejSHLaqym9ShrNRcx+fiv4P8mICx45bAHqz4gMf3kO4K+daPQNow6f
ovaucGB/m9RUmn9qF0lC+o7okTXH2bhb1SpcHh7ikYBb79j7VTiLjIRDuZfRG0Hv
lxf3q1pYJQRXC2qvBQkEt3h9LsQ9uxPvbswNn743rVIk0OeIWG7/fFlKQW4kQSzs
sBnWMge/gjnsrnc+gVM0DTwiV/eEtylUgEudioClFmS+VUctYpbR9ccwVa+iu9D6
4BEs4UMjwZQKoALNgiTE87xOhKTGCNU6/wG/bOlRwVdgQOt1av5zDtlOpWpirg0e
RQaPsD8QNk31ehQpU+tmqJMU4ZE+nF2zBaWZ7N7XCtdkfuwIZP1Uq3KfO51NH0sb
SO+19pnDYr/WKeT2/c5DQ0FkFjKrADbftUPtb5enH5xvDcwqSL80t+HlD6KhDTOl
mVLJaJk53bCt6Kuva117q3A3DyjjK2lHieHWD2b71nuxl16vgZsII/8v/1iByOlS
LyQWhiyx3xgV68Sf+g5t5jnoPwjtyxCoFZMrSX6CuPOnTKXDt9NErM3P5vbNMnfP
4VpV6g913uIsMZx1+6zmS+c6gUaGv4PTIyYjuQqaN3Bn98/9EOqJLBb3IuStzqoO
i4dI+YXqGaUgh1BftmoAi5+749N45COW5hLiOlbT/abw0vdBs3Ojyr/E0/Z47bZ5
FFmq+j6VfdB3GXzcx4vtmvWcxe3VmGrYOIqWuBuvcfriy06vpHzA+KOOnoGZ298T
+L/ml2/9KNQqKME9Z76cVq1PiiNcKWGUORzG5xlJUaYeSq7PCidKPTVMTeQG2Bj5
JOe7ze6vo+Drah8f0Zh3kHo1T6Fw21e/H3XCxLjjWQXON4PKML5Pqf3zZtCFomLu
GwdFjFGsl+iaHbNRlZZr8kVh50P7ku/sHLuJ0G34HN36shxSnWihv6m0RSD0wABT
H3mSqT+B+WRn5nElCq0lN4QjYmLLm5QOzVZDxD+cx0aS7h+wRANxhBi5gD8dpqBW
oWQTX7+iP37GrrBRNyDN66Ox+McykuacfvPJEmXfca9CpPxwu0xL/Ar7+RT+Q/fs
yicJ2h48AwxCANYtXB9oZhJldoln1+cD0EM/pCAJg4eQW6gnifAy6+2H5xC1qW/G
8u/MYI0SJ3/qUwMj4bMdpTZL20ESnqcF5/ZXEN9/DxtOWYVTddRRLkMLwmQkrycO
MLQdhqxrBLcYhOVopgux7oSWmL3uAd5mxkzrQ15Vwa9k+PCs4M5iTyrttHlZM+oW
mxg2cl38cZL+76c7CiNdBpd8pS6s+zbC/ZfRG0xgFrLhVc2lhssgpNIZKagXUd3o
ok2rj7/UnzLYFYQ5OF1bULcw4bdk1BLk+YzjrlXENKih7T8DdSiNEvIbwmrspNjk
HPtRRv/DuRj8Xo6dx3J9gfKERLcun2GmbwFIOq6t0TlIJtKQjZl+0fMBX3Vv0oAR
HTJMla0ixTM7vrIIMUBvjXvlpQBQLX+MW3rVmOcdTnyl4+2YA2HmO71mAYACpT3S
UDw8g4ChBK7iqyIb0sNq46reetWHtPrWxJ6oE748CA39CX8FBMV/AYFQbN2euSZA
hpwnnzS1azQDOj2OOIwgPqx5oqx4pK8t0MH7hy4+JrQK66wJotXpAtuS4zQfgsMF
joGlREXyNsxNzbV++tofygHH411mtUlic9YRnjQ5TPmMQMfQtfmkp95GRECFDFR/
Z81F0blDymdh/biXQzvh6BrTDNU5QD/ySCig20o6Le3JKbC36EUjK1b1iUBFC6QY
fnSLzKVc3CNrdCFZTE2DU6lvNkPpS1RGYjCoNVUwXVdAE5zvw3bq2+osYmc2Ojob
N356BxzFIFqhnG8ErmXrB8cf3t5EnYNchxTJ8hINE0xADGgVYOVj6ZIva6h8IcOK
ytPOG8BEWBs8Vtrq13Vanm27K/fRtkwh2dvMWYrZcCfsfM9DDWB9+ckHw3xwJ8/6
neZjX5KGzUZYg8u5gNB0kyWKUs/gjGD0Yi071w5vOWyKKt28Shqhi1ncg29z3cyX
k+vxtZeT/UDIRZ7wZDkEWWAagQQa351++hN2Sx4Xzd7FUrZQn8SBPhCc1qfpw/41
4P6ofRQFg1KLgrZcNaIMwzDEEZWCpBYMKhl82GycocwI1vCvyjmITpoFYNFBPViz
9Dqs7kSF/fe75cbIt1UTlA0t8K6ZsMEUcHYnZWzb+9XwvCH++kqs7tkKdsOCvt2A
cAtHEdCJSLlcXCJ44yJBwPP2aaufjE5eE5sHru8VKQNgfjbslVlazTEq+K1oNLdj
eDG/z293uNWpfsPR4O10thcNQpOXU934KEaghB/yCKm58p2d0DShjeCk801tu91C
1n3xJiRVQKM/ToOAA1bbN1DMk96WZXYxw2JUhXsdrrj/c7bldvUF/WYIbqX5pw7e
ylfkWm7C5Lz/Oj5Jz/OenARgaIbf6NVhYZVhCEbrS1aLbHwT7qPtdZUYSgU/9WlV
ZaCZ58gXVLR/Zd5V4HVHDrOfrRtORwOXfRa6PURWcixI0Q+7/JlOFCMLiFA0DwAr
jkBcIFEwwrfQPqT+P3vFd71nHdLkjKF536uSiNqtFhqb1XVcWvxQcjmfCX2K8Oux
FAsdALGMNaxTjICj6OXC1kvti20z0+CYZqpme/YF/gN17iwOf/dS5DTni4O0q0Tq
pfY59as0PviGo9hPILVgazbPRT7UwdZWGur5L7+ApL23TXd4u+/Nh2dix891SvYI
wUr9voD+sLNdOxWv5ARdmctCVBgJ0dMK8cbewN/TKf4z46oNpVdWYC0et2sXFm4D
Ekoe6elZRs/E+am0pbNCCkBc6f6uaVoWePdQPRS1rZeCs1D3xklx8LvNQS7tgpWW
wm80WU83PMH1cUdWWKtHZp1KvLHtRhPruM/NFhXOUE900SxZ7VZ7t6YTkxWLU0LC
wkH1HpEinFrlJx/YP1yL++xZAdmBHtgBDh3//kVjaX+Jn0h1RVsqVT2QctVUvHnF
TXweTnqZHJJMqqlPHloSFk1NaLZ57maCMx0GOXDm5yRknu1qba3IkwjQ4G+mz4OG
YnB/Dc/BYsNJFfdatA3X63cq8r5cInaAj5T4U2DvbCMBua7fBU/SA0ax9tFd4bn6
W8PL3NpPurc/bRYBAgvjlPupLNC7HYKbHTMXZbQdUdnwLB8dWLTCBzvth6vC9Uwp
LlVXXyEdNnvSYWTk7BdWC3Gkfu1ygCxS5tK2OA10PCjuI4ePUYcQnQoQ+qRZH2Td
8CFSfK6iEuoE7OrfXRpaavgvTmlhM2HQbRo9rmmRvE2DwdUXj+Z573SkftPcMgyy
BrrA22yjiDXCjh7RAdRnAiSu9rYLqCuJq+gooRGafGNpuGQPRLd+IoYip54tsZYD
GAof8/NJcFuY9ljwo+P4szpPqYdIdO6nDOKJJLCwYUfMrVgVL6qU8hE/7TP3j26v
MwaGbX+WODSBKajDgiXAmcHraVbShFgKHpMojnivxqicyP5yc7uVxyyBUGGMs0nS
fgsgq/BPtYLQlOalt9WXaB4L952dQSbWqM/QCVpT0vYhKGU6dANNNjYzym7Esjh1
264hNzJ12rGIb1U59/nTvCBDD/QXqoWd++thLZ5ciQe6wKnTpCJJWAEMN5NwcHHC
kN50ob0BrZTJmUmaq7pGLOG1PRKokCG1giclA930bkkeIXoFBxET3XXgkJ+BmLi1
0V8gIxgmN+qffgEPbWy5MSpgfRW8u4a1p9p955k2OP9Fz4UTw+X5pdxq65Cneq7/
Ru+qEAVySsLINuN5VE3l+6FjdXxiQ0blOjcTd0yqpZfVtV3RDUKZP4KfWSrlsinh
RUz/DUV75978MFWEfa4PdFZ8GObEsv1Z4du/S/DmnCoXINVFlmN30G7ZNAxCj8Iw
ecgbwC/cTd7GVLKVb7+htFnHvUjo3p8QbtV4IqfGhv13f/fTXFiXXBNnoucDNdvR
Te8FNzyquKIPtWR5GweXxj5Hjl4haw22WYT2cpZQuGagUhaR8ku2IZF2hcmthw51
fCAxGnalf1KS4KOlTwbYhfNsabA2+WQpI1aIxj00ye0DnlmYLgL6ZIIzQWFa8+al
6KmJ67WtBKdUBFPnmFEVTKHQCQ64mjgl5Nkhrrfuhig7JHrFBvnKPuL6OFgv5I75
wPgDR7jzOdg9O4RyFXceHnjWi9Dk34TpWXAd5iOC/aZDVfaoNux0d6Ot/E+/zQwH
KrsiwTlQ71QrGPvpRf/5BF+VlgkKA6Bol19zn3x3tI8mPZ6oFDLgwFfr+HgMj4BW
6e9/5BzTyfhYYYdgvb2F5OdrOCdS0JLsTSxdYsYJbFPAoA/BeHa7RojmoQUtjoSQ
6X5YnMDDVzseKM2wEY7WiEKg0BrYW1QSZjmoqb7iy1+E+Eq9ujRDZwK04sGWOr3r
ClhJUAh0V7qAKXWhK+clTFNf/DVjyEef5WEhLB90jKV30DOCtCHVgm6th11xdFAb
oxYi1BKiKxRr3yGKoJH7qm8pSBAPbhLHE+6TG0aFOj7OfUgNqOb5Y1FxzEWvYyZZ
iKGya9O4QkWLPCo2C6V7z4mojeQQarCv/sSZSnwhfVRgX3T84FhdZMZ8pbgkRBmA
uyBV4ytaGbi1J20DyzQsphV3jkIu5tGpH+Tdy6m1pt05sWzYnRffqhuKm7ZbqJRM
IZ0YU15U30FxaKsgs/jQEz37u3wM8LWXgjz6AzHMzCUhmLs3oXAOjUXzjyCMm2nn
hIXXtXobseyTc8SDfL2/bQsJIZI3/pQoF53kyg3csM+3yj0+zrAbG45A63Yp6d6C
EnpO79ko8R/fyPfGHDy4kBQmbLIrxZZMDcAC+mTeXJ8AjU0d9ctJGJsSpeGM1Idu
pVvFxTGBAtlToszGbQ6ds02ZpjMQqxyHT4YK+VJ4KaeigtneanI1blQOIhMNqEro
rQ+ujWulZ/3LX8b6B04J0Y3p5+eUipaS1BUOOXYtsGJ28jz2rSoD4uNhuxwP0FRu
ujV2f79il4ogKaPpg6ju8lWVSUyhYH32CVF+cOs7h5pcVVGV2b/p/mOtnTw3u0Ry
gmPeCcFwPqMSaPN1GMmEW4kmOdBFZL64xCMKCyaCy+9lzAvMHplsQi+FUWUO8Kdl
XWV1mzomYUz3Hi+Xmm9Pey+apQxgSwKBqDAcdFD3m2M5fUGZOkJ0pwUYBKjomBOq
+EMbpyHvh8M8+LrgdsZ60nbAHFC26gsNx5wS702MMSbGJ9T9L5d2xSLtIqCeF6Zk
P840aqO+x8VTi8N3phBBod9IX1H4Ea15F2D96359jdSUxbuMJLtrxoydgjC6zxRG
yazQUN/Abkvyqq44oN15CPMIwWG/1BlXYB419Si0odaugNM3V2B8QOYvanv+HFEp
fT0AvgYWz/OluzJkZHajUSyGltA0iIxsQ2Kne92Xy3/cHLA/VpNN2ZiTiKLLVz8t
4Ix5goBASQ1GQOpxYbInigR7qPSOutwYUBYhpt72gviqawhIjHF1n1E/VoULtIHk
9UjfzA+Ckab3MriqO8GhKwqqbc3DjjGLiJZjpJP4a2NVCCrIbTS2MV2x8vf1WIXr
Hvd0g/Lq8VhV4OyXitFSvgOKZaIbwCQHQORnMCfc4+S2mVL8f6hfE5PSonwnyEg3
ijBzt2W08Pg9LeR6ZW2SvN3JvooyHBOghSsgHDbh0oENPbtZal9UUJFniFx6sFrr
ESVy+l23yFyHWQD8ncCq3DAKefo3h8oiRsQKTRFHTQHwcN495i/C0HRKWTPJhctf
bxzU528DA3ec5HVvXM+jFlnU28QE/umD+pl3zgjjD6LrxkosbTc6rNKeKSAVRIq1
7uq2xTUsKWLLsfjgXOdc/NH4fEufL1Whsof4OL5ObnobWnAUTLtawS3Jh6G4dSFM
LdriYXSsmsmWdzCqUtf+cozluK4Xg/W+//0T9TdPyRXdjKOszcGypL9Dm1WSAH6Q
DHjB4mVq8uzwHepueFqwTlCX2YjzoQl8X/kMoTpsu4SF2+P0bJ3s7Sa9fX80m3PO
B65r9//YLvVz9kWuXELH/g2yifVAVmZyflAAHAp7eiNLCjqgeUWGs7V4tOAb6iUW
Pf8XL9W2+FtKDdWeRmejzBaOjgxZKG9GOZzNwil4lIU0Fv0JBoUb/NFZPU53tliZ
eO/4Rj/WQCHqhDzb1unrWU7qM/JQLJQ9MkZpR5KLIJn3S7h9g1qMy1HKc200eWae
NpIvpagkeLSKAFd3Vd/ZyCk5vv6hOsJ4tX0IHQPmdm0oYVRhsjiOGuU7vh0NEuAZ
tMpB5d/6sB74qpXwZwrorHC2cSd3+Ya68UtCL7KhJBBMsF/47HalZtDc4ZIbnQ/2
xHF5nXIdnaCWHwpb+WFiHOkfMo6c3njxEPdJ1CQY1BFfK/9ieSoNTpaBQiIJrwS3
skJqh9trh95geSOohQnb97EQwSHP5WDSm2bLA9x1TKwn0bB5DbBetUbp5Y8P7KvD
UK0jIxLkMOrGZsMHxqf+JQ96iLla3UwEIt/CkzLZqbR/9F5ajydTSzMYtHFZs546
58aqS9GAmYk1ZDNRbHr+yzwjHYVt1DHXehC9ZtzI2GlhUXKKWGnUrXpXbOEbo2Ea
+m2ll4Ia1TdrzV0cLqc2Njt/KJc+f1PFokG+1ZmwnOhg64/IrSRp5VYQgcyOgeK/
12Efp0vH6AcT1/A8rMSaI1MiMP9+x+vwOsDPkbjx/xMvifJo2brVubBfA9bdcghi
7XN5oC63aR8fE03zFlplpNxii3apeYRfSCC/mmp3To3d0jnmYmfT9tWv0Bfge2nr
tApQoQDbroNUIut1nh/y8GJG2+s14p5OtAOKOXSCqSUGEBqZ0viWU2lfpfsFnOqt
L/SasnEFbBuEFtK95WZoMJtuE6e8oGlH5bcf1SFRfuIiXVfsjilIjskbNe1Naolo
2IYZqeanNErIEdjilwiizWBM36gJgzkdQUKLRef0w2S/RLY4+2+5n3XqRBMK3MFs
AuxgqHguenUCthxa8ZJiBLWFMd2HzGCUDlmk+zB98AUsNzui98fWV6LHqkXV8V20
8gbhb8KRIcBK932Wr/x7+korbCt4te3J4QzaUVRP1d+a+4asN9kLkQekK3suY2F9
iTH8jJkrFHkVV0JSjL8YCPEg3+3cwjIf3iuY4HIum2a6eOZdaSIbWyaE/xgAO9IC
JOWXUmXp/CIjpPB2kI7k/mz5oXVr1hhN1/XwGSVVTzOoh+Vr+k11Xu67yVGzP/H1
8YAlhQ3STvKar4YSvZ0xZ6tF0ZC3VsEOlqiwTKhdLDVB0stDCA6mZCe8XSgiPevr
0y/gRyrr5vBNGwsX6CJ2EyANYa8/fCW+MgKkk37w7fMCKbXDymKoONJQt1M/Vug5
jZhvDs3/525opKQfvAp0L6m7ct0FhFTQorhMvDdaZ/4XH1vdbvDuxYiiKUEKdkef
+N0tXCe5XOxtJQA9w+3xj3e+qr9MtFKzVNJ+7oRZHgqXO3CsL+QW39WEv+FA0dBb
J63udIxBELWcQJ8By9TcYYCMC4WH/38jIG6dJVkmoOhStWbcBVkVPLfYFCiHVKpv
XkOqOVZ48W8/aReDYZHaJAhx+DEqrHSgYHOmz7SeeuSy+6lGavijjZbwCAU5pIx8
+2u65CrP0VShil98RHJT+oLWIQQ92ax7o+1ebgzl3Mwb3Zx+yvz92/mRTfq/cVeA
QnVGApsPER3MgCW8+1okSP6Hw7ayrg3gDhzJcnAZn36JVYn1/T2+LTfJI7dISlLP
fmGHf+WxFGWEAgF3PhVHJ/gFPvvFWTFxC5dqE3Wm4o+i3JyW9lPPfC07XjqYXZ/Z
1XZ+0I9IqRadBs4/K+NHJ4UbSBlR/vI1JIaHOdVtwngY20O2s9LhfZLW06qj/2mj
7xOTzy1P8/RaZ3DafTj2DSPbVTUHOw2eHXJjqGurnLz57reszO5Tv1wcjToNC/G9
brJAHQBscZ7/yFW80ZD/3TUX1PSt6FuqojXVOrAEh38NCATaNmRIariXTimaWb6B
Q8IKBJq1GqHzMWEq7EU8sN+Ygcm2M57fHNIOTt+8NiOQAmsENGCqJNiC/Rg5TkHo
BzXgI746tR4v17hnoxyiWboVeLCppMbmoSBGvnVIxduMAfgNrCJqkr4QYGtSLB/k
RYTXIoVax4Xx4lUcxoBSEh4zpMUqtcIz1i4fCyLJjn87xmXeTK9tbr7Ox8nK4rFZ
IYnmzi7zPXNMcs4fbK0yL1zH1+YUmybNCzEUs0wqXjDFQoUbvdC4kopKXkC16cMy
ABEvDt2WKtBndqnnHAgaaZ7vyMZX6cVIzxQ0wRaSW2yY1jzGBYHu0IhAq37XKgNg
4bg92SztNQWp/Zaeco+ahkeEzQ6JnO54KVkH0B43dA6p92oiPkLoUzW0Sd1hbchB
utAaiCT8ZgXSlS9SSFPjRrM3eT/d8UloXAd/iqzWM4chcAg+F3ddvYDdUal8ncu2
ZDb6ksrZNP6WJEynfeq7dU7+XJa3tlznvIyq/GRxlVKONzjKtHxRuFaURf8/eEo+
4WkUNJLhcoRDL9t73FliEk+gExAKGi1NH44R8OXQwZu4Fohkek7vwe/dplg4ktsE
k0+FSQoRZ6uh1WTxk97qWl231pKGZGazsB3OnGFHjBX4G9YjSL2sZUjDPw2uPEQi
30VWKazy/rwwahfcAl9LTxbNhySZJAVp7fTjeRQF9d56Bbk+YkUladFHVhzpXoWh
pkf5ENo3f7GQUH7MpU7spaR4iRxmSWGit5LqqDEQQjsBSph9gnRSgivS0nUv3QnR
4a02p7YV2qba+avySiQGPnd516z9K4ECihnZqc4yGIqTZNjhDkX07L9ME2aGkUf7
lhN4BP72veRvgF2Bls7vrLwHv/pBjcAFQNljXAqziDYOpq/CcJ/7NjtTenQLfSK3
kbRSz71obtPXeLM0hQ1lAKMAWcfxXMPtRG7xXlW0mWeCFA9p9M+HOqIWYwTSphGy
9nrhZpNsAXU5aUmvRxWHp5X1iSCoss7nAd0KCjNQBmATOks7d+8I9aMhN5NjZrTP
Jg0/NG+1CeyWRFlo0EodkI/GVj8UDmItiB5ZCruuqV7FA2Tb7gQUVsk/95oIFTBK
MjEwXwz1RejvO7ddbbvtROdyTTlOxf+BelIizX8blMs3zEIKm8egGtvsuxf2NFm8
4ckijzK72imi+DbfXCoH0jmztwsGbxlB76PplzjdZ0TMIZoGCVaOpH1D3DGSSx8F
6K6w8UnramwaMN0YQbZ5+8EaWuwP8b1oCxp4u96pErsAqFQmu582ul2aFkjNbN6H
TUswsQm9IFu0tay2FFNN72CUGQY8zkibqnzS+jcbGx3YAApxkeQZiDyn4t2ttkYB
CuFdfdG5swzWHVM5optSOoSkjrVc80tOZr/uXHqT0q3B7gGUeBlHtETgD/VrVA0k
ToY/i7uXTIo9y02pAnAr6mKDWyBBBLVXVKn4qqrVgMX0zKRsQ53+xSq05/IvXnnV
7ToFywx72y3LNYU2J2/bRG/nXn56QzDpzvqCN87jYGPm0JOO3FgdRnNbNYeNvm/K
fui5m68ypHcP666LBkf5JjPEIv+tbr4/GoDKX+UfTF30OVRMEL+Z7/0wngylGDXI
egFytkMS3YdHNG10oP2lzf4/YPm5WgBumS0Owk7gPmF3zY8ryi0URpwuJ/PKRcy7
Zo35GiPjuQD7Ptvmt+m53IqpE9Ych37khd041cKdP0isBhKYmP5mR41AacVv4INp
ifOnnD1C1MONEWEVs259EWZkLqaGRsm71Nf1y7xARdPVShGNUwtvxvxPFTmnyyck
14ZvrzHPm/Hck3S+Gt1/6hFiMfVKARhwgBcH9YBl6cb7lkztgS7P3bfbhVDBRku/
qtj6y0n1PDI6U9FXMRVBVfzp1Se70BV9DxY0zG4tvz0IjSyPOoxNJM+BOhO+ly15
DB0gRVSHSU/nUPK1rIhcIw2kS3HDuzWI7noRQeIlPD+eCWFSXnBa2a7FE4FdYuyZ
Z+NhDLOV/wyhwUxIQexYMn/fNobRdIWcTFZeMSYAkcmJTxwwBWcT8bEW0HQxr0F2
WOlLiiW7MopxLDBL0nDgHigiGADDuJu/Rf3NUnLN1kpDGYvDSAn8pIWQKpWIIKWA
vKDQTjCWcz4ftf+Giqmu3xyrhmACtahVxE7C3fe+k1OMo2Q38eD1OagP9laJlPt6
SVlcsY91qHcL1N9op7L7t9+7kMGUq43akh0uyYeM44d8heirw/LNsuqwissZuSyF
ZSYf1kAbjwfowb4TxpWtw1zMolRMa561WA7JFm6X98mF6VX6LknIkJEWJBaiE1N3
2TMjK33Z7hD/w50hWFQ+GTF65djf21r8/eCIu3wlXIDVUmzqkiLIQerpLjK9RVGs
SDW9FktZLwpU9VLcprNxerp6PanaknNGeVLoW7jmGRtOYQL+7uGg6DFqGH3Zb+Pt
jlcIm8WIS5EdVsTn2TI/mQ8SGQpWL9FVJBbbiHomuLhDfEJQudmvJxdFU+8u3f8K
ZzX6a5FiHmNa6oLVYFYuMkTl1vN0Xr4znjA2aT7lRoUBCv7+HksDwUdEadzFxQ/h
7DgX4iwSWCUY6bAAqm4IiyQRnDwxLfwiaB5FMy585iaI4BPpx843fb4hUbvkegyx
r4CuKyWBhGUkzrfqxaP8twL6I+qLQvGPPk1Auje+CPxvnHsVmpW68hKRh4NH8lCJ
Zq2bwVPEU4czwR84h15u7JhOams/O0ZL8nzMeNkRKsSXbTBaPyWNUPh/6nYJzENI
FfuWCX9Tm2PFq9P56FnQrE5WtskfmPvmqhcV2OfH+vP87WERj6mnF8LFb2HC40L8
UdCO59dRI7HEeEmDOgBbAl8woAAR5l1qKWTINzAX33GUP6VjNSUaxD5qmzi1tMYf
VpAWzfwd2vWbdQcBA4fglfUwL+VPPGlMJQm++Ua310Nmi8d+qtctebdGqRy6s1h8
ZLaTfLUZMXNsPHqcThDSaxkTFsp9I768pMjzGS1dotriVlcPgoHwDhngbeKNQZpK
prxX9pPh7HeUNf/WRb+2q/gV3HIQxyJV9aGuU01M2c4zB2bl90M0breYub27I0uD
5nicMz3r2wvKVJnySL+ahLNhll0OffuMm3WihiSm4Gq6PhDwyh2mTjuNaDo7l/zh
LtitCkpLMFtJL12S9tyCmAn6+ArVlMBgz+yDUkorH55gA6+Tnhseu6OOc1iD96Wm
55lGOKeW2ROZtnRHq/pODmpp5876F/TLS0POs902Npg33kTE+sXR/v8mWIotvJn3
An9ZLFyCvbI5z62ChZm9MIBM6wNdiWUJexn1WXQVZVtUO1FPTG/J7n+7n4T4VhJc
j5SV+WrAPcBWok62Q3MMY+qcJ25biySgoBYxsuJ6wOhwkOCHvDwFern+ZFDVJbmR
fEF8RwNN3+YNHoXkwriXskfarrwNuC6jAt2WRs8y7G340GlvgHwXb3DRn8LLzfYa
jt8c/+T4khVj+RUL1WtHYAp3hoFkvZWh/taoOOK12TZic93g2RHjBULyF/kXdsV5
Cv63H5pD1mQVE6Ow1rdwTgF4EIsCR9cTsi4EtZODChRJaYVb2gtVGplgmyLtRkf+
2t3gLnl7knU7oQVM0R+Th0tY+7Jdf/lub3wI1R8YKHCWjgmmo9nJXtMPRUtIS6r/
niiXhHgz3b9KL/14ZvKAk76ABU30jaXI2nk48COFdHG4UrGi6drseRGCR1Vf7GG2
B1i+hnd8PF26rGv9jFvzg64maG4ig8VffgMTy78D7mVpheqjdF9A6e10SmAOa8Bm
0qWLJAs/jwawRzwmDeqdg0MqrTLDrCri0Vren4yKOgpD1MmeKi0u2rHoihyv6vD8
5jgUHES9qd9EKAtHtDJ/PxV3pZnFdOzSdJuEqN6BCOmPlmyVHxM7Tu3vV888oTRj
9ubIcGGDeDCkb+6AZ/Hqpu4u6l9lF962fOBMYye2qUrD+QkWGJGEFM45LVMPyjqs
vQHBurYSllaIr1K1a33d5PBuiI4kouQj7z5dfscoX4Nj9vflCc9JlkhS7cCNpP61
RxwAP7yWlAbFsJYd0aPVDXmPf61eBx7lWrXyLUe1zzE8NwP64hgF0KgubdGFJUNc
kJ64rVwakTzPHn6rWHUTiuUg9zhktP2CFcSXIHozg7uJHiy7xLxgLgDdipzf3qG6
rI0R6EKTXe7uZTiJpzUL25vTq9VW0omwXePC/3W3ddIfQ2jEeNP/0sCrP06crsnj
t7sEvp1np+xSbkrMXLDKLbCt6Ebj/ieOJHhhz/vxXkpLiRl8VPOEWpWOa5cx7LJe
5e714mfyaOrrRxSWYuA9k1cBVkOYAcybXCJpneSygzVF0w2nMpX0OIOOM/jDIrut
SpkZCJD7gAR6uYK8r1VgSXS4jMpstqko2USmz0yTTqqx7OyXp1kSw5WlD5oyp1i6
beulQwKcPuqatRht6YtLCe36jWU9dpuLjplfRBJ7khSQ2AFI8Pz49hD2tWZjE3E7
Er3BP0TbIHDFVXg70iuu2utDS3UZ/CO6r8X7vonjmtHTz7GX7+ELFUfchKV1Q0Go
oKU3xMxZAd07DKBfX/qvfZiWIqvif//Xc5NSq6i/0S9QvMVFNLKMsBYm4YKq41ol
P8R4VEKUhDfztI+Uq+01kOA6Z+41Q3+prr3qRfANw57DDMavWbNCaYWRk3jEkhdQ
GwCeyifGBs+6JGILLeN2v+dbLQuZjtZNg3QbOcinv9+MiqN6RXKg6wOzkiJlPfIp
MpebQNKYjAFn5rzzAbjy7aj8vnkbYGhe4/rmLi741FpHENm0nz8O+26xcVbVZ81O
+Zu+/cRkvyg4k79hLgQrTP3zSJ53H3PgEUQzHrLVRK+3jydHugLC1E5/7vb0mbNb
Glxo+4QbCHWRK0dbxsz8mTz/TW+/rwS1sTF3AH+HNlJqX1LVIOr4SquAWil1jftj
B9mg53ttB9Nx957fO5wdhzc/8ZmpfOb5oY8yGNuCSxoHTI0wFgX0NZevU+fxhHJ2
Ok/8OHSfAxIIqWkvI6GuQa0ZChcbGMiZzq9ZNHpQJsgpsJKg8v/zVMgxPgyVq6iO
aAedJRxC22xZ8JJDqlurhZ/c9aqndnWaY0lYdzN6CuFeOyEJo0LFTqA4/FBD/rxx
D1PcIktmdR3CcHxrOWJiwWrydXypgIzUKOjqw0Sbua+u8cMxgH/Fxc7hsWiNEfiU
1ecmUqL9Dgjs+hzImOVTkApn3hzouIXvvk5mshY1Sgyc/PCkblCxz91OvAgnmxBb
g8f8cAKFv3jSo7pqaA9Cyr1hmQxkbLGGNxHYFupfCvlrMHpDoySW8uLJF10xY93U
mCglRPtRVToAXmX1KsOh7qx3xBSaouLdmYRvaZ47cjDxEe/x/VmEzdAjHX2fNuEh
wlbLNRuVnWr+D6F1VrfBXo+Xul4W9dZYE2jBOdc/BbMB1uczOLUlsNRxUh7cipJP
rQFE6ooEmCPgXwdBvED1m08uBPMVLv81rVJG92qeEnazRsu9gdApiEA1uo8WqdwX
QA+SwnclIaAw1dxLGeQk69Lktt4eFavmrcgHy+JU1O7UzIQMVEvL/Kv3RDnLWV58
PfvYU4VlHdmY1e+0Mg+nhYKYwjzB6tElGTwPnI/gHtBMtl7eU4w+mwx5Ycd8sIKp
LKo8CPys47kmYrQI2qimmGT0OB44FjsVNEEbMf/AXSAPvv6J9Rbo8WQ3xInNyeev
+a+XhJpxmMyPhOcergL5IUAdIry3AUBq41HJcUnDL+z+llxZvTLFgBAvioE5wjt7
M8OK68tUmQNl2qreepNCX/fVhK9XSQdXgH4RWNTGLd7eexXSPouOo7UpXgsYR31E
/HT+IMOC8RfVbjxl78g5yf5sF4JNX+/vVpJRWdSJfchz9feqdx87tU76XraU2oxp
au3PhoDnHmZzLQ5NGfcIlwnNnPqcIXf2wcCD13iEhqQYuZmzs8K39Zgd6IKJMYpb
VYzy++YGuttKI9Ki1WiA4SURVl3n+lLZ8FV/71A8hXSHFwKzb4TKiMGALtNUnQ+0
MpnVrVsZve1t+XYNiIkjqcRzOdRDxsV60aspOXraTzQ4j7wVo1pPYjH5JHHSnELW
QFFGXRP4DRtTBmICPl8syo+sUpRous0Jw3x+xsK5+fR+aC29K2u7JQBtKlUvS5tW
XASrFVJg+s3vXJoI75pM+vGSds969bXfTYMqBqhxDbg4eGbRESVtx9occC9uAaJG
xJGsJ+iaCC1B46KvFIWp//ic2oaAiE250E7AAmSl/XQGiHZfyGRZZnA3KwHwQ6XX
NY+N1EX/iUytGTTLGjS2oHFAdjH94LBDVO8aadINUb4NdiL3pB+mHUeFKSc+ywoS
GGrDiGrY41MaCmL4htTR8Je78Ax2izMLPTKFSW4Nka6T9Fw53rKADB+QdYXietFR
VFiLUsfD29hBnzezSKa7PiTkFMPmQc0eWddFoihFbZwrTOqL0Yul7OvUQdi4R2c4
Z2AsJLiM40JkE+aACe3ife/wWM9uLZxv6IwosGs27KT1oti2xW9CiAl2BTLZzK41
JWBJCnq4UH0Ag+2kNYRTFuyMI4qjIkH8/mENSJrBaDQPBzjrDWtDLAOdk14o+Unt
Q73LZD0Xbg9IDAocT1gD0Y4VoOragGveKzLzpKoj5N8A4KBRkOoKhJJ46hkhwoMI
46H4SYiFBLSspRqYd2WxfxrfTgWEMIuMLa780hzm7jo6VVkamMoeugDNe4TijX9a
NcMblKEI64CkS/4P78DVFEuc0i0Rn/vmNwuYhEn4JqpBj9OrcVHduEqwOSYT7Un3
EyuRuUwssHmx6VhCe0FfW0jcybjFMuxscqCvyfDw2W/vK0lD5pJcg2LsDb9ZH0Rt
M5jiQj5Nxinv6deD1VcwbB170UY8nRL8KlqKME46NemjLBmqxd6DYow7w2NiOr7C
50hSENb+zoPC3SioPcE9/0//p/fCeqjFXtONOI1YkeG+wGj020TM8pQ+xrs24iHN
1kdsEmlxmwADpeMJX66SiqfdiyB0ZJFzaxARugbp25rfjtt3bvsE/NL+32fH5REM
u6l4TloUdxC/dwbB/8XJ58jJKdRRWpstkkm+cmsTdX4e0YTgJpttogn8FjLYM7Zd
ObPQbGJqEXOkqFISkCPQRI4K0scdiTa9UdC4FRQ6GzB3GsdhD2HDnTOmp3WyopRm
aZMSW27+Ue8B7Z9o0pHh/cG5j9BQq9jXgz6R4rYNrKwFcrcnu8CA1EmGEehcM72g
MDgxph2gm9IOqyaVzxabtCglYBfIAnQhFl9qMeYUnf+3B7KT6ZxR5YZWkzlOOYbX
R3zqisBFyACe6eSXjBJWkj49dW2Na/i2SRLiCaeXH3htqwFsRb4Gh9zUaQoXLFt/
guNIkvk8GKxyrXtKCKWSTaSJWDDsCYBU9Whmwz/q9mCdIMJmdci1O9lGZcjZrPU6
+3rkQz5rhwrvMg9vT7s6OMabdbwvO4dXEXQXaa7gGv1vw7+Eu23Z1RkHjuo0uRao
8rP/GA9C2sAbxo5YkZm4OQKAyBi1cCZBIWSveoxMhQ0MyVIONAsH/DPZhAZCKSp+
LB7JEpc69umxgMmX/vC7Zv8Dg8vfhGvLuIzpnsZR7mUTcwaEkmmMz0PTu4/11oi4
wVdE7WhR7zFkNaj2Fid/69nPEVSXuSGwv/JYn46QMy7A1FrNZhZpnyKAWxRp8Gq2
7JT8zTD78Jo8+py9vn6mv3qFs8BZdB9Dh7q/4ymkZlxXCrzDpvbpEv1CJBpTSgq+
T+F8S7bL+GTgP+nWxUYLM5ZiYVRkqKRlgSP129b2luUqjdV0TPwUk1DBe2p4HyqJ
U9X8ty66oPo+r4gsUDo72HPbUSiEqemICsK0RVElvSIUGESH0zrG+XbHwvVXGFXD
xh2F4UYDsEkueGXYS99O5L9dduhTX+xGY1yWlvHd6dD+5YlAHdyC5Lbj1pCbvmnd
nRKnpcH/xb9INRWjn8YzDkaLuLasNhjoTbEUhBuD6vKD4aSEzlfnVWnsgtMWYgnr
82K8BJnhFa9cAS9t5q3n9CDUcvEaAkGc5n/jaquzM/S3rsaDyLmT7wOvrsaCkZIs
/oll6YE9Z/0J85C+c//YK7qe9q+FDaR8xPpSld5ShfAq2LEb25YXrJaouwoB3Y/2
1rcGUJRoHSj4EGwKoq2O+oKT65eUeC0AS1gdEwEzXBbAKofPRY+8rK4kUmnDp6H3
Xmx5ivV1ueK3bPrHtUxW0FMKdGYW4MuoxptuBnar+PhGE2VC+wLCg9wforyf3zx6
ib1sNZdbUYly797tnJKsBbJH2J32ldiqzpFp9WJ+MHG111Nl91WuNqGZsWKnugay
XdC5GbDvFv4yfZ5inX526ImXhLEpBrlJXsLfkwDhOTWOMuqoV2j3Vuivja5VIx/t
mS6utSSBQXG0/GZ6a/41vTb+fipbZwUF7vftjTzwD1ABXdkM3985jP+DqFRq1nbu
jxOvXI8dDXbf9rUo3XqAq5BCtFjst6s8728UsnmqIP528eaiq9W9qlwPtQR3VYmj
XvL7xu1aQtb6kc2ZE7owx2FNZZL9ORSsOwOvpI0Lxbz0IYe1gvpBg4yasfaL5ktl
MT+sBTDLoYW7k/pe3ZpkVvebvHCi3vVuagxzhS1JO0Lcs9RnOEWpJbXxLXU0bNbT
xtvhXPTN9Bh7myhJFRCFmPsFDOyDa9Zx5JWmHFVkbEg91ETiNcg7Czj93b2xR0eT
pzXssQpK67JU4pdr3CEGg5v6yM7JjLQz6UTg13JgvQmFeCcUNbATOH7gUh5sXHdM
CubPKHT9DpGJVMVQcY9pdUBhkwnZ9suHZCU02cClmDDvJRSe37pINC0jjS+1JM3q
0LvWG7HU5DOt7miZ8UOoEXkuDvs6wF9nQzCoeULJ1/CsTmQmL0fZ7L7tqNLxVmDs
zPeB7NcQmAVPWpGoBHCepE/+VNPyaFSpyDZA4mvbQUrk6PIrmd9fRGJPKXUf6Hug
57FsAvkJoRtNs0OYoOc/H3V8eYN415lGqfcAiM+CFOdUsw3yX2r1FZwd7gqEohZR
/tA0v5GWf4nWdiR8bNr4ZySpowsYkSPPb9haekhepQJnjzquLWCTpVFyf5qp0IuW
KgSYf2/KGvQEKrHmjuqIGE/Xd8a1rggq/pqPKGdQ4f4EUxtRg+f1mJdVjEml/bC9
SDSd73jT6EhKjKk1+mNmVjShaFmzyhN7C7kifUpmmvxkP9ZrazjvGwc2tIdoUP/Y
GtgLtetzHEZRM3IWOUfhQ+ZED6fRCuXGJ3wFxhG0xmruPVUOZknvH64T9RTHjD4X
Ub7AkhHr3MRoq8i16zOPo0mAw4lCPalQWzVB0PHspdqCHJx6RByWy58aJd54uJe6
1VQd1qPYsIoKOmoL8su7dBO61IOa2XD/JH0TzMFaWrFqisevDsSzI/h3W5J+y+RS
ue8bG6xhlh8b0C8m5fOBrAIeMhtmfv5Lek62b4vo8rRVKC6Aro1+Y5NCzoRjyre/
XCxQLhapMlelTiR88sIqGrNxSQFHXNXZcMPvUrPFE3eJE9LmiWCz+73P9DE05iPT
Ps7Rup9mDRbDpO+LMJtomDdsaZOyU6y06pGryQTPI73Sf0vp84Q0zUaLOitXfqq1
tc4SGJuz+8b1JsIUBBwhpqPIp+b8hKW5yEAkOcHizIwcZyEydIoL1xVRHHKov/zU
IyoMhsBwKPgPmT8HtLR7dDsfTL/Gi3iS9QBrbMvHyR/Pjhdsy50nUXoHfU7lyuFG
OtlZBOfrncScY8Fa9X0USQl7oPfmWIr6jxs7Oxufp4LHM6TPXzeKqtGVAuLc4EGy
J7QGuwWXTtgS8tMK+Meqtb5vZm0HDn82ub61rn48J56qGnI+sGcmSFWUSCw5/K/H
fkFwMoAc56mCnLhipD1ZbdMx/9igugey/InMKJsfYf8KXS8f5hY6blMGADK7T16N
SAsrF5DudFP0tmXU6Io2yxJlMidS0vFnPjsD7YweYjKghvIKPH9Zu3wu0ymxuGOT
WfHczKHCt/d5ZC+A6jUkhxFuCxYitjWxCoobD4LBzjbmpw8mw5tIf72Dlm7NqtXf
drojAgctABV6HespoNoGveEM7eEFvAyYhL/FR8ESTSQR83wPMDWDqR/4LM/qjMER
ZQnk/2QtWLKrpB8lAICwIPk3++syVy/y11+5h9RsIhc2ogsCygv5GrxWzeizvG/3
DICdbuyrCgvVrhdg1m9kvGzC6mql9SEqugQpq995C1glaSMC1r2RLtR9jldQUwk2
tXmpGD8hOSxu8RCAvbNtptvRjaa6q1UIRMT8QSCnTa0N4kyVVfBvZ0Kt8PB8NYwC
TTjJZA61LgQMLSJ2dYRiSYY+piwiYVJT9kngssQwyDSLGqoqSMGpzmaahF26lIWY
5ZX3xoD6B7G/IJJoXLi3KxrBj0fi/H0RJytA8cIzEhYTQcLwuX6fh08DLeU8ksdM
zqAvNxskNN7ZbBC3Bth+uATl6g7JPb7saCQGs6eQxvnriCFPZR4bumEb7EdYFAym
tz5XYLZcieVTBqxwaJv7AA8/2wnmXeYP1BSshYzYQyXPbj9uLgGyOMd7bY/tyd0E
Plwip3rReq63zWrJZH0t7CqhkoREUvxUV836QgylL7Sx1VMrrWReQhIcJ/BhlmHh
icPifcj0sjXR1BxXw36NqzJPQngjACmDsDHryxDsNK0BbeUwtTB629YoS7XUeTxJ
5Q7WzLC8oOjXI23l5WLUZ66U8U3PlCn+I86uxGl1iM8Man+7i4H3dEDskOidP0oX
ni+dJzijzGlqG3pEjBiFOA8XOMDduamxCzBDmrqamNCGYjw2B7qCJQA8hB6jpMn5
p6buJc1SSaS9png1A2vMK97POmePVxR/m4bOVal48qVxpkhMNdC0skNp0JT166aw
vwdLcdBN2iirtvaeYm+vZ3OgwuZLcRgFJCEw5cNuDei/C1VAWemQ97YmfYWasQwz
IL7XWli49s673kvf3VV5JgGQbuCsVSe/waWncdz8KM8It46cbbBkXLdbDoK+sEcG
uwQ+Mu5wvv3/jjsl+o7fJoJKGpfWrKj/Gs7HY5aQ2Om9V+B8psey6HqtUsK4gomD
ws4emuuB14kVl7WnVorHeAjDdMq5CFj6YyAWFwrUDWE9haFns/+jcV22DHUrEIKu
uGVBgJeC3U1MaqilZFimgvT/lLhbiV8AoCbRV3gyT8q91gSxF+iICQDSEyb7sMLm
AkOB/PD50eineucr4lsaLkuoXnnhkZKPKeELatYf/glUi0HxPiLeBrB4Ql1zr4P0
VD3N6dSm+M56e3JmAIPz8HsT8fhzQdCZpCQ5q12+8ILX+/sjzIhsSEqH7V02BjFq
PbvCnlHzdseAK9xFJ7QP6HXXOloD4IXINu5vZtZvrNP1fcQzfBC4d1uBE8czeg8M
8diHk9MdxDbULz2xmxh1rFV8afV60rgmWvNNOyMp79kCjOAQjhwg6JXJ0K6iiWGT
9sURtHoP00CAfpT3cZAeVkC86mC52UigMAXJOyZyyuDm3JGQfbmzRBapFYLbx+hB
wkBpLyFbKFCPepGhb22B88S4mlMfR/BqZRWZqYKcIujn8e5DdGWGGY5zFyzOpz6F
iOr0aEYrdVfRL+YtWKXhy1o0mu5hmsUb+30tgr3SfPP8K1ww0g/St3JmdUQ9cvQI
Y6aGQ20BLOFFcx8opi9vPD31IiinJTXl82sbzrbORNlWoPfvxTiTND6Drg/gvhgf
e6INRuTUgZWNjbm9LABcJMxn4YxyqXevv4MEEfdnG4P+Z1eTuTfPp2g1UVUuWz7s
wM05UaEH9Ymkth0vZipDQlg/esuCYmALJ8Fb65/YaXKfuM3nFUlceHoPcEi48N5r
gdem/bbhhwl83x5u4t6isUjz9r3kGGRciQ/Gu107VOI4CMfrdeJmtKxFTfkcRiH1
qxur0u3fSioFRw2oXn2nxE8n9pNnDfw+HWiGYaWvULj5YRdkcg9w6rJ+PAQNd3S5
PMtmwaauL3AV4577IAhpgNyCdpuFvcgZY28QP7Gm8ZpLvWW+N5TU7abLYv4R6Vn4
K3XDMG7sD4hRGxeKeYdJhGdoXkzYHxTPYsGZBXCfXn/KKEUgG3BOIEoNyqZ4opEs
/qusAdGWYajIIAXmM1TM+0vSvejBZRXUXTqubcDNyCsxZ4gOsr2Kqi82GmE1vYl7
QFwJ1Dqph7n5FHZi9ywhguwdWAK3PF4nV2vp0y4KkiGE91N4+YB14VaXJVdcmmmm
ZNthpp28pyXpMnq/7y/mXkk1zWm77s4Y7GZ2QmD6SaHsOC2F+B1Hfr6Z/ExND1D6
I66t6+5hiFDws4v5Z83GRwL04LEcZ08JpTBj8w7i+bIf5Yfo+YLkIYtRsa0aNqtn
66AHoVdHLjngCJaxhZRAxuuXqVxbwPhyyiLN3LoM2/FmCNlHKfRzBnuAMvfT9MMc
JaVSVlXCiqjfE3GpPBzu+fRJtelAI+u0IYHNPXeN5dkq0XirWGXj11VXszRewTp9
tiuYdV/qN873Y2+VhHqEaSgEuVOoZE+n5q7FzSewlxj630eZmh+uADSQLr91UxNb
j2hYFChwTVsysL6DpZvGnRaYUop8ejWGsFbDl8aSctgLiK/uaL+Oi6nw95TVCiGB
mfWca8d96TPobytE24jaBrlmZwi70vx+5Us7hrsm2QhS9BHVOg9Pm1s+hh42Nv6/
CQSn061q/Ld5HQC52zJg/2PXqKau8VqlQhL81MqdkhNDNP/ATyS7M7x0b8fcldJW
GPFdr23HbmXgI/eGNB9tg8nYGZw902r3q06WHSDCtBCEJIEN+Y8GbfBMXS4PMFve
PeAF0FhO846VeycLZf90H7GNnlRHj/vUGC5YQQYvtdmPTNN/xblum35KrsTC1+/B
5e+tuZQSCKR0NtbQl0CUmYfDSNit4dCaAvEOhvEtbBnktBH/yQGauCD3S1HuAaAq
fAk88V4+GhBZvHS5vUy22p6r7zrhtkCDLehs6d7+I+wzf4HSbpdlp9WnaLgRYrvE
JtaaK9pPD51t3R3e+9cyxaQRnhUGtuTQaUcH/KtIeCvIX/HUmxTosp2ZT2V5Lsa+
aEYo8vX+LP5s/IKjvYpPwwveZ2GzP1B6wxb62+Ogz5UbRrEnwwMJfNB7HNqNrtYx
+L+8K1F8EKW21Z5ou+cHFs1WuFRMeJ5Fb2cZktmrHHeARSZwUX79Pu3ATJX72O7A
ACHFmJDqlFDOti4qNgCaZyiPfMjb4JhEwX9ACvX43MSktzo2GTM8BsQHU4ZsNeeA
CIosHXNCjYR52pqZa4HnxqwzOqMAthYgPjN2W8PJ+ppVGq2gMbUoxNLyKPnSSPsd
bvrIowXWfkUw4pqj96VW9dUThOkuxIB98bugtA6CFkrqCe8MGjILQDChR0fz5lSI
H4MmWsOxAhYRozSKaN7l5wcaifkWnIwYgcKEGkg8V0zmpCobg80C+sBseNzHl+Mb
KrRKSRf5UeLThw2P411lCqM28BzINKSdafWOtwOalLst3eLtn55iojpZcrd/FOw3
cJ8HQtv9fryANb1ZBRxWhMkTG+19AqqYsPgr5VdwnEzoppRIKVLJXysdVIhY2iml
SOFTxhiCR73GleS3k2ZQjTZ4sUXhkZEJmuQZ4N7fqp5fpv5gtpoVd9KLQlGLg2+S
DczG9gdX6OT6s/jRCE0japYbd0+mRrR4/1anTrg2F8o9CoCMfu17D97XycyUAgme
eb+ZcCIzno+SVF/eXKlCYzQ2jXp+IFjjrLbNgKZZki07HuTaan/5IIf6PH08Yee5
Lu5TzsVunk4qc+tDmz1t4pKT6zc0zL+RpBuQfg8gIY35VIGSYxJ0TipOrKw0+5P9
3m7IB3BEKp0aTVCGmb1+irDNdG6snBoQqBa7GKyQ5gBqNSwBZfj7PbQ0rNxuDHdP
3lWRzoC6WnSldRabv7Wtyp47X4CUel5aYuAiwcj+BHmUYLRx4FI94vZO3PDZSMX8
T4caiW5AN5Cy2LrHiXxC5qhQKGncj/yngOfOnLocdPVA+/QbRcBz5j6CuNhgg8eP
8AEeZhUFjnKeWolWRwcQii2/e5VPqt4utatPTgirLOHDt7Yby8Jj4NJL3lta0vv9
l+8GRhvS8hiNpTzSawVyUge2Gf3A7PzStFzwP5pV5fKzSraqKgt7Gv9fpCNP/+UQ
mLsyQZwKWu5c/COzwQilMLHXfOIYdf/2GBQ2Vq24isiyleWxYorBBAtECDjDjqCP
uWJjc5LRsS8rm2EWLh7lPECHEhpVjU/f3m3Ga0qcPd+docyxXWp8fbTIJxOcAf/E
OOuKn0DQmb+BLA7x3UQuSTqasfMNq6Lq5TiPRoOgDNlqFOBW3jMLq0C2YTdj9qP/
Hl8uEmG5i8pDqjOk1/RQns2Ta4b09wnaoSSK51JMK8SJj/gVtr+0MZTN07AuGAEy
GGSECm/cUh3aX7sNXCb5yRvyjCXcFplRXYajfH1+78VVRVoAoexl2a+els7/Foq6
rE25N3GXJgFtMmTjQY9jwnybOqCZgEPZz4yim2vOsVL2X6SDHXeCVyM8BUXHBcPR
ed3xvdrLQs6dzUpYBGvE1Od0yjaNsOSfNNI4Sr+vkMlwMYjLhBDl38p/mZj+d9h9
GWVWIQoKT1g6HWrXlNXI6SmiAlFnZPGSOydqd8jOzqJqgioK7D7BzzF32Tq+aHsy
PdHljNhvZ2MYA+3qb49FNlbfU/9luKkeCxjYAF/BnJGzYJCPQ1qhnGnYRjfJmFJb
CW+rf39BL+5XcnQ5UlGb31ifxL8UuUCVzznqB68w+zoIRIs2ZVeAIA9sqCDE4x+x
vyEaa9WYUsKi9f8EaCxPBwAOkkC+a602sK2nlGRM/aMiOWreP7ukK1oT0Ao/2RVD
sOiXduiiZW7x4xfamAoG7/ZrW4c6hfc6KRcmGO0oZmcfOEWW+ym34XUGlYeM8W/5
rxxwyRTg67XQHmYNP8lQfgB3Psot7oYh3JnMyOykOUmaok63ZgZAUHGcp75aisUk
UN2OLWWsVI22yD0tj7abKjEaiCa0vco9c5DjkioqInvz+7wT5+HbnJyfIYLEIh3J
SvmNqm1kWG4/pYSIBRu48HsEwkS9t0zyrJJPdVc+BkCjm/3lcad0w+6PHM3HW6QG
aNFhKXMgxxYg6QxoODQnNLABoqECSCavP4rv695afqaVffrPqjpZ4lrY2C1B9gkH
QlauXU3c8RtNe8+HASuaQPFnMom6koahTIs2cUS+bXpb/z6Y33gtE3pQ3mRv34Dv
8upBYnQUOwpJV9p2bRBXUw3EJGwqd1dh2VID7ZSM40FFkxTgQEG7+uRk1EdRgeOC
Er4DmGdq3Tww2XN16CwvakkBIMxI2m2BIKCr6dl+KGE7FW0AEEVmoy01olgstmAr
ZryMx6COMbb2wixltko+OADYacvhzcqoAsvHAJEanvxcu36DWv7hcGlozia77vCK
9r1cUCwYT23VeQaqw35WfwJZiRr3XpJet6phK47mDzcVirxpf/7kTxY0OFwerTTa
GXGl8JxdSezbVzGmS85V/xLRHgpjVFirCMPbeFeEM+glDgBB70HgXiR7zKg0MPhx
AnWt70JeGKLOGYlOTTi0o/H2HRVJzFQ+sWp1Q5XIvj6L5Dn+AQyuwzPmlyfPonVB
+/T224aPiHJ1oFq8kslU5usbOiCWzQALCc95fDNM2pgCMnQuiEezYi7nbduBJerN
IRJqyHVV3tct/oXTOC72N0pSilEcu2IKzMb39o1wn379HnUWhLKw6QCTuASeGsrQ
kg5pzdVJzOXBs/LSS1HLBUosSHIJIWok4/ccY9lodo6dgzDqrVZrmRNA00eMq0jV
H/nBHjCyVEy0G7s0ovRIauGKwnBmcM6B+pF26L3smjQSITFm55aq+d0kvyNTkDKw
gv5nf2qhTJpdCrl2cOZ4/37V5sK7bXzPCZl25+zU6VZT+2rSpbSGzg5l4AuySOIs
+3CMztItnq9Tjhzd56jpovphsg0ekfNSqZSAib6rbnuHCIEvkU86cZRNVOJAlcpC
7IlW/BfturpUf6x9Cnkoo/kb9rnluVAi1kRNwx42fRfudiw4mCux/VHcrD7VZ1EP
s0O7aGXy/CMkkHJNUS9a4YivSxGSea9cEI9DUjiDMfN0+lzZAaSwqVF8tiF9S4kS
/fo9xLAv7O5HOdAUbRh8mfyFTYSSiLR0Ce8+wa12ewfRPPMw65yg5KIy7YhCF2GZ
OpyMMgnXnLC1cpbnT9+oJU909ZWI8qtWMX97Il4p/+NptOIB14XIJpIUYvWxlMhb
BKk4xgDcYMlJ+esslubwHa9vz6bqxqP8ZwIXfDGU0TikQcuRsPseIt6WH4TfnKxo
IMHqUEWyYrP2QjQf0/WGu/Jxk0nDKDEdVoQyhtsfQqfSFmdghryWgtuIHrWaqVgO
MxJd/fG+k7kpUyXKjsE1pSly1TKIrcfJGyr7SGuEQNZPgiOp5SwZWyhs0JrAPjYm
gmcnwlrw3JPvn8/ut3eCtYkisK64qfA+fLSLGkBCkm1ceN+J4jFMefYAaPzGWk9A
3BCRT3tY5Am9EtdJPTpYVz+yPtQQdoz1J9vdASBINJ5VDXbznYFeHMql3o74Y6GQ
607qqGci0JR4sjDmjRum9eQ+uCLVj8uvLYXtKq+zzmAQTfMhPzKAHsil6wG3vHJT
b6mEyidB9ITU+vgR8/iEFrfeskf0NEtmYo3HFpZ+nkyb/fRIiFcgi0ByuTCEMjzS
GCYjD149uCQ21Kbrvty+q8m3GltiHylacZT4C+57JZYF/n9P1qc0rWPduZPwp7HW
IRwsFQn7thRkxqlWzuRUDJO5Ua/SIimo6T/czdWwQWFQv4I8Qj2UQc+Q1sFGSAc3
8MJgjGXYXtbR7vQYjL1bik1dcF6x5bDEmqh6DqLn3D2SI7eNVaYSrWfzxxal1uwt
oUfECvEXrHlXsc8z5OMwpjV3xvnBkwUV935hYW/fjUf79xCqSdoYs9RzYYlrtvgs
dTlo51SL2N3m4GauuwqLgef3gMCOXxUBFHas1wBwdlN5xfw7N2JiYRLu/E27dUNT
Qpi62ePgyeCtcmoZWE8rzPg0JmRIFaNWUuVRTBTloF0RLY5RezfYcZPVzhPIK6cF
tBVaX9g8ADEI4F77xm3dFoc0LX2z1fJBEymCPNsr7dgf3WywWWjZRSesQtGN8TX6
yedKCxCj6G+tgLKIXw5Hb/o2Mknl74v/GS+dokR2sjFtrwbwoD7H7riCCfaZL74R
mse6CIcTebmOoJwZxBkrRg1Wwv0ddaIhwGT8adMM6AxgQAbxur13X54MqbRJBjmh
zVb7Aq5832/XZrnlS+t7tFc23aJDFY3h1KkaQW1lCIkUZ/Uu7qOF9X1jjWp4Bj+0
ULP4WA92X4XJmNM4SjMAN56pU11aeStqk+qkP0edQxPnkO73WinIm1tLB6ZWgPyl
OY4Qy5rz3QTVXo4i8yZrWg6w4P3GCnEZ4uUp0TvTiRssY6YrrIK1g/MIKhDX2Zd4
P2QJV4TUiO5bnPe4l7QNJHkX72trodAsrbZD6ujr1YJ7Lyjcr/nyTkuaRZLM0imv
OU6bjheOtuFCf9uwGoYnQbtepTOHHyogP1xW+PqITkwjIV/BgCGD/5nOuXjA092W
uQG2fCkie3uZfhk3xiMSjMpX5rvfLm9Qri0x69eSXqaI6Q3I3A8Q/em2hCsxnxPU
VJ8Gv1eXkQd31Aza8l3MNir0hM3qpwVoy0IXlUp79/zSP0Gso2906//oy0fYoxIr
Gn6QB5AezkPWcYw8VuU8zpkK4ka205X35tNdTZO5AzgXDIxHueHfB1F4Ixa0MqCU
Sik4sxXr0uCLCWzyZTqYhqqU7WlYnQC/r7lmXW0F/CfSEioxMeEs2rUqXVFhGX7N
qTWdB0z93hRqcfSpBmMID4ygZet73etZlYxssleP1yRMhQ3PpWRbs1h8Ys9mR/2K
OxzePlMh+Rql2fH9zAiI1jd+BW5GsUWb7IZ9Wfe9hfKwASPlyF+PUOlG7ip1AJ5z
6PDp+ffmHfcegkv5GRTengEpZEfr2oUJEJfjHU+QGMV3Km74RjMU4J2dQNt7FApS
CAvoD2G5Is5oEa6dkY9mBCkDMSRtNfl0CAsTKZ5oa2DsneBOmJavY2rS+DueNGUG
hoeWJsIbPqmEshKXG6MNgLxSSOTVmUw7gq8rX+llrjoUj3ROUgjhpWJAZFUd64fT
AaANBpAC1ZZUSMHIrEXyf+S79cWuYRn6mTZEWvX4Ad5/E8K+wJZCjutDllyGAHq2
G/EDoEToFgfP5r9DeimYcH+r3d8sXLLJKU9A9fAXpsSrwBtzuGHJskLTIxakKtYP
2ixdM5rQByeVqIXo8OIt9Uz3M9yDVYhw6dyh0FvB3c8PameGlzo8nCvVXDwp0DXc
w2T2XKD1abnYLB3PwkuYss1eacQKMQWFy3nN9swMGlGX2ATaZKnSOczx20mp05Oc
r35OKCq7ZUTy5VvbQKu9qmgXEfucYNewt5dMFhbx6bkhVfatr1/vLNK94dndNW98
dJynvHg6YQvW7SwgWjQ4zzjgc3eIZlqR9UWiIoi6rYYmtTjOGSlpwiz/fxMa2kBu
/ICrN0qPcCigKiLQTmmCSAonDlj6psDH+jlRSc0Yuc/GPnDWQ0yPCfVCMnA1t2qV
REShXjanHhG61HhthEVASJcUHSToFgcfQHDsyxahjxbbmj+KB8LlXvKH3hYxD4re
O67v3oH/yfOVR14LhsxWrzG352lKTQfg3hWOkhlcRUTWeUgLGLc0DVgfieKAvUx4
98zXLUpNYnN73WtWCNn+hfdhiFE4KuaETPA0cwj/UknWf1g0DAGthyzaCGENuw+r
+da6Ha+jfCi+VK70FIRHQtfDOQYdy2h7TS731qafZ0aFspmqNCeXmf77tCWFRjLp
yMS7N1QTVNz21MSDrXWf9QvMoTRAk4HPwjzVfRpdFyVm1fa+KPigHSaUzfteQUSu
sZIcORT7xJ5l6DJvCD4BxM8xB5TRyyjnaQ23AaLQsnms7pxffPAHhqRLRzWOO93z
J3Y0863+efqpFjXBmM3GYi0yC8XyyTxvseOU2n0KzV9W6K6u+JkN6VXA99cbr0gU
SpUGBSWDr7EvjZuCp2gY5PNmBumqgCTmSDS4iCrFlgibiGDPSE9RyJx1xRJuxPbG
xe8fbNKdtUizTzj8HHB40FLmvdoTsQI2yH0El7VI7A9l0LTI7/u4XJK5ccYgP5CN
54wPqxhnfJ/QuWokKxtHrKzo7J5X1R8O3f6pnjyttAx8s8+ALUM06fClaOeVuiF0
eB5y2VynJSabA5sw7FqjkcvRCqMwbOBO/NLzaQihS2DxUw63ZYtfcOIf6VN0p6Zc
j45HN69cuoOOwklAHX6ahNnpAgE1jxbRjcYnoIEHfZlWwPtO5aYGd6/uPg/AI8ZM
vAmNX7hKahIXLiY4WOf2ITMmpxzitPhOWRaKHFkL/NcsaYpgFjp4fshkuGh3aKkg
we9AbpNpEKJ2s7ROemXQPiWUgJd7pmLfaPIMpEXZYlHBA71T2u89b/lavRY3PJVm
+jmGuDoTn4rlU5uBbJHB+CY3YdxagKZMWPF9MZib7GF5osoXlA1O/vXKO48MW5s+
q0kD4/dy/eYCaQzU77zPs2wgaWpUx7PIT2qKA9MFeLVRqINWDPqf3bVdIAaxGwTe
rPhtWmG9KqoHcSZTOox62st9MSursWDaWVOFVXXcXK4Pc5W8jo0WB4UrnaFiDdDi
UkJ5hQtc/1D1BqR7VQ9i8VUdGbM7vhx9fpJPtUCoizU1sJQWl0ICw9h2pDzN1E7R
t0o3OkZnlu9n7ZMXMfNOtoldxwg6+ayIpyCRXEGuwwKtO04kGSxrIvYDT/7JqnYp
uRDkUAaYwnyKyL6d5N0jsk3/++yG4jqp+sxpEJLfkxFQ8ROw/OV+JyHV+Gyy7TBF
jgQ1xz8bVI9LbHIGO2XgyeAQpKFE8zuc5CbnsRfVcpZCJ/MlhLefpx5j6FaPnY2B
t3H9TvjAR7B+BXNiiFjqItjXqO14ZE6EAF4QcyPdRjS8HnBzkILSS+twmDZekqrC
zcSHgadbMc6HNfW2sjoQci/iE5evHV8n5YcVq++9xs4DPz3N4ZM5OSrwvI1nd+46
D50MlblEYvhPTOtwGVKf4nQBJZh0ngNipmVbF6oGPQPpvbvyPIcZAQUXUbh3UZdg
E63kKa+Uczp2hvSga5pNDO/YHPPcJtjBy836lBYrtClCI4aa7T5H1g3xcbZYdUOt
B3mOCH4kESp0TkjTksj/4+MsW5lyXz+HPrFipK9Evgnxt3Jm06abOV7bSW8v42uj
s4lSKM8xEEjJXzo+AsUtgv7srnTfTEIto3L/rw+SfEhRSAYNyxPq+peIx0nNgv55
s7kOAs1hqWvyrrSrphVvagJQmquXSgwT0oGx5MVHbWWeLxQE2LLJwqtRx0u0G6Sc
wgRiOvzzQsuhCQp4Gf2qZHgd5K2uMbP6+DftepjKQZt7OsXKeyqBM1v1VwDe541u
sAlvel7K1sLJaqtMkWrtBHHXszdd/9l3/HAFfYtEaHteTxup34CHhxOBTErnpkgX
DFhIcbG9L3pXdEBcVjfrs5lTsjjyovgeNSMdhY88ASLGXwTwLUb29k2LnG8i8Chv
P/hbKtZN4/oZwQj1Q5OiIn51ZodpH1XkjY9OSDqbRKcv5W5wu1RfCULeT1MvpZL8
SZMKq+kW9PIpxLlKCn+9vzmMnB8B9YfEHQO13mH5x5lBRL7FuncLuBU+oumRTeQT
fjOzO7zz6SvGvrHCEbO/R+gHUt19yJ7bdzxlv8rtHdk96MMplGSKHx8z7Jbcfpl7
5HwBiEF0mFSjiv6K753/GYYBWizY8DwcBn1xudzeu7XhB369VTX0mtzM49hpEIJT
gzc5NhT/ekTyzL9Uhvm0JE0dgCEcDj9VghTYhbtcR0NvjUX/MnQLcsC6AxEgUbgC
6qDqeARK9E343LjVUVqsliH1Kcnj74pyAD1T3DseExDq3M/BfdRsGEqF3nQVmUCx
6D0h2beRv8IfYbi8WF/h95h/g3uCgNUCXKwUnPDUCLmnFm15i8QddON1wIF1XMn+
nkgg7ODlUuZ9Dc3rB0KZJVQ5lPe40m/Y/ugUULy3w7QtU1rSUpS38DutJvsJwspi
kSO6osfuUO62+rtLxLMoKy1Z/2JEGXb/KffpucVtBo4u2UJBHAgpURD2PMNPLnLP
6xRhPoTYJ+iNNUuP9WCB3x0b8H6zbxF4RVfrPkR3bq4eWokwS3SKl7EA2D++otzG
QoLPCo1AylEtFploMv5lR1ymiQU4pXhIN6AU9KiySwJj0ojd+8pNTBKgaymJg9JW
eHDwUxaOKJT69IXWaBYUbb7vkuvY1ruK2NMsp7yrK4LrS3ScsyttvlggJbCk6jLd
YCA2oL4MBl1lGJLSvNBTmqPJjktSjlTmvIqRwO751zof7V8c+2riLf/F8QIMFBbu
WwtCY1YMZ3C1QIWMxCOslGl5q9cuW8KMAgX9Tp+nIn4aaNHLx04wN73leCXI1s4K
fijf4VbUdcMGgTEH1sEjpzrnaim3xcDPgrUMnApJ5y8hwZC4h24ZaufClJv/3mOc
3mKzHfYUGifVeQuWE2BNeB+ADr6z8ODXsG3RXzVHKm3gsn6R9F1GgOfEReBwFkXJ
NzLFswJfeW7tb9ZKPha6DOCKnU/XYTkPQv0TtgLJc7rbDyH9GpzV3R4mPJB8PIO9
FF88/TxjKnpldcqS4vNDe/LUMJsELeEtSFCIOD40WUolZkf3F+hc6JDVg38WI9Me
HUoQjjNJaa+R5OOKuXZh62sZ/HQ0UkNdrLbKrqn2EuhkndRmtTQ1uj2iVqVB8e6L
GdS3kAUbJZ/eWXEifJIeSaZzljWWaCmlqt+jlLWWFeke6c9Lyw2uz+r7PSumL/Hz
MpmYPrUX1Xu/v/WO+Ela8GUlWb/D5GbwAxNJnOnHfZK0XJW4EPiFixRpAyepfiD8
hdHFgaCF6vIxXo1votZmM8+OzZ02lW6unSR378Nuk+Ccw3hZPVpON8KMBBq5kWfA
sRmPsy9wmhxHc1Zqd8+h10TS56v9EMX93IPN+P/uE3NFsdTvtKVs3uXMsKlo2Sul
8oq/co2ClV9PkCRq8hApN7eqQPsT/7LPRKAcU7DU15YU/gnt9EOCePMDkZeXgZb/
odA7DxcBHmC1420aHH7rFK4psjaLoUg2b+PK2tCkCkmNqkj4AfCxlhhgLjA/LbaL
j8LjLGJ3/otaR2nQjzQHLthzZtrB495DNx31X8OalnnV20+wruG2LOCloEt7VYDb
JJlVD+AWzgrzZOPFZbub73WdEa9IMeCRPyFG+cNFXMllKmXAvjO4mdvrUHYhqD5A
2v+QnoNXZ0jnmmK51Jl6akarmN0FTwYMah0rA+3rg1yZuQyQCcRvHIgrVTVN3mmG
5jst0ctsT5bMrF9S4DkqSt0G2cLb2XaKrOOgmRcmJn2y1ni0Gc0H0GOj+7SQhXYX
+JIhhZuSe5vB6d6WeoenCHzcm+Shgqfl8w19Rp1yfzU4HaskCFaafXYp8LGB4+qr
aeeRSxkSavGVFsfUlp1u8HgsjxlV+xQ1maC9Itrry7gsJNSB4244gqUftCp4K6su
07kmrcfO8Qgcl+UpztpDLMzllpRSqzK2ukgk9kk4tHEhYnZrRgQt+3sIKnv1qTIr
XC5id+BnNF/wV1nXUGCxup7PE/joQbyWrOt2DT83efSCAya2pQzUn9LRn2Axlqn4
VhHa4WLy5qI1SOsX9AA4uyDKioS6NoYeoQXd02trU7fAP4nPow8YvOslV7Zk95Xr
l/jV8p0rQcbkn8aoKOP/iLPRzMS4lAPpUBMuC3gkBu/LJPU71t9znqG7gNk4z9+4
SDHFxIJ90pw+lEHh7WlgN8mCN47HWRsh7F1/HYK4D0bklsLtaI4L5cHKGY4ginNE
swNPVhgosJXzq/QkRsVDANhhi/7JH9V3Fe0zKq5p1ELcdcuf0cprhPKl5bh8fCzp
ikPzFXlT14DD1mbUM3uPrz4oXAojd3T3GQ479HXzCOLJB+2iT/vEfrZUrWKkEomH
4ipsSJqdSrx7DpuLc+FQcabZ2zVdOB30BxGglUu+xiqyTVNg+ka2kXRg4tJWX1SL
pI14hWBAfQxLZF8SlkHI7Z1qCHV8WQo9zGolEiJt/gj14iCQjh6OcBxeGSkoTK27
1MpheFPgwQcq8vQxFW4vuR3l68z+F3lv5tN5EnFYusu1k9drxa91AH3xR2Ewj+iw
hEdGB175vPVaY/dF3FrMOXFHvjX5z6JpHE8ZGSnuppx/Z9CJl2a/5vCPcClf6SxX
tvrQL1cdr+qk8ZVGF/IvFkD8D0KjITMEF05sV7yPkXk0DtzN5a8qasnvmNtlgTM9
FDsDdxsKbJgOJMtqz6r/9/QYSH8ZuRabOx2M/gKx1CfKyQaK4FIKVnMh1W4oEaox
26z/zRM+VWrWLNnQTOfFpv3w9+RzNFdMfDbWWAn86ojjH0xTYuf54n9M6Cg2/oJP
HQYVOb3AHNOkUjx/X/UnrGxB0EM2qozp8hbQn7ZKXpGnHOMgVkCc/PzZgQ0/j5cL
9rOmgfsiznj01brFvS12x8AxKF6DIZ6qdOFSaHucQzjXqgGs8Wwdfvuz8zVdPPib
YYGMps2dTVeWBGQ4wVl02U1TYRZK5b8Pi9FXmhVuASI+GLx+VGFw3Aa2JyJxOsCv
X6JdKeBVQGmvIa4HT5/HppDn7SX0LtEHRflk9FkjAtZzen45Lir8GAZs2X9GFxiD
wBmrstSxTKteI2ZjEoK6bhrCFUSdhiG8pvVSx+VXxtiJS8mohii7zrZmJ9nkAvMJ
j7Zz+OHzUiFx5htQG5jUSlg/gR9Ky3et7J3pkeQhTLkUJcgDtseVl8sHMCoP6kqO
Fpz0xzmLQu1x6sWgrFf5SjdqBVw3VPm00Rm0IIMFavykPEwdyLDLJICWbZsy/1Wi
kgqE1oSOzEeVFD9tgA0oWdl6bqdC3bqcyuFhxDgXZpwMqP89QfSKj92hP+AvieAI
aYZyEyTeyQ3xttSXse2rl2E8YZvB9gNvYLxE/o99wpxW+FB63ncUFyfd4aU/pph6
yY/T6oJ86FeeZLcR0H31BqHc3ny5S+3brilLeYPq5Tcg2eQW98BP8CFPsh2iWS7H
YkR3HHKgwv0lBZ4GsngJFTYbXVgpsrAT1eCUAR7JZykUmRFHQhX+n50JZMlBowhD
/hJ1+501VyqktKCbOj91+ewRFaD20B1D5AZuNXjQl6ARGLjWRcxnlLytfa8erWLj
0AJIIJAlDrGKayVxRQHc+gBj/6CGCxPFEHiJqsdKjrn7pfBBTYE8//FW51tIbi5c
Yi9bikL4lBQC0NYLJR6Av/g1WpKGagrEN9SB/Ro+IsDqpkID5cgkqhZU3wp1D40E
7HDiJzVIZlcD6855DrV8ebY9j+H1a+GKsH9BaaIemgF4+rKz2es8Oj4+RnKk0TeV
CY2KmBQND3rvkme0YAOgEA1oY+aZcYUPuTNWsNOZv7C7+XpVmnzDXGI4yUlfk9G0
Gpf2RbG4VqPevKecBsSLnhCjFu3Nl95AwU6qAoLbvKwDy58tQtwR9NSGV+pcc9QR
WvYtzHs7bJqpI/wuHnc27sntPJa64oIzteUUe7jh+J6X/3bRD3ZAv255HLHcA4xv
aJbOHycO55AZFCVjsn73TALYVpxfYUzVyyrczhxX1KxG1/04hhKPNb/ljpnhOTd2
/SrbGZPD4RbMn/bk3uSdZ+J/SUaBAD/5aX71pQwX9cQxG8HTTkj+yan1eBrF0WEO
qrBRanGkpQWxRPwP7KOmaesLJ/MDhX5bV7RbecLvfsGK6JZBjANTYlfWYuLShNge
YBeWSOeuU0q4Yp+7y+TTxAbx24YjK5XJ5LNxmRNW9UWMaimq8qjsfjimDzP7Y6BW
HMth/IsepMvLV0Gmqu1bLHe53pBN4HM6WCGK7Am9bEEiIb0sdMLpnFiwGPmoGplc
1EHzB3uAwaYyXozgUWxGWsldNKhSk0jxBHzyhaWhJYsV9GV4fD2lVSZPGmUyRDKb
mblwTdyblpcUOQWrxz6o7JE0BwGJaHzw7vigm05AW/89HbLV7fbCIrjnUCIExSFd
CQ1FlOIZFpaGm76PKnx1KJGlK1N+PDupDtSR80ufZ8dN/U2HuUuF2DEHPt2iJP3W
NBJRRfSaZRWTASp1bAgXLalksplBdCa6RbvUlHYi82+8aP7F9I1ngIleCcli3dHa
R7ltZ7qZEtY71h5CB1EjZFdtCOlwO+l3bC4gUh8OHj0dgJsvRsQwhM4kYfnIyEpN
ez/0ovkFGJx6RUR8nDU6K0JO2QhAZv9/2TSSV7rBeOemKUC6quJ/cC1v4hQQkbMs
r1Jk1nSUA8O3NMQ1S41rMZfPClA2x+4JcZzfDty0BtvMSNYzFcryUwki+/EGCau7
7oznFv1xbcJeIp9J0gy7jagVGI59ix6E2kzKyYuZr5ryVh4xCGPOMG0rrxUSL0RF
mkEw0dhqHv9cq0oFETRO8t/fL9ede8igLF3K7JMe6tZX9w0NtAlyEhmyO0nCtaAq
hn+BXKDHkNqZ5CYaSoo6FkEdaBAH90ernigeY1y0+pwo3riFMbY5PCZugFSdWhV8
f20ywfZ5Gf8W/OW4sIiaj6OmzqeW/phcO24wUpxcn0pyDNXmVxellggnfZEFilBH
2osD0iOl1aoA+twW+vokMtlwuWTFksk7k6Ob/sPIlVhl/KjzTpO1yTufdeT+Sy/n
Y2rMPy1kgtnb0/ME3zMoSDbPbVHHP2oT9Vg9Ou60gmvHDxoEmInEDDPoGGTpWuPc
3w8KjYkH1j9PhUrAo44V6oLlb6WjkSfIcScpSNb4oBzp2WahpDSWd9KL9lPWiBZd
oHNJLDB/IgYNRr6TriWiCVy5p7uuctqdMIhRqAOWZjCy2pzcKKZ7ByafYdO/5hG8
KxBseXYdkziEz1cITugs/4pihjzv3PmxgqSoh8avjtQMX9iE+6dWQFVLSER94KQx
JkV7Az4XOKGdNzsqSaPg4Jz27zrnprp1HFmMXKSYKeChZgcClIGUqcB1p6uW2EtZ
onPNamNSHWRigbAz8GN7JtMgxYg1ELk2odTQvccyh88o/6obXUUGkSZYGhm9aA7N
fc17W97I25Hmq9eBVx97cKRLyrteXZCd5gV9oeqv5PhDy00EABQEEEn1kVZdyOFZ
AuFJJAakJkXMxF8DiiED9y7SXn6treX55xkl/L68InQrUCiQSa+k/P+HIE0Sg0o+
iiR1ZTIROPxvYGtkibS2wjEvEGUpnpv0dagvvvAmJIaz3eTX4GKJxmA3+vhzx7wr
rQw56+kYr4MZoNgSDbDqjn/SCVmNYrEa9+YumaKECYbgnfKEEK28oJzPlYdQuGTD
IrR8UroL51tPRVSYOnUI+RVH9OfVujpVUDE38WKvu8xmmUNooUeLo8y+qSiqtulh
bOi2Lmllre/pL4YtUm9X5UjAggGZlcan9/aSjWNn13RGgKyrDUrGDOIkqWkebJ7f
a4YT9r9ItLU6/KWxgHOy1tCoEy7+orIBhgEvW1eXopvzXY83XxED93UvRanyQ3pa
t2LNy2qqruSuqTGXWl7C4Yr8mZGmYLZxorRlsf8kwuChC8EzcjJ1vtAZEvE6g1T7
mqLoywZKRa/xBFeTCV9fU9uCByDDexPKcDrz/GviQOK0tKtMch05v2biulOf+V1D
UXX+rr8lNbWPYRVWYG3Oj1GFAGE7I3xt4IuYv9CNO/VXyBRANMCMQGdpF8N9iupK
loeM9KADJABpUNbaaH3NKdGtJnhBcCMQJVRx37kkfmIROmEVXwETnGz9mchkLHKh
2JTPiIOb5Hi4Pcn41lpfCGn9SsKNcxM0xxnDjwFnkFaaxdnalhMf4R7+zLBIiYwD
HGpQD9EzrhRqCKqMxO26cUnOm/SUChtZOoh9hRp2DrK5WmXvlm9EeyRXYxZC728D
V/fwEznwlQfAKONO4EFReVWnFCkt75hvwhCsUTv99XGBjAham9lbY9s/8jl4gKt7
3WA2cGGy4amVm7+CHDvU7By3aP4C0H5PDexfSr350+MBVCcRQ7u3O9HEx+F/X3oW
Jp+DV0rpFL+HnMxB+f7Uw8f2MqO7dPQdgcX8/3lquoR8y4aezgssGu6fdm6oqejk
QafD5zlOV84K2uUM2McGMMOi633h7UEI4IPI6aSDK9iMG6AqEy+6nhF6GumPtFGX
yTuS9+aQHRGDXsnB1lC10+Tago38KFsjz78O0Pqij65DF7jXFXRUmj8pTe9Djtf0
djEDme2zKMdNuNXuGvvg//KHrgoCEQwVmpQboUPBQ8PZACUnIEmS/xTL1bKt8hMJ
ELUkopahIJpHkFyWV55rT5N5xsNU1b0f9/CphVzFvv8cJdH3ocxmUrNhykFZmCez
XqGmOvWtaRwYPbRvyG2StILMX2usvqkmK1GvoN9XGd7wQzfvFKPE6u66FIxtBbtO
6lKvTdFvYs0XchiuW1KTvM5biNhN1u7DBqavjdfIer1pRzSqN3JJrEKQcULZAixZ
pnP9lYF15TZzDNbfrSqducm21U6GmvbU87GZTp5BX2QuuCNPfbScomM33DxZp8UD
oBizXG5sLQp3zpdhPhs3D1vqFa5x+6+MOn+rWilwSXaRJQWbfbA6otAP+m2Am7Mj
lrTHh6emxuY46zvF4FFb2UTSLSGCMDlrnRNjPwHUKQfV3UQRP9Az0z71B/7PoVMs
CfSfu+5/RHLBUVzDQ/yo02MQBZHrg8Yw5sCwfVeUZ6ZrkEDYqfOi6j4rPFOfrfIt
1jpshZNOxq4Jf/xgVJQtH7jCPGi2/69Kr9gHcVsFMaFu/A4N3YEjDpFz2u/wUyXC
yvF3GmJZsoo1ufeFqilNVyxX1JDU0trfBkITVyJM361+4iICGVNz8Pl2xalsPReA
abqvbdHciSsChJSYBtai49xVp45Ol3YnWi7PI8yna2DRsjMk+tdxU1zyinzuMhwR
3oEoZbD3Oz1DskxH9/7KdNql0f4f1kmYmJK/WkQLC0RVLwFNkCqFRKGCF3Xtxo3F
LPK8E98wJI7aE92i9DFoBqUfLVIS7aOxecsXB4xy6u4nI+9Iv2g7Js0U0hXlE7VC
//NSiLBsuSCN0ZhSj7ma9XSZPFlr1Zh4x4dAcVgRYMMN/Ai/5xOIXUOIg4YgBNIs
UypE0tZE8f6Uzzsnn3jAmJYsSKc9gQjhyJVxK31aZ/fmnx/pWuOwMlEsgGa2z5Hy
TBCPLXZdREQunmbh4VCst4mmNAfmJROD95+ARyqIr1/vmZywQgN0d4zWw5F+809R
PcIxKk8G4hcn6OD3IQZqg9qhlLOgbW7i7wMOW3qaY7wpQlksD9E+4YFAB446ih8n
AYHF7+9GMjNAxO9Bomw50+TvM/CGAZ0y9LYOEa+R/EIjZFZsEMhGruW02+sQWKHL
5OQiu5DlV8HIzoVCWxvZatoTPVsbd1RK24VROBKI3+FsGTljTfdLFClSEKYIx7hQ
YFMS0qoxcA5D9HNYlD3tJLVurE/GV/AWgIAxX9dW8Aq6nvT3swaOjdDbi7HLBiBw
940uiJshuKf2nyDZSYbs/Ulv9SDHlxfc5jHWcc9a6Q0C6nFHIhstCrAIYctNhDMW
sfwsGmyHd9W7vFzqmGK2zIUcs78MWVfN1JiQ6g6g2qMwvC4aUryHv4JZtTjC3rvp
XaSswkpL8RKwap7JTrHOLbH24PtjwmfvX/UKK4h/mYbaOYzkjxl09C+cPhUgbaoL
kBMMb0x3zB/s5FonrkhAsCSwhFrW8Acv5aott8TEYrsBg8mxy9hrNcDRZJKUXmqL
erfoVeiz284CKUYPQltJI6pG5rgHJ4obpHTwCWXBVrwz7uMtEFdNZQGkCDSHVHt1
w2RhPVQ0lmTn2FxCSxGevy7SSUaRqHBG6I5+WXMnjcp4WWG0t7/MNyzty3s+LREW
Y/QAUN9mZ3xbnYQoMfEf2uuJKTGd47pvP/lPJDeelcCH9Xg47SCGjmhK9nUMHiIG
y6c0PBjdoRbsWvWdjP5lSWGr3E83OZxgzGiXka8YvGBoKpLWVqveODushQVxG8JG
zbZo2zjdI4ArZlvTf7i2hUU2qC2kJ4zW+lCDt58Pjj4ltW92g8WwNOOxR9uaIWaN
FFi+2tA1qi8YAHdU23CETBzd+AS6glKqSxOC/GKmi73In4weEFSOKYqqF7CfHZVt
sN30//SHygF8NXNQvQisVbxPpmHyC5Zjdf7b6CiY6LPtteABKzhRjC/yEKjzxZIB
tysDa2/tYnv/j8nZD/j1ZGRXukQghg/Lx/4/axaCAEV0HOnkV2WLjLKHCQeMhKli
6GMlzm8BZUFsTulRJyljEGnG1GmJlgBBRFoQbOcrQOpLosdsKhf3WKT8aqaTHkVc
d+JGvYHzZrqhKn1RHJc0o5MT3HbedpWIZZYATKWAb6T/BPIXZe6ojzTO3nqe5DPd
J7b6KGpdt5wr92AAVjs7eAUTs9Fb8n9wxo2fuk4h79Lm5jn8JEgQRg0qhPDDYaRG
5DqutKpDhk98ELKOt7fh2mN3hQCnq051DegoMTLAo/LAEi6aws8RLZxJskbbyVon
sgWQHGkJaMSDNuf7Ad4zO3a3cPwrEsM4GxjIxxz5yFCqiCH7uxf0UHCJf+CzPETa
HUUWajHtNliU5WoNQmtLvGCdF2Tfcnk/GCnrPvsQ4HXflPNqtK0PeEXFwlzIyTkP
KAclLq/oS4LPDcvVKh4eLHZCHF/hlbZXBgEzDZEb4V8kmrC3gEoqTJNokfFDQhiw
/WN7WgLGH0DqfO3GBPTtCZgHv14/bsVmAIlUjoZIDPdTNjzvxhlvkffbvzWjQs5v
iIk6Jr+GFCPfRUY9R4BD/PkRO089OIyzWLvkorbxF4gOEvU4GjfQJWvI6dAb54lJ
VSimexT4KPOvwUFsiPO9Xj3sKUFHKraikmr0y5qkjseMvVMO7gkWGFkEd+PsJCNf
GnoAjvYwDfXzybMOw5o+lcGUXFHN1FTHdLEZkqOaBhXuCUIxV0c0QQN6vgjpLNlV
BdblEBXSJ2PEl/w+/kvG/IsSJByfiMJSwVTWXEEkUQqQPMp2ElBq86yOq0J40LiS
gKJ/+SHb+hYgV3qZn6OS9yHFUN2IN89tQxS3t0vVqN7egojN5EDliuNU7JMd03In
mIFChzLE2uT0G7rjaZTUPWF+LsxXXiUVQGWBo2tmSAPzJzi/TCw5QKUdquFQGT6I
GPiQ0OPU2a3E3lbAuZYJeBfh4SRlDm+XI2FUWmL63K9d1CUcyab2wnNKO7dc9VcI
YGMdUwmWTRr9w7l222h2lwwz9dr78JpZdvpqRn9I0dbSO+OilxtJwSXk9CV0EpMF
muH4qjQBIZCm52qaBquu5rqaWHrwjjVHfbg0wxZ+MJ5vQ7k87AVAelAT5WhE4FX9
ByFUQwfmSiz5RoGTEwKAGrVzyDr5wF2L3hnMaWYvqt64ZEyIMVdgn0mhPYTaAkyf
6T20n55IyXeyKXmVacm7QHgL8IbZHSNMdmWIfMg+zhJ+RFmQDbkGdzhEzoAiPe30
OpWbCAxCPIhAEBqHImSb9XrKwmvrCpm882Llwo1rMB5Tso8qU3ztMJednMgRtokZ
q9+Sk9uNIY+wkqizHxvgXzwGbBy5p3bJqdbyYCnsZ8DkyCw12cVrTS7jEGXtb95Q
kUD4wKNGHAidSn4GlMkYLt/pcqV42bw2PZKoAlcfR3lBww4jrZTpToi52NlIidem
wOdQX8/WxzoiF3lTGlljL9fRM/5uGIIxMh8zgGF62X2EJxN3ah4dVUDxzWBZLhfh
Ncah/OAHErtwN1Hp4Hy+uzpQzFCQUpQVojzU9YZgSPIlU9hq5es/uFK1YcYpkuZQ
TO2jBAS2vptp/0cbulCuemrpNS7eQmVFR/AtXPiCjde0aiLSGvf10up/leEdstco
uMAHyapa+CPx2v7TnYqBfRzAXrs2p2RkFc3h121rPPGOfk6PUsfhlyhT9ZZ4bsL7
wSP2REQe5rwehreVPW716JB04zYnSHggwK36Yj3irbOEuTjRbkkl1PIhKM6xarrV
nyWCu3e45phipuTYewKBu8Gkyn9JNesnM/x7jZs7P3vJQv6BorAYfdM22mqdJBWp
P6NvsvtUjJRt5XDVt58Zf+FK1Rf2NUgkWGjHwChhTiDh4PXwU57XM2B0JvoY1cqx
yFJLBFwpWNXt1lhr7n+QL2j0CNWgAyuVv0zRaHNMyXE1vgWC5ArpJ7eqVNWsM9JJ
8YADH5mtWf2HgF0qwmEv0h+KfopoWxVtpQIszm1b3lczBTss7KO56jr8FJ1U3P9Y
dwaBbV4Q890Fmz3IHnjun1VzOa5hUzgEj9z14Pwo7mH1N73StHXbsvx4TlVVQ2cF
WwX4J0+LAHX325EuuDMW3FQIhgIh6bLzQhReRJltrdmP51qc0BQ/Gz4NxW/pRp2u
tGQy6Cb/dGZEg9At9+UASZppbVLmuyBRFgxzGQWF95dXsfRu/uZSJmx0/3WXkf/R
HIXXorf5A4EIO3v2glGxRd347OIFlaDJkDhmmub3f/WMTTAYAweemu4TBOnTgW9J
Pg1WnmkzokHg0pUDaGJ34pK2pJA/DMxswpEhm02WswRXKXOr0AkKrxxga6jt1/UW
Y4Nb9skJoseYLqtlVWjH3ine027K+cCZ9fnn6tnntU3D4menx4eIo3ydrRnbu7rP
OvumPUrlDgOMeoXntMwgRVu105d3YP8en3huUIi2FeUo3EbM/FslWWZ3+SI2xYvL
wVaNKBf7sqVIdBo3j34uFPi7hBRjKpGwrNzXjnRM86adcdoDqH/6nFj35SPfhy5N
t9h5z9OwEdIlgyCHUCWUc7+UWmdoupZFg3OGHsuK7M1tvc6tDKPTcxjkQ9RXR0r0
aSQVlMNiAH02GtUAyx+K4GiDAr3Uu3fPmQhKgssnlY01us+zWfZnUHv6B1xHeqDj
RQQQuP7NC7X3Npr8k+0HTAiPMdiiXAIttWtN61nZaxJ+/0eLwlSJWDU8mzT4gA8I
dy86v5FrqiqXRWdWe97MikJTov24TQZryINr609Dt4a4WfGyJbErY5Ho03GOiUe7
Bs9OwLyBXjtHxT58uJZl6WYaY6fg489+0JlxObanu3mSp5RmZ5jplfkjSqoWUNRr
5eoVFGZbWGuBHsveZwR+27ORMQ3j6zeBXMkO/xa0lfil6/vMX0wPJEzeMDnw2oQt
7MhSlZcgpKQwwkx4YEvyigvGVqoDMrsB2bMBGDsRFjr2DmLRAySHQ2FX/CI3MoGY
z/y6A10GGvavgcjg4ynx6iMReWwA0m+pEaxAFnCyfCmwhaQ4YxwoIHKAu7x53OqB
BJUTEx7OaaaN/sFCNn08kiaVj8QHpQ3HUvtPAgDSV8OpDkHgnKpngzI99YJQlwPB
Ta0Vo1fT5lq3TlL/9h+d0H1wySI4MeNSb1aZ3qwSuvQ9jZ3GiHOBzIwRBEvPmhcD
x5ps5SYfbbfaeMkNGtvc5nAeJKWeSxC9C2B6L9BvGBWnP1rXHHODeSmbVxRpkMM7
8fvbs3CJm+/s9gTd13hbh6EaIQ2Z+6PhyET83hFxX7YKtpvMEIkI+CjcHA2XYSCP
S5ZFG6OHfE+tvBzZQP3eFJufEdPW+AENRchLdGOGVGJMLbomVLVtJN0xn7vkEINj
L2VQl9ntsFcAT/YgvUUZNs4sw+suEvr7zNN81xmpF5frnyAXjVxfj/Ngm7FeuOSx
u/K7aiPCq4pLNd7Xwkdr863O6FaZX9dUkvBqDdM41BQWSv/XdEjENmLFSrXUQZyh
zg07BEXUCcy1LcHP9QOlJxyXcdoYCe7UTMFqH+r/YVE63xEWyuA5Kokldoein6yw
SupgQhhf3rlmw39Z39upmCE2EzXeuLJUCp2Vwmg1Ie++h1OpdlMEyiZhC5me3bjV
oRpSDSHDbRmnY02IpeOFSWIIvvNeM+gE0EWYTygXFlxEd4faOLpimbLalV5a0Lml
T5i2CAcRq8ie8WMNipKU6nNo50zx84hat3rpcl6ro5VY6jStTSFdrXOB69e84dMz
PwjlyNTN4yBTJRbRCJKiZJ4HETYLhzaUovC/FJSYHp/QSyVZ1tsXflWKN9p+SfTD
NKfdIo/OU9v9E7RuwGn6EQa8IWvdM5RPIivo+xXf2aX7kf5cE295IMPtrgTZDPpK
BsFBfJwI98Q2io2ytkK+Cj5ql17PmLQ/r6AaMeYpZ3zF/aggH6FPpZavs4lt6jP8
/R4gX6Jl8gVDRm7ZXZqUR2Xk8/Bx1wmsVX9uGapno7xLTXcLG+qcwqWDuMCOlJvk
LiJfjuHqoLw1Cy48c2v7Z5dteWzdSIulMn81JHBH/3Rbosilma6JOgeaRPU9xDoi
DWDC/TnYreNAtEPXfh9wsqOGkowqAlSD/e+hG5ZKP2jZ8kt4uPleAVGh+tDzuzX2
JK6NWc6fpsgxg7W6SWM2M0mgNbyarH6wo0KipGaCggKx8Wi8nhB+fYJ828gSwa7w
2yNL5v/rHndceydWRdtCJrc3NCAY+VklUmZAw5ouw7Tv+6o7EgkMbSxwxRW5Qf0d
SQ6wIS1+qyifB7KAdgO4t8lUXaUpJdKXr8E2vzcpHdn5oOKQ1HNDLUJ4sWxwEhJD
7K8pkhR2Ebvvfx9r9OrhxBK7Pos5vvWJJpRq9plBTGsAJcVAih3iqQojheoiR8Y4
7BEjs67toL13invMyO7BdOweffbEx8sfsWza3JvLNY+BDUPkm4BKB7ZuIpzvXjw6
brKtycodtUhyE3MRpisKuV7X6Ufn0qvfJdLc7KZyFfTH/lZirsQ9fjSBaw2qK7Wt
t5FNOQJF8ghSe928RzbiUQFwGbfeSVV9UCAsDBFnNDJrYI36NLc396d2B0gtGERe
k/eT01MD71BTBJRRwK7zWOr/aW98Ny/yiXf61rVCbb8fZrBXn8948HWDe69EaJdW
fvpg73J2A2OUfigc/6mijdFEhBFmlLBt9ve6YWwOWLt04Q4USmZUCJdaS8ptNJpP
rZbjmdZu+6tTaJJBGWdezfF0idfGatItmI4td9r4QBIbmZaDgkzV8E3/cvTFs+MF
+mK6hd5uN6q55jKmQlWYtOl0Kv1y0v16LpFLW8mDSwizYQvfVGv5U+pT0cdYexw0
rgSj8k1Nr9Lacnm5MZTxjVx/iTOi6Z4HdVzEwqZAw/VwlYLgIjS1IFLG4ZDv2ngZ
YeUwy9ur5TTyYFZZle0D6WP0xOJ2bS5o4VQEJWcJ3h5EF7Tj/fAodri/DcvUHmTL
9isioFfw8G2LBRvasIQJbTQbPdB0OMgeFJynOcwc7Rc/u7MisZcia2XwkpGzHlJg
jqfT7xkqI67zLFuK1d8mcl5DBRfSeRsHJ1jmPncx7cIRyhhX3jxc8RgEeIbkCIoQ
3iZ7oH8qk0z808pm2jkCslyt5bIc2h57pWlgXu3XvSSgKbp7191STX6sVyaCTkCc
6owVYLtR4chqRkAxTDgoJtdPkTbnpv6yDkhCCFrhC92yHvy2OSyGhfn8gYtb3gwS
6ddZZH5gJNsJwIV4ihE1+TTquuDfHjDSHfrrBiZXE3E3WWW5f0ON2wERNvuy3COL
EGdbz8zpeaM+JKldX8o6twhfBuZd9rN2JgY99jtQpW/5YsR+QlGoSkd8q24oKlvE
bUUcaHmL1RTSDXZRFWvo9Zbv7Us6ZJBUeEVJ9G1YhAQ2sQ1SNKxop51Z8U8ULWAZ
W9jPUf75/pHMCzVxKuy7qFIlKhG41BFNiE5ps4nrh+xmnMvAzVMKhI7CDDBnh9Wv
2zokR2bbyhhmpqow1rLU70HmFgofVTnoVtknuvih8L7lW3OVuptQ084st98zFI2V
O9y4NQZAazGVNoxY1SJJIjztohhwNkEgHqg1e9/WPa5LVVyowndekyWT2WhGLaGn
jWouEisEKdC52vtRYYPewu7TvcxVRm9yNaRiKcRc8Isq5PpXU1jqV9CdL2audDFv
dnEorjY9nBOlLLKbnSvc/QQJfEhXppKR5Bk9SzI+Ud3kaKAwy+5pVFXO7ykGa7Mz
S/AHn3ips5nsd9KMdnDM2XF5VVCFYLy1MZFGE3woE4nqydOxU+zLEfPluCVI+Hds
AI0lX7RtAXX6LJZ4naa0feROGEIlt0PwEDto78O+YF9sszNIgPAGMJ6+7QQE71lQ
b1h/I6axZlwOVt3gB5ydGT1xCGznYbFIGxJLQfMY2yOR3mIBKs/ImDaMzTQS/Uk/
dGTTzWA9h+kDUzZJUdRzy8mOibR3qbVIIpAOVEq9G9NvMOK/UOnhP9Iht0/u+q40
sDfbV69JRw3dQYMMCyRVqVaJwzYPJzJ2WFGZl9re1bg++PFlh4m23W9Pos2G7W1H
ziF59ComsFeKomW+IUUyOo18TKniR2mvHq1igfmGlKhyKa7+DwcEIe+Hk+o7FHpg
KDAbg5pMl/MyWsLJqr73JTl+ucFCccuKzwzN8w+Cc18Y3Io14uej2zC9H1fQhPYF
G8BUskskIR++lOkj2KbTE7jUeWZpZ5bo6TVUQnvi6FC3D/tRdHOD3zk7KWstUIA9
N6aZUpAnmHz3jQvxl91QU2UE/vwceEYAlJgrxd2ZdTfD0kqYaYonem3JmFT86xOO
G6tGshKE8B3J+ZFjkAX/WPkjRXTIHeXaVywuqx6i7ilktY1GUpLp0Lo2SPTq78EN
wcUD6LHhAjZigxLGSH8xXLNbpxf770BSBmZf1rIRRP50hhatq/8jtygkJR7+arLg
U2ebHVKHA5M58yybmT+iBgKOeCT5tgc4/Tf6ZG21JqOxPei+MrJEKqLXSCCjVUie
CY3ub2SihGVCsfBZgia3xaW+ieCdv+uId888E6WEsslHqqNCDKh57pLIixlgaIlB
RQLttjjG8eHD6XmfrYfhvSrRbZRMAhg83JBXQEI7aTLf9FTtj2JjLGt4lnh8xp9o
HKQzo0ajnzbKvpIrEQdwR5fJoCG4aNDdvEEFo4D6P/uZb91aCwRP+RIr43wbH88+
X1347FlyIT6/MeU5bwGqJSuDXnm59Gdz2tw8Rc+ARJzV400OGEINTYR7zvV3Pe5i
Lpdflv08dM7IzjbvWN3x+j8mfXpijYDI7+PQLtm8MahOgv8wtOEmmg6WDsrgsEv4
rTICAmRxUXvp6VkuHZ6EDL1CcgohknVdmZmgVn4S9f2K4UtuJ/z167Di7EKqqDVM
uVSzxhCWRJQ3S5ds1Ds2dlPLg5iSzBLHKqQLYZidcu6k10d3Pu8DlCJ7P443wVhn
S1YgeVFWeZEPnaPb29quek/zyQIpTJnD7VnlLyMA0CZovrtIuHBnP5y37YOmrjRa
VChUlENmsZGq4Eea8oC2XiS7aFNyau4TXOszirP8iIuQ64LrRo8ktIQcZg6td7OD
azfxu7zAYsVMrIEQFpYGwGGL7z9ZGvQTWZn1ZxoHb9vHko32oxzO3RhEbxArBuwm
H21ZoETmgSuPL5Wtya1KHgiYwto9PgvPmcX/0Ww1Yqnyrk7J3/zMOOceR6xWUUu7
DTOJmN97NgqQ63H0T2qsMp/C7YW64ngOEsf8O+vHHGaH7fS4K1a94XUbMEmKlO1J
DMr5LTVPw4Y4ZwXn/Q7odQqI0zQDb63v6QVqzzkboANq4jEx0cVR1N0R9gXNLmVR
HS/Cf+ovrLgKD1cEyrZ27OJMmJsrXQKGpCt+8CI5FSKU6Nifga3PjBLUKPsMUq3c
gerpkFc7d47zmo57kFR5jOHugyuwA5T3jhwjF7cJlPIY6AEbpgJCAL1O3pc9mSCB
Qk9zxA1EJ0pauWAv7HpGXSh1s7FtP+HJjQ5oXMgn0RdtEW87Q+hk202A+DYFcX+W
x4mULs6M9hLevqahMOqcZb0ZJAW+QlDY8oma88ovXwqS7/YcPooqSvWzveOvs7iX
NpfPLACamsM+IfvANPb6B9awczX39gJFpEmXuWlDZgwhNQLaU/uMzOVQaNFVZj71
15AOxgzqu2J8RIvtlUKI49m4RytDV+SY8KccKAnYlnD0Z2MC2C/00huE07OdRz7+
liNqP9tgINAlce4XttOmLrhBhVLskcV+mDxQOcrxM01OnfKJlWJouz6wDvhTPFeZ
GjEvEpWOtkPP6/63G2syjSbZ7cXM9/eUXwZxMGn0zt4NMK5K5W7UEbgSSlnlxU4J
3kjjvaif7KEsxPAzJoW2GFv9KMYu3xaOqFOzapFMxyLS8FELCvKs4wXi6PeCATKr
huI7T78K1tMU4xhooPxNxR7oLTayXqGni2I5EJC5v+oWJPEXYCCx+caTs+f0ro0D
EHqr8QfEqTbbQmqdV/xKcCiBR9bP8LP5H4OjxDuAHAJHZyOquTEDxAi4LOyColo8
Ihj6YvFovqWcDGGkxSz8lmYmgDQXAG/jw4XNgReFjDQFoOiHXbzVsNvyNQ2VopRB
EoFa9rJ9q5omcBuxjNL3PVuTu6B5mcDAQJLde5qLUFN4mKCIep147pmQ59t6sdgq
D7Aqx8Zxh12XzcX5P70vfAGQJf5CuMqorjBA1d62tG9T94S49weGHpZow4+rwGzK
jigWwgNd0fjUBZ5inCZzhlOL46XQRTLjft5QS3I3RmYaJ9Uu7pUuUXv+u1mS+Ywa
N3NC4qF0PoUG6pOfE2w7DIjV8QCFDR9GGV0wH8w0n0B4wQiNQWnW4R48GkyEScbo
QF1Is8lmjOH8nUsM8muoz/Mz7ZLJmuGk6kllcGxzBDbI6hQAHSYoovyzoPB0WgTh
e4NiVOB69MpFz22Cq3w+mQwvjwcgrUuDEg394BU0Yfu3GcEDxMT8iv7CgNCFfzs1
Sg2CvmOOqU7SITM/sDcIa0MDQFw6QdlnZU1jSxZUhzaPDZh/XyoWz9L8XUObCWli
fIis4U7yzX9gQiWNlWQsSkGXHMT7h1gOGIUiZZN4GaOPLMeybrGT8yv80UxFoYCZ
7tdmFhoVbEUReYq36UJxRMt1L/Vsq3MLbCXwIluFnAAwsmh2m736J/sPuvxZjzm6
mAqJd9Zl5HhmksFfdmje9nxtDOdDNIHMEgh7sSlSoorz0zq0HRIfvZg3pxP0NwUR
+fkkuAWu/f39bZBkWlZfy9im3E+R5LRSYr9JF8mOJIrI6sfYwiP5tD0VilZVIEt5
K1X66Idm1KI03eiZMs2XwfiPGs8vXHqGh5qEWYT84StB1YQq0nuwf+xmXh6WkTiJ
Csqe8+e/iMKghBtc4MN4L+wQZgUUxOI3BrhJBhPwLDUmxyzo/IdwAgvv6bn6zU9T
g8XIk5sZUAKAyl2/vsZCRxoJ+fGY3wivqaHFylEIxK8ZitQvZyVg5Ggi0W4C1uJj
OLqW8FvlbiQkEYj/nHojSo1SbbF432BE/OuLKeh+mdXI2r5xrDuZPh1A0sY+PzE+
brw6etUdQBlDxNNXIpW7KJbZkXTcxwI7tNHk7y/Xi1cYzEvPdx61FwxkOTS7vyA4
Fwv08xzXIxeFFeiR6Q8xrE7wIp0AqKaMSHFuaaKnBYWN4j5XlLiPWOIfwenjhkGD
32DAYCgTltCgz5rO/XaFxwyuRdedNgJ2vZZyOQaTC0E4tmqWINPp5fMiWLSLK6fH
kyjp94qwkL0myh2MkqbaTinzPQC64Rrt3Xts5LVO3HVTxdNSWvA72xaAIy3gBlYt
JbofNnphzx5DKzLKfnOer2hzM/ER02JdxbLn3TswD4xvCvirDcPrFblQhwwD/oye
ag+MoE14lsKLDuBM9jiB7wTDI4KS1btUgkjpD1OacNz3V7ovHXKwtWplBsPx1Pos
EvRg5ERwhPeM15lYWr2Rj5IPu+KWU0jIKofc9UeLX5SKz6zsSKpF21rmQeWaKtKg
yGjzSI5NETqNyRk2l46CpP3iD/1QRiThS9Yy/r28pvN8ONXtUIi4ASR9Wh3vIYvx
g37HZfu1fzUtl4YKmghVexAxrhkKdVL1NgWIr+3j3W7Waq4lEzZ68efxgpk1rfB0
UJarpo+i+ePjlol0Vh7A2nV2fewecwvFVNFMe2+csnHR7i9mhhq1JagyGTY0ZpjG
mDWMvSdaccMR1WoOyrImpTpvDoljkAsh3sTfBpQR0cqI/QRuZeJBsLrDw2xd1cTs
hRmgu6rL7U3QX4WnauEo8IJcogl3076JWBiDAK7Vkcr7Xe3hTW0TrJbjEYCdZPdn
HEccBTD2eBPgBfxBRtyHUFTs9F6JihYnqIrgNR5yCAm9279fU4WjYNKPAAoUidlF
1yaaE2xo7Nn8Wp5ZVRsicyHf1hLig4BArNYym/yCge8fwO+2hoPULB56fXlrH51Y
A363V6wKFWUing3ECIom/ovpxOBk6s/6aJ/m7EtBuul253Svaczfih4BL/Bi3iyE
JOrL1C35Xe/uN5QToIi7J29v5ybi/ukIJF0uC19qcNXq/z+6YtexAsX22KbqsxyJ
kyhzQasoRoD6VQYy2d+bGQUKtsKh1XXRsIvZqLpn6aL10FcCpk34nnrwXUKAy7Ak
NjV6v3MKwYnXCFGs/7HAfuSYklYw6G75qw1wt1eOXGNZL8VhjMXI1gMZF//EPIfz
9eiLfuHQbY3IAZihvAJb9WNyxvBJC2DvrNr2NRQtbVv5lgVS4UM6SQn+S+bK6jad
aX+0mH1k/Zu/zu0Fz+IDo2Z4jbTDDrh3110nlFAqxwO7EXvuDiQYteWXQrlNFB8P
zd2UIvhzqPZ52OLAcsaIqqO+cxD2/W2PSJH1Du5SqUA3d9Q53sjOyB/CrTv50U73
0Rx5PH5GvYYakYDDMzqb/8YaZuh1wPPKJtvpI0rESqt2YHd++SUjbQ9DOn4nnkvH
dzcsTpZakTKxr1Le/2ZfpPM/DWzIQilxKJZAoKnRwAoX4ItIT2pKlqgg0K8D1yac
X3hyx3kKSLu0hL/sHHcsPA49QXdy9RilpKDvJtXYt3Xknr6abiBs0lO22VfF+mJU
gnNXtdrP1beGoZZoHINlWRUA1qkD8KD/9kNN1M19VIv5svfbIBRxqruyQxqe+t13
fzFwtmr0zvWN05lCOarYzCuRWWHu5hGJq09u9KWe7cVvXLdxU1RUjFO3MHOzDUSZ
y04voDzceB0gWYfGHdIf1jtdeqM+dbOjhgWDoqM+BnvzGn0CjDXZzoRtJbCs8JxE
6Nnwo3EJCPS5FfOBkIrf0RefUZLk/9PntxwK19hAu1eD3V1aVJkRrNH1F2sVx4+h
ioL50zM7OLrmWC23tUXoAxzY9PgPFwWKMUxD4kdfQoaV9P0ckHto9G50UK2Fnncw
dDW1eqemIcr/bLRpi9P1h/hKPbz8+dChOAaMDO571yb9C8RWa1XqHzvFS5avLjk0
n7hrBPa897HhejrTTIwu33IhVku5AheqpxqUiXMGKllgnC1LwXwINrjHI2Iiu7Rz
oan59/PfIjx/nvk6yV4XhWBSszHET3Fip+uzcOweWIXYlSirKmCj0C261O2LAnKM
KoyPWxUpYUEJ0C1pxHlLtY7gl/re56XQ+GABGpMoblgzR3rcc8yADrAejlZ/iyNi
h5kQRBPjDu0XDUpE5ffcCYcs987gxaFIgTUs7jSWmVOkPBXt3jFUsstWE0KrygAd
opmvyFq826A8/ZsoydToPA8ZGgIEn9PSAmMSDkzreXnZ8f01MRQ5DkfZMpehMmy1
crGq3h/r9/DE+tLdWg7VhK8D1pgBD6t8ZIwNHfWJ95TCYM7k5OR44TP76FCIYl7X
yohitEhv/XUg7NShORhozc7LlO7oW0BE7RbmNw1/it0g3SHr1e5d+ka38HwFgrit
26ITClfAKGUQUT4axA/R0BDNkZZ+KbjA1E8iMZFcMwH0AS+zMUjlD/N6Is7iJDZ6
Ks8af8EbJL6HFM4E8eWGFyVKc9eSkGtpE8/qWYqks4dOMzBChWqbac5uicqQvXcf
BtsS7oJLLXgnr6M2U5ROcHmv8DabwlUcOYrYhhBumNTPDwezN6WWg2C1K95016hP
5zDrTP0gTM/GOFFejANMZ5eMgWxNMgHQVDjmaUXqRnowQL0yqWP2xCKvZYvqk8Ty
zIPau0cMtn2AL769LT0wg6edeL8aacfOlfY+VR7mQEjdVpLUXiBIEHPDpw+Pp+Bd
p7yWLIsr/QY/1gcT2T0qqZ4zDHeCvIUETWC4BpKqKfqnIMPcaWlKdtkX+oLFH02A
2Nb+tuZXa1MH4fnU3XMzC0Msk2cmKp9qH9Q3dhIfb+hLp+GlpI/29hM5b+6neUDT
/JZN1Zf9VG2HnymALki/xb/Lj56+rc0kRpYxhfefgR0JTK9SdWwjI3K8Oa/Yl1Im
6Mesaoo+r8oV+vIz7gmcsbEkfga2tDhK6WbeX9xdWS+o5EOpmF3UZd77+OdZKlpG
TQxSGQ4Vbo04uQ5tBtF/YKjG20z5OSOk1qJ+141LK2Tkzdv3uKyvthazOiycCm8P
M/fLU+AEBrhvB4iNiPhC/y0yNgB7XlBubEf+wfh+yb6LQMrSY1aCaOSzC3hy1EVn
w/sGOm+NyyWUHaKO3sHXEvFhV9MiqnlVrCbgs+bf59JbBdo1rRHhTCccN5fRiQ9z
RhGeTPG27fakOa1k10H7QvPMpc8sVyRVbWyyqOvCdsWvBTudZ6TSkjm36QrZyox+
4vS5POlJkxF/epKDuF+YS3q1NNoeJBymDFL7oeCPGRymffKsNJLghGNEC2YLneQK
vzHpuOKTDn6U6ZJ32otij4SHd0Q3T+lXMDc+GFT+wBvVr8SHNBlTF3mO6qoAmvwF
24YXFreLHvqPCUPol7TwX9pU/LmU8Ok5FgNXup85cIe1LesW01+tFtWGE7RGPQpV
ajTqKPjY7jVxS9gTy+WpzkuNlNcJcVHAAlyAo1yYCKWYM4ivtCwLiH7bSDK+MxZd
uWXPt/edY29cP2G5klbx3eXzhIwvk5r4e5UkkqfB6V8EDe6Z9DI3DBy0zJnrQ70+
dcbiSiKLVovujD2GfWZ8ho9ox1h8xx8xHm4RdbJvlq2fSJ1YmwH2XrZTgCumh0XB
RZy0EvtGrkP7b0YwNXyJfMiY29kEdFio+CTWWSITksd8erXDw7pW+jWXjMrIZfGG
4BjcwA0jNweERdK6yVwhiQE2yDoFgQKGQQ2kz8+NF9/Z9R5t9uk3zzJFv5VpbWg4
JN2/DEU1J6798FF3DiqrhbPUIn3uFpD63w5DaW1EF7RtPeytvufCfzh+XhIbi2Y6
GJ1CMPnwM7QAyGWYRstPQgtKj8Y6RqP+qW/PLRwRXWGUH7FJzqZHBlpXS57+uHYl
SpdYKfSJZaeTaVaLX85gbK/mu4j8knAJNTzelN5MbPWhDAT3n6gVHMCq8Vwf6dch
TCMbydxtSA7lYujab7FSEDsOZnM4/Rk2h/qTkL23J4RrJGUx19AuwJFZsOPUrKCo
fbbtuB3PKJ+PsaLsIizRUJzX6JIB1wE7QoT3ZSAqk2WYAQYeYg80fdXQPuP/e202
bixGSkd0qkxPgzYjsHF/PVhyztIg11vijtdjeIAdWKwnS8rVuZI/IuSPFwBsrFUY
0OdCegn3hrGW5kZKoQh78JUmGIcH6f2b7gN3YSdRjeXiZ3QXrf0CDemryP0+RbrX
B1DQ279IWyZKmuLJOYBpxy6kylbkCSz5lxwU89i6XmPWvLb6tD/4ksx1g6cmzDHw
amcuYZvog2Vt67QjDtLXzHRHtT4S2opwnS3ooo546OdmesC3tb/LxtkLSZf5fBxL
00OyZaAIYPPAwUuw8xeBzVOeUpOlPhjZnXSKcTwzngnavSPRxR+r6bVKgEbGPP/C
DGgT3i+s+DhMvyD4zVVnPYoPGwNmCbD1GMAmPriytMXB9Xufuvp8JwKUJdFRSFcA
J2INzTjHG8a7U3ew7setzk/fV8MXJmKTRJMICxmy4GNDSAyQVn4c+IOcxFa0xhd9
kKSz4Lng5ziSGquSaGPeisrwZkLDcmeA/P/S67oZoHCJibab1gIQ9P1xf6ahSpfL
KucUsONlW/Jz9qcpGVu3q0tEE1fUuOm0wzex3P69dpfoERaS8EMQJrfTRI3ivVY8
DAr3cQI1yHie2dNzT1GxdmaEtN5VxzhncAjmSDSeqFqx6j60xx1i9DNCwBH5M/iD
fhiDuLQoWqJkkAchWkxE2eZG1aG/PHfXxmJ95XeqkqS3X+QtHYMrah4aJXmKvm6r
eriNlJUdpdlJLs+/otyOGqEhQYLJpk8dbt5ifAFx/XpFbUuBisxkNSdXeXGhaadD
achcHUFQXAsk6i16eU1BoUMHLInvp5D4a1R1gvqv9QypFLW1Vl3hm4lrM103Uo/u
1U5cXwKY82xpnwy3LcASj/QFdMgfQ5RRsN2BGxPK2m7B97AWqJunmo0JUBMC0Gy0
Tp4mtM8rODLnPN++0MuUNZUPHhAbaHBONb6Zyy4KeuygPJe72M3lNsIbm1WPpAkW
yZHO1V+ZJIbPhlrmzfZCHpQKqPesEF+DET+X2JW5+o2DTR5C9NMGosT7e8lSFM6n
w1bob4C51ifK30x74wG/xvvOmAkJzSitUI3iOauxXvQ47TcDAWuGK98aNI1OCMqE
gEgPwD00gjgi4aB7LwZP6ua7VhgKZ5c2eJtELfYHMy8d7K+L2C3JlUZvJW9XyXnO
FuaB1VRFiUc1HRGMckuXKPM7dKHYgIkJI2CuFx/0Hgll4gOr1ca21YwK9k0LjyZx
188S/gGkgwUoWW0Zrq4uIm9ycky6+xfvJyXqyHgbKwZ1EIECwGmbyr4Sn5L0dpBp
2qz7m5rzNXZavLgpNOi7UwTWRUSPiwatWWCUvD7YtZr9uL3PhA8GKh91d/ekGGYL
UYrjeDo8UU9zPsa4bWrzrR5Gf0oez4ZeuVM/Ah9tc5FgrtA9Rh+eK5bEtbgUHdDQ
6uUSc1maDH16ZDOXwgnZnfyh+cCDMyMLZkd+EjWP8u+QQRz0fy8JRlfJDzM3gLdw
BkWjZVBQmoyK1mblLpGwGs7RuFqI/MYtLNV1lBuXRC7Pq1xbjSg0++yHXYU8Ivof
iWJDZOItaypSWrw/Yzl2jCq1by+aVQGaTNcGf5FWdOYigtNwJwsbkoyZEcwSMP43
/gTan3k6ajPo5J4yIjWsCSlkNRRHhz9CrOKQP/Uz5d9M/zmKMMSCeuN89cN/daPU
BXd39ddJ3AHzFfMsqyh88/Yct14nxO1Wj40odTF+1W2JD/xfNorMi6mIxomnTwN8
gVjfTOLIb1eKnmkegsnq/bZL/EVxyQlshssGAimPAx5es2UBJPv5DR7r8BeftW0Z
YjzsCPnV305WIg9l2NyUwbFsD0fqWXF3iGa9BY/tSWqTd1ZJQpeL7m8+NNIWSvFA
SsjCe2gYzvoZgOw9TyxcisJdF3Cc5y/Mgfsji8Xznuj2m4WlRP84AjXwhu3rzDUF
o0+BfaLVQFhO7tWTIpMEoYba1pQYvGt7kJ07tfdfDAgcKxnqpkaEsZGGwxXmxlmz
aGSYKRixkO5SgIl37IA/I/Etnu2Rx/0SQzdqK7BoPety4Jy0chhnadOjEBHE+/aG
QOFK+Es6xdb7WbSLXhtlmSj39t0/X5GE3BhXm34DcKaCCeCwlHFJBdjEyAxwHVE5
HjjKPt3HZ8t66IMSjyd8GT9qm0Tx/t2rJy06lExygs43hXpb6JkaEou3rKqfCKOa
LDG6YRIY4gW8DrVvwYxTmtCes8IXFdcmc7Eqx+QvQHnrwMLPdSdwT+cinj8uekeE
hjYsDjf+Wqxu9PSG8qmf2zjZR+ctfm4Nimrm4VBW4Yt3lRzosMh2lMo6P7Go2+vS
DZPI4cdynYYfycz/GPq17SC99gx+3KH7JGx2V3bPkMx209q+r0wWSC4J0bj4GO89
ZXuFOB5yCNE6WL+7fyuz0J0y/fpS0R8yNf5oqW2gbSGaRSUFzB+z+RVbSfup8xUK
ePdd3ZusQxwykEHfqqehz5Dif1ZUC2hnwzmba1wJ+O06MlS0Jz/VG8vIYUNLjdDk
oquzf7gxlNwa79kCwCYaJafJSclFQZDVbEg+y+BW8byQLjFT1nBzuCA95QsHy7Y6
f8IesYMdKRQpWxwwNgC706HAK8j/mWZxKLQgJdGUZLLFCciKTdJz2AKUxKAKsseL
TZ4pa0EmicRZPo6w0vpHBTz1lZNB76yN6QJHedXOU0FhIPmmjFMKWU9niWkWV9wc
cBqkoaXhMI2X2l8f5Nst78mf60xvJ87mLfTGWtNEH3jLNnm4pNtQwH+JOCG72YEl
PMPKqb+5OS7ceBLGxH8rQKk83SpX72qcO0XoKVGHEyvfBo7EAduDAZMNAJgZ56do
omGPFiYSScN/V+Fv+wYacl4KbqbZGSDDLydCX+qtYPKkEYMmgUC3pfZUALtFzTsA
Kst8df7fg3BzuEA1i63fXQGnAtRWdu/f3jHQgki4U5aq04oKtk/+q/C5gmAtBQ2G
2svZL5QP4nbrqPNB8NgbDnUyL/OERCoapP+5q1BezbcmLXSuCIyaH+VxwdXjzBDJ
Hf8tCTm7sObwQBxe4p1aJd2lIHzRvf/DeI03EeljS82soKUqa8d0joxG66ZYh4/g
n2mbfuMr1A1Mt1aeDWoEQ3/q/aVAZW4oVPOpIrv5BbcpDTIZvmnNnrlAGBztK8nH
CtQ27wuP4zPiWjAiuIjB5rq3P17xUbdGivDWESyZB9+7sas2UofquoNtVaiVRLQW
1jHW0AT7CSzSvvHsMgE6hGPDY3YHtS6HiFRlTLCBf9xTnmOwyDylvSixE31lB7ce
Lgdlt31VTrpf6a80JTRQDZDSNfUFle4BYPiLdzgWAIY18xbVr1EQZmWzZcAHzyjY
Y0wiOY13GU6zM+QjF9XcmHOpMzFf5HrBYDJFge3SJKe8QQ67zUg9hbMKA4tdY+Hy
MZ0dTHo8ckNegfZdHZY8Ae6Bjtz8GcD8AjoxN6OQOdtzPMn+/rJgaoTD513/ALit
vQ9Oa+BAU/6JzsnXy8uy10+4Hha5HqT8mjkynRQhYLkahuestcVO35djB9z/Kuhe
QI7Lfl0FUpLnu4VZ5A56cQ8xqfvnsyvikPZt6BKuSXBw3PetB4duInLX5hvJx/NV
dfVSRuIjKyVkDXso1j8fZ3qk5kmbw2tvzblyinq4ms73fu6gofny+01B4iVftS9B
qGXupaCNoE8m07POPwogU0KKV/1mJJTnoZYpBKwfF+Ijez3QYQs7gV+aP7sdVJCH
PkN7gKKdbREYy4R65O9jtesRoL4oO3BYgTZFfUnAcAI4/iIR6A9gT4rELdDQ4a4V
DpGtvQzFDwm49ogxxQ0Au6yE+sK37BUYzQfSNDFX2L6KunKm3yvEqI5SM7mY+BVT
A9qqV/8GrLVNm3qOKOza065tyzpLVJttVPPCZVPloLuzsKUvs2Phc+YZkxTz1a0T
vifOoXAQZF8gfY59fdaaO5mtSvj3fJNIvltdqqzGJ2V8d5z5ZNYIhfVNVsJL38t6
djPX+HE1kK83yJgT+D96vMlxK7Il3mYcLHqvdDTnVwn5OpR4YwzRLRWvvMp9brFV
AZCbJBywK/uVPa0ZfUUB6aVeuqERd25wSEgEr1ond5sGZ6h4Q9COYuHt4xsYADCO
JueG6K9HNa42qjsMXg1OMY55ujaWBkmSUoxcBqWc5AKcSlFkd7Xu9gEM9kzByBHC
6LohJosIziMjyPIFz8RpII+pUxOZDe2Kv2k140ELnUz8OV3/Et3NdwS6rFpxuhe3
iFbeSSqvOW6MRj3n4j3Tus6p9f9XGXC6+g13CSis/NkEP7iene8FRrtyPwJQ9aiZ
MRU76jlCRiXVzo1DAMPdN/PpzvbT64S5HDWB+DZLAMcDJJtLshHgmXJvHV3kg6d9
nj4Y0AsFOK/PTfN0tmpM3U0mf6vQvYO5YJv1H57ucUx3AyNltauNqHKBn7WWy6nQ
m8rBYofr8CFeoD3zR8hOs5bQtJlpki2enXyIOQbmd0DSTH2P84gUYMc7qnPXmFIX
A2VpDN6ksJaQbx00DVx24MoLcH2dj/NmttvYO2aCmXdvkuXnP7AwJkIcsFCM/DqY
WhjJ2pRWGkR3WVohEK6v4Xymb6tZprRFib9L2VDod0EkYhV1+/24Q5hEBRKGRgTc
61+6Z8UVqUR41dh+X9fKhxo2HdvHhuJ6puDyFhxowNNtS/5IV4R7HAOX26LBQELF
HG8SIqULomhHp7pjkPC8jD4bfeUsKFRFx0L4F/rraJxCxrONXFHKBCeaYZgiXtcS
HYCK0uViK+TDYTQdY/nviYfVJ9q477eKS45ChWc/wPFwrdKXJHUCNnTOgrMkZcBX
mO4iwHTPSJ7JbfDCuw7MGbEpUPOhl043i4iBfMpsSLSpi3l8D40gI4ftorDoL1Te
3HGXo4qx05TYlObOkEaS149EZMtGBnmSCDyU2im/jEKdR2DnZn1FCQiU5x136QAe
2WQoY/DfbAB6m0y+LfG4QTMAytHDhOPY9LuG55QJgX2qKDT6RD/n6orDTA2teVNq
pwYAeU0zkHdlRbtZEsaQGn5XhleCH3n4DVx3AU8gVWWlUQbbqsynTPQlMh4r9F4s
y6ge/BMFl41ubo1CES36noi6x2eGdI1eSW2m3P4hq43sXUw6Lf7xFGxQHkXHq9jj
6VyAsPQ5YsTV+WF0Pxb4kdTATpAZ6OoMwwOOE6mY7iIrbpBLOV7OCilJbPQf2sHj
/b8JjtwaFx3yZypGecZfyUGW3XiYtvPgTPUM4QSoUhaLyQtoUGI/FfRSkO+u3j8r
BwKIgPhdbg4tOjPIg+yeVC7D/4K41SGOc7Q1DLSKQGOkqImJMdS63CJSCVOlBmxe
qjQtk+UJyxucKRHKl9H7YWdO05OgRVn8sWjvPcbxjlxzi7ovj2QRwe3+g9H7siPB
bRUwWxkA/HH4c34U6rCwhBA2YupsBa1gJ4aBcYlDyn+007X/54oa6hVtfRztJgQW
u6iChOGPYiPCE+sX+SKw441+tk+2mAH0zrYIa19W5ihJs3dsLLpOKnVoMB7hYk78
kH99i/nZNl9YaGnii/V9kqxEmqpBZ1K+TEeF3BIVMRoDNAQHhuZXavNcdIsJ/+YZ
BMTJ3yWfGO1oz2ud7nM3dN07Z0vPT14K7GEXjH8AcgcDtISt/XAat9R/0p+N7RlB
4YfkPuiXFchDPhBUYIBuxKpSl5cc+pskS52NxO/SznVWkFSqFCBglNooTQ3HZl3+
f+jSKHpc71mlVrZAbnIb3ABC3C373XPHKvX7oydn08R+OQ8HUIlD3g19PgEjTrDS
bWoV7mZlqi+qGhryGlxRCFriGVamI3v+23azCq5G2qmMUtnbGW/ApowtnvRQ7LiV
sksEzz3+XG1+QfM+mzcqaIx8PI05XA8cjTdYq5MFFAbok9KN3uZv9dhTNgDgzzGP
cAqpnR9iHwzTMdbkH1mwP1oMDnYEtYoKq8Rm0FhLIGRGW+TPPVemCguVOX0lYmPa
mpSs+s7guWJJyJx5isTxL/ZFxmpT9pZz8jtcCXRMtJVU2yPozAvU5i7bnctTOukU
83qTP4SiKnFwmtvCZdVf+ztoONt4DnlorV0g+dBH/JzSbPGZ4S1z4Uee1FQyXE+I
7BVhz4ndAkx//c9oKU+QFMTi4PBQuNB1ZJtd+8VQIlg1MveasHGxNsnWmRfJpXg0
DCy2hxv9//ZjTXlzqnmwy+SvOnnGivLI0n2etu2WWKuofUTYYBwS5bdZfHmKJ0G0
UfxyJXHu0QRr2KUAcgeejaFks1kmQzW4t+LCvfvC1qky794ah1w1AXcTCEprep28
yelJeLqsL9NG+kSqFBxeaQ8MHmAtjkykRjHhWtow6OJnSKIwkEUC4gTZGfPxc0UG
cyuReKFwcNcXSX29KyGevR2lY090Lje3IjSWkUkukghOySJsSTUb122MUTKr9nRU
295MSdG7XQjLhu0tCm0eY9E4BAp3AWcrui1fGRFdSXTET/OlLGFU3AQ69G2iNhWp
HFbrJJGy5n9+Fv0RVs7EVkoeNd5Mesq/3mlNrqukelHLiBlqJfA0CubP/i4chHOL
xNsGDQWGhIFo7Wvf8N+lyKItfhHffWm5RL1U5vSRfqHUPL0ro3MlqGOQdRmOeCfZ
Rs6CTySVpbiV5I5ZbUXDBRCZ/vw3pJX2uAxjCbj5BQCpoyvHSqUPm8OpsXeXWNzf
5n4K5oTQJd+p9SN9xLby/yXswGuAp/5KaK6CL0I6gp7ejGJvtmMA3MdMSHS/EaS4
w2dAfMnJf742gdpvyqZC2e8mXHviPZ2sDqwl+jzOfdssPLkNxRuYNH0qOiAECWR/
FUmrbk0sw7HSlr9+fUYz6ostLCcl1AMWhQAAwVvB1D0p1LEIacQnkTo0sAl2HNu8
UwGCEmMEq6pA1iVNJvqDZZPC1EtsOd0rZsy+Mk8KFoAm4Vo2xHKd55nc6qNPxjy7
ZStTC3N8qE6QnQRuWXkiU6u1uaB+QzDC7ck4N2tGryGF2x4XdDnsUt4Wh/qVwG7L
fFCvYCGxeHj0qg7YZzQBh6QQAy0qCCz5+7Up+MTruwfL/Vu5qZuGQXqRIIuGTIuu
X1NvyK0n5du9VgWWAfhqVMCYZjZ6W1usgX/9f/0Bx/EsH2BibjDB98z0f3Im2iIQ
mzk1kw08AkDv8ZXO36Df02C16FKrTQc7hG8dIPi0o4AgzT4fOZA2F4/YOmkUJfHr
vKace4zrn9Rf2u41oC9hXws2bMnIrHAfroVd8kbaw3/aL8B9bEpKBfWDq3v7JMes
3adZAkVnq2oHKX5w8KYIvP7w293Xz59y605HIvBFRKi0aNpflh3oGHxdB1BOw0Ov
QhzYNsNcx5D//AJqysqZP3MOlqpo0lReywe4eLNRWWUdki6vF+pk8GhOKpDif/3c
3TMGWKcumpPOM9KNIdWTqM4oQslj09qQmmO6qdOv2OP9rdjKn8FSb/9eXKvmQfeW
4mW2dwYd9PARYJPyymqcqs2JcfpWyWj/MtHnCAmdTkKXcSF3lytJLImHPi/F7qDu
qWLd7QBwmIxB56vRdiihop9AizmJtkavHix2gIY90pEzUrHmMMF5RZVOo7vlnbl9
7+Afx+Ym/e1lG8Pzl19PL48CTCCna3CMctBMgW+oNtMG43F9TFE+5+xVSJQhV6F3
Y4/1RimVFTdyxyhHLbE7uR0q7NBSOwBwYaCKTLX2pjZZz76KQbRpKuWv444fv5sH
NE7hcixQrrsNe0wh5yc2zZACaojtxuOqepr6fXesZIlquCmn9UMoq34uh+XQMkuv
n2hVw3OhMSNdKLrHnKlP+KOk2xVKckfumkjaSJcEVbVs6orTIsMENHu08Mdkm2TA
dnCzMZ9gWBWrGiuYjZDgo41FRtBlIX+AFQPuQlL1Nmkk4DLx8dBejALKoUQdm8WV
xJUVCL5lwSgVO1JdS2+6vg0OooO95kP6I+bcMETQXD+9DgpFq9DOf3tDWxRM28sX
HfY877y+lYFUZgwafdnbjmYrLRzZvPO6u8SnL74t9ygNg6KaVsgm7/Wr/J7ibKaA
pB4mICEAjUlaH1OzZAFu8q3/WANU10B2M11ZAaNK83Wsxed/ClchyYan6fpudPc2
dpwQnoNNkSj85PINYGw/3TtjNiOzzcokHy27FABrmjIAm25Rk2ukqjESrdlxWGeb
u19DQkequ1pWlcP3S1Xksk4H5q6pQBMv2Z0qGYF8IFGG7RAZUFVU/UsUlWvNigPq
Q0jQjvBwWyGGZ6Sgf0CzL4IoYtMqTwxYSlZ/Ai6X4Sne5pmZ96vfAC6k29VZFwrr
KAFMB4Rir9CAMoavzs36gshN1xxLjIit77dfzwUKmhkgQxguthvdj6WA2N7hH9iv
WcXwRZ1lJJsfarpeZxmDU4ci9oKOEcHNKon3EsMPSbVFSydfDRKtil10vfcItNd7
wW0lRddyU12oiRrnAMDolxyHqRZ8Q+8zVjaAd7HfB4afL9S4QZZrKCaWw17frWO/
H5cCeHaNX3fNQOr0bXThDzI1Uy6Zi8sRKtpSP9NNZAvfhWrq3QBtM1sRoBjVDs3K
Njfva11vSj9nLUhhSH8yEBaqdMX5CIi9oGzFbi2m/8AG3uXo2rU1tBwFut5oJzZ/
i7TafmOIPMQarO7BMj0/BcQxa7op0SUnPfpse/nsKOssdqxQEmJUpt9cIzJzj/N8
9sEg5ExnPUwDPiPUpp2GFWbpbAnUmpJzCGf2foJsEb666QOsqHms6r/VVVstW4f0
Fi1IEMoLkpEtiEh4UG2+jKSXmJSMzUiJmfKFiiMV4+vToHIOAizeizOa6yfRjbYD
vV9TF9bqr1QMwTrS2VDTnU3a4hMKxpfDo9jezM4dY8YMSDLs4lRY6GOtUbJMxmsp
wzLn81LN5/7DQLsUfnqureqdlFwyHNgnopDRKBaI8XZV1RbV49gGee++iqW//XBo
5278HKumD50OmyAR1lU84kyyGeG40ZhAYHfo/laTpKJs+5sJ6KZ61XjPijXZI1Oh
DtlouGyKR1jKgn2NlRFQpLYigRAlLQF854icufk7hiPhldEi6BvNgE1+aibmn9zT
LzssFtao2NItfR8sClx7ZodX0/LZJAMiJf1ZzCAASh4OwDL2AYHk1m+6pZhIZ+xW
n7YeFHyuxtV4AAi6vso+wRqJ4aPRMdsxZn+DTkPYksJdjGCehy6c5CHDSM1FbHsz
pt2ObY4KiHpH+pCtwsA7qXCyo3mXLDStM8q5Jh4EIZw3a7ITswpL9z7lUNvOO3Rm
5Ls98gOoTslEMi6R3s0o4znOJrfibp6iNhrohN0p1BlZIhsW6hzTCriwbmF/lmte
9/RZImXS8kmN+DuHxMYVLjk4/5F38A+7QoSjDs93WUjKrqp+7UsXaye4sZncq8DR
/YTJ33WOMLbn9wrgnguNf3SUW3FzWpMqK5yjCsAcu36gn/vqu35HMeusecsLxGFM
7U6fa8jONVJx9qoUn/2DVO2NnuoyVemaVgUFfMJNJkKTJqPGYm+GH7wVVEiwWj+2
SmT8GMkhqbNFBeXE0DV3sC2shTl+RwLvi9vzWoRjZVTe4gtXgQARah56ovqlUrng
OvOZSsp/EctxZsb3af3DILZF1yf1JTo19yX3hs0ra92nD1RU+LJT5FcM7afXp8Nl
yvmKoP5hKX95wH1yegJHPjD40xGVS42dfm14EUfhBNw1FlooMNODroklNK9/cGP6
ZNXWLVdy93LCawNTSMyfaGwcJ65DshvDFDD3oIUBd9BgjupeUCywxDw6aMUz47ex
O44dnNIDCjcKJiDZUmcYa16/GLPDHi+qMOm6o7z2UJZlvcjXZLzPvywJpJXbZR+o
/tOEaFXel9GOLGQL+4H0ytS85nx+wO0Aq0hDAwo0/6hcAA5MRXTXIzW0PE3MD9nl
Mcgh1bJFqG2in9EfyyTE4nrd6uSUuPKNJwhH5i/EVjrnBsEG/X9RTozY5eptIns/
St778nVj26hC8VM+1dM5MtnDTcNPRdE+R2Xi0vrBPH63pKGWviBigSNJ5vakDsOT
CfIViznPThbii8+dxb+c4FFZ011JGB4ry4OFaYI2+bwxbVj2i0dQSxrAO0AHRSSy
AywEmW3QQVSVKE2pRGp79n14ls+UBJOK38itFpKHyQsZQg9mfNwTtmxkjWKWHBS/
FPfemkJd8ag1dc0A1Xv4/7xds6hMmehK5KXucg/Sd4pqL0diehS6KkYQ/HP62E6e
3Bo8yRZlYBVPBg5wkhZDJgGviLI4thIvW0LLeNCPuK1uRXsaVJUKM17MivuWfaDC
EIBd8kTLLjTwkC8HV7xgMTZ3dxul25Q7av7z22+1roEZvTpbNbPU5TOTlAaVOfzy
2wT97JngSiiyBPgFEDiRB+RAPi9EJrbUgTDfa3tHnA1NKokuIvhDAT1Wfj3GkJue
NZo2xd47Lokx+WH8aRxEtykdnPB+a/F3X5u8Dfb1eRV9WNa1X/IMiEkSWEWOsVma
AkdkgGCIzb9d3v/o8++r52wLHiIBMwoB14UhWMaR83yoPgIi4oijzq2kDSJun1BU
WCKabgCFMk2zSE52pqc2NqdWudZujhkJTBEAA9xSOxJYb0J7ocm1VVR3t0swke+e
rRhNGyAjBebgJs3EM/HDv/2JyX+YPKbKKy8dB3iOIDNBPrHjFHcZ2Sjx7q4JQzdz
FCpf9B9yjH/0W/OTOJWSWJ7jBzNzxvUCqbBxqkpLlLXVMq/+lWriNyYS2qALpxnE
+VuN4EuSx7b66pJnb9HKGFqyvIJxq5Wh0YgSRJkrLlg2wzKke11sHDVunhydWrLC
9sAXf/Dw956gR9TOzU04jPT0VL9kwGZuwgq2E+ucilYTEDlUaDnF+crvvBP46Gqd
+/I+ESo/OvTgQQn1A+gsRER41K3AKZ3mTokN7RDkiiRI0ygm/5CdhGv9YIy4Fr53
Gx3fy9rNSW1cKTWCf5rr/vh91gOodRNGPejAAOoxLXVvkOB5zyKYPwk9UlhWzGPJ
dw5aLjxc3ISWhe+7uuRuiytlh9ETSGpWVh5gXyXPHBQEzmHD51HMynDAfFFb6iWJ
mNEJD3ip4YZzBu7paYx7lq6S47j7yEjVx+O8eUNTkSPL/2xpOQcsC2YG7J+c+kgf
4jyYuEt4712L/X6f4eiz70rxD6dIPG01+n6ky6IWJfL7qRtg/fBm94Trs1DUCLtw
57U+WZJPQK+X2R1Df7ISK6XUS9iFfcv6jNblTprhi/GzdBFxd6PxvaF5+Lpc5Q7o
htR2tNEsyPY0CQlOGM72k2B0yDNIVbeCQQqhzOsNU9QWOyfjRQSAUIH1ZFLcHbK8
sCG5/5i65zomjReHIDj1BI7JPi40ENhVhQch2amns9XGYe8BN0CwuZvTPPtLuT0h
Rdl4ocBKjoRksDA/kqOe95lDl5Ypt3oGMbGuUmlhOPuM9csv3ekPF96IQDnvxXUE
oUL7nxYnLVOop5jwhGl/X8v9HPkYnamj5i97bKp5uzXy4ucWI2dfAIWJbvs7CxBy
HAd8X0etlZciU9m+puYcv+7BUCqXDXUZq2M3/+Tv7Rw4q8JHQFcIdlBOam6QBrO8
gjCv9vt3EKP/I7XWCLvFXYfGcwCCjZeulVyK53mmjg4j7QgGGi/wtx+lZaJt5aah
t3++yI9DL+UpgiE34Svv3B6q70V+VPJpZV4jUSvb4qUZP/q0rH5FOhpALiLvA/XS
lg4Uzd7HR0cC59DEnNHiLUyS9rEC1/QrP1TnPbbPEQB0CMUprq1Y51FelTN8NIgg
8mr+njQsjsO+yS/lz2j6nvYGORwn/QQDoE8+RdFJj1R9i25Qz0hTC8DOlPuwmVz7
FaliSkcZO3HZOQLXS3X4aZut/r90QYltZ1vTL/sG8EuS7WSC5XBnYZPQQc+ZwlBl
yv6qlmV1CP801Dv2UM2W5Io2QQHHyiKEAZAPnW51iOUGz76nOXQMstZslPhsAs6E
/NINh1slNZ/pdVjYMIuJGI7keQp6iV24KaOTztZIY7trdisVPeZTnREU9FQMdiMW
PB5YqduRCZgvkYPOGZcHXjgZOsu3puYmw3bg+Gkczm9YZzbJoUUg8U7A3RzyFp/u
8UL8b/szyzIQ4C8aCtXm9OFJtrFxe9vNroVipEwiCrQnYjG16ng3Cedo7qSOrgNH
XtS0FuiK79OwgbE//UVboUYs2dTUaw85mO2uli4YGvqJVJTx9yy+XXQBZWl6gs4o
uF6BZyQ6oqSsV/dJkYtJYJnyiMP9fQvVZOFz7k3M0FI4cSWb/tBQQpE/JMgMgf0e
4jpfqNjsDLWWs5BqTXyrAT9i5FOYx2BBHs/bAJSKz3WnkAw3To0dElFAI7tOm60v
L2bhYDax5ZF5lpulWbm9O78KdppxN4h2Tb4YvuN1F6zpCoxJcmRf5CrYwAAb/EAo
LO3Bf/RYpTERyqYRAoexx7C+jm3pOLbGr1hMm3WdPwgtNWh0N7pgFMCVNJIW7V68
HMAtpXYOhQ6LIHPqcLXC7vQ5d2PwmWOn2J9hbQXQuJQ/G+06dC6+27mfLeXZh/Wr
kObcl6a19tkxuPKPapYT0ojRzVbrtkWfUunwwY1kFfzG3sUJkNMKxKeD/POd1zf7
PQDcZTXzM4bx545k1+yeBAsmZDoWggj1FnyZuY591d9Vt9/CU7BRP5bwfbYudoPx
WhZrMn19U0DebK0BnC3pYFUsIjmuJ5W2bKf/20ldPnZj4T8PowQIHHdbGvZekrci
lxb8XH65CWXIeXA1h9yy14xsAFPji64W/lm1EzHvF+KuJ9kAUqB2Sj+4FwImmOjH
Gdvbie+eYIKPd61c1H1rf1Oi+HSniV9q5AtMXmVZwqrIK40Q2wu8TYjmszK5IF92
1WBT0KxqBxVmyj63E+f6uY0LTJsPTEGgNfX4uFNm8Ba2T9aiVfcMPiuffnhUjHa+
nMIfX1mrqfPdkhR5FLvURmKbXwD3d/4kJAacnNuqxKA69K8IzY9vzcAbvoGNbA0v
zNDhw9mhKH0/hiReCNvjhchJq8Pl6KcM9/JkFVgl6jeHI2IqBuwctSRXbQtK7tgR
4wp3bSpz0mwRkn/FBGSIOLQJSwua9FVlx8Y6k+Wd9+yOa4IVQ9Dyhva6Z32d2/HR
Bq7ZiaSQHXn3636FyC+A6N8WGZVLUW/+U4AERO1Um+QGNJF+MbVuNvCduQCRY+lp
PuPrcSESkP+yoq9el5aS9TDoEZ90OOjbScT8ywyLjtzBTQrG0Fqj8gUq6RhaER9z
PBG8e7HKFZbGAre+6pxAEEtzTOEtfMh7kKqYFNTp/UcKTKRcyd5KgBvOCZuPB1oP
pVyGLD/XWCufTIdvFnpKVk96N9UaEvWV08IRctpFw0fZ6oh+GFoj2S/v/W87LmHy
u6m+uVSHagnhM+KtiapbYraIf2kZXsFGDut91azTvr1oLWbLMfz3SK9uhiXjLa2c
vhnsjgM8lLXh6JG86mU+Vb/L0ydjEDyThgDGlqdA0SzA9+0m+ZZ686uph4Md4SEz
Uhqje1UveXiJ/fx8g5A7+yZTOeZwi8Mr2XHZ+5nv4/J9+oZ2MTrhmqN0WVOo5Nls
s4fe5t5Qc9nGykey83qv4wEm7AcBGFMPhITAKkC28PAgWQkMeeEW/o2/a3X0kjsr
BcO0sKWspKnoYkxEKGOA7X7HctJ/4JOejsvBb/GIkwSzGeV5ipiz9KLULgm7Vsgu
2x2dG/J6EHA2UoSFLSHTODMfrDp+x4HtO0ivu+qvocJU7RVEFPFby1DbSrneseJ+
CoAsPzMX91L8nd7My87riHD0UEJAzyy/GfSHR59UNAKH7sENrLb7IiB21aUHk6j6
Dj9RcYxbdMzs6gYSg/2xE5ab8dzbt6ZjecHZwyTszdvycK+3Uc1Aa3IXr0J4euvX
iCmQ+gN4E46c70wxd/+5C+7F+9fozmTVpTJ+0gVPrYoNfnvk6t60GgsMGtuWsejz
SST7W8ePnflVg4wM1ZRNwR6tLv4uy69xVrSEC6b05V+YaNFHaHbVQDYY2WctMO95
jqukAUvfc4OtynrVcnpGJoDip6ypIkqywSkONnicp/OCm0GXWWmZBBwhP5AXzKBl
L+TQGi5w71QwXlSqls0NMkmQSimGpqjfcU/jp/83G3ZKf5cjpv652AKQBfUhuySe
GhIOv4RXi3EelpKNdN22+dN01LCOjBG1UqtU18rzGkM0C9CEuWqWkiWkpHQA5GXg
/f0D3S7A+W1uU756vkcr2zKmVRKNvEzOP2sTr4aAbTYXZb4D+/ILNQ7hBj8Be4M7
uG3wjTLkLZQji31r2VoEId1ywZduT+ivfB9hpoKQJSnucKUmMHYiTaX6S9DP8Nwk
2ZQYVGvFKc1IQU9Y/msqqzKgbEda+WIhMzCCzSCVDZw3I59aZspfJuUEBosV2ULt
bjYd8y4HqZAQwePGTjGltuRZMwkUqF9Dy/fdYte5BoF3WR23U+74o/osFeu9gTnM
pkB4GUNgfNDpvZHJ5zA7Z9rjeds5ivhmbqkm6RkerHCkkSEVsgPI6LVFqpa/Nk/8
E17L8N9i099pinZVVnioCkvT4lyLGBy7qhrcY/4YlfmdScrgJXSyb3it0HxpN70v
SGRQoFLRM0bWAI631laJjhDt+D+edJyXwgUZbBH5KA86XYP5GI5sRXQ+XZ+pNZ74
QUOHb7gfEzWlgfv052DmTA+AAaZeiQQsjAm3/S6+uAIQfLBt18WOlJY67q/Y818s
yydeT58hAkNu5wCkO8nkiBVZ3L+f9shyfzwmqKDid0QFyO5vTclm8DnJALdAPedi
Wj4ZedDXRoqfdkRPivfP5os+l9N8ZKz6IbS5EowVmEE93YNoviuF8l1c5tiuVtkN
wC/nBvahxG+Vtp/FKAyAT9gAmG8zdFtu7u/Ir92fEJCcN+ef8j9z14QBhqPZAQKK
nI5cXHR4dh9KOoWfQGmpMfcMOq5LHQz6krQDNK+cg6p/Z/02Hwo7+RU5A7rmEdk9
9mOPRidXWrdbvnYq/zihoZJwinHjN0hKO3v40SGx31l9zDSxxnW4RCv5lBQdySyh
QqWNN9ORUcHXpfkssA87IYi8pD+DJ7GuqfS2nInDKTesomN1f1c5RoX5nm3aNX6E
8Ubluk2retXAbnTgKImTm63cF7hG1rV+AO/kCb5T3uhshbAMQh9Zwx+0uORgPJWS
8qaUS5K/jedRzw+h5Uv/PFKhkwWVGAP3Ad6OYCOUth1sV43iE/WISRcSfbbwEzKa
TM83uO0VnBwDq1GmVdjDV0aCYgvMB08Yv3nAEl5SP4gzegHaHco10BBXKMZEzdK6
tf43zP1Jyy42fi5t+OyBWJiV9kQES50xE7Eus8hhVeMeG4hu/jEvQ/9lrJk1lbSb
lb52OzZVk97P1tNspsSL2GG59SFYS4xKgYXlpDx8WbOBSWxteFKtosteVb+USQQg
1LBGNFX0tfOYN44akxjM17cy1NvQhPOBxbIhthRp6es3XH6+32s65LjDJX57GmAr
aXDhalTzyE5eR+NNAJXMNnxkBmrEvPIl4EZ+3G60ARWYun8Bn1QOFnKtxdvgCfzF
UQsXhwpAGuek4bgjXQfvevoYt7j3fF040D5YTDtdKWf+r9BeLTfcm8rv1pWHlyXM
Umgv32W/Li+uajBrRX5EKPmeUBdojclhX1igbgpUThjs1K9m+31YsejP6cmnTlaj
g/t1l84DZHoOw5EM5ro9DVix3PVCUcbNZp8XZ11BONvGd1EHSSzT1DjaqflnVQwJ
0zq/DoVDdANkJmrwe4rvdPQBi+h15fRwISByX+4Bje8iwTJthrCXdAEBGFD0AcIb
Ageu6xsWjbvVqQpe99EhpGRuZYae5PQiUcb00CVkpogKWemnsP4vrxARMUbQOqVq
5RqhLvEIfWGyqjq4ve0DMMyk+0ctmC/gMhVOo29o+NQT2I9l36vCrQUh1hspfqm8
XM91FjUkWVdt7Ee8IO1eXGuJeDTEbIeHrAV+3wBfV2CZce9vbn7qG35VYTdFeuT4
/tKS8WbALhmJrsSMovIM+tGfUyx29oETpT9vPmbBLAdUYMIguyvgpQ9eYXjRMUN5
ELpKwRXUZlpnCZcvseqHjg3sxL5VSzIy7JJXWqJ3Xp3f8l9nuQIMJll1Zl7DInp9
K6k3XHxC2qjpi4ltlJnwMePEwKUchg0GmHZ6yeFDy6Q5U3b4Ao0KA52w66ZF872z
QTkwV9oD3sz3zO98TKk6i1Z+ExHw8UjZUMPyYgJ8jxLWL4wITJiRev9UE/ARD82v
LUAYlms1IM0n9o//fj+KrfuFbmVSZF7NT6ZiOx/9/MVIlT5/qjMxxxhFjV1nlUqu
YLXQH3t3ifrHF8OssKh/FcFQGkH1SnJcTJhc0s+4mREmjCZHLFmfuUhhio3eNMjk
gjzwhK5ffC6lV9PeOTV+x3Gq3mlEWjQDMXS1oVWfRZJj4AJtqUwBuOCmSpRZJqtk
c4eTobu/0ZEX7BbRGUD7gnFDoap21kqFYS8DXHIuhg9awseSnm3uc7zCyG6MJUt9
TMz7uKgYDyEYAhM68JmQJCVmJUZ82yEhiYTqX0KSHHAZqPiAnTOnXCHSvCd18vo2
Nmi8yY9Rty4MRjTZOcbQs6bNaZbPfF7nkObyt2VkSfYPCs4Q5Zs3ADfHn9M3c7sN
ce4NOAyIz5U3O9Ubv08go0p8IMWCnMBxCbtmrPV+TSEYsKoN2yzZrEqlFxZ2kTZs
UZF/hNvH5mvK2hc4212B7huxxg+e2KYTXgELXresD5aa/txw+bZL/qMHGwQ2q6FR
DRlnsDEIBl5hmnHQsGfUR874jdD1PgaTT6BYfNnv5/CnAdzhNl77RQck/L447RwX
lUmevBhbF0QChxitQPoR72w2j4duoswTHdmzLS2xXXLqnu9vs3+9+NZFykYm2W5C
N7gAYb82hQpBKOy6m7QG/IR0kgA7gBuLDnlJgZsYFYvUksCJiHC8HtgnDiaCeDvZ
hkZtX+xIaIq4mJz/3lOuK5o4Jnuo8zs2ike992HxlG0VwMy7bpGjWn+FME/3rCB5
Ykg39j0NMEPLbjkMeEd1IdKld98gvHWgQfGbTommIJ9SGXVxtlXN47KQo7l/ay8k
xB+EXHblqvArxakGM8uC4GEiKLwV1gf+U0d43P3h03pfg5RD0o+B8sRgt4oWQRqn
ZL+HZu9q6mCy9BfmuUVwGH/jLpMQ5kDHdgeLQTvUeWdYfJZ1ujhKlY96ImTb9Ms6
NOSM+bT+8ZtFqu3O3sfxpMp2r7hYPVem/XMmPgyOyWvIewt+fYWPyd2RVcIjH5wO
Ub2BTHvvUU5cPrGUNgmbIj+PMpXYNlm+zA9R1S/njZOSrTmlu55QR9oGApyvbmXS
X7BE9xS+S/cR6hSZmBMxJ9SrqsXqjy0C4IUL2VKIEYmUuiy90xTXIAkKW+0FSMzy
Vd8Fp5mEVXBu0VK/GLj31uby9YbOraRjCcYK05fvh1rC/z0M5VmPnoVJI6bTsSkN
120BvkhSd0NTgSO+IgH27pKiIf5LqzCx5/yExtR8XkiejqfE6G6pyBnARHFpMeHU
bf4a5g4LsT8fGqxdgHcTOZbUPXkUXSjWti1a7eB8PW3DJe3zwZ6VgrWI3HABOXEA
XQOvuW4Ff3Tl+a2BBsm/kpY6+t3nHCov2eJJDWf+E4ueoUTZTLeaxd3RBODCRc9S
jvZpsDF1PCL1HiHP9Zvd0EPJ3b9NpEnPJYZk9o4u4DQBPd/gX4tY06VKc2LBzJqs
3LEbKBNKd/xFa8hGf/BVxZqM5C6aX5xYZJI++mtIuhsxUo1bakYIcLZiT3PhRobo
psp4zkwK2CCRXHtHOnbS7sfbkzUodYlgfJU69z9mJC/JN3DYqvh2tM+QzZbStPC8
cxqYi3dakLPEQSk3Eiq60oeuebX3x1yMC8wX1MjzM8s3mO1mgip6MoolOobpPmDK
hGZxduTMbt8LuTSn+JgacB3ca69hxuOtcRKPdl7PttqL3xkeCtkeAzSYrM2U1Wm8
aaWVZdaaJ4AoMlKG3YMK6h7RhcefEKdgWaYe3/TMFZsKN6O8uM6iebHT9JHT/wDt
2HpLIy4A8QVYf3MOlUKKpb0Otdu4QR2j7DjlLsRwNBv5Yizur6ftOXzNrL9RjI5h
J5SP8nN19DnoAxsM/jh46IyGfn/5pMT+etw3Jbuie8P5NzeGaSwiunhvS8gON0r9
5G7IVGj5Wgzpr/cTtJn/Hc+dHGkB7JMHbDTmFMRjbpyk42zFGDS421AFUJUhiF4O
2DMINwkJqEN8uov3LfNX7ELq/Y43I1oRNoL3Z0WBmYsBpkkfR9zQvevrN0O/rS4M
uLtQE6+0uXk4DwUl1cPyC+j95WPlvqdpzaijURsxh01ZoU0csMzdP+JIywIl7Jl5
Tmx3ZLHkSVd3sEDHHB9nBVM8oaYc+Zucaa7UIxQ0dmEZTwn0I7zaJDfrtqBK+3CL
dgHrs0vV79LX/IgBA+4zVG66Be7xQUrxAbke0CqbpfQGRx9S1xjKVm0AHhxm0aYj
6A3yyh/ZBVBkvnN15lOTzYYVvHlU6pMbsa/bsx8ksw7PYd/ZAg0hnVLT/zCq0H8W
D0UI/6coXRIs26SOCORwQtWwbhvBqcZSgNu8EwVUY6JPA4ZfMM+3AiBO5uOWDPAM
he78rQ9BeHDRgUiN1MClJib72mLDBaG/6Wt1w6ubjEi5RTkUQZpaT0u+3NRKx286
545ty3AIGT8o4l/8QUeyWGzTM/9yQfUCKqUGXBVQ9mN3RQQ2kKx44AIL73wWaVEn
GJeqzZyPEyxIXe4rB8JW/w+ju11sDJL/pMtWpGot0BiGx0Dub8Pl3Yf/DgfVPjOV
dj0ANi3Ra5mo90Et4nUJ7CPYRZVIT307m8BzcjZNChieWXZFViZDljgwHSEUiV9c
TB/rEVgmnUcyZfrCNxUhy7QG3X6L9cdy8kZU8GCFugRmnJwKcq8PvR0h0aORC8Nz
BuVpQ36c1ZIH8g/2CFBItz4RjineKpTSWFy/7I1rE45dFsK3vsQbANTpdpGIh2H7
ZBCjaJqT1zd1AZdsPmYf+Vd3ZAADgUwtVYGdZ4qiNDpZ607BsIfmkkMOzCIv6xqd
gyiPTGBhElvq1JXfD5QbfHbmDtYpaj8Vft/BhmwvmbpVN/Zv24H2kDR0UbjndxRd
KtfEZ8RpkbN9+PfyIZsr9dj7eqhHNOnYzSmT2HTpXItLBJfjqJ10MnvTOAG99N4j
lsXyn63KBPvEeAf4adIoGQymUZkVQ7fPyxlNgbGAHaAw3DOObtlpIZFMH4ahh3FB
W/xsO+5jOqtmgDSBxMCZQXLEG1LSOSA/x67DvUguVoVWRTC0lsLJABrFl1YRfPjm
+6dPaLZNfkJkCit1ZLAumTQ+sw7afoDHHZGhZZRH1mFupztvff5R+5xnpP9pI2CI
IIXGsakXEE/MzDWoSemP9mM45Xgwi3ahTAXVEq9VCLdxNRLJeyT3OYnEhahnIBPy
Cuqg/mw4k882ulXNMYZChyvRVG99dWgx0hN8B8QK1eNUEGkGGBLjoeZth6As7wc/
QOZ6XGbxnXVdWRnHVcrKDKYiOny9Qspst+94R2ScFDEAxtdw/BFJ8uUriHjrCR17
sL5xLLhrPHxl+xECidVuKvsdH/W8KadhAaE7PtUVIqMYlhhvYtA5e3zUtX0BZhD4
n86bliH8Qt6fD5nXirvnjt1VMPQqsLm2Fdf4Z1WSmq2Xz/Coa6e4Pkb6+TP5mk8o
2771/z2+BmOmLIYKhcTgXy8Uj0qzI7vIwTVicmOY3hGCkR5USHL3SP+VuA3ncyK5
3nWuv59W1bxAqZN40BLl7+50SO31fnxuwozEJzyRxFYrF1i5D4Ghtrbg31QKp8WU
XOqVQb6uRZrBlS3MZZAx3zUEdXrYUb1U11YbPvmTt+W3zWx1lE6FwJZTLmWnGabt
9Oi6S2q+FZEj7hRTdN+TpSIs9NPgt860fN0cssuEts9M6YkIkVpNhe6gHmieTuLi
ZJ9nVLV+mz3LdNiKfM0EM8lLWnDssCye0JxNaG/oMHSA/+UT05aINsMM0vTwZ4z7
50Ml7WjN8i7/L8KRkGw7WP6+GzfXRBXbRvCvqoPIyVW4y75wXvGlmGHBkMCIWA4o
2Z1vxALh7ZgXNUA6HmcyV8c6sfmiquIPLYpxfuwmna7zP6abSL7eZ9CdZfdeN2gt
WyGB9Fc/GC0665ZW6+ReaZClSsM8sbCi7pfieCtIjwTivZiFWQv71CzeDywzzxZH
zLPE2Adkh37qeekvuPlaL/E/8mFkXaXMIAwWayK1j7ryGhf3x4TgppGmugfSLE2i
+Q/9p/8drbmYep+1pldBpY4TEy0owmOcxTVIlW/RLqBCWst7byuoYkPmVwwd+CcG
wlW/5u4DYbSzK58opRJ9iuKZTf0YW8qPZSoiaP93/ddPj7TUgGM5qIzwk0GPgBJt
nCq5gwpCUR6c74jCiQ/kZvSgFwVBaoEpsFRexBqHM73qYjMnJ4plIp5Jf6MyXDcs
ee57je1kEmkfM3KJylCyfJp56Qg7LUQJtEvgJ9+i+OpklWOb94toC1YTnQ4KJMVa
bMwDBWYveG3lyQOR6XGF3LRRHV9bZ7S9IdTNwGiNuiDtboKHr3oFK1nwKF5xcfdA
17rgQnN7C9eEHBa5Zi3ZzNp+SZcuxkYtBljldVXO26u+t/nkN4qR1QbWUV9eU+wR
NP7o2M+8Fa+o9ucpr/JkY7BNLo56l4A+D0I4qGsBFycrC/cIepZRv+zXmE9mj6F4
CUqvsY9VDYIQ/eClj4Umpsmz70YRriwB8QktwDVISKgCbAkfgydhm6zvKoVT112P
yygvNw8b2J87+g3eQDkImuWb2epRkEch9BUNt7AhuriOHiuEeEH82ywCMJfNX99C
q5ByuelY5QNgjq8MSLKum2Ek+s7V5JsJzb7n7JO5saOQPY6p7casO0sRGl5KGfKQ
25E0BMmtpE1UQa1+py+0Fu3hb8gRcWo4X8kI4oMJ9dVyhLeOIw50YvvfvR0jRxwU
i8oEjxaCJB9w3JAtK4MkDe/iKQH6onEnUbjw7/2PqbiZn4OT2lEigtOxhtQ9K0D2
FH3i0SoAH3ufao2Ekxy0z1GL6Qgya04m7h0riJAUcKdwDhBt39TJb5pxkDW2rSAr
vA9v2MVLJqVJ1WtoVq8X9urMJ5VuDrTG57OqebZik6yrB8jiChS/hgjzFnRD942u
YPi9JZ3HdxphIp0wyed4MXYd0y/5l+DqcSSl6jYOHG0NFEAjol6Vvhop/H/dY8rX
VqSVjEE/+Ssp+r8qv2miqiYxQS2bQ5EFBcvlxP/4wQDooFnNNa84rsZrdbN86sm6
GhXtuS3wDC+uts84Ce5rRhgsKbeB7ZxkEqa8miww31jAG1V/q2vluqv3VTcLrtvA
EP/n/NvELyfLZaBiKx7bWO+ZduYVlOwuJAVMY/7e5T67SoYULPtDJelGCP/2BGnk
3SnRsBDPRzrkk8F1Zn7IHVX2fHSOo7aToSQ0vzAxrohzABTrrCnEiNk/hAMwuTU8
h/vTx/SMZzpNDwEEqqNGtbNXCgdm0AfrQIO2DccK0ITuB+pvJ3HY6u9zqzJ0XqyO
XodCemjICg1liGb5pEMD3uinv/sCc7n6GnHhb/N22ogF6SzOEYI3ek+N+a/T7CxC
Vf5ezafUI71nglGbsdHDd8XnxN6H8DMZIjVVKUN+1nDvKoeBUD6dduPdWxKwl3q7
eQXRiaa4ypMk04F5GPd4Rft8lrsNUbL2t6Jjn/Y9vX9dtgFnFWLTN/5WPGrkL+5m
vTTRkj98jH9aC6VC3GsC0BwP+mc2/iQff2a/skPlceNpGg86j4D4topOj+kyRk5T
iCb9nYBCNkdQPkz4fKAdhNMc0th8rG4ZHLOv24Jt/fhbuE7XJnJhAkHD/80eXcoM
LzMd4qvtwr5w92SKujc3HF1i6/JQjdXXfc9IQNawMznTUj0eCvw9TcGNIa6XmSQl
mbKoBq9fuVI4hNiNAjyERDUhyip61wb7Gsb8fZSZE287nYToWLIJ+zzQHx2EU4D1
mn1qMj1efZoez8wufO8srdPbkrocLpqyvSOg96pM5cIwJUDQ56eV5+mqS1vejhI4
RiYj1pMr8VBotq4byVUXBtsVSJWdv5k52pwyVquzKRNYKpY84h7Px3sDhv01PXy9
Mz2XS8SHi4nT1+p3poIkscBScWgUMZy+ZQU4PeNrSMokh8A+JrDOdfNHqbXm4Sw+
GfHLC6xo19PJ8pqLqb4S0yRgDOrrk2cGHhgtrGgj2X0Xq4lJoOa9+lhxGW+AD0dq
ji/lb/1MUcfDODf7QlyvfK4srB3e1M6M72mVfkQ7IXMjnAtcz5uMkEhmohzmn2xE
j4qkmFP1wSiLZ6QoCIvjm/FHDN4CdAcVKNtSO8NTvlX4qslXRV4RE8KhlH7y21NV
gxc10n1fYgoG28cqIxYyNYr8SWolgg/1fgHptfSOHSbc54Aq4EOBQAOG4DrVI17N
EsfOKrqS30OV3Psv/FSoPey/+uzsvSzOAAuTEWINIZxmTwsBEu9zNftiiAr3zV6e
hxI5h9J5ANvRe0rKnN4HfBZ7u0spftq1bFAQ2pWFTFI0FmnVgn42KhyNWaqqHeHs
pZp/uLojxUA+r3+TFe4BPfYB2GFGk8AZYMGzFSo1U4UabHPoDfnCM+FAvalCueln
MXPaa2MFGJx1MOuosfb7ypi44A+UuWSkDucAClk8g48pEBKqJKaWaWSpjzrIYol4
iR5KxW7dtoddRnr2EfCqdzXcUbMw4rfURSD0DZ+F1JyDyBcxbJLMgBxo6SUEtyAa
Qf5NfvcTELDV3K6huQEh50hxEcowOwuWUBSB+6SYzVogITsvky5PiUAoc+frUM63
iwa4leRZAJ54xO1Eocma8KiI70cTXP5zqdn3TvxOc03e09h+XSIYCZ8bTS8TzbyT
5/Zp7qSmawY7c4ekoOtT1kz6/L76ZDmJTY0//7FrHOeljo2AxF3A7oHWJwJ7/+Wy
K6KiCqhuSGXsuPz8Xkegp+0A/7N4xzNNzC4RRbQdPBhrXBqkxPVR2vzDQajaSln3
xqrdNhfsCnCMvWpUpTbfWqN0+Zo0kbBiqoJZJXBN+cs7A2LiR47BUc1cgzwJ7z8D
CDDx0j0d7B1Yr+BUzdoGGz4iaCYVxv7yJf3noV6SBfrvktwHPACo7PVMFacOBieZ
XdKSmqQGxk4rf7BaIFYCNsnKkrLrQqdlSVTWl1U/htVa6jK5pAA7XUvZ7TmPCVf/
GkCwXUmO9vDZcTItJtBLCSGBZHQuI9odkn7HNUlWWufN9Uv1+M3oemXMhF/e2MaQ
Tm41xG1aaz4TQwHpbCEGDJumozf1JOBlkgJFxL9AZvEjJPxQL0Z+cLucyA9HhRd4
jOiPDmvCv2WfkxxZ/42ChRV88fz7mbdoDuiHufGIQHziQ2zBZC1/A4HB4TUvYWN1
gFC7CqYT8/HuY0Y2lF/gTGV9RB+hM/+U7fIrN7bKx2v8D52YAGo0BBKej2uDwOmR
dK09vGO3OWDKYnOCrkEXCYLIrvY48YJjy/GD9TanxJhKW378PgJpsBfy3glwV5U8
jPQs9dGH0PBblHQIwJ4BdfW7BaXu/y3iKych+dOCtnwT2Zb8ckUpc4BPePOqHBT/
uQKG275NRJC4R5yvpFkzMShXBmY1H0cRmkq1KTRjLdrJIY0d1OUU5HkHa6Q78APa
7gxfrb/hjzzdnnFyg0VGk9eaKAStOt4LhQxB38Ui+ZXE0mS8zGlX0+OA+B6bS/LE
X0rxWuXsn7io7eaVfJPBwW7vz6MnsPb3B+gemx5Z1ccmI61OS1uoyQX2gjUwBFUW
ISA74rFddQjBK4TE9tYFR3s+HtXGTJJiswHT2QEGFLDQkKabXFFhLv6pCazK4ITm
KqsxGPkePdkb3Z8TS+h9en7NLSdw91+FoKCPfpRliMDpzJx2wz6iuQP85Z+IGx1n
gK/iEXlGJws7QbF6QK8vQzQgTi8f/nWgbihvf8k+fuzXMpnfd59MnPN1wS/ccPck
QX7GKwmoL6SF12Fmm752H2UBOkdPdyPJHs5WEowiYus0OLXwQCFCgBUcqk2LpU9O
i+61LpDdLWQF60TPnhZl1GMREjuhnv1vrQMVOzKU5IVCVBeLp0yaqXKmckxJRt3z
wj1ZE1XijyMiF/Mm9C9Or3+EwoOm3CDewljwPqfBYJqEuFDXMslNZfZkJG8vGR4K
s2gKHQs0QyV9EGa4jFysxB3GiJ69M+O/Et4Nf5zSdoR5AmyEJIrnKJ+NgLA7/FVe
CeKiqyh0r5b3tUqOG8MkopxZy4aAL4if+ApbSKOPyXqZxEbcRc6aY04SjDyAIHj8
EWDz6KP5Y+v5uBVRKuQcyLGYh0m8RBf5RAPcdR+nVEhqGw3PU0sRnSEOv4nhyhAp
SpPy0qai7jHtvgHX1226wuUNfwjhr4te/79Ohned4yYqJpeQP965QJdWmdFxd4vX
69gPaWYEX74EcVD5T5UIsDc6UH4gJdvQTyM+HJ0KG0AVThNfdPmnhU+1fQeqL4nx
2XyKBzAc81UpZJw2OvfjUox3B/n0U64IsJ5C0CvTk2U0jVWxGLNBpSayQykeClyJ
a7H0E755+AowzTS4JjNHplv1dHsu9S0hpcBlHgDYEU/wFAHw/t/3wnmFqI1cubLF
EmVBxUEfNtTfkFsCZxZqqOax7wlOKA8XPxieBAl6SPCUDfSq/QVEQPPJLCxl9eHL
ANisqfxy7FdLjdNPxiteXdewPjRKqlswLsfn8mRvG67ODZeo2vwYojxFkSmZaUZf
OgzbprSEpiqinpKoVyXuznUwxD22J04vuvyJ5YBzFzmZn3T9P+r13j9GKOd7rnIT
RpTOrJok1qiAw157nAMawCRXH1vi9wNqTHiVwESz6DmYCW4fdlc6FMryUch2/0A9
uSV4fTwWTDQ0xAzTyEY4cjDrphjB3WT0YxbrrtaS1GLdVIJHdGpGWgyJfP0wdHTy
CBVtNjzQYjivQPn7cQRMlb1vOmqOpxDVk4sE6+Rxoj5P5oRSdxNh0JKirPt8el12
JlygOgXY5kWUwseJ48HRZVlDYfuslslUA/eeWhe1of0iz+bjcn37MY7gPUbeVN53
x9p4qEUAFu4FRcNZBYlZ5+AnmxOIiXvu90YIVdp890eSEbeYd7AHE33rr1jGAXl8
My6J7WPI00MGN+9+KGu5Bg6zsLWuTtHUx5ECSzplZH4r5+oftBn2Zahpud5qvHvT
YWPEwV+jmuNgHpA8T/cITlUKYLKv8D0dUdpy6iGVF+Qcp2J1uW9WSti4r8FNSnNO
2mXKgGOwVt5a1wrpuxIb/UGHD9bpKJASWn7J7aLwa9541Lf0cJeu6iRC41B0HwPt
FDdM7Q+W8kFBZxxKU7i83+peMy3P32ZH5OPPmp3M4aC6SgGACReREtgYUGqGAC06
X36R13z8i0MwhiofmjGRgoCwyvByUWxq9TfSZaMt9p9xGaDM1qMZVJEMHlAcLri1
OSAwSMzDnGhC2hHiXXZtEjmu2NmZEeLZ74Y3w5acbxMjIdgbSVv8pg8PIV85J9av
rc8TGTTGXRMhrB5UKz4FT/4NyH0IKXyX7DOv+KGW0wvKGGGIqxDIBPHENm2M5RoD
9IB2dNsehbH7Huqw/eJV4uxylL4dMWAtj6o8ld6cgW1fRnUZJjyP0seyFwIURdHG
gV+tGemJT7Oo0sL8xo6JOsc8tRl+0LZT19Badz93PTT2srSc2+5ur1mACkX8hCIt
AnBA56akk2ed0HWiz5RsFTCMZApZP+MZXPOQxpeZjYEhA758NS0uFyrBIwiyMqpu
1MX398ANFblLJRxjvMojNLDT6Zt/zVorMdakv9vw5nGsNtBNehvpuEQNCZGQ5pU+
jZxJPsUbHR2vTcvc6yaTEXW/sMU7DzbySGNpvGbqi9N8H91kmBMZUx2DqIDENcIA
zvRag/nR5chxAJRmElrk8GEnBtE+su8u1cRlLjiEkyeTp0SChL7B/iTU5iiHViqY
Pk9Yb9VEq12abA52gFRiqTIRgciJ2rTIecdla+/L2GYrpYcQrhBBkARmZqTGZBuU
G53LfeAPzuLpTTB/X+sJfGER6SUZ1NiLg/BTKUB6q1Avd+FxsMQIr7Ftoi9ub3FF
WNSesmAi4ab5Y5HnHcywPiIwgtj8bHv3jBRSIs8AFxCiHvJqU8VFT9QRwUbfe6Vm
nAg5H0U5N13+o9i5PGfNbFAOYsgpw0G5eOCSO50uHS8L1/J4SG8AvQTGMhdZu9Rq
KYKjRacDeFjtRU/uM/F6LK0CsjhQZoh6A99k1/Ykbq73UwPhlP0vTTb/Mib91ACl
QUwn8Li++hdnXveNoPNeYDbKa86RWd595GXttLD57EHHZuqLPdozvrjiRlLwVGMb
mIsL1c8KmlO+GKbt0Pd8lgZaxSqV4fruYNH/xiE4WmIQCWgUH5rCF5Aj4PG31g4A
RJA9kQ6bGB+ZRiahiUC4DyEqpn/Z3FQpf5H6TyrEgFsSkekAyvjoQ6FKiaYAXprj
f/CyFJnLMMfvHAYMmV0VxDOsHxocP/1C4T5rfzVP/2PIVTPDOwi9u5ryv9Z03i/O
Df+uqUFrTv62W58kXTYL/+PmybQCS0uQU6hr/zfKK4RYAAmjnyhDleLUK0X915XW
fol5K6Of/Fc8TiVeWtzHf6MmEx7VjdrqUXPidRINJz8f+oODKo1kHq4HNfV5E/tF
F4cqM7fMF0zV7PeLuD6UEOadO+uv1Woy2xw24GlYkte0G4Mj9OP0kF4STFZ8Zr+S
GuI7WCwPz6su2Ro08Z7JtWOImkU39J1LI3njBka7AXePBxhvQ61ycSz6aAopll9T
kxDPrv+5FAJhYQToqzrtE3yq3L7HbTMgvQgSzsT5sj0oqXaNrN1q+41/5mxOHMQb
CQNGlboi/Pjm2muUK5dbUn+lsBuUTkfnTZ2NmT/j8kYTLPhwhrZ/JXRSsPQNdBSf
Skd5KhhIs7tJkC0eI8oZB5Fw0iHoKElnzdPJcpfMOytgG69j9yHU8fNfCniq3D7C
0FDrpzL374Pi2dmOlcMZcc3EoA/4Tg69EB1sSkZ2DHeDpvgvasQW/OsfeM1MTgQz
cnpOxPfyHH3tphqmga06HqJW8XJBRJ7H7hF2EovfRddyOvBp6F5wkwjM8sz0cxWZ
kD2sCqjJXGQg+MYSK8hpvnenO5BTxutzzZXojotp7g9FbMB0ng4ZySVwOP2swt2y
q0Niw7alQ6KUJdRp2iSWJ63TpKJE3VaH0jZU3Fp3YfGT6339rYGeezKOOt3vjbnt
woEkwP/oX9UgpGcQy9StkRVyy+XyhX0HB9M8zgI15Alui3MxE+9itCJajBoG/6aW
DA/EDKKv7gkQvDbzrJx1S8sh5fz2QWHqbNiDAL2v2o2EfwIbzbsT2gLL2fqMMOSl
RE57l3vOAOnn513wO2BQL2iLAJlClVCZWAb86zvrpH0Ph+WC6tdcvG3fuWKo8OmY
0TlT2cciPfZ47tIPF36k3WI0Z31irYZzt85eTyjkJqi2gjpTem1ZqL8VeQsEoPKJ
q17lLRB7/y6s0uq+6H8w1T77r1Q4m1YauwqPdHFRxbxuKczhgL6hJaI7e+LTI7MU
NBFvqzFHVQ12mWcTUWq03eoMxMeIwKKdQLhA/zUxMO/AcEs4HCtWG8+m4g/f+LVT
i2No3ydVGfQyeiE4Hun0KRDIhShCgAFjC8dgmiH/RHZcECK8A1MIaYIVql8fOtjb
4RyowYG/eMBDOqwjEDcn+0sygxHQgIWTaO8RPv3aWEb5PBOphTOJeapD3BuvpJyt
IaiHwprp5q53sex/yUVvkQkGFQifcvCcNayZeRE4XiazZjdTpXIc2HaGZWKl3soS
wvGQV7r1ry36FdZUvZGp3+WfM1oDXuoVwVEyl9lXM8N03rJ4aEjNJI4gmGEj97uZ
h4eDg2OAlbJtI3d+XUVWo5SKqxwm8pjJuVQBAdhMz9gu3Sy9VEgjJ7Gw3YJ/oQS9
G9QIXj+07lpmpE9jjGj1FSJirAbYS+bqANiMG1tFUN5gNCpAI/2QrFBA2k/ozVat
AHXkeKycELqZ53h67CyuM2Iv1Pbz1RaPTa0CP7Wy+rvFaz8PfI9qXXCI7Wg8/r2c
3K8ih0FAQa/hSBHU8XVxtU1K0Tk/t7hV+ckzTQ226ZWB43XAIj4kRsJIqEUEzoFA
T4zcfPSaLidVSzkXtbvcsS98QtaANKOKf8/thpWjNd0IY1NM/HEkKrVCuwICYXZp
WXkgajMcSOtK72lJAmXqW8rkQAOxEz+XaaoDd+NroAuRBdjX2VsNnSvQJRA73Ku5
lX8NTvB/uI8BwewAWdTzQOECCYs+pNSEvOQhy0BPI5EMy5KLW2l0p5aS05yIgFVg
k2IDmgEY33lKwXRLoELW95gh0wzykRsMMTKktJHGAoIYXVVSc5fqIQTHFgvg4+mK
+rvJs1FbbUjkKqwEOeee+GSKClJ2R9KDEoilSbsXkxpxU1lAYJ1+OjWt7rrjnHYz
7h4hd0D7T6am9wW6of+Txn3Sq8zX92i+MgxNaKaZIhwXutTux08qY7BUGNJVMcwF
Wgpu5x2FsmTCGEudO+n9hhAvZ57YZj1Ckvt7rast3ZFrm69I5jfFUQnPlfB/76pT
OFYzePy3Yy9clUI3q/+F9WPgHLRZRn3hOmFAw8pR85/wk7G5INa5Eff515Vbl5tY
NukCpOw/oD81oJb7xW4jfnmlN5xWVIOHTvIygJilcGFKHY24LmRWnIi9DXSu5dt1
8dq9vZr2BUi3ARcz/yGI7hQYv3Sv1YR0QI3jKER/Fgppy1XP/5Vu/EJcXOKPD5sg
xsBXn5oN/5Mxsp0JIB+aUZkSi+JD9EXw55ARYH2hjiwsGdpSyN1wsxTaGV2lym4r
F5gR29tgIhCKiEIXjx4yyhgUg1ItmncGIHTG365hN/zXoYt5YLo7fYGyTCpO7r2d
TEHFtW5EIeX+PU+xZU3K2en6GsySP/ADV/9w7s/WtoXFL/phOgGQzgXEm+ZDcBWo
+4Zz/LM5ryEoL1/ef5OvnYdOglxoSliTiPPYI8kpAC3AXGttPcGJPk0Y5VyJDrq1
UYFBn3LWfEtMK8yapunk493tveDApv+dr0Am9mtTHFXk7H7mngt0cr6/pNjj/CWo
NOrnrakuvb+TcHKyryqBDf01kwnmz/tyRB33auMsJC1VtzF9egByWZ5VGIohIDPu
Y4yhowSHR6AFrOWj+Cfdwfeglln8WS4GVHBNQhC9yf8W4njFPXXAHIQtJRVM/g5k
qC85GUfnY6mEzQizGAZFCn3DDiERPhgSHApdZV5A5ktRckBUZixV2K8gU4/nmrs2
CZvY2skZzHdTIlRReBSfLZ5gP1Ogt+MRVgzFjIWvruaFKNTZCB1s5INBuUXcqWql
r+6UzG004TGZvho4ot2CrUkYOAj2YZt4Sxh0f9Xz5Uytv6d45WxYJ7YT2rMDruZz
pfTj1s6QJzcjR2U/flfr2Soit/Y4P0UwjC2W1CE2sOod3j5rBYFU/3UVPCD5hS6/
XSnyEMVcOkzAwz4UbP8nDreuGvCPXP6zjooyyIiYdWS6VCIetKuBpEdJ7qCsmp79
R123Ns4hEG5xB1pd0VMI+e25EflifGeO9b9yNR+rZcexTqXetNhy9FFcbG5G4MRK
iblXESbKcn4Dr0qFDj37yg9sqxAqTERMTsH1HjR2IdIIO5bYz0IDpE92rlc1hccB
NxzNEawu+gQ76g0lqp3XSj8PXXURdWKrM238IlRHo/lrw2eeG2kSbusTto5p+DfJ
D9QE5I7syQ5zxosDxiiE2qwpsmnjeGStIuYDcK7paX7trYdIWuEKt5hyUAQ2n8m4
GvqmohSGvpM8vGMQuIiWsFk/5cdkuj0kVbmdKxLd30oxEFi6XuMqQaTQsuvm8boI
nCp83+dHPkEE9/YLpIcwWk8x6tFaSKnbGZCpD/6Iu+BHUbfrKO+7Se5/2Q/nrivp
CnExyJMggO8mygQiYq/PP8XY7luxCb2lmN9rfvAVOphIO7YkKAmQjjw2G0vPean8
lBOYe9ZOOOQeKG8Iaxhn62xf1QW0i3hzslD7SV5xTQ050s+IHIw9zvLiP8dbtpWY
ak43nGTRcD5lqrARt8b6kaYCn5eapiNsVdD84oBAAWBhRcUIpyKU3bscn0wtH3v2
85Lobozv2zb0lgEyDnCgtoUWPlhpmKrYYjHPid5zFDKTVZZZwlhhnz7M53LdarMb
dd+qRELR6AN9lPqvndSfHv6aslSb72XY2yk7pPmm29CI4SHxPOUbz6gdrK3I+Ux+
0+im8ihqm+YCopUkVIqUmzsAjrDp1P0i2JfbV34oPricMnsI1rRGX52EGt8U733H
QJB/LcQWJTrMFa7ykyhhGw1Ut36gxAO/R0CISm0OhGIck98Xka/6geY1TkDGiIZV
E4AeLKDuw6s0wqfTx27ouqp8DUwcevPLEq+0pArhrN8kHuiC/8JVPvYTsGcAoV0n
mHwUGMCBZ/AzGcY09tEXg+Dbd5EmQeLinC/eQza7aij9zJ2qKOOkR0357mch+Kiy
Xv8Es5qJSxAb9htMCKW1EcKI8ktVXrHJ3P46H1XYtGnG/vmRWVr3kpz3E+tcPsYL
Y0ezC4Hfr6Soo6XmwxmmA4kM+wyqvafBIv7MdCTlHxfCixhg3bSlIwMeLBFybyuA
aW6+oszNm2IYSN3X9/GZf+5XC2pmnBUBJHol5mQJ39+80/+xDlDoqiDebh51xzTR
xv+wuUm4dIaEgqTL0tUDlCk8b0fBjDudMeklo+mJPgmwfNE7dQifnGzHOYrDxecn
sDvdPSASEO2HDoaaWRdMjO7hmKs/C+9DCNKzi07d/WjuRagk4yPKj4Q0yJgnkb+l
bg9DnQqKWwOFVjfAPMdIlJ6sG8EzFs7b4+EUkHzdy4tQlu/TMAL8i0GYc6+2xSMc
nOLyLa/vNoNM9dHwq4vcohvcAVXJEet+FoI1ZKNc9AcCtC3IBHvt6SUnCgSjwidG
Lcoycyq1JXNRqWwmS51lsJProAWdhNVavG1gS2xm8Y2Pzkv4K6pucShxzRVvAgOq
NcdA7nJMSNv68J64lCc0/V8Ryqsbr6ZaBQn4a2v3DaTE+ATEXLLxmjZbF7BXhQcf
2xbekt0bNuRWlWQ9AqS1XwD2diSR/la2IZUB9YHJbx5fcnc/A/Pb1MTovpmTwZNQ
oUoyKdxqkVN7nX+hFWoo8U/4ngZypn0uWtKUTiNEEw+85avsI+nVX6ki2G2thmGO
/DCVgU3cpFS4ZwUnQ8JoBiIMHep5EZAgCIsZxr0nDsgVdtxBjYURL4i4G48jALuU
LJ6IxPvXDk0sStc+wgibU4Y4L61pkYM3M7L1CPBzBWRjwrBB5d+XcC6YndG23Bmj
M92t06ekezA3RKFy7ayZm88Jdep4gYl8gfJAqNHlITfjw1jxtw2aeaFlhM16qbX+
FUI/cdtjtbZavqL8zubTPdTfcntC/aFWm76iFLzs7bPxRTP5RaE5XlkGtQ6DocMp
WMFOBXP6PMmOShgt6EzTuXUMyn3+tSlFvem93yg2K5zhol3AOjXqHv0m/vXD0QnJ
sWVLsmDBRLNrdraRgUL/NueNwxoChoNcJb6bd3ql6CrEml8X9FtqjjQv4mIf86ih
VWxfoa5d8zwPW4qX8eG3m4OcWaUuAYeqwuuQL77rgaLCkkby/UJc/b8F1wpPWOWT
EYQcLNHQSNOjPoUeEv82RvU6Swrwv2MqbxY0orWztgC/qOXUMoNdg5x+GnM7CAL8
syOg/ufKbD3VwP21WmVsEPzfyHn3kCn4/WOv+39wNzqT9T/xFRdv6pwEDGNiiVLK
XjC+HsNaFgpPZgWe9fmqAKPRQqz2E1sID7zF/Fsbo57hqI7O5t+bMxZDM5+oRqke
O4uixtXZACsvkchq5V4UvMHfcYosVTrsk4vyimRBHzf1M0ObQRFK7ebwydH+RGlH
1kmlr8WKRDTXr+ZorqcRjA2ppPA9QV32U6+M/cbo/ERDB4ELCt/1ELGPqy8EX89D
Sd1D8PVVL9FyZJHqOnPxtfHyA1ZN3bo36cgP8zzZtTyqjjL31HXRYjXngRH/I3hh
+QZFwN4QefdnOX7oNEAs/J0UEAVyRBCMMsZhQWXFRZqVgA3N2UAamnHOBtrx5HWz
JT3pwm4aCj6EYLwqwIjONbu+0Eq7wW3IgDfkEloIR2/3/C1BSc2lMk9g9A4wBP/U
YSOVn+PCT3VfDP+aKF4OQ7x47PlJm2d+KYJboj2jD2a0KD0vKTgyoELcEKjVbYrT
qyxKwQv0cy7BwxsCmyfSWsJEAC7DTZtI7PPhNaMjIwrloLussF5aUx5/KZ70XA0f
u8rovjID4gPYcpBlWEnxAPCSCONotJmpsTUIgRyvSoE1HY7l0CS6nPrG4ftJwu5P
GyxOif7jb7WyxVpNaCtvoDOIUyV7JhYtvZ7tkaxq5ylAZzc0M0hut78joQ4PHzNa
1LBRwq96fanBqC67CFqPk6jseSktjwNX3N09aFPDBA0fdWrtTtshFpkcvlonMzx4
L5m1+SCZcq1ytjL9qdElJCAB6mpllArZBS6zjU1MNepa+XuIanr/i6NExTdOWmIC
me7MM7cuojwQNX6rFMokHCCEzticzFwHigLcnmZnQ2mAtd5TvrPXPVhOp4Ii/jCT
sLEkO+e7BG0a7bFeTGZNk7iSzcqVHWbYPwGXr7pF7h1h0JQMYMcN1LU/LB3V6ZJp
2gkvDqIluRWGrYNGLsmBH7Lp6jyksLcW3eIG/vDUNoYCugUNbczgDQ8cOBxVSh/u
eVyt4vFU2F2+ZeYW9jwJG8emntWzyiEumAERqjfqCHCDkHR04UhHehnovUFGMAn0
dPDcNUyeUABlsYSWK/H+Yp09I/18j+5lE5Pb0xoGDz9qjT8D+XV5IymGWDH4aCar
Ywma6ZDFnRpxiKgGuuwW7AfZGoqRcVSP68K3SHMkIPz3Zi3P6H3teqw2YwGrk9CY
sG+z4v47jSDmVTfW45+JI5woE9R10BdNjXKzgpvnY35+6ydFuNM3IANIxpKyAZLf
JHNkfnRIjmQ/Ms1BhaO3H3df3AJGAQjfR0IAbig/vgGxfNLW+jEUH357JzZmssSP
uvRvgfeQy336MJFHzizXIBM3BRb1lL9xMXnmLUrtuCoo78SL24Eg4uUR0mMWGchn
wcUsaUQsxpmRKs0iPAt2/c5+3WjVzTpdGic7qdUdO/+bwK9paechttDB+wORQ7Zl
McL1H7whZDlaVPbjBkFTIY+gwB7LcRytCSIYTDBnRwFdKUlTRAtRMeMffy5q0NuM
n8DNVINGpP0OX+f7yL6veOTlvXD++eT1/0vdfiW/5f7QecDgbMtofUAhY5DD1WVC
6OSbMZQTeKKjfZ21sepL+G7cOdDVMFnfBwkEV/FEcP1hbnIvuOnXjeRL0KPkKOmi
OjOv9PyCuT4XeiIo48sKVdq5htHVqK00B82xjfOZI8dpXwf3dwZwapmB/bc+qshz
LC8g76vwPqdXB81c4IGaw3OnA1TwkaL18JLGod8nIiqbaSDft1Ov/ATOX0yEalaE
pYJEPH81J+BlJ/+hH6d1ZOULHmWsNU1NQ+0HFUkc49x01V5HyO66UKWoq6r89JBj
hK7r1ScmitzrmRHfvHJps7sJ0VX++XPq5L9hfU4t4ue4v+KRjtAdZPSYtco8nhnf
1R05ZeKhdW3wl/PbkqOIxnk9SmW/LXNtxjC+qI0l1bqJv6tQ6+BWM6pWNr2tRSS1
2l0v5kl9SOTpNSl1NmqOxrLOgJE9kjfyxMBiRnCjA3pNdXMcUB7nxB0YO+Q62snA
c9QRCAC1EvzAiULiG4y0dHxKB+QP0PcvQ9EJ42+NKEFPg/LgV3Iq0MIWSWjQkF+D
dy6JS4B+7E2q0Xj/WX+mTo77hmg7+MRTMHH7yPkPH5Z30AeQl0Be2hXFH2kNH/BO
B0t/vEt4BGxlgAvh/mRLmRBn0NARlHD2U3xI5nCyfbZ0lqwf0UPjQwiRKxteorEu
7pnM7koxLyDHPusgoXDQvwlxwVM0/sU3AlZPzQ7nt7AJ8BhxK+lol0nlwJXr5G+N
3SJQRRqLQUV1HDrtFtkKl979qnDgWFkn5y++pAC71QQUWKHtFNWTOX6k80SVsjTi
vtrUWWw30yFPac5TUVwd8YA/eXnXV205VQyylifUKDjGLtpCH5iT5qClulB0x6JB
VtyOBvhlSqwReIy2Yy0IF5JKcZ6IO52Zt20kKNeTwmaSfvJkepXjsGhUZmq7Li0c
/m3xNEP+0ni4x8sCN/as2BMtl4TG/f+qITDB0c2Wepb9jlYie33xpIJRs0rjfXF3
iYdUwfQArAecsqdEc3EX1xitWktyXTvYaz+ydQZ6D45R8sTsrUfK9ybell5AV/zs
Kk08RoP8f68+iDK20tuslRVmNRAaXipTEWL3psIhFEJsW9EUbEN/x6IQwRKjQsjz
5r2u+f/F5kiIHHJGe8/fDjw0OT4fLiLedebl421AnG71ewBu4uU2mKSyPEsDHPdU
XG/ldHDXfOcr+ihpDmNKm68ILZluq4HQqyHxYzplfLAWCKsVzbjQtPYiWJBnrVaI
pSiUXexqrcU+UO//cqAm2HgHe9Ib8BHm56wnISOI1X+4ztV9zZZ1nj+V1dtGEMkS
uLJIie4dRIiFOhBuVLId7A0UZtNSD5ihHQZVHw+/UQ7MlxaajvVZqGlFXRIUPbhb
AZUmSC47stbRIJ7+D77qQofwUWXTYRK5ACX2xziuU10VGfU93AwosD04JE8nc9hr
FCps9/QS1XrtMTqFrg2+it8bkFgRywpwIigqO1/O2D4a7HCsXAKqATMK2HbaGl8U
01sRsE+8W+uPdrhH7sr3EGJyGtYxz8uRpAfaMVj/3HgGeVGl2won52WDGop9S8hp
dTd2H942K6Za+RWWO1Ger6zzd6nyFsBTpPlhwkW1hPgUBn23/sGcpXC9g/ffbOeb
9Nlwb05uBIPO1V0w/Ks8FZVOlxMB4A2A+vGESRbQvI0oarkDxKj+O8P9BG27cOVE
DZPL6OCxFIWhTxF9bXMbegIO5c+nMM1NnUXucRP9pi2SKWmyvP4Pj+7r2kTvergR
D4+CXBuSxgPWatcmpxQUompy6IYap52P5wK0G5CQevCosQmVB/SgEi/ec9e26rII
wEM0VQHwZBMccQJuvssbPiaOq1WD6vQc9RPDEivfSd67JOMOe5Q0zwXE4Pqi4Q/F
TSezRW85dsaEx9baET9dJ67983hhucYcmcovALcyJSZFZal0dCnlBiwMV72WjRz3
vEJ9du6Fwy4RaiTZcTTRfaX/ex795vkBh2tqx5+eF4CiCtl24wNdnZtRCYl0F2rs
FMpQUiCrV2wDk15ZDWCrDtjZyB+RU/LzT8HOI/ygKXFcqW7xSKKU0doEVAngWFvq
t+0r5OcaFo5UNt868YlOe9fdPcfjPuTfPURMgFj80AKbFL5kq1n+Lfd+B/zkUwOX
9XgrWLivkRbP9pHbjwzFbgyUXiC+C4jkeCLGzj4YSjZDzY/TjQyrK5xZ/W9Qy7Zj
OsAecZrdt4jlfYpLsl6aqFBVNnVP+1IgygNNYztDnlafdOvraQb1AECVsGPQtX39
gp+CyCQE/H5ZJ8DuS6Bkv9GfyVCAg5G5Op+cSGzUPj8dTivJN/G76qQKG3UqxclQ
wVCUlykItbc8ytD7MXYx3SGAEe8XDXxn/CtI3qSRpN9VeuAzrBWIO0bztPzTfLYm
i0EhH5+PwUHXrycDnV9TcylfeiBdPIr62metGXebbflEzRGT3EGNs7gGTnCok/fG
BMmtZYw7GmX/SpfQs+f8eAez0BtXyOefyafHqFPIN5YPxlZKNl2ktmTHMOznSoNw
SJkPczmTPQyR+V/AlS3dJlzSWvLPgL+3eFFHGLJh76tN3apc82CLzfvr8zjz8Tg5
3BLn2fF+htxGP3tCO9tjjR3GtRkOYpoSYKViRj89GcAorzLXz/o3ccBQ6Y0WVwLU
nrXWJgF182Xc9cCPCMOn6KgMqcj4Drpq2Onj2sUdHmtXGdb0C+Osk5/RxOen8BdB
f2hezcokMKHksefqDzY91G7bNJsT6QFLZFwj28evfEOer9AErrG8fyuALHcdmXUX
8yMIyXs0HwHw/Wq56GngY3KpAdt1/TE3uzYbEatMf/mxES193Lx+Fy9c8bDCbusW
4iX+16eEZ8ZdWdZLus9CunZgduGms/Cce1vDc3kgCR+JCQ2IU6cUE535kfk2v10e
Fd9KN1DGRKowGW117S1CqXI+UydhLXcQyNnBDte4Yy0DVVkVLa1iR+fAmZiX53uJ
ouBCVnhjHzc1kOAG+LgNOnwKmDovy+W2NIv308dCDiEUt9W5Mrma83pDTrn6ROGv
5Ru9LdTZ4Xk7psLUa0txC15WidTqNyRd26s5kNkFcDMjMNa0Z2IB0txSNaEeVj5i
Jb6gLKGVIAOrpPo4TNhgnQZVpy/1QjGBP4Lbk5mNMTA9i+vU5eyur6eKilK/rfKK
HR31/R/n76wuEZ3tJWE08y81W9LBj/Ke0fUi51FBSDFZFNTH4N8BBG91V/NCXyom
q5zicFSpvtXHueadjkIx4wnnYCErcfZRO/wvTqgBmEMio/kbWJtuhfmkaN+EObWj
5GhWtgBd1sRTiGQQkRhLbBZZK1Htt97mH+tq36mrtjzKJFDElCTSsIvkvMu+ynZw
9McrokaRwrFi4xfseIwl+zYPL4LmcgW16fozJ99ghj2KT1EqexVikwxG1Pl2Y/sP
97rEkM/Bjg4LL06rVn7t8ioVNfASjX+grI6K2nEbjGCZm9BZcFOz/EtBBWYDlbdL
EwcZmh9k4vU+PX9TJVt11Ybv52gasI/tRRWTaPgz7j5GGORHWnlC324fqj9A8N8D
TbhcMIENtqq9431e0luPOMbXAjTpvlminSz2ZISssK1fNrt9tOY0mOfxROM8oFWn
JtNlWmJdooAQXq0YlYYO1wJPMEjIVr3mrKuaKwiEgC1QkHCE3lsAthdPGw7EuiFT
s6cKESz7KlKvOCmsLXpDpwxJRlFsFC0tZowQOBoSRNtszayBlBCtHmsJPJvMp+3b
RPoDtvYSG8FO3ybYt0f/21qbhX4ttrL96x/2GkZjydEE24GGvI4yXFyMh14wTeOe
gl7sD32I6c8WPp4Ytw5KpK9XsdvdmwxXXMJWg6+05YkEViBus9K8rEqEsimd7Ws7
ZWHYqqTjaOKPa/NG6lqrt50zgPEYbsa4wucP8byVPteuZBsOMt8x/YHd0ZDUYExx
tLfjBZ7qijCmgUPB3xSWWx/5Jo/2eBHtYdIFKgKXrO4bQR/Ed0y1+RfrXJx3/ZOd
0vLsxIoB8GT9eopM/Sgu91VpuDtAJTMexTgYWTd0tCPd04HOGoIxcovSsGhcTElb
ipC0WOcU46ki9Qx6K7E4BqLyj/fOLh020HBBVoYFtNYpeL2q6Grq9jIg7g4v4flr
nZ3O0mCgBsTuAOkIdpPQjZu3ZaXbN+o1GNksAnosXSoa0fgDl6YdrWpfkrOJmBoj
9MIZFw54SI0PYs+1H/BBQDCKZ3kyDVntkSKEtsnL9hesC3fk4SwpvX9fAs9/BMSn
JfbUdQaBaG7BqQCZBlhBmXyYN+ap6tyEO8iCzJSeB0Em1rtVwaJ+v09D5P3igI64
i2Rh0bGmyF5ZS7X6qjGPy/wWvbsqijsa4keHoqbXp7NbxIYLGhI59QV5oBAUhOWE
NmKgXwnsX0ratu7ySgA0UgycsMZP/ExcuSNM3crYcYQMvZX7Wtgx6KMqi+9Q60zR
bLSD/1Y95UZXRADTc0HWiTfgrFLvBV8tsVRxGmN/pVR+TiqOtul6JASwGEsRlJtL
4ylcQNhrVm0yC9LciCXbx9iFoLdhKuaDILqUU3Lu0TdSmWMBmw6swztti9JVOSxI
3EX3HvqfhrtjFwbGm37s/P2O9DuCIcdeL9SVd5PAcPKDYlzgNkDzWMJbf48Z9k2q
zYri1EKaMwXzzs6zWCIcUKg4qjmGxuxoymJh4VQTf49IZ9mvE4wNQ0/re5ukj1lh
si+DCNtTyji0DwvdUUwZtIWSyMCZUO2qUgGcV9JbahKcJgIrTbCpaAi5XtWr0p/H
0P23GjMw16+LHegGBCwjzZmsshUVKUo3z9bV6yeC+WNy5IZ2lwivkzhxASRy+xN/
3bp9OGGdbJPrpNHEb92Z7mtsFoJk9kRZAnTV8v1oMRUZPiojx7yQXyKQOwSLetjh
jvUAzOYrbnTHme0yE9muxyCDuCa/HunWSFbvw+npwBM37qqar23//xdsFw0ZlLCG
VguovwV72e3+Kp6aI9x1TNoV4Ase3gnzRJGFnLOagfw5w5BX/XhNFMtcAiKik2jC
O8K8Dnx/hGPe4yVcwUQf10GDDl6V4QuWma3OfgV3UMPXW5qUB1p91wg3KKZknOOn
j5C/5wIns4quluoU5oc8TQV/09hoYy3yRRuU8dcJebZxtuDhPeBnVDjuSGEC4g1b
HxNtNN2hAc/mEU30KvyPwJr3AytWIiplfgI6jUmrAAc49ULId8DSr2I539TGMnUJ
sxjExuVtHrxxGEnRHXA1sILIofZnOG3aDjMaEIN2tUae6h0wcliKPJdGsI8Z95My
/29PmbJZA/4ScD+RpFsAuJzJLFdyeAuRFicwdTfHWRmfdxs2yqSCyuMP/0Fz6jt3
xmWj88n99WMhCEdK25Zyn17Hja3a+2krFnahURmLITO0MioFgPD0vOiyaxGdYJhE
EylVyEqMXk3W4R9bLlgNpANt9NOQZFnIRNEUkO0FRbrl8g2en8AkeEE2Scp4UO7I
a+PngF0HaZQ68XJwHXRM0sjooyuVhXVfFmTPNG35JFRGKXBy1e+9A3P4XYb+BZHu
XjrQ95eK1pGb6cREzyUpSwoDehbLruQ4LIBget/LoVbOt1tMwswmMEqOXNUsINS4
VZGvisvNbr7HpuAipRjBiFk01Dq19Gid0q1o8PequvbnX0mkRhRqd6owSgd94onR
WrdtiJkixr6Ff4Acxd8zHYqGa3msqNVXIw4NM6eS2Bt9YotH4FghSzZw3ywZr4DJ
USV1kMhsVHk47+CDgMHbRft08s4sfWAGiTcHMbFVBLfJTWvZyeXup+VhrFXJwcG8
az9uPM1Dg+FEEmm4xILg0D0tkWrZdkqiM0vkI2tiivqxF91c6ziqMJkd/bCWRIrV
h3yvBpVM6zlgZzXk8qfSUxpiev+sLkKANaWTfjy1rrWiKbWHBBAloKPegUHsh9QX
ajMaaaXVoGtu45vkaVEh2TUSHTjwH0Xlyim8qdSmkXWTVb5homSdUuIBa6kESpr6
xR3O9Qf3pQOKWMR1rdHU0cyXH3QtVcLS/UBUJg/ImUFhWOh3u6echEooRsyFCMXZ
Lr1bV0eNJs/zAVN802cQKVYtqRob2ms3Qd4Pk/YnuR4y4Y3GRdTz48TXDPfZw8I0
HwTxyHPWTRm/u8o3MIyqSlkVVeHYo9Rb6Vyweu69wQd2hy1VNX8lTuWV4eAgiDCX
+0+5LnybpiBhAChlvZ78FrhM2BaalssKgfYSsTm8xwBFcv9iGELXbYC8miMysGRR
6UF85hzoY/DZAYe+s/xuuRnLgcgs1L43sC4aRVEpfzQilfbwXtVSw9G3IfhShS5W
z1+CGfqumiJEia+GILEMPnYVkPMxKehLy4usdBzWAtcRNPDE5flu/CpZSn102r6j
fmJvCqBZiDovCb4qG2FCo58G3UaY7Q/5xjvNNeg8mZsYPKSr7tkgjSawb7+G0jmf
rN9bUyGq/LzaTB+uke2aAOqfiSvJL2tm0h0QvHXqBPeBxQ8msWyi2maa3GAZt0tY
yJSifvAMJYUqdqNTYRCK2nq+qOivc+AgaOmTz91kJSfnEzFHmqO4cVdq340g0CqC
U+/kAhbZvUvfpDsqd9J/lRf363ATjj6Ln819HCo7HsArbgNNMZmbY85GyjosXh9U
22Z637/ydqX2t0iDslJ2zEjeruqW/ZWJnsGFOYjz7yaovabshu7wq/f9pVHRF/A7
MtKKvfrrAo9L45l5o3YbSAzK8XyY8zpZv1kSHfiyS+CB/WFCNv/2qT1qw3LayFZD
sSb5TyOsz25JD0Acd/XdxQjtYhBNVa1tkOXFOUmc6RwBO+rqmcHWDcZmn1FJjRr1
3k6VtKghq/ctHbL1V3EKc9ZVAtLeYdpGJMCtzEJ1fDu83jI8IpAlTQPttD/5EYpU
q4fuxmZ9AaTo+VapYqMnzZkg56Qf/jM4jQPTnqrH10Rr26xr9w54Ckoo1odAJX01
uStHnj4af7XnfQgJ0g5cEmHhBHJtR0m0mj5VbWFXR08MzXLie28n4KL/OZukCdSF
vm+YrN2cPUnviannVOY6Bg+OL8kC3zo8ajBcaTQYZZ5+SjxeRU69KUCsWn2uby/z
b1DYVs3+73GgxE0dVV/8bPSJQabL+SLXKMDgFrqTND2LRN7Zz0/bIIoqaZLmgUJY
ilW0bF6bbbP1ytMTVaXRuGfqcMfejyNmeyGVGczvbkt5GU+7Jsu50UtM8lWcakQj
aNq+5alu7it830bW06478EQk7cNpJ9bak7d64QCCepUIOrR9ZwGwM2l8fKTTkFd5
SkW9dPZmbvigNO5NBzTyAqjDwbvxX41idz7MwmXyz9wix/+ef1Oux236kJ+wptyC
tNpHKFCMI957XJkzgdlWmr1gYiEV9OXxCpRSW50FQ9RJlv0ooGKB29RasAEf1EFd
8qNN+Q4yOsrHiIRJ4kngJLkugPeLZ9lELlfWl550esLdyda3FqevFcQ0gBFsVt76
zP3APBTjvzINkvNk2TwlnHmPu+WU/AzIJ+aFSgExUS+PLjo/zgI9KsfKeDZqF9xn
/jqjY/EHu9ilSQgC+ogXA123VQlFOK0k74RKzrgCY1RGNENXstrJdN0/KHxP8Bfd
Rw9hB4REwFgjfUzHD9DhtCZU0Uzm4qs4BrmJl5BmBBT35F5Sk+b2iAYbYC0IeG3M
ImXbf+vncw0KEAm9cnkfOtZgbiWpNmHUBLtrAZrg/wSLCm4C5TzHdB95KB3CFUfd
TezAb+aNe9Pj22KAo1DROVXlSezwY8uDlczW4PenNFV6pe+lEPt8AoFarlF16HEA
JsYthHoJUqWSOp3a5N8fLsVhdPdY0Os2pCrCBHUHVatwN7l0xZv7wbbcpyuYclMM
zQI/iG5fo7kdjIMFRRvq/7caKHqORJhdiJiAETu+4olMCz1noUcZpO1ulrvXUQtW
23d65PYFZfzamCLF1BV4H2Vprnt/U8WawbxNxh1Ws2O4c2l9/MeEOkQTIb9Nv49f
xTbkiwQ13mz2CVHwQSrt0Y4HJH/dBi18w/ERLbCM0r/Plv6f9m6wtKSw3E/FhwJT
Hitbip0klveikBl9hXrk3YTogQtBoGU/Xke02smL2UWeenqaMrbNkr92j2JJRpay
3ODPsv1Eifu64IKRg5xpi6sI5jERESlyDcvUYtwgHZhWW/Z4ThRE2hauj+EQU1Ts
Tud32KjE/HnQslv98KM0zb+D4pO/kSSOBdFnI2wjMGGqyolGS4QQ5V8X3dhdLYMM
sXlCc/e2zR2I8zZOKPm/lnuFOhPvw6zsZOAqvIbeDRXXyiGSH6ATk1JvO9H25KJR
27HS99eFq6chRVuK1SXbnOJW3y7gz4bcHQn2TdRC8auWaGbwKUZeK5A1WAtDo6Ic
pncXX3Ci/Bnl1vUElwkIikC9jKqjMc2lJZjV8ltt2XYWdGqTABzy7fqg5m+SFUr6
+oo9cxFTQ1LXjPrjcv78ocOBrOiUtJpZcn6O3EDgsaagph+xSJOCDaFKFkizG3fl
DUJ5mtpn3eyDAwo/Mctz3Wv3eWadQwqMmrAR5xB74bihh6laKaHPcxzPBkbrPAod
nusnSwn9OYwmbHPiPA2SdBZdwxCtDzSbNvMdBzPXB4xv6al9tiMh4w7zM6oVXMBs
urPYkHXDZBJMS9R576fAShraOFjsuzD8yLAdTrP546/IS4BtOjEweWXmSQANAJ+f
8YWXfEDXaC7Hg9RMYdGiyijVYXwM16Qv/JLza8Bj93eItqpfn+fOMW/3u7wwyn4o
GMVcWia0rN5p2iOVctvtYfPvcpOd7HA/8+Sw/JDGH+LwVQJiYVYLuv12HNSpi2nx
64v5H28x8r/M9mB8i2hE5O35ZdMe3A+H/d+SZJBpUjVhjksHUAsNCLuVzLeKvPyo
XLOemCj716Dy604kY6C1FWKk8ZHfBI0b9V0IFdgzQtndceiqDacJXDukpaLpeANu
qCpFguucopa5tQqOiOL3IC+exzHuksZBCcPBvwwJv69xn9g7P2xRkxklbFgwQHF3
wVsmgFPf2LUIbpnCuyOKBKf9mI2aJGL17YsrkuLWpjcK2bqequIhGMk7IlJGqChJ
kCqKmkp1ZI+wEPj1HUwxiB75xGXgy6cna1E9++Klr1ACNHQ0eGPpVTCJWl/Sq3qB
CxFXuLXOv4q/sHYz946TUvLuord/YIgSxLeDqNM5YYjxPozXSH04j6ssT6RhxUcU
26da3Qg8X55jXYP14Hu1d7cY9EAx/sxa6pvV7HYUinojpxZUeM7/zIM10cVzuPrA
qSgemzd6j2U51TsjG/nZhOOAYHpdrE5JwwQtKcVyoSONTgAh8BJyyiMLP2Eov1wN
g63GZgvMWbkZ9yFrktmDP1FgsPPnQ1E4aJVvnEWW5Lew+fN/603U6kwnx0G/WF3i
gsyOzWTwe3iCNA1TXQb2OFMFBE8iAId8fD985scfGQua0X/nUiEP+p4c5S4noqYk
NEFRwXx4ZVfKkQ7lBdcrgDVRpTzlkU0a+j6jROHjH7jbevyFcQfdT0P+WIMf8uFz
6lGxeprxZyqw7UVHdJX2JEiGty7xhZWseV4HoOs6lwYmh3K0J1ha4C6gyPJWOrDx
bMNAB9UGPet8yKIxXbXZlCSGK1Phq81iQje+unsdyvzmee//bKJEIG2hXKRD5u8S
wQPuLNyGJzZmeNJuI42Jd6KFKIjtIjovZNxL7Tqjx4JKROO6pLCwyFlsYNMZw86V
kXdY7WjYqfIQBKAnuNd3wqgtcnIeVSfLVbtspi0JbCJ6i0joQx1NVkTRIiukjIdu
VaYPjJZNbewr/cV5lH1BuJ/BPTCr2UCvp4305vLpb7QD6zMhqCvFfhPWzRjsrMoS
ohZzRPlCX8bpAiAO56VZihA4ZZXUS+DnqYHymn5lm7wH7bKrlkLhAhBU/p5+OzIf
H0T1ao75jMlURkGxGmpmUJeUmf+msjjw5sToXQxyzHueBxCk1ZGoICcC3L34Tpwt
iVeNmBecncm1Zp+75Ptr8Sr4llrl5OBJD4FLACn8NRF8yQEYM/gPPQd2n9HO7tFP
H321phvJaP9IMpnqHEFnLZam/yro1RMLM1pyklKEXQwcMaci8l3vpO0zA6X3npy6
PD686Y3r3x2HH7kXs3XzrmqSAPqH9j/0OkFaP5MKLWO+IFnuJYRVsXfuKEEbNJtc
7RWOtD0thc/GrZaD2dEoXJn+3wmQELj6/XEvmMQin7ACZBeh8RWdttXlRo1sNKe/
odSToJn/hAXlPUxFf5itnYHaXytQeRZyXWtsaWy5+07uRI9RZFkB+u+9Z0g1ih6f
SAmVP4W0BVNE4uzXo5MsE3c+KEU7FnLt3OKPZpsMq0tQS2VE8IQ20+mxKRGlkSAm
v/+1SSWO8LY+UERqBJMobQwWr5A8NQUltmVL6yQmuNITJhCLTxI5LaFo86McLgMG
gPkC0J/W9vBMS9PtqnnnA6Oel9xCT2qjmCTuHmcBbmQkqpnG7DmrRupwyhoTQluE
Jv0X/QyVcrq+ocysVAoXJJCgrApYraZ/1F8ttRfYwNi6vdFJXTYau4uFdSqWYiSS
G8s8o6+vIg0aNMSaBBoV4Z7G2Cdn6cN+AVv3QWWLB/rohfCzl3mVQIiwMrweMoSk
cY2accHCPboGo9jgyk8Ig6LhOVnTQUbEkpB1y3O2Wuk/xGyViOip3zpWHOkS+sVe
fgDwNa2EgVK4poWswDoxMJYuEbk25GM9pHBSiL7886/hQ5l1vq/0I9qLuLLPuikw
PPkEn4bAfAM7aL4oQUflf48x7R8pVtKk/xBmTdAKLU9+62QM1RU6Zkvwyz3LKkEi
RFPLEfSB9/ua+VEOHYZ6pCP7zDF7RcPg1WjIf9HfTAahroSA8iTYUeCiXLZ1Y4Lm
DoOubWJxSdNSv9NlCWg7jfGgP+h9cSldyOHUjv7PoQInIiR5Imuu4woMSwrj4G/N
A06K/2lohr61A8/32HiO0pJubtfy9N/mN74l7dz+trOCNJqQqHC3N50V0LJ+VKgh
nFQWs0gjzHWjV5ebL1oRbIJ+1i6B7JzkzcQEy5OVLK6eHsDoz8zeVEyRNQWWgk1/
T90t7g9WRRo34hmXRb3kuuyR3CtlqYym6xsCyNLUmtl43iZktRRSluT4C3xB1fJb
IpK1e/t0feW3NonX+UDIpcAX8spsF7irMkG98n+SNBuISNCCdKBk1J2dVFNKfaFn
UYn79H7GbwtfXkiqD+6XwDPcOnG9u1b3BwJIi5y6qnKJJqmHWOI6YQdqBorf9iOx
YroR2Ty/IgoMsW2m9eWbzCSc6NKsC6t6QsNrFmobZ2Lvo7tB/n/qTqE1S86nu8xB
IFJCQsI9XFYFmpVklESvyYM2cLlhy4aDXu56Dx1zA76JnRiWCOPkNensC/vS79e1
BWRuY0diBeELKegUr3JuYuvSNQ25Yx8mrZ1W/rMWBo0foouQEr1HLgnG+O8AGziX
grtWBuWSxRigR0vzxrNamf1+BojssXLKP+UAz80whAWhs1CrAImRtLmM0p8R8yaG
YsjwhIPc9BRTNH8C+mXplHnAzD9LAva/WVTnWzfHYKvc+DFOWkJzbhNgKyko409O
Xj3LsIPNwq4sp4bRCQIDP0YK6XmQFnzAw/FbZ7NqDEATn9C7wmachwsAoYY3zWWc
czPRBhmtmP3A8m8co1l2Yu66RXwfVYu3dnYSjGa3gsi3gKJie76Gz7k9zgwlrn7a
aRg2vfGXsTF/x/tE6JlDLVVJY6CBCE3gB4dok3HvJCGDVHmLp363WzffeNWgNxZU
stM4W7Rzf7RpVVHAD4AVX+R7Zz7/0T81eVZSPXoBBrR3zj/FRTQM7wJ5hVMFzfXz
Axoi7d+fJKGjQD0QTBaCMrKoO9hO2R3GkKeH5E2TA3lz529Kaf4SLSIk1I67b03E
GhlAwtymZm35Dsw88/Og6Jf+6AqJpsZOLMKHWJ3za1MpHLWxetdIwbRmAooauWND
nwKzXIcw9ZW+0jr+qU5Q7Xk2FMqaBtU3GfmZCKxV0qX4bY2CSeacjf5QV+Mh+gTE
QtcHAWiISB5fcYVRIEhIreCUk87UKWVjRWp08AfLJQxmwBj1sXQCW7norMh6l5RS
YxMqofRD3D1hU92XP3sA8ewZo5q0Y/JhsoOk5dxjlPZSCQQ39Lms9wu2hJp/9U6C
qVQE7pY6PzhKVmhKqLNDPMfKPBvryqlvBo0oIXswxvqhGW01yPNYU1K3L/fbR1AO
ljbahcG+oBqZSNDjx5Jurgs6nJeO3RHXFvOLZcI6W1NEaM8q2243wl8BxvKHJ1g8
lExxdmHAFHbMhTogbDQfb2PCCKnJ6E66x91iVX7u0q2OyaIVs184zpkui3sMVL63
qE2fUC2uM9ZtsQGynQMoj/Rzx56OkWP5UcJ1PD4+xx1W7GncWW6+8Rxkeg3KA+6H
o/Fv3K2Qf0kG9r1n5k1BjyaWD2JQZepGila2LwfS2igXHvwCrZAXj5FK3WQsmFw9
s4BtA5Cr5y2hWi/1xhvt7eOzy3WUKYgyebFa/S41o1OIpxo2Qg79OyVuo4Q+UxPp
404XRVMaxVJ+0XWFSyFeYbTOllVigenzp9jcf0g5x8DBKiB4LWDvqiNT9A9SHDJI
T/KJixNe99UmgJBN0NhWh2ZggEhB6RJd5CMAl4NKpljlZg7sCtTAI0ociBPw1IAh
rsJzqle9lN8qLWdEHhsT+nWTbiG35NqpEvW4MueTQrKWaopg+eVKbuDZGpJ1ACd2
RBREavH9YK4YfKnel53Qm9kvKICmlNmZDRfIfyjq8aU9HeNb4r+EcmxvLI8yJFmB
QuFpJ9feblDMMOgRMEwxYtphbrOpWt6nIquG/5VCegWyTe9RDNKJuAeE+sk0I+ni
EHTGFM9BAqJgOE8s8laJOZgvUYTwU76BZdsnw4Hg3O/VWaXrOhzujEYbch4/pzyW
R9i2Aaw/lWl4BVlkhITjO307FK+Dsy/bavWEby3Qb8xaHgvJTHNM5Q5iVrcwsaPT
IIDk6Hmgn4CG5hcdTcJV4EG4mhJa4Xer1q+gzyNmlj4ydpT+LDmg3EU5Lm+WnEnJ
ipnMfhdc++M1Sa+NReKtr5wBvzY7dLkQcRdDZd1dqwwlUM/k4W2PsVZqX4mPPeGT
nTqvytub3DGo6ZjXFAyLg/9GfTWVsSWFmmaCjivSqpwRlYNnsJ1asq19yEjZ9lyb
+JkztpF1dv+lKP2zpLZYV+ZE5cRpEVXqU6nBLK9+vWo4HN8NAPI3Fzw9PVHSBVv4
axGo+S07K8bGoP2F7hrXUmu2NxUB31JahXhMPqiGtZGP3TkCbafUTtR6CYh1Kkcq
P2nnRJJA56vjuMu7RuuMcbnNtd0HXPPMyrFPdqKtsTV7uZqGF3Y47c0FY6sSZEsW
Vu8a714Exzh0vRVQjn6PMo7gKIGdwHGWyn/zwwfk1iwu4oG/2A9jC79NNOsQKw1A
KXQbubttrbdxo/arYSIiIjogzqQ3HZl3tSiG0IWOTMBARsd8Dz23bkznSfK/pFDN
p0so12PnnDJS979dl6cSAYBaoHlr5HhrR1SnQw6mSvEmOjG4mwV09YNWfEmsarNs
HaUK7LZDVCmQd+lAbWaP2wmYFu7f1UoFZgTZ0FqR9w+l/8Hzj1e2Y+XPkVZ52eST
s1nGQwHMjyIINhjupMdoZguA1WIxhoaGgT4cSdZ7SFAa8UeGcTYcbXuBcyunwiQc
RaSiqEoydG/3RnSlowppUrzA/Ka2PpUy1MqZh0e1cmGL+rwDMS29S2oF6HMkWAqF
cti5MX5wJ0m3bsNbAhX8iaSgyXZzC+C2zn96yg/XXurwiZG/mn5LS9aq00HHyim2
3EhxfYbW6Iu3rUMbJ/0Kky+gbT+Q9FirehOGJ8rZd+kLcsivV6AEzpYf4VAJRSk9
ZFmRugwzeWn71ux5SMzQ0i7V6RSNrc0+s5rmZvh/0jjUbZxw/h0IsAmdOA5Ky3fB
aO1ZHZqLC7rLNR08gHUwuiln/P6IytUEQfi8WedlwI4QpKLsCHJoVk6mBVX1Lecc
+sOjUIbS4GrktNYwKOZo8+12qcFxpNCfH4u5UoBIF3KXdNefOCCt2AIEXWdad4IX
kRzedKIQ8aswU3E4+OZytDTGtTejr6wyNC7zwIXjRp/e4NZr0PlTyPrOQJ3HaFvG
XqlT6Op9qKfFQvFfBG0bOHX05rcGyYClLtCSQe4WhSN/UzO+PhDaa3O+HwGvo6vO
MQyvf+w8sJ/QCPjbmm5rDRCaQuVDch6ocAASjpSPNiwGcqPrw7zXvBl4WPIdDTxJ
/A6+BW9FHX1cIr3tnpBIV2zEiXYMyFqrnms4TsNE7j5pDCYr8g6SjJFUPAna9cIZ
9l1EZwA2oTPzAGN2mG/dwq/5Xaz4gaUcG0L3tmqdoy/8oSpHUkcOQbY1NToXhvV0
MQhfPFcbsVFrMsvNMvUQ6riWDmFvie3gQf1Z238YkGOW+JrZ4x2zkLVWZF0rBgVa
G/Ba3ZCzwlHxCWOvjdBIWaknDpx2gEErsKQkyQeAN96Gp8VO6i1gP+2+p2l9i9nz
YYVM6YBfKwIlAGEyOqV6AI1mgwHIazHOjbOhvOevWEimbyoiV/xqpFEQhGHPG2cT
C1JUvRobuXFPGmXI+wyDOpOSbhp5VOQlt/F7Az2dYcq1rx39pG6EyY+PDyOB+2I1
otOxlCSsu8Zm6S7Y21qwu/KAG0v3WgMS2RMDtI4cp5hgEW4vNkGM5QtpFuwhNH6p
QJb6OYdCLEICCbOTFA94MAnijlYcUfl44I3ms++t5XLtb05RM4lImnuDXj4vpnzo
p6uyJX8iXfVMDIU3zrE8GRRBJ5ew3ETKxZx2hrt2TEWVM3tHnr0J6Vc+py1DUa2y
iTimnR5qs95HdcCmY6ZyynYXhcBRP+SJeO1b8jL8U+iTNRxwGfeIxq9pqbpFCYiO
rMVXI7aOMq4Tmiy3fj+sswS+xJXRoPqqz/eRrsuNuV9Ruc2jsBdzXDZmPgeHVOr+
c+gwavUgTTA0l2MJ8BB1FsB1JWRnAbppJz74cj9xpVjZQ6/m9lwft52MbXiUGMu0
/N5X14JkLzIyfM1eYD0LoWvkjM2KyouAQAvBCsGnraD/1/y2c+GJBQfRnBoi8CpV
eaL79kDFNYEgL285uQ3IUknytw7V+36FhYvcU+kra6Hu8mdO5yYC+Dx1opI3bZE9
JShaTvvXEwO3E8gQwI8ecKkIJgSd2AoD50wFU8iLhoPHABaX30tZmUfstvBpfM4e
tOg4xT8CM5AxMWXNwVdwO+PcYXB105WWccIfy8hn0KXhosOLZUJKFe6MJcYTPtKE
ILHTOYHqja5ZSOnFmabGjckUJiij+mZPKcXG6Dk8Ui4eE6Kh7ToizrfNywm4CJkG
iGQB68xTVCRaroHyP1cUrYqyQb72WC8is8/xtt9R7c7gFwDaB5TwVTtYASmkBhFZ
87zwIU3vdZwVPk8+xqcEOms3hX8+hO0b42HE8+vHp2WTxUTJgSDZRIYCdkG1exfx
FiSoOJOlKPxux8TYjQpVjqZya04GVA6z839uxgt1wop6M+9Dn/ynZOkI9pmcjzhG
SH8cJ5c74NqWz7mM0SEc9zSMzIVETUX7XzRZlI8fxQ0FJ0MdS4kzPpIQQwRTpU+e
jWIWQlATilWJUIkz6/ZRgPkkf9CiK837ugKmc0WgpqEh/P2LVO7NcrDHCx4//Li7
SoWlLk3hu0wccvlDYg2VKvULG0BE3xyQ8UTBYLz83Q0g2LeFNfy0Co4EOUNUcAT/
Yru2R5CMnQr9Npu/FralHlehqkY5bIPvFJp/Y3xJOxX0/3KgURD8lSYO5qwEUAVf
eFCtKWE8BwP+myh3Ys0uj25dzTPj6GQgr+T7cRvfBc2vaETHATCJEZUzqgR/Zlzj
LexBmeFYv+H4pV1JGc7/LfFHNYw6CHMe8xNqiqGcqGoQxQZsFGfkx5P8LxDjet4y
5PEFgbPcFZH62YuV3LU8c1X8NkEkuhs70ILAvOdwz4usQisVNwMxqXTWA22ra1kA
JHyXqM6YMTDU/xOLeU6DnoAZUEA4cRgn9hO5qvrvsKeoNc8o+w4FqUruGP46Iul+
Hj4ehhoa6YHYxQQL/vP8miynSNyI+KrxRGFkWMaTo08tOrV5li7Xdrp0hv/aThFO
8qrmXUdnpIkV1HZhvt7EjS4C03bYDTR0Y7QyI7PGGNOxqIX9lHiIx81sYaNtTrnN
SWlkrx9f/cnYf5sAeOLMkuKNC3ST7VLlBFnklgtErX/VmhXBrlcl+myqFTomiKDn
tYDcDaaDi5wYWGQQ5cDUnBKpB7WJKR5TEEgWT443ZEVaL5HS4ueZ3+0kAHwIrGNa
rzI1WYVN9I2IpFDOihrRnYaJ9aoReWfIZvGCJiOvP2B8ySfwdPxZQqfXZ6+HEQlh
sIl71XxeZHjdkUTTvHVEHe8KIBYtnbn9ZLkdwstM34T3my9DSmRTd16ngZouNIg8
PMY29vmUMzbI15l7EiIDsfiRLtnztY7v9IxvTnCqkbTtqCJUHAOBglrs2ZwXK4j7
BkC+Q/dwmzTqIxjPtavEvjNF0GeiJmXRK6BeoPbjtC5Zk3TEAIpB+HsH0GwQiqnu
SWJNqAxupH1C9emcJxPWaLVQKNZF4ZXNh4Hmg8WNABir5gCDnK1EEWNdVy+PgZk9
F4IsikPCVE1jhAsB9TIf2ZL7g3pvhSr1hvf5mDVrC8Su8IPSbHQLCr0MJrMg+VYm
2xmqYXMe6juGvMOoD7aciEgI2FcNYLt39vcem0KT5O9+15WsVKuBe7tY5S+T4wfA
+SaJysU+KvjR49qb33l1DV50MYAzDhOsq8R3K77eK/kqG0EAplAO287XyoV2ssPC
+EFYSFYTezM7dFUCI0XeTW8ksdnE4A3vQqeDwJLdghXIxZa7duUGknastvjDRVRd
UP0eCqXgprMYMyIbKYFexWvxjTLYoLN/D806ftSBvAwYnlduyh6MgAzi4iPqLJRN
wt1cuaVpaGQdAbnO5rqU7oa1b8pN/t+hXEaE//N/p+gLCj8ODQbrWZqzKbPQPejX
zF9RHUrJ9EBtRjLq+zhEinvvzDf7j4zDJtVfpuFnvyD4kry4HpizV6k7AqFAFD5l
z4okVc328rrk841oeahaFLds8qGj0++ahcE/kYYZBtJfYRfFYCthk6NHRDLQ4qrE
ZjxRvgj88vhyMGkcZAtdg1bUp+0Pbs77Bcq0vbKCE+8QcprPM5JDtkuHLpn8LXgX
1qMScE/c2H04eGVvLme/h4SMKzFJld5wz4ZPZMUVbwGiguZPHROMDzXND2UbeOTC
yon+A/ccQd6rTQA9GxguCvK+w/ZsXJiXImOgPuu32ekXgNv+i3tJxy3ILSOYMSrz
6Qg07I5QfOakTSgQXYq9x1f9uo424gEp6B6B4QKfdbB+kEMZO4k94JK/lpQq20Gc
q/2QdfoDdHRQQvQBRIhxXRdeTdYz4zkZovJ9FMd/HG+pdIipIw05CRsLx9gRioKN
s5kp1XLGew19ERHznqSDq+dD09Muk0kQPnb18+ynlCD/RdHZp+BZW1MAv5RXXKxV
ETYYJ8ZAsPfX7v7nv+mZT9LnqmtuWn4+zlYEUOfP/L4O1tOeZLGzvMwN3twEuzAg
RDeQs80QSuasI0b5SQM/EKWuF3M495RpJsB+FwRoKkoDtvI/d6xFhHX93MTgM3ki
+u876Qlu/xoOoUFnx3Z0PUX6Hb0PtsRTC7hoLhF77IyqQpDNqlFIyzTCXoXYA8KN
nH2XhhkUFCr24PLs8EYFCcIN0U8dgHVWMLeqzBF/DUbe0EYob8EP57g1hEg9bYsN
FeulkVL/ew+0QJCyWET2m7ij+Zhdiln2qXUYSSbAcviHvZmg6QK0p3G1Pg+UDpHP
G7Vukk/NiGC1jWA22JGQCGBGIj5j9sKPTsfgNp9HjrXexfvJyl+DVrCEBiKmut0H
3JhY4i3T6GcJnu4wf7CGFsJr0M/Qzx1SV3mK+0IHsIOjio82K+ZjeBkJZcBkHIPq
uW7ZypXRjY5tDa/m7iEeK09jAQf5cfyQKeNBou8OQ5ZoCAnRW0UDGWNFKQiiZzjA
zFonm976V/CzFbohe0Qwsp1cu7OIIx2tdZa9uvC4DI4+I2KtDHZyhe8FV9N4UHL8
HvfB+jzQaCkZGw0I3sKzuzCARQ0IQkNX5QaLi+EThJhamcwAWgYSarhgHtmEENtv
YMixE2OK40xyhua3qEi/URzXhruJNCXWOGEzOpqFN7O4IeVpIttaxWAi+ykICBBU
r36CF9oylamQAc4hTopUj3327Bmtgs5YcCmdRmX9EwIKkiwrYCQQ+kmUk2bI0n+y
8Srn54So4bKDGWRVy3C7V2xqfBZgQ/PBtFcMpYVUs9ActhG79qZJ0DAq/yoqcYAk
sZoYvQm+axUezLnbtNlTx3LDFPLvtxVpeKNcBB14+3DhJdA3+xvvi6kTQsPhmIlF
G8m2DKFQcSiFD8TrcTjW8r0CoNiuSEB0wSsJjG80aNpcGacAFah0Z/QLDpupPEBy
P5J9jnqGwxv6Sq0PxJXjzqp2bNT/lxIh0J5haVviKTo5vUIs75nGkjC5SkpLdbHI
ARA7E4uwD75Fdu8B4HYbd6jBF8JoRHrtkurwb+Z9poLzGM+lXtBYrwZP4WIceu4Z
KxcjaxaIR6gByREKqpr+QzHh/jkjVXl2lhBz/GXEb5JlusYodT4KuPWlXbKqCHQR
QNIbKZbZj6WrXCLrslXEUViBrGYYml6UDfVPEpY3Qh32rwze5Y2nWD6nmBaKHsO0
JUd/9XYkoZpTs9F24qvYnBKSAI3/udgCOtMbvJD/adg/f7cdqKyjoK3cqIEUKLJ0
q5Porwff9EJDQkprztWANaOwTuX+V1BbWcl+RQbXAcW8oim4iHuH7xnBSO8C8Wxl
poE56JNbzXhHtvzO65/Fv3+c0ntnt4TUQek484xFgBXFuMOW65ROMZwIKdrL7fjb
x91Vznq4pZ3ct5k5Dbw3gjIN3cBRZa6EDv7ZJKRfy+rWgf0KaOaNlWgfg7xp2BTN
iFCbDEkNiUhfS7CdpK/bVRMEoyaGDU8GUMMpHgPwMstmeKTWWTYKRcbm26/WydtI
dhZxDWpdPhFEC6s2EoRhtoCHl0SVKub++yn42y8N262VS6WOStvRuPMq/7stWK3K
h5QDtVjXbP+/sb2sn5EiwGmVU4TFBZoJt6y+6J+dn7mvn4HgV+ASMfiz8L8m196G
Xb2Yp98sqHbIkjDQk1v6d0aLrfV8aLzurtFvx/TKSKFn/3ux8WJXgOudCOYtu4YE
8H3HS8S/VkDHA1OIIXQU3enL2WCfn6DC0ykARBXOCiL8KCXWv+ORqDvNQcLb3Wv3
WF71SAGviFEG3RdBO97+PylgKGVeRLgMD8MXuF5az8zNvnR13xf0r3ovkyNc17Nd
NFuEltbU2IGVVenZb7ZoFsJLVfrz2QEvkqn0AFCFZBTq56x+3SwHU0N9bam+ILgt
3p+G1nxaFVAzdgECU20p12qwDcJd0KB4DxJ1cHgX5vkgcdVXasz1olivM5FkySma
VidEJP1ufj8XV9/1+O6XbMtTZ3CLyUl9bH2n5AvB8inAaQCq3OqeSk/us27GQ160
9CXvT0RZjK+oPBFbbEG9OucBqBdm6Fy+km6U9vpIdgpBZ8npSMqxC70sM0igTh9m
oT9aDOIySBIEU/UTvlyUBQAlVgTchT89ktSBrSvklxZsvv5s0BpZyFHplc4pFC4r
FhLzs8koTFW6OvjKWOKuZ+l7Z30bZKJrusHkO8ZdH0949bE45LrI9v8r/AinxZlp
d6Ppy8Ei8aVVbtx1Jx8fl9YQv3FULTTDv6oi7RePdAmIBQV9rQBu0DGkbbDkVxaF
J6/dvju3XX9vFzYJ034lILl1qNW1JOqzP4gWaNsk8eNM+N32dKAXxzmkrja3TTOS
pxOFyBtsWVCsZ3vQbqxwm5LfS/jEqjlUJqwoCASDlfrGHHiZwJrGZGFi/04hxBHr
Z4EQDbKMOOtNUrqX99QVbYrsBtAiCYWtKt3eeJVijA7J30Y6sAo8ZMyADLxFyob+
du7BTjk/ld57Py57MbHfdk2vf/2SBUO8xoUD4V13gOWZ+YcyPjk+zKU5QXWYNfIH
m0FeCkfsQ6NstC/vAf1j846e3NQxoRiUrvUYj0lcgswAsFTC/iekIekojP2sFyGk
ZkLfwkyxuunW3Rng3NwB9lk6OAky1uem+iEfWr7R/XqSozIX/Ehmn39FyLniNLBg
EUUWDDLrrcvUL8AJwVAhmV7YAJTVjzEniCdQC9MAkpQzi1jo+OtDcwL2g1ZPuHSa
V1xEeBeRjc+jybnRLnfzlYoHBaMRc5fbiLDS4b2hMLnFgB7QNAqtCl4Gl+zcpyDd
PaKpF3qddU738kQA1kFsRfz+xjDDpmVMTp+iw1RLEW4niRhu9yJhkt7Wv/F38Skm
Ha+N8LIgpdyWob1wJLHk9sfw46RYFZhherN+C2NucZdBhc6ea89awTTV8/A6VIck
lW0Shxp5+B64ZrMKtCp8ARirNQFpo8LIY/wRFqdgsXCm3dMj0jLa9BrB9FGeHIRf
A8L4XQ5Vs2BgsVEgyLJdg7hl9wTFLKbfKlsZZ3bSh6WWC1ir8ANlaqyeTX5Fcl7i
SxhF/GWaP0uFhfmL4yfr7HhkLUOms/RP4eg/zyp+scIS8G0rtoghFQCoR78ZhYh4
02dJrGZfnSV5ttH2B7ULR9UikW1ublBlWBG3Ahc4ctFUR8/4FPZA4VU977Yqiykc
i7rftrY2Pkug3vHE+QyJC/4Hi77sfQvDPCjTSQfUjSTaXVvyZ5QvoSplTTce9XGR
jb7VfTCt1OezUN4vLBWQ7KYnx/KpQwZ7TftYyQYlgWPPsthjdwTxr8e0CoOQst9g
OzsKpW8+UawOy6WiGh2mtiKwgr9sDjQJjQqM2q9KaMBB0qkZbE3nxIY6yEDvtpJv
VGYs+cTNnvVUmDhZe72vam99tJkxUqoVQbZf+3/Lep8FtW2x6ZlFO8iZpe1C3usX
pwdMpm2yZ5QI9cFSiKgp8oOCaHe8/ZUYseD3/dLms6ImyfYLhXdKGf3Ka4o8GeMT
1ru5vi9R2TDVpAGN8JigWbs/xFEWAPc7zr5+ruIKsV5pHKas44anpPnjg00c3rdU
QYNNugPRLR7VASHPK3np2vBzSojq3qLvO/SO4elhrIZ8KVvMDzLCd6vITvKE/41r
GCeyD8Fz/rxWmxxFsgFbV4otoejHbXScpsojbjxb3SqAhvvSOPxcuSbrHWgTV/ly
yA7HcmZyQc8WT/vz8UYDiFq7LkLwoq/aaiRFS1T0BUBdMLDt8JlMQnKtVHOhTabz
0gTgoGIHJ65SDYOD8lwUcDCb5M4P47aE51doPJ3muK2n/L44/0AJ0u/8KVbxmYdw
ZllufQAZfqz08HVOnL34owi3UmJPju8kmmCHT5u/zyT1m8m+r/tuzmrMDCMsFND6
I6AAB79KB/oqDlLUqHj5EIIuy+gPFEuIS0IL8qSFYe4P3CjhTaBoOez3z1Vm+DgD
bjXvncIu/cvg/ADnv8VpXoz50hN/s0xcS6B+TrEKOXwUf8gwZvIv/0q5Qwhwf0Dm
fa4uzCdrupiJ3Swdi012yKVHhXNVgg7Xj/BbHE4Hhyvuf84m6+yQBcrbpRFgR13a
BA30BkKzqMTCv+HF6MEECgjLNF4G/SNZBUtpk/neMHJvBOia64/WnMWCN+8eTr2S
YjYk14MN2WeFqGFn7rMbqhNekRYg4LpLmWL61k+59HsAqvCHixjbRMq3B1eAsFYw
2GxxUM+B4F4ZoYK+U22EJMM6yv2HnwYiJAGscu5ERqcGfGWD8HKJdTFDUH71A0VZ
JzjIu3C4dPKm9CDTQFnxtPHQT/706nN/e08QtQlWoIDIcBUmZxy7NKtr6KT3gbZX
c6ILgrbuX8kMHrEw13d0Fo23pmanzdrlR3xDTsxn2uBNTrXwpgHhCp7L9/UCHwdb
qTYVrXH2S86U40kTDpV2oNbLqoDKUCCqKakAASw8wkyrMG+U3N2LkUGoIXtxJk6R
AbMW6QHNTgaRjBMrWhIBaowTtBne8pDkxCJ3jBQHeBCi6w8YQSzpArfOqCDjOqoO
l3bXumg9KVMSJbNWAHRPOBorS3AQtinvppdK/IoGh9NjDQlzIfRA0Q5bCnsyG9Xh
B9711zI/noiYjLM6xu3DsA6ATP4LkAAzMpp+4S4Yt8FMfJfv/auqxRBd9ROjVRrm
iG1HIC0IyKzUBB3hB7hRdTFyT2TC1fL4xydxySEDKumzF2evR8QcQmM1HvQmo8CT
hLCrw82S0SAFeQg8dSb0hFNjboCq7+p5dmbjqmjOWjbufwo9gmz690EHDSW9fnGp
lSBXrMg7QUe9eMTCAmeta7d5+HP34arsVvmA4h/aDdPfrcjjRhUDMvWOp4UX0dkD
jsLYltJMh7VZgQYruY1dWxL75BzS/EtDdMtaE/x1Nkrd268KqO/eH0ra5g9uz/qu
Kw1FpQ0Mk50J4MQvy1ZTAeQzPtiNy9jjKY1BKfeOxhhM+6FhKcNLf49mmJlHkpJ6
TR2oy7izwF1tjuVutt0NSrLFBGqCwBsSoOKEmRXIljvuTyBQnlhehrR+XDV+Z9XK
Aj5nD1hBEskiqusXHMRNb8o7s7LxYZ5vAVA2Ei0LfFiqDvOv6o4kjZqZV1ESD4Xt
xVP2VQ8VadpI8dnA2kg9dcfckK1FrtTNZcDrxuuJMnsXlub7Dnz3MVZTf1vytJm/
kWuwEWjrW27vBPXR/25T5ACDnVNUBKGYVF/DkSSSOiLbBMdq+aFNM/RWr/YpApcv
BKGE1wIS/rkt58ignjDxexkf2Zvz4dLcFzi3NdYzXWT0rp4GTKAOmjZgtjAWcLG6
O6b5B29PR1Dp6Szd8F3YhxQsl4uzB8ws8c0wqytBl3n/umcYydUQmsXISUq529Pn
Uewv2ZvK3u7ixNyOiXLasV75V0g8ID6IzblZSJ/CV/FoAVMhRgsghEMUgMf70j7r
IYDMukKP7UJK49VhAKNTLdrEc+EE3j/Qnd/xJctXESnU3dac1SQTDkSEZd1b2pJj
E5LEdszCkPRc3lkicHidLvfiElYFC4avRj2uy53wFbaQWNxeW6ef0+HpsN0TE7a0
StSDpDq8sT726j8QhFKJ5z3J8vYC5q/dEg59Fn1b6f7B3LUoJoUhvLZ5PX8tmGlg
gQK1pVn79PEfNJ2k29tHRXEKKWeDigDuEWQ0fOd/4mqOh0AmdXQ5L/DHrs/cy2Dg
qVq8JQHibJC2EM0mD1SIE9s4UuOFXzCRZpLNw69lvxIMiCTA0/cqyoX3ZPg7l9jk
8dVsWojVKh7AA8JzdRgJz6kVghVW/gJo2ZlIcHo4x9mJAEH2IXG4Ni/g4HjHg3ep
Iyt7SrlBLCWfDgED6YbJvJUywUJ25ZKS5Bffu55HxXogcnJaOwVJrzHqmxiFvJlA
ARh05mcF0kzBT9qjUfqvdVmOW5awNEzh/+zO+/mFJkmbiWQ4isUqwTdOa/1vQ/LH
zBOBn27dBoDmMSbfnDe6IfCiEPF10NBzSrlESozpBBjyfoUc91rE7vl5XJlWqDsf
m+353hZBD4YyD918i3RhNP+o8fQL+Xb9lofcmnfRNW5eTeFWVgZ4irIyodeKxRBF
ez3ZnDSZQkjPiRWodXoeaJGDfIhBKANiHGtCr95uyxXmvp5aqZc9aznbuSR7AMf5
7ANK6bAUVKaQdfKJdf/oTLcqJorb/UGegICB0Pcc0f1+T4ztBSBdLtvlzBH7KENI
ozuOCK6y0UnV47y0CmhVTN1qELEvynlBSU6gGlv++JvOUvb8WubT3V8qGKZ7+sSa
Irt8E7LS0+i+SWW8BxmUmP2RDIGomMuiIcEXIN7To1SMl0QBOZ4Ppc+57Pfmgcdn
KcUced7J53NL9YthHO/f9XzI0rddFGpzxudRulJj2VwMeB+bUxI8nGKKC4PM74Oj
k7SkATIxHJGxMxvltBCsMR6aKChGy5KFt5GPNIrni3wfKQTnziAEp+Pe+Z0lYUwI
52W2zWv4FaKi+KjFOX/7iBqhzR1lr6kiTHoeV0NJGa4Ua7dgMelOvzumwES6crKn
KFsSbDP7Kw0Oy9rkY+dib/OEyXR616vAb9EF/MJ8SFi8Z7wEaxR4TCQNA3WhdN3E
ydcRzq/m0itUEKARct3wczPkuNga5rrDZQpaxDMvn7xUc+Jedo9WyzXag6b+CC9q
LwXf2ScfzYqvC12kSPDLZKVtSsTa4I+lWKzHigQE5ctbA/zGc4gBgFjNY9d3l00/
qwmZVsNryIIMCYO7Mdgnc9cvTC3pzoUYPoSZg7RwNGla5gNHm+e4qzNyL9YgTG+u
gIMdP/bOpDGokjjTrCKAR3VFPEM6xJTlA/rdqvMuEq0u2QwoIsPQ10kNXlYfcL2O
X/XjTRO50PPYeUepjQdu5LfKZdBYmeXKi9QiXKUcl4gZvhHLp1Px6fpHnnggb0tV
dVqcOoS5mz4aJAbviTmXQn45DOtzSRZMpIy8hdGCiFewJ6njQibVZkIAU9tWT9Xf
t6R1PU5MC0izNPY/pxlxxU0RUz54lGjS6gXQr49ILFDlUPygkgDKZsICqfQFK3n9
pjagXEmwuCNXb/6hQhKdKCC+K0p0J5cdF5ynCoAsvOk2FMrjV0GiQdk/0NVSufoR
n6OM52unFrRiermEC2vkq5FIZgMGYcxSJ+6sGpAxxU0NfftdJf8v5+e4g93M7zOX
5hjmYdqJlYXoURte1dsJt2HousdmxHR80kOQONH2r60MxN59c0GbUuwI/lcondlJ
O04UgXuXXIrWjfI2whq9Ka7k4UxmKcV4tbpLwvr/WKr9GGYsHd7w4E75wXdvgTSe
AbMwOzCTEmweBH6htOBwkiOmWWMYNug/yF4ePyK1/I5ZQbsBIK9QCEB1a7T9uZzV
nmcZrD+QCMLGSSs92pVTZuk7+EmuV690UeivJF8DD8i2GCtNS2o18iymcZXUn46b
LF92UARtpNchL1FsZiaxFz0zYhzcSyIL/OcqEQKaeaAMfOCyI4P7A6B5HM5KUTCw
M/FVZ8kox1qzNUSB3/aouKllsa67jtgVvr892HN3OZbP8mR+wNWhkqNnILDGw/yU
MgJHcqo9aIp5+ewMg7BnlMaOX/7N3pS93cgmSix3Wub5NSFfqEfJhqXC6xESSrwr
16tuo3QrQRDR+uLgfetWgB7BlXK2MkTeARPagcgxrmCFDOD5Cr02/4/T4h0Mf4Fd
L2F1bZkSWrU1hdyVNPnISh871jiorgleYZH6GJq7fTQZ1G8j4yn+JQ1WLOUgd7ti
VVgwYNZy8n0o9vBDuLpBLoQW0/fJF3OxZg/kOmxIvL/sP23Xlq1pNpksZ2lp9ANg
Q/T2bKqtjagtar7pLFbLSKTjULingDYFzZVPe2tKu+wfFqMBXOfx7jgsTGFsWlfC
YM0Ftg770fd+FX7U1aiAMFP2kQpkpj5jHHCloDjA6MkKyVtfUeotIS9nFGFFU4lD
blrfkXMJUBRNU1OXZFT+BQCTrleOV+89EnWzRuEhEncpZPhPOn+2v0FWXrNLYNzz
FDQLaRepbixeO3VgbYtu9hPGPOKOIsh0JhDPSqrijmoa8oikdrVB/or+7ZHN3s80
AYRC8bCcIQ99uTijyIqTks0/BAsCM61UnLSY6g+38pgJeWWIaAxs0vWu1s15QBSW
jKLBN7QLELUM4BysWUbF+RugHppS2lU5d7E4w6Bo+ep6F2EBeL8ErOM2OUFxSE7U
AwYviNctz28eGTaMRE0/h5oFtRjJDM5RKj+d2Dq+Xuz9Alc1jSyAcUuLby6a8igF
rr7ADe13d7uXSx9Eo4mWW5Kqyr1qwaN66QAigwonjAQjXCdwbTNzkOTyWCrCPifA
YoVID60dAkPdBC6o8tu424EwwhLA/DGWUtFv5akSMhZvHSCA7XajgdNOHeYI/zWZ
xJKxJ0x6ndE1drmkKGUxLGKK62SduvqVfE9/JCS9Q98qeApqkqxiFoBbdpcTpuN8
7U4WLRc45bZd3tdHzkyydH/gyJ54at8Jw5iOxNwKImxQLplMoNfOxXAqp8SD5t58
CMCNgL5NTh4F7zLKKSGa2/eXCwxPYhkbCJ4D79raajV2r9hI/ovd5toJXCE6Rjk+
fbu7C3wIFvUa/e5P2tDgu5a9kwF/pHClbR1n9unmMzEvvFHlyd2Ep0sLI0gzcLCj
AjifCM0ngSMAB/tMSdZeXeUqCE2rOuZ9eHdEM/47Sqi6/ky8CrWtdquVwbJdMc01
S2ysnpvUDEd1XtKEpjappi13DTI6wveZWnzyeh7wbaWtZLHBtKYK8CN02nw7PLIv
1jeL47VhfgjjROz66dWboEpslvajjPYAg3O9R8s88Zca2HTLutgMW5TBwLdO2Xd8
WyEIjCTg9w9FEse7LCZ/AQK3KIGpntPpEU7Vxt1E1QsyrxLaw9jCvZSPOuXMHJQQ
dzxdFTFZFjWjPRw2yDWX+Rc0aotqghDaFnTrWwFB4ikJzI69RyWkLQTRE/NHMuFk
hFyDfTfNsU4HQveffkuQp8cRxTQljIUrD7VTGaM2w6SEGVHQDPZHvlEPEZnlXzlw
jXVI2Agui0nL4jz33XNOYs28xphvyYi4gcJ/S9/uHsjDwj7FCZXXm1SQ4446QCCV
hbFmshAv/s/yNXWPrYF3LdZGhEhSICWO6fmHNZailx7fhMubjzTkY7iuzHXmC0hx
nZ0VkGXUpt2JJkceYEF6PgTcChNwbuknKjzkc4D+5PnAP1eZpZZd6S3G8FPB1giK
sUuF8emGcs5prdaKo35D0D7w2+WjWUy+Cwsj3s2HQxbn8T4gp4bhV2WWe0PjOSqa
ABDxX+OBtWPFpdk651JyvAm0PQTYktzxKfq7PTXvXruJXXkO286teRTISsCOxGxU
sjz3CylADkwas7FTN1prT2SfgNCuu+AuMhCP9Hq312kmoA1r2WnrktiJblVQO7rd
gN4BiCQaeVZ+ehN5+HZ2viGKzobebmYYeDqHdYgfkL+aozrLNiSQb+m+0B+orltX
tcEzcoGU2mmqIGgn2nx4rItHhkx7ePKcDkH3IfMm2y6LfpzNxWbC0paNRGZwpKYp
q5XXnj5ndC9Lmv17s/tXqqBJ1k/uIMgQzVMnhNqwRC+EksRQ60zPcDnX1REJeMEk
kyiMH93zfl06aWiEFu8tdJwsGgnMdz2pgja/g/IMPU+v25/sFjcqmUexAk73Tt7h
8GHoYDRXS+tzQUnhiEqz26grv2K/CG1hgM5pwf++bkEkKMblnNjBxi4bFQI05TGQ
8AATpGnkOKQhIxhA4fu/c5DfM8JOj8JGBV+CFboLmvvI7Jgad+AGSLsGV5p3xjY/
JKd/JCD/X2cewKvXsbc8gNNOI8OIrIxaJwgCq3DTu0orvLqBLaiJV3c68nyswBCM
AmV/YJgoLlGWlTqUHn/hdV4SW6Gp4wqUCLNf7meAN+rutSpHqXNbQcMrlwXIzfGh
VG5L9wJYKK+66Q0W64h/qAZOL0uqA87dkMlpAo2X0X1POcDHz6/kIo7Db/nera/c
uWIOMK80U/UuRtSxRzuGVGrOZyYWTuLLMS2/Fwgf5ZgLxeiLh+JyW/dJMy2LX0ii
eU2YuNPVc/Ji7VGaJEuOvBCA+J497Egztr7gRfV4B1+Ij/vk9YG321DSL2XU0Fob
xEoxKAwUwdd9tt0ynb5c3jGfnyfINY85X4BkL7ckrfKeIumpXUp5PfLpUzjWpdLN
WAThgOHiMO9OxCEDFzTEavx1rIHAWmMSWxElssTV1T51Yqb/ivg/gBoqwqCsPIRH
h7gU9bGVrvMzp3bkCgthIf7K+PpgRi9BWCcfe4sqOf3f79+rwDGzP8cbY0DluhwD
JaEnpQzUSgahlS0MTPg01mlG6vWTLmQwAHW8aTTp5YsyKTt3SsCTlXDSlYowT94W
mpcnu/fL9QKDznpxmmK1O6Stxc4A/tc0CaH/DJ3CNs+jbgDbAgMxrySd2iu2GeQl
Jw4HcHwlin03XaJf/ACd1HhwFZZ2Mv6Drdez9IuIOdF1sNafASDrjhaT46yNfqKJ
d3veTHJDKg8TrYIyI5mQZ0MHeVSEeVnFQjjqlARQrfBZHpy5wi/2x2MPt0f3yV9o
vF4LXtopLgSCpTNgrqwdTMmgMJoyqjV2zh+EwkuVj9xkyeb9KhlZdoWEf2NFMRXs
yye+23/KEv9FS+4z05MY4cqghiaxR8pGn+ugbbiDqkoLbII2pk3SgTqeB2HQj8km
8wQUoS4neIW4kQ10CITITHrsUvgpgZ0j/I4pV1oA2iZmM6yQSbUqwBBCYdb3TwrD
/iDVQjXJFdXZgVQAT8xPPPATN1O+kJH6y2t3om/lcCJT4TXtnuqve83MUQySPg65
hmX6pL5ZEslZFMVNSvaiR6Utx1xnWqF2mI6WV5OZN1yOtf6Y2K1DxWaw9P3AOsvK
CofSWDtxVD5LUDqDmd7vszYiZgn+5+Ub4kphA7JRrE5Y75SZWe3wsAKHp7Yj26O0
SoYpf5kzD/DqciAcaG2XF68UFXw25i9YiLKQu7G0r/6t/A7S+OY82PdquTeV9gOP
6yjn/Ou0QK6xMOaQiAiK+0iMfSHfh9osSiN777bLR4wiwaLApNzicMjfsa23ilPt
X+W9KI3rh49Z7hRW+c4Zex2XN0ZD7vNwVuZ0ew+Q5Uj6PheVs5wnWcx958Yn4V8L
8dkpKVQCMjb/gA6fiKDemnmhG0XBFcPXojesL2dGix2ZlIQ0hIGkKwxMLWNG7bWK
XKKyOgOlZb8niY0Mo8hSN37GgIrvpegTka6RxPjzq0JkCQD39jJ0JbZNpQkN/ds/
XLGaFhvzLZXvaQmjxYd1Qo//nPBwmWjSvHvdv2LdQkumaMhrnpuP63CerEUCzaYb
vVQUjEh0Y/X2I9xaHc7CZEJg4as65smdeKHxHeXrgphl7CXKQAQuZLFgEwsOiDEP
ytzin6IPOSfQaCFXwc223BNu4C4lR1+/CxVgqe9mPPCtxSMGAx6nn7CqSR6ZYLvj
mgF51n/z0zoC/4cpLqvxpjJKCZUCnjOcOoKcUYtTwwDzDlFqTx/HqJel7F3YFTnC
3nusRIcIX0bAMv+R4fqe+oe6WS6BUb8YIP/MuFSST2cWg2MS1RTYuSj3OqFw8yyG
dqW2+VTQb4z8chuwWKOzqA42R4ejEZlzB1CBd2Vup9vppOEUSb6TwTUtixgLsk8n
hjctH5LFKrBWnM71i1o1LNhXBY8Tgyth5/8hDqckDXXG3jW/DxGD54eO6PWy5hx8
RpxSpBFqVygbjsBr44ryZpTwEAWg7s1ClMDYiSpcjoDYiKo8bSMfTn87IBVsOlkh
kYxfyZ1fZgcZf596WdZOKPEfwMbYcdwF5X3SALJig2z8OQTP4uwFGMPnTpw/BCR6
UY9E62/piTJkxA5N3YM/0xMwYZ75J5iyqEOdet9iJo2SlcL9BaRr+dliFgVPca6Z
XYvQtnH2uKeFKLjz5u9ixYUchXXOgKyBLkdvbGsjnQvlGAbg2rxUmzetnbDAJ5HA
byc8oJpsyWhqQjfcI2XtsOqNUgFDXeCMjsn8OTuAdDRr7WJSsH/6stWOwiUKM0ry
MmXf9IrVI3zfewEwX6pU1nBMRBm0U2lOujywd9bI5/f0u5d++UmPv7fv3LJuehWD
LXuP0GtAVQ4z4Ye2hMXE+YQ8DB8wvIXAjSb0nAB9XCD5ZXZvQMrNM16cyCOtDzOg
tU5WnWq3wTmEOgjDxcZu59IgKBnQqtgJiqTIlHwpI44E81si4u0DwxLKg5btOxll
ESAEj6WILA4BAW1p6V4XFoZztoa39O9OeaCZ/FNaYiI/rJmbpz4g6wcdSfnB2c/E
XbhzcrcIQwVSF5FEd50la0+Kl2Jth6fDTSzYdwpBRZdXdjw2Z7MGCEmGbxSxit9L
JBNqUJqI1o8Oy9UuEBDkv9RvULHi4Vd0m1RGp4/SfU5Zp4TwH2g9C768FI8QcVb0
Ees6knoGOOPGWnzEbr8Mm9DwyopgG4wO/XVwqV2CA4r0wf35xMjcGttlRJs6gtQE
KDEiE/E36h8tjnCoKziHyiXNWXZKB7Y9Bghn/wQYqwo3xJqowm1wSZEufz1TWogs
XeZdlthcwQ6nCi3D3GWzT+eiTe5RqLMzvgrrpRVYnpcs7uQBWh9eH5BL4nupGIJb
oPxfbHSkeveq635cjGCl2VIWh0OgfcXEoXlFngFB81bco/TLbupqq0BbXWpqEnYv
YXjhDaDH7eDq2ItlbJXlvIqs+MxWd59r0yytMmgCyiqCRXoj758EKr3H3dLHGnfw
I1L61wksY0WHl6zoEf4bMLj2B+fM5TUZlhOvPBuA6UDowBIy0QxEUWQc2crEzBQx
lIOCqrLL5gvB18XfHf72Jiw4sHjytU552UVsL4UA9zwaKIA4xSEUh8HHsrhJyuf7
AvkJqDaCeeUXckmRf+fRdlu/um02DqG2YeV3k3L1A/HLyhqpUS3XfP48XiBLjMmG
V1iqPYZFM7eW5jLwVQOW35GxzlfppS26t2wptAWZPY+0jd2i4LRpdCapbceIM7ij
sQR+B15HipBxQ9jUyBusqKkoi8C2xuJf+mCr9JeMgB1KXIjq+NZJG1UVH2PxI+Ur
ltUsUZ5itIxuvpuYvDySZhDhlgq9izOr5HyU/qFGtulkPXKKaDxEEeIc5KZ/5JmX
vI3+yGMDfVF32dLrLFk3S6f0ZVRXfZaTyQL9lZroRTirUGqrpa36aCibONA7Ex6j
tct2JQZDg/T9iMExuv1TO0rjlpC83nIn48fAHZtyzKw4Cp6MLyXCpGOWsg/bH+fo
7BH/Mc+NWc/nAEx1eZAtncq3Xto6zNKVwBeXjbb42Au5VqRd6iGk04SX11k3gGhB
U2hxmwINAI0JTYj3H+RCvsf91Kq2kSHN9XBqpRRX1KrlQrbv3STDo8veoaVUnXhh
OZfdChSjc9l20V2V+zynhee2LNowQ+IgT6z+VVZ51JbMLs4GWuERWNeqmk3x+mC9
8ofFoc6wZM8HYvsP0naNVmP3y0oTzb21THU5LtenW4o0nVA1pV7w8//I+I4ThfSJ
igT1k4FE4GGUtXGicsHZkbR0qNAnIEDAZSFlPb/HNKn9/0X8yqENWfTzmtEfmLW8
j6Voq47+hW6T8WtoyYFp0Cc4AM+caR+hjUnCN3KgXVE2LMvOTEQezQmInK/tWlBW
RV8fqTTKkP1ZakyScYdzqauIeXOsx1ocCXHuvVGI6sZRMEUllxcGaSMkTtOFnsNF
twIp/mk5D3be6RMCdnPK8g5VmMRNecFhvdvHBijmNNpCIgq4TZ6ikxo81qay2C3S
d4tc9qSj5HjCkiMNKeRDRQblCXt8mSwcCQZTiYso/4n/xMtMfnNtnSCfS9Ztcpca
/ZAwy7y7TKECeGwcWwVbvRbLjRhVCs/DYYPSqjfsNgSsXKaOmRKFwDR6bZWrWZvi
b3SirmOv1wIAZeVqsZ10Ylf+vBWPn2Vb3xUiVeK1Y7Rgg3wopUVWPO9EpRxn0gru
Ke1e87osK8W05blGXwzR7uNl2vqnFdvtFBI17N6l5D7+2tYkumHlRn+omu7+RueN
DZYYK5q/Q46Qes4VrT7nSD6B/frHSJeQPUHaf2SdZeRTTTscaLylA5GlJ9F0WgCD
N2Kshcmq6Qh5i3ANajGu/h/aw7R0rD+duCTPeh56dH8TpZRT6Y+XUVOgxAIqlAIv
7vPjzUQ5Uz2O1JN7P8Y5r3UOSFA9NYD9z3TbRPAhtQdPVJ3vlGi2//5V0yVaWj2i
NTjV9xVJ+ad9N2ufVzlDVinRJSq797VGcMbzpcjASx5v5hGw86KQcNqAn6nKdoih
Uuy57SptxiVR1F4cKAZZkReEhx1IdKc5MR21Nnnbz57EKkmQ93H2j75T6c47Ebeu
0v3I0j53A8l9odqxqRE1bydsfjTazFJYxxJKkWWnSJIUgaAu6bVk5VxJZSia3wlm
3fe7vjg5oFaYswIfcwVbmWqpgUqdOU+knLrc5aqXZ4s3ab/LRXpIjocqn/sUoY5g
43m9j3R/tWVJD0C5PzI4IYmcchaORrtvvkhAk6EgLUIvDr0okkJmIvyGzHtX3sEv
aU1zGWlOWC/Opr7DVJY0PBKFdtp0p6n8NL2fxmw+VK6R0RPw+cLoRnXUS1+EdZPT
5X+QXujQdjmR9qmILwN1jj4o8g+XgFsppd8292xOEn6/2RGwRJ8h1tRFKdigQ5KH
B+2nZAZ8MiQm+wVw41MFpXrq0Fr67kpiNIVfk1G0Av+r2/BH2r4KKrzV4VdDYyY7
zq1urzTuh1Qu8yMvnHML99H3Pu+DHqfK3rDun140dBo9yUo4s+jjf8DzhTFH5czr
8Ln2DgNVyUiEjs7D4letWT5rgMYrV90oAk7rXpkq31NWubb2zdV3FqQGsMhRy+ct
7v4rqXtXzpRW6Armts5O6AV8FLyoSRbST59tqb+qSAja0dqtIbcNRSu1Y+SOOLAZ
CjuqgJEBlq8alpwmK3zkcZMDa2Nfhg7Poxa2vjmuz3EDmw4tLpilwn7luw9T+UCJ
xUDbYSS/h4AcelOyfmKhSz6m+PMnW1qhKLo1ZXpirDFdwlu8qo4YaZYyJ9qAGbOs
dlz/nGLU4/Foe2/+hECGfhV0OWE0bkHfcAfZhdTBrB2AQ+KJOCFXhfrUv+MCXUcl
rVJjrUiY3lWjMdNPO1Ixpn5xnOmEDdcuFRrMxIAS539jpI2p8U8lh719zfziLmf6
sn/HihAECUZOUp4x8wD9or5sH/LMNdtvXvAvryuNg+ntBm665GC2XgMDgnSkrLtX
nCnpYgqx2IDDX0Br6AsMwDtqA3vqz8bBSzC4v+i7cWxbh1TmEjqgJ/vfUFPNBdBV
bBQgp0ImiUS3/AzoFy9h6LYRAAGEYYk5aU3pxuiHWJgpgbvBb0CoPiBvqAGp+Lc2
S+hJfK77Mk0bnuIaFNuo6jPnqteBs5P5JJGMD5qYJCEP7ap8fQ7/9ocxAexi4flj
b/xHHvGkzBZtALtDRuF4IX66/lwe3OHAhj1KVud+WC8eY5BktsjHhv93IewjCpn/
9yQF0lZiBcqVPQXVKZnSTkXYbNjJ55PWB4xJQ1+DjgT0+KEYtrrJyiO5o2G8VyKF
Is+2jYHMs1OdAHpBNNJ9XbXGNPF6cbAJOGOClxsVwjsRDlcVk8G0IE2YT2tyiMzV
hflWTfzMz5sT2wB0g18lyt/iwfypDYRhlGpDAAzKGlXOIDF0UAJX0Jj9wO+RiYH6
RxW0PZsTM/5PX52taVSKtLxveewqIWcAJaYEI9OPXBJhfA00IE38Oolm6BeUBNR6
l/NP30R4xG34OyfypsRuhhHbeaakmYBHvi2T9xO9OSBrKqWeT9g3PjCt2bwf/YZa
WNo/sT6LBaCWNrcxYzjxa9QQOIZvVgv+9KpryOe8WIRuEte6W0+WV6wFIcEC4YZP
L8AkEr/EuM8A0dXbtY2Qtbj65hM6eYVJbpS77miAUA5rWoV8cueEdd7gAMJQOfCf
Lt7d2swZQOLp2poIW5Ghbo71iRqAQBozfKaVhr5FTvAFfU/DVuh3IA0TU5Ii8qOU
JohSSyjaKgv+0IUBwvHwn9RKOmbq4f7fNGb5VYsebfXGel5P2PJBxo3Tw2cGyUCH
94d83XUx7GMpKxJ65Q9s1tOX0KTCmpB92EpyzSI5LuOCAueBx7AfG6lcBZq3OwoT
sb7nVZwdu+/dxOwxxIPNi7Z5ohG0ONxvwF1S4+jxC96Zhm5Dsgnphzn2XCciY0BF
4MQJCCW9XJ3c2Yv6cIPgvK0B3vcdU1nfXEQFmyCr7+tvddI/LKxPfATmJA54kX8K
UJJJUTvLjmq85NGxscRPSWsaRVymcng2heJ2JmlUeoIE9ChUe4/vplxPMO2WFbLi
rMnYj0I8QkRDea7zBXkvfjv2QjS0QqPojNxvWTkNxUwlYaBh0lmmRlSzUm7WahJs
XCO8L9L6Pwi0rUy60Yn+vtFI0jVm/ggaOd/TATS5a0z4/kXBYekDU8Aih1Y2/2F2
xr6AbdO6uC9FTQqVUIXvCP3d2nRNDShaWzNIHCyBRqm742XYU+q5wPfyB2DXvObe
H6jH66bATkjuiFPto3bVGnwv7jehBCiav3B6MNys4qALQJ2VF5/LW+zffrBdCR7m
9hoMNVSswVW1Sx0RaY1+NXHCPh3+ta9GxtuzpFVHBHFCJ7OyoGzxR7/vQIZNwZGZ
uGqBeq/nfCbbYTV5RmLDFcovCZW/ohjJW8whcdmgkZdckGFjP8EKpuBylDwYuXG7
YcQd9ZuUKK5st+YQlmGzeAQ77D7dBzo03dtQQvLx/PfiXFcckiWCs/TrWijdgtiy
z6k2EZMy0EErq0nfZBiryyShQcNdePfy6nx9+DEnEZXnzpouEpTHChpXPRKiM+D/
fUop4zjj4locbulOvFJPzAc6jlvGM8yFJZzqf5SCjr1JFVjB599vcUy7oszvJ+Lj
lUi5x0YzP0koey8s+0tCOPp87MY/WUjGk4jzNicBki5YSpqHhxfPz8lxzB1LOWA3
R//MXC368U8ikeUyAsHQmQlxkxMq5s+e2fiQ6JYALCQptOeYkubtkjzBWrW/wY0+
odgX4sF0oisvLo6sCU8B+qyQSpAuQqQC/ShTEpd3c+lAOeYmVwsie8L/eLethh3Q
ZPWZspSDwqJ5Y9AaM+d5n1sSNeBS+k3ZJ9XpZAtjPrXZcrmEm1FVolj6LvuvlyXS
tRawiXdSUS8jBxvUco2DFO9glXyBf3sTFdpZOTxmCAfTzFHHkV/KN+6a8zn2htyw
2JjW+czRIcaLqB9ILtcFSI143SADucuNj8HiZAoPJMd0LJy7oKVRSUXbvQCvo8qJ
Ya+MD0WOjmdx31JjPYM5/uacwGnQCAMAUi9r4TPOCKTji1XFwuK5T1tELeOb5/oy
VbiQncczcNefLYDCZaQ/1GvhnirzdD4vVBZGgL14X/XXQ395ZlcZPXKJmxebR9F/
dAZEktvbm3CpSL4f6qTWzGfqpoe6jPRfjsk9k+eDQb9KsyOIEvcx8sp+4Lf4x3bb
agCzGF9JeDeKZes13IE23kshD5Vkmbs87n7VCpdqK56Ods1Y6IWR4tUY7B3FwbMU
CwP89OpucM6oXIZaCHf6+yQybi4A2Poa4jPzhPVuWZyJ8wdBzNm+JzapEr9XHD73
cx3XJgmruqD2PLPUSaBj1WfmNASY7SVmc5OSjOsvgJnYRuLBlNYnaZfUMqL/xep3
rHV73C/LWHe6nfhuGtWd8d/WWTK2Jf4EUO1ufTbQNFi/M3CFzU6N7UQO+f91pfDU
0SRiESdz/ry87lSc7bZI5owkaVkzsqrdDTbAsBz/UMJ4YP0gYZe+NTB3lDSJXRhL
KsflPkgVPVwFWYWINEP4Z4z27WqSIsXi2oadTFlpSj7PP5nik04pJsVV12KoHpRL
N1a8Pp4gu9Z0ZDKM78i80qUl6Z/plgP0wt7r2Ay6E8x7tG5eHrmoUcuHNwGK4vFQ
JCXrHTLnzP+8IrvtKTBia4EfPV/LfcmPRS5KbnJLZR8yeHiMvAt3IgG2v7bs8/+Z
6q2qhge/iWh8v/ANdCtkTFqMIrrV5tarhid/YrXY7MRFvHtJHtU6lcPvqrGWnw83
DP5A/Tdo335FL8S+5DadthqmBgl/bJBiHXymiL5JUTOvp172j6nIIKXZIc9QgahT
hO+ryX4WmW+s+1oStkovTgNQD/Ui/LHjKtR9CZXozRT09LP8WAV1NzoQ6jCGwXUC
wt7I5Vt56TW8qLV/RJS3Su3A7CO/5Pt6K1gAoxR6vmn6zPPaE3ZPDcMJPZZ8mia7
3TWrXxVve8cK59CxVLvI63xagGt0nOMLCm8jGTC8zrP4LFA6IG17p7Qq59C5E3p6
/6Yz+TirzQAUwUC9ez+DhWLCiPT8VbDHGh/MagsZEUEQA6odLnwuoEjywAkA9V9V
reZJK1skjueTM+K39ZZQg6YRZes2A4m1h5e5MHBpVD30N4LXYVtcja+sqUr8vft8
AqIbJZkyOpFxhGn2Ugy/PvTacI8TkP6r7o12Bkwv/KnyUVCQqxdCZWb9csK6EAew
NxzsjbK+DheCZ76HyZaBqX9xfhufSlrra22suTv6zdTPgB8R9dKn66Z8OQqiT2be
cfPu29vtle6al4eQbLbHR1nRkOL2RwDkPMkoDL0UaSb+X5ImHq/uGbveWhqV6Le+
pI4qbz/nW1LxbrZ5Gf/YFYJg9sjjHbSv3YXD3ahm+/RLaYXjCPk0cp+amTM+8MYS
2McMhR1MJ/EJF9F2BuwHbOlxuTmC3y4cXTgep7wLSbBf4kzmM/D3mCNX36WNOekQ
hyVARi+NXrRg00hz+is+RCNEsWahlyS5qnuQZv+PLNDwPHhQaZnvZN8Fa+CH6Kv6
bu26vXycUL+P2hvdvTUX4gWpZaDHH6FkuNXvBcEzhyj50hxSNZIY6cuw9TF8XnFV
zq7Awwt+08SbRQ9xo7oNCD6dr4po4G4Tuz4BopVONAxeQu9rornxG1vqRJNWG6g/
MFzGpy/nUmgc8/VYoW4pzvAk7eGePOFLS0xy+WhSah/CDFweAHJ7ThEmrkYKFVcy
DxoA61wDzS+WrAcsQxYQomhIQsFKHwvSxfEE5I8mWnzKdGbgAdImAMz2MY9byBCY
2RVxKI8X5w4mQdsuigqbzBglTxjOQHgfSbqBnC5AbKCHWXsV1za9fKEX4hg01OkA
xkj3vAMtNs3uIO+GFijlp/88/Kl17OHY6OUdmXMLHOtG4y1F1hrWjPMj0okMkGnJ
PgAmm+pWqBWAxv8ymEuThkXNvxL+HeJF0HOCqAo0W2TExXnM86Z0bXpIvHirG1Cf
b2aGx2ZcXVGNCgna2bBVGV54Ret+h7cwIDSNTsS17zENSnthfSg5bVWnkCU/oOjH
nCsZbYXBFp5Jr2YZh0YIyeC5BKscHilI6pzzhF13BUk=
`protect END_PROTECTED
