`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZyaYEIeWUliIhUozk4vEo1sPEvgPXo3KcwvhBvPDZ/3e495IvHlkkkfv8fP/Brrq
AexrP4+sr+xt9TFc94AFN/w1PS0Yxd/cWz+zQ+An2Mb83Wg1hISafBjqBWzqUUjY
Cy8qJHSzoGnzbp1cWvODbFCxNXKBZGyDwwckneJTiUaJ1QgyzJXOoeZGjSQl+eoL
kZ49A2LotCuEWpQ5So8MMWo2PRpqmpRgDFnXgur8RwFM+Up2WCENfagRSitaCY3d
vZXLU8JJc/jtSDsnE7Jv4WRPSR48v5gMhgp6X8+Y3h56NK6ENF791bCzzF3zA1JJ
JlA21i/OvtPlbRR7DHLLTE7WGgC2BDQzy+riRL+tHYzpAqvwcRijESaQyT1ZpFjK
bLO/xmb9Q/mUXO1cgXRMtR6Pn6LUHEd73+rzHoy/ALP78DhSRvF+B0VbMzJg6BWo
kXtr3AsZqO0uF+nBtlI6CrrlDHcOcfePoJr7Wa9TMJo5ElS3ohshqUyTKb2Onu/q
f5MBS9WkVCviSvTH5lM57ozj6OhsfQuLpkXRhxVvf8NtLuI2TN8Hosp5mOh7cVXp
59RY4onqZLoCKGeZyHFuesUw9o2hvb8b+/CC2Ubk1KwEToNjlWcsKhvEYbQIkZsO
wMFEa7K1vIhxQlzbxoZJJaBHbeiQkg7Z5u9c5rJr+rGyx6+COML0Fxbb3tnhNqAe
8Q79zLWS2qsbY1IwQYIGxgnoLsecK2SAmEsA37pSN3PsVDanpvLkIdMpjz4znQzv
uEEY4p4RsRXuSnTO+0C4JuMfGEvKP7+4xL6nPkVfCUObrLNfyqVRSeNyy6oXbp8D
Bp4OXLMu9bqbqb3LUnWPlagsffxxSFWBWiVA27446IyhEqPYvLzS9gtjlfC4fjgq
DUV/qNEcmCtMQWfiIOpoqjKM5iyHq0faLp2uu+JYoeXH3OMr4sRkEM+O2dkiSmTR
bruKH1QZA5p5KEswgQ35AAxCxgIV6nt0YfwD4gJIfphpLbuzRsjuL7J+U0aMFRmh
kLqR/hHjYXTnP2Q5e6EWmnUGkLeEGmpTzs2I8xgw4speqgrNKRpddveNweSgwNDV
fxBywLQV4Tezyz5wVsrbZ8hvN6rhb0UYqMxmQEZKSzCTIPyRAHOGZuM6IS8EMco5
ewglAuD5gNW1eJJUnUJHhyHyAIq3HkVwFnCj7rS0lLA98wbXxkrhX7Cz2kUJbSTh
BhRxwAt7CbaDbAKINpfIPOZkTYaLHKdUKWnBMvIVEG/zazxgJz+ScI4cnN+5/Sdl
gsGyn0lTmj5aTNvjadCoCfD7IuahDEi3tilbqsjjaM3KCfNrhhYdBU76w3t9Bcoz
eR5N9RrXqqMGoP4hTXBmahXuZDHmhyui8QTqR1NQzUrzdkfBiPjTE60qikIWWjQg
zkHKnS10kkEdV8gw/jytJ3TR629OXGriJlUTLdi6ck+/p9ap2V2nONKc4JVLVZTN
HLiL0cq1pF8ckiO/Ve+vKhGWL87NQiqX6GZd6CzgtCfb2mllYj9SGwwbSdZdTt3D
qhapTcufTWhNOdc33EPSQedmzO8aUQ9MIVJSVEx5rhuvwwX/4Uv8RniXCRzggUCT
ALQm285lHoVFzl83ZOm6aIzuqBNqbjfahE2+p/+ki5zcyYoWaXlc+RNCP+HdwX2C
6vS0rx7xec3MtYI9FLq8hxJxEsh10/oQILATTN8yF9e9G8qP5GO++ykU7cgFsERA
AOujqIyTr4ZW+oKMvAYdV2DNe7Ul/x++HOSue7B8bdm04mL1J86FWZlgCQQqcNDF
x5cG2m7Cp8A6Dt4HAqj4LVrwE/xsU1cSDus2QYUUd2f+EIT10VZ51qD1lChm7R6h
n6kbZ+mdU03J1h9a9R+SOUFbJSLEk1cokvxpv1noY2tWw0pPDbLq/MzGr0SPQj9F
a3uqBitIDcPY71/HRkS5umHeyJEgyU0sxkLkA2qwNS9cGCKqUcaYyqa8l33Rw36l
CEUz0f5/bJxby96Tm5zPos810J6rp2df2pSRugv9YbivLIf/TosmxzgcPu57x7WV
p88I7CjFe5H/mp7gac0sAOFin6RozijeQ37y07cR/UpVxlYFLGRpUyl4kj7rNVAi
AmQ/jcUHP+AgUIOX42ZdvQ6qxQ05+XsunIm5QNnX3IgpsRH8MN3W+bQJHa6jvMQB
TtrB/7/QoOsRVm8ptaqOZzumvlrILOCTMxdXowOEk4o7vx2iMUgP8GYPAjvtPZyy
XhM/88LMUvfnbKEQTa8QkZzWLLND151DKhblYLeqJmRevP9FLWj7cQEGcQXqEEZL
Fl0SQYtfoeRfxLh0L2Mvkh1aCwxcoOVJIqkVjLND8TSh09zggj3dpm1MCaCkZEC4
RruMl8/UcS9WtDbm5QMXvgfnqi8CXQaNudNLpDMjSPLOPrwIr2sfUOgVjoFIPKAE
ALpRTSQ+Ez+c+qz34mft0vOC+Rp+HxBoOapJ7LpLSp/+jutZpICw+n9ia4JvBW51
C8LjDVuEFyDVTvWZ4ljpVB+M8RvSfUL2bf1EyXndl1MzMNYF8vSy47b16Q88aVmc
V8ZH9N9qHAAWYhK3BADLR7Brp4j4xV4c7GvARVSEwriD2DajWD6csTvwm1GTWbv7
JhV1keOeK/Etm+DcW3wxdUvQWQ8oB9Sr9+ucYwz/7sGwRccygHtLA/fn4eTOsLYy
vZa6NOSOhXymvJXO2bXXeMCupPqH5mNsgMwSoh2pbd30Hc1cpstGOJc66XRb7RH5
Mqmx0MwyaiifjWBBjrfAVIa0QNBcXcSL7it0lpZDw31v071OEmW7UZ4XpJSJf/KB
WtP91bUDRaBTNzbS6wUfDY/U6RwGMRkDcM/Qe8iLaVktWl2DpK0IzWzsmBlQJHjB
SqsVjOX2tcTuPpd5i+F02pvnRkqSXVzIx883vzjtvaiZcuOpfDXPowp5S/x69RPy
BkEz4qrbV8SRwralXrUTKNWXBgMq5nQfoLprz5j4e3D1ZNRYEDNZPYOrX04A1F8O
W6LSVVKuX8XMYZ5ih3ZjD8ECEnJ8eYmLTgJVr4m6LEqLI879fGErngZujoV/gt5v
Dgir9USxRx6z/yjyT8bAqWNgspsluQs4FAAelKQpDP/azQ6mcEC7qWIpuX0tAUEI
WRQvF+ei70cic78xsPOjl8ZWoU+oz2gdAQiqK45+kwU4a+2PwjjpId2U5myj+Uj1
hMvrJ1dS2541s/ppybdDBtvkG/uInz7kS3blbLeZ4Wns2ku/mOZ1Plc3gtbxmkdk
lM6u1drWk5O4ECf4rs3LilTn+DiiNyvsoJlmJkQhkXAuTg2e4KRIuGbJ7PpSDA/3
rgZu0mbZVgsarAg4/fhxBklkaRt9oUzbhtzSr7V8QGtgy4H2QYp/NK0FqhJYABBb
4rbR8h0xvk0Vm4tuXbLxEimuN8sQRNOz28u03U2s1cd0MY+dzoRFhJm9yOLCieUs
V0PcPLJX73eiHhMGP10OjNzZf1qqnKK0j9MZC28wbdjGunA8XVNuvZ9l6Q8RfMgf
WUEG+Ewo+USvN30E10qKfhn8EWN3mGQiaKCIEuKIJpZE6W1qxiZqDiUPwVf8ub5O
FBEQuGBKIxlRfqhk5TouTeUXD4Zy9cvN38ug44ydQ7c3VdAQTy2UlhQ93cLVoGbz
XiwjDR/QnGnDlE3CUK7kD8lyIiMotVCTZmpi9FOgVFqMkwbqc8cpUrqcYrhCjIxX
rk4j9NwxsW/PbParAJgzH3ZJUrlz2QdI5qoQ0Gdc4TVlHanlrps0hCoJQbDKA1tx
zH5UcOj/aJsGlhA/5ymGqrXk+RAgif4a/acDnlM/gBrkrjCpgAfNycmJ0GghAdes
Vf80IbZhJRK4TVk7vkhFpntGlTrtvSlo5g2qYKbwEUdXdYatnaT9kaKaC8uRZBp2
88slVXmZSvMQEUUbaLiySMWz7GeZxSSt5730JHGZG+++wE9aZ/IjY2z3LEecezTb
SPEwtBsUqUkkhRVHNifsIt4u0yJET8YrOKKmlOawh6VCQX2QlPxCoYDNqo81n7uU
CG4989qeILBdT0h7pU9y5WdxuePhmzxWWOFQVQYZjGjTYC/wQhTT/zQYQJ1QEdNB
9cCbDPDzwocwbqeQXNROt4a1gpuSVqReSH6Pp6b0R/tnkcAw05fDmJ0GIy964niH
A+nBXgCZiGVdBUlZ8XYwvPkhYAcZJocQ8XZeYdmmyEs0lXGWKTdvehU9zphdjH+T
3OSw59ByEKrlCZQ6UhHyRfbY6w32QlGblDJsTD2t/lDtwqgrnRnUObuBuXHV/XC4
IFbYE6OV3ZhoCdbNdqyW2zvTNel5LKB60jjEqClUXbB0GMyf3mQqWGqXPxePUSDQ
IPkmddv1Ar27jjEhmmsObHmZip5G6izFJBbUFWkfuv1uwm8vOdMlLS77H56OzLO6
GvKFbVAKGTIhhNHx73KgYfpTjgTvorYMn5uuCMBlA4bPHuxp/V58lxV1XZPBA0MK
/CYo+q5xlkKPpf/b45fuolvjJ/UdcG+3lICzGb0+XIhQpnBwrSVbvD8b/eCkPZkK
lMkly08vLiA27MYDUofRioXRNovtBCn/I0/Vej7Abhr7W/TFA2JgcYLloGaFaL6/
mV5LH+tGSYAx6oVZn5N5sxsrWqsqJhi91w/jw6iYmbIjaabwtnNO5NN5H8TnvoXX
RvqmH2Lt6mX5V1hudibsOxfxYAGbjaBQILcxxX5JNYotVp88ib01hGn3DMSOV6/S
BTb8nhne1OJIlZDFe9hFpUiDUA3Nu/ttqemb4Wnx9ze/nZeijxegaHmV+11KEVv1
Ls5pR+s+r1ClumkzK/GMykH5aqaI5qc3nm8qHw4Pf0pKUaU/E/cXd/kHMwLuKBkf
m0PGTr02mXoGb6PFf16ZqhkHY2xUen1EkJZLlOvKll2kFKugYZX+6WP8ZA9v9nFm
1p6YlXeDCOc3qCMxfuUEuHVW8C+Xz8P54V4yY4I9YUTfr8qwMQ0JQEYW7fCyjiPg
yzX6OmnPurov4ivro+Mm2TEPRYTKS2subBOswIhjFwHEPrARGYbZEozPErzfJGVA
nsC2z53ZI5s8lnFyd4l+FrKplJbpm+FjLJrEYT9gQT+kAASeWKz9YXbyev3M4OSx
dzBmU8gNud93pe5WVdoUgoH05TIUY0K62uqgZ2be7WuDOF0LH7PRUbjzTKGu+WgR
CMGOxu1HSrDJGX9rNvLYo4zFW1q0sPNTvAUTolg/wRGFUT8O7vPlBJfS6RYd0aXj
nGIkZji0J/rMpvSRG7PjKnAT90ojl9uRJv9ymNdIF3On0jDmXFuXWDUqUcgJo5qF
C3MEvskLqsczPdEknX37aGkRWIbXlnhZADtPr6+r7WmVXXvIzBYuFnjfbi89ZuZP
o/KDj1Y7rkumXBfNqAlff1e1XW+aa6+qvcJvBfh65i6UfkBOIeIoNSftQsE7d113
ZrTdyu1MIsQ7I2WPucCLMmOr/nqawu1noSQKxitrY+5620Ayr81samwrDcxATDFP
Ruc86rEf3P2B3SXDnj/S168+T6Vq3VzKIyTHJMsleUyYLVMRee7L3CuMO4wObCPf
/0jWV3aqJd1+UyjLV8XQ89sLnW/odnIkbRbsQVxnfMXQDS5cyc1xXHPBI9kSMest
6ZFebMiQv/ZYmAF9c9jbR5AaNRa3YUcsTILU3TlXeKQYaKssXrD04fLkpSZwAIEE
8Af1C+N+JO/r1fu8rxDGRTQTGs/TojECFtPxECaW1dOX5n645honY3fXOLY9VT4H
sdmPKcW7b5v94TLSVhppSbE8DV4YhBrBPdUzoM+Wtio2tcMDjpaWmvwse9XQQOWn
n/zl3np2krTBaPY4wUmAq8YSjTZ1Wg5TGonMDZFgaL3Iq9GtYqV5DoXmRbfKOJEO
2B8/e/0y7IGYoTho+hM1dyq7P9RKg/9hUImtMX+XKPRh+Vl4wTIzVaoTf4uxoalf
np3hf7ZDM+7l5GW3wZk+G+plA8RTY0KkkrHSRJrZs+eRg2TdPNGfTOU71cAfktGa
s4QqQC58/SeIhNGnCu4e1n5kuurJLbtK+AMK0iyda5PoVT2JZPpnfxcxJw3fZR+D
Bag1EvD61YAdLEPZwIKLdmUTXjz9SxjNISfoAZL/5r89vcD1UmjYscCqoJ5/JT2D
8kzoCuc5g1Hunqg6R5wxiHN02H3VIsdh7eOGsqyiKcoapMSzi3XLBKDH40fbntIC
OjJJ9QyfXomTIXn3XBHxKZcVLT8fJ0OaXq/Iz0H/Uu6XUDsy09iTgj9/LCvk36Mc
sYPQgNmkCx4FHYJzNIqRMATiRJq4Iiqy69YZn8cSSMNznuZ1P34aRMVTzqMU0Eg6
w0f/T0I/THYtQdKdDzDgmriUV02ik1ZZT7rAmTC2XUjklxLdOivx9aXxCoIUIfiS
2E9Hpr5DdBm1H1MPqgG0YP03qlbXQ0glgEbub6pmfy0Myf8aFnWWiOQ0SRA9sq6K
oCNbtRwV3p92WeuIQywSxXzEofG5imGQKFgTB9Yh6fx1/Qduw+eDGf1oW/LsdMgm
Emm5hsZLq3FQNP7Y0hxcRyJdPhubgxQAYO7Hz3IFi+61HQyPv/AUp9mzmeUuDre1
WTyapPouXHCGQSp+RUtB74kFwFpV4T84O5q9RktKZMR9+IceVZZIeznn5ah+4KHP
TTtKol6tq/mzrt48VynXfT4lIxwkZAZaDZdsrcgf4zT8bT1Tov+We+1pf+zl5nyt
fdfPyPLjv3ha+Dg0KTF3G2YE35DjHqg9JDpt5REoC+lrK3IzKWf3a5bNRVBBsRzw
BLUPIQqyBrG0lwnMVKRk4obqOKsLr5uTJABOQogJzWaX8IHHUMZ0FIViR2EKzcRR
5AeBqRFttfjuA7vOsz9doREiyfaBr4mGdieKjGBWpeaaYcsWaKx+/XktiIWfk+ej
d4KGbC3Yrj40oirOW/zyVHU0K3d2PettF+tAYWeVLasb4Mwth9ec8ehMv0RkLUe/
3t1i0W89yO186lnbR5XT0tVnxpY8XGMjQEuEGCY4a6CMyoUtaJnaf69H2H4ABZRy
EHou9V76bNwOMBgx6JX8ntovVW1Z9pzQv6GYXWX6YuMf5KcQFXZSVA8Q5VAaLqlb
5IxCPeoxrhQCgLtR6/Hk73GxySb1xtfie60PUEtPGjeYiuUefRbyDT4zMMK8SuK8
lnrCxsMa2nE5NRVgZmcsBPEGpsPVBEJKK/yXRXPgiSmPJvT/C+9TAWpXFBWLFp9Q
02PAz8BCKaF2T0Nzz/zLlikq0BQZwenFIpmBcUY88wqsAQHDy4ddi56wNakFmIEg
pNiTuUsyRA/YUGGPkXz5byGi0sbUmexo300OAsT3fN0L2zL3C87iljDBb+SMdwtr
vwZcCZbUzZQwI+rfXMsH/9N3telRmgs+YnOodQa1Ht5KucEmODc9r54QiTP3yId+
qSxnr9kOgZv7tyfe2jFQOAEhdQ4xXXTTt5ajcrIwtk7xhNsrnk8U5vtuIU4jR/y7
QOaeU2ev3SBdXcfcyOfT5olV/AACqv68jxXHr61fHuvoE8n6U+CijFXhFOSBO5x0
zPEq21E4ByJBLJWt9ydo/7jmq4emaWtWm8sCoC2my7VJsThA0BEWpCz8yroUlxHz
45Te8u3eHJoHvLX4uGwDc1/Eab7ErMh+yNLEWm7ammKtrYGdegz5kOSfb23ZbxIR
RT/cl3mbAMiJP/Ac/PBXxJmvE07kfrNQxfDPz5ZY1xqx6D9Y5tZ8GTYDyNM0OLm9
aw/43otTWZFurkgWfJ36FvALPWKzs8Xk9U9MNvJXMRbA6dbLYPOtfyNUoFLJraj9
ORgharpWaiPt3KHQovD8+lF+KzCuD0sH8N/CXGrW+JwMwC6oD+bMd5hStGioyZ5W
DvbpzH8f1n3fH0H9Oli+5BBFPZWwVyLsmdjPylvpXeExXLt9mWpxJ+ss0ae72CRn
dVuDFBcFq8nb0B/R5Nk1dBztrX8VxtnSy+sBc8WGAIlcadduoCXXHBm56Zxh3D7I
Ta6oKdnc0L4oMl5vy4/7A6NlpVGW7EyoK4DiK8pjGRZ46i6IojCmsVuSsMiHGnei
PZk3p86s5FUjTnV82l4uHW1tvAtcE/qxao6xq6AWUpLRTQ4t8ybeJphHSVPTKxYy
yyq0lmse7mvhf2/SXddgToUhQx6yLzewJ+8FO2Xilf6leFz3r//+2Rrew7ey0m66
MZviO+dfSPhEKMhFWlLCA2M5iEvhfSFlPMW79cdnJDHYQCUsCcfEDotuDwluoOZf
aZS5iIlaS1JWJwgQF9f8wuPiM7XHZpEc3x9NNELnGjw9yK6FyxxdbWDA6rSdigaf
/ZicKQHqaAItVXMv4tFNGnirbsrKaYlhURl22jmsRgRUIq97qYvOjr4apxQNhXcF
KPf/AkIBdRYeYsBZ4WO9HADVjaVnJ5hGWia0WPShsqzYYi/GLAFEFWCmDGnPJyQG
Qho9Ufp37EymQldp6M9yPJGu37bc0HJzePwaxDoxlnrzJZ4h5a9hOge8wC2szERx
BsTf05cfxoZIVK0wRTJCYKEYoEGsx8oGlnLOZ7Uxp8AQDEJ6L54JKtnJ1OHIem3W
byvgZtTGrkWm/+gNIm+GaoEbYe5qkhn3hZaO/E19KxUgz4HBgNesJziA1658H5V6
SOyF4503awVmlaU4ia17GhYt61yCO30lUKh61XEt0IDSqygw/KsRIp0HhnzTcz4I
h6iTmVRJGs/SeYZ0HxN1DWjCXh6E7sQ+umCuByn5DM1qyVy4upbG7Wi3wAlugKi4
ZHMuyOv/Jso3eFYsORxUveflzb9ly9ZcDkZiwOKqY9WeTdH+onyi+x8vTk6mf2R/
BWE6yBgr49Qa0uei78kmDQ==
`protect END_PROTECTED
