`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kNOZWtde55RWt5OKMkLBaw6Qzt77yVHNMa0+IvF222jRNLMWkMt6HecLLQM7deE5
/A/Grw6k+2HDxElbRsG7LxWHX/4OhDCir+BFlriLsd24gWRNpD6UHCpsP9fTpyvW
8qEVp9Hpq7tpPyfIchYd7SkSIBQzThCySizHNRzBcd25W0TgiQ9Si2tFKDP8aE7s
3bjJC0DiMztda07xUKg72diNuXKTVpv0kSGWBH1CBsLNmHHju/GaQhMab+HtGLrX
ui/e9kAo9WMQzdz7WN/B5aQULOo5CKDWwpexZfxbOQv+pewAcbfOmq4d4jzeelMV
t9M4gTReQNHhDg29URXmQLOmQ0m0qHzdMF7UVTD3JdhPct3okSF4yh/1a6IuzhoU
R4HDmvqv9cVZTb7+sfi13SNE96MTpDCgvaFNru8mTAFRZMNgFOSQHP3FsMUY1EV7
zXfxdBj+BznAnbj0w0mLQvcFK2jtEd333iIvpkSzlBn7P/2/jtD8HoQHYo1dwrO7
rFA0PkkmOMJG89LfJObGNb79ADWNfEPWK3Lwea0o80Ty8HDrWbYvt67tLzqh4LP+
6SjBoLEAgB1lh92cbjt+ylqgcl98i5bBcUQaFzWR84mjpPvWeoKnPDEAy3bOW27X
RNxxb1+nYlb/69U7goAZq1IeCuf3pc6lzxtRS/Sl+OO97Wg9S3xavaSBjjh2ru82
sXoNd+XndqtbelxhVJBqQaIVolaYAgBMA+wGehYZX2oPwPqvRrmGSmNHwi3vbVBz
4F3Yql10ph48ZEQp+g2/EABNAKXfoDXpOEHVyGqOfol89944yr8o5CE+PVH6Ka+4
JM2bV/LDi6KHYrnFcz9pphw4JOk9kTOGtFOKMqiKs72HAzy97rns4XJgelNS4B6J
9MtuSd6q+ad9O1NOq/e470PTLB8vfqGsMdNBKzVXjc9hnSa4dCWhtQazcjAHxLqq
gE0BeuYhioQcX0h//zslYBU8tjAeTNLjRzc4GHkHnAyLOJCvWd8mEGOU2tiiKCb1
75EhbdtbM8b5bEcVN+fvoLkbjsPFuLygKafRl1PzJO6pt8SySJcfy+G8Oah8G0VE
0FzswIwQwsPnU8BX8AxByH3EqjB2eoWq5oC3zQ6CZfDhOIDY9KiMJK2R7fuGimpF
RxJL3OGUKadXccsmF3DXgzpk+cyowFtUkmc1RUb4mAA=
`protect END_PROTECTED
