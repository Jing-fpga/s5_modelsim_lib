`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nIz2C5CKhAufVpK4bxIPHlQhACsAd7IUsz51lURN5hnStzmwy6wHSWmDqxdM4RJI
9hOPno5kI4s0tSIUjhrZXeoR/Q3rLQrx/RIoKzNvtMjiEotfqMocogz/R3VofAKl
4KbNZv7aEwVzOmNPJo6Sq9O8NrwYdPhQNdejKZkMSTxGQ75pKredGNUR4itRMt+d
KIyOY7TrHIWUoYArpv2DLRWee3pvyDO71UEpwy6sJdfWjvB9YBK7oaALGBxBGaD3
PWWC4b98eb9I5NbHf0DzswUMeUp4T7H+mStBiiNCtlg+5TUuOJbwyf2BvT4v1QCn
BJdbRrE5RYqdCr0Hx9X4uKraEbRd1PAF9d0149Fs1ZlvypDbbsA8/Qx7C7vNSbED
mBlJev7dHObfFqxN467SxcVGTjtSRHtgRDXdoF7cGD1RFBSpLg/J36J5JFO6XnzB
pF3BfkEhvdpaK0xY55opDbyawFK3wgL5vtAM+iChgbsrcxKxgta2MqEIJS88anGy
trNeXL9VXzYEOrgJhrY1EGIsbPXbhnBmkTXyCvpDgrfIuBSzXUrQgfWsVHFT/VF5
jlf8rl5BbYD2qvoZrIFBqr9MWzjzZQljLRUA8PxWoPo=
`protect END_PROTECTED
