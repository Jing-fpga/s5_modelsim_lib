`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hw/0NJCWQFqCdReT9iIqWL81v2qSEKasWXqhVfmKBEX4Fcl+stqcWHm5cMRycEJA
yq026MlDTfydKwsSwaPN5osDy88pLDHQxQsR0J71p8LxB7XDsdq83n52owVYBPol
sz3i6TTyrFcSh1NoCmPOM7K+jSjiNYdTzaMP5MbZEFJHq9+FbuyucSoTMBn5pDet
tjg1RSkIdnelz3VBV5z2b7IC7dPU2ZI9bQVRPenLTsVQGbOQG2GBa+Ft4EZfVxUz
hzswS+rKTG60mJqJ0KpgXmoI3JJ3nltqjHWGkxwfNb2r2ypXeujxLDtOpGeesuxv
Mvn1C4BzKqD5YGvGblRmJhqvSB76JRE72FnvYOUTsp9o3B8stt6MZ2749OjBI5tf
mumBHCfjN2fbV8nm1QdHVIf/xthb2Rr+OfqMj14kC6/JMORwJeukSi8WK93HxpGX
sHIf+VZO7p7PvrionEukmPHipkxM4pH0bVeBVaiCg1mCctuukWUz/5RZEX41s8Ed
T2T3gU6MT+RysJjOrsg/UVsaim84YTcyJEC4YT635uy8APQ3K6nBUbBoqfneVag2
Bc0RK6n1agjleZ5thcC1AD/tcru0+xOw3leAyoBUJSyz5CmL4Lp8VcHsZT+3Xqd3
9n9NaR+4GNkqnyXjZ1frIoKSGlVhTeYupPGZgJsW4OBYp3Q0iWQ0zcAXFXr46C4V
YR67/2LvHGb8U7mhPxjGB9n9zQ60o4B1LpaOOzjqnWOp45OThaErJVSknDkjdGDX
y+WSi4QF9b6xZcJhOqh1xGQnRq52yiH6gDLQtgL0dPnoSj7vTpPJqns3m/QdrW3C
GPZiUD1F0qKYftcxzDn7e/NGLcpbKqxk6PSOaWaTu6saGSmkoqK8sB2Z5X5jGwmQ
uU2rOyp7gUoFzW6KOEomEwL4vKfhdJlP5HmKw1MT18x8wBFWQmIc5D9t89TIjFmi
ajsblyhOc/bAhqNEj9iooHdAJzWYVHjAPHxUrp88ywBJQ1vMPnawqeumNSr048Tu
gQIpPpAitlLMU/ThBMkSSZfWszdbEnFbA1k5Al9wwdhm3oqng+9ZxjnXCu1Yhm8/
x93RYMj1dOXs8d24+MNoEFqZNcPtgV5upIoXIMFt2XR0AEu3K2TvzIawkXAtGVnj
NlI+50ohg2CJ4/8fC6SEkW6ygtN9C3YEnbF/wnB7MoAGeFu2YEQpktjGVr3lRF76
Vh+X2kypfQE0EyHm8qLE9y9taSiXYhZ39ilbOFelLM1ezQ0375b0xI70/+kVb1Dp
iD5e+0CD8NQDf6gJ37zZEX0qebc4zTCP2dwu6uBt9gbN+bUVO+KqQOn7khpvmdWA
FKLzUrOKj9jtfX/FwTP/LLh5TUjWc1mtqZWuPDPgHSasGu/Ys8uiUKbrYCAZ5as5
CI8cWOku1EfcxNu85yq7as9LiTUctfyUww+KMzSgDxJvnYt9Zj1v34JG40SwL6lU
ybokccOzDT5KzAF2dSBaq4lyFiNJzHMQOrPRCSPW19z3vlEwhip9uaAm4Yds3HA7
jZ/iLNduWWK4Ni+ke0nhM1JqzODHM1xyMgnqUmNlxqUnCcp1UrAngzAvjVJ4we9J
+KRe2I30t7WbUdq0UqshEVwtPXczK+CkU/Edhev0HmSr/zxbARGn18fnxL9amgZW
loEGvnMtI/c4240PV05TQP9RaVzFcdhgehlabEi+NmxhlsQtc6eDD1gtk3NfsxrC
b19NMEBFYxM8f9YDzqkBBqd2IPhvs4UXgWEx4equjEzoGF/9eBdipjj76fwdws2v
F1xJLQGW8vl0qF2jFWX24zOlQ0eV0991zaPsLw/vBNioWv0lj9TN34BHdq8kGLZ9
Ma55zuOz6KCYKRbZAVZaAGikOZcvwCQXLpZbhZPoUQbqGj6099X8YBS+kEdFOWvd
7gg2fy6OjIMnzaKEJLyUmCwuFRghaw4KjU4Hxpf2NaF4RlMQqsBj/CnOf/tUlO3x
g6TwbFo8OvAd62mxTnG5XcKu+xvww7INmBOSVAXCUmuIPMGGn1bfJFaAa8bVH5QT
X99IseBnTXmxeFmuIewNLdobfD4NfPN9rzWam1cWeToI2QRTobyadAYqmThylN08
J24KX9ofWgvwz09xMJOI1/M0W1xXV5pys6FvaNbsM9Rzfw9Xl9EAdO/k4dIoutxu
o9Ezoz0VCIp/dYWoJJ0XY3xJkOrKXMw27ZFuboAyJThnjq3VCv0YfkA44dYOwL08
qYGDm2mn/K6i21SsnSL33my0aOpVvsRtPMKR+4SnLpOXLzukbESTWiGvPt/VjlgV
jNRIBZ6tb5zEL1XvxL9vtm4G0/778x4BYn3/s/6IXKZgXkcMK+efAK9oXvav3yEL
DkixjsT98BfcLhQtj9OPRaBEWunhmK+9wSQ8qzH7jLv3+0XFrllFNYQeidbx12mi
RTWJYClArIMkrGnhqQ6dxVVYsQYx1z+za4Bux8kmtTQ9At1lL6OVCs1T02O3J4Bt
gutftb3E+wYlQBHx3b+Af4tslfHDMWMb6Hfps74a0Hfaf3qr0Rfd14W7awnJgTqz
GpJsYhBp/g9ZvFp/YVUF51reX7wN+hRzImJJlKhMdNPCsdH+uozthBNa2IPrCZSd
ni7f4xxcDBX3FKSeRq1FjD+e1ZjP+mWMOwg8TgGFS8G9lPm8tmDBW2i8yl/32w1o
2Q7T6AbLBnlCWOs7QcovxAX/WwpIGR6puetAXvh+zkyexeVCToUbOYRuGTR4bICw
/2AaO4I+SW/xiuxqnieK2K9NsXUhkuqQG97eL+AgykgfTWhRp2wvfVBI0T1zxema
ZHYsyGrJ5DVRtUwRGwRfkDLS/FLVZ4pcBuE2X5XYEbBH05S5ff9xK5HC9A2RBO1C
UC2S155qD5mPSAcsMkIHTYtbsbKkRhqeGpOV7y/f15GopZlu2s8IIasRYKZuqW+2
6DCf5NehvhenhnCumpKn7lMh0B/tubX+e2ClRv2tTd0UMQ69pSJL+gvMRkZMVmBV
a37lqz85XmHkENC5rPbmPjhjow4M+W9glvHUE69ZQp0KOa8ymoOVTf2pyGlbrrom
+h+uN8bIREhHx3LmEZHa1yOimx5zCo8tfTlO7I0RP6UVF4NjRiN+j29z8cqWS8Gd
RZwYcuXkZtsf9JDaqe9DxOvbpxDXkc4Ang0eQyHVoa6BMgA9Aple/TxpwLVUlGY9
MOPmOJCRujcy9f/G58a0x6cLqPdWBWLphbdnFVWGWKzIUrulkJ9u24GCbdXsKgke
UjqUd7HGe667wvwK55SfBVgtrBeXwe7QKAi0eW4gfZblCsMENFq0hhSW5JSDhDb3
fmvMXBNDgXVcvDAl4GMSQcWZPhZ5Q9koFwiYYWpsxA2pNOJABge62Vw9rVgm4CAa
k7kIUtVGEVUxEdSYLTqpiuKW4JwkbeqtwFTXLNMy039+8lD458zC/K7TlDCbXTRC
2CKFqAlOeB/enDb5u5W5ykNYqJVZvmhL5h2fZPt1rUxG2vs7SULjuY+O0q/hkfRl
XZzrMK8XCQykMqdNCtKR1iTDi8q+mBGOmMhwHvNbi02sTG1prLYsy121b9INGeRN
GSQ8BF7311ee9aOJAfmc0yVV9ynrcb6WsdkX0oAIGl2CTwyAq/dSZNVtehwlOnpk
kw83oF1YWL7lqVOMK0BEspwl/MwBPFEtm5xMrJlKt4isDYn8PIrvRtjyLJhCyIFm
q663TsuInpDcf87AiUdG14tUdxwTSSer3u77N3ClOWk4Yq1Vs1kXfMGcAJkb4ckQ
6x3c/pYujjhK3WLkJgYFDv+3JvBHcxiGF2eyziz9Xn9gM1rh3Dzcm/15rpFfF/R+
uTKOVjF+or1x5cDaJI+pT8L97uKhSdaSyOQY4tIuRZ6ko+2yctUg30Sgc/Mb+aYe
qDNmbtD4t/EwTmxOS0ZtWHQ2izl7/ZpSeEPQt3VkiIRlIUCcjAGhyboX7ZJ38Sb9
fuX0lIAl21MJo0j0DjNrhFhFmt7p8A7Y+roGSrwwI+5IKVq7Dbsflhjx020JCmVO
p9ew45tlrAAV19F5GFQc2BNQbV6/YZ7P+hawIbfZOZWcoe2z1VSwjT32VG0SPx2D
ipod0W24d+CpLia2Kc8rvckRJcJSPeBXbVnPRBOVL9lDaP+q2QjqX7wRaiJH09bt
tNZ6yYcwTXnOmN+s9hgqoUV/NmCwrKVYJys6zebDP0W25CQWPoAL5SvUID5VP3YQ
1/0R9MQ/Dol1xV9Q6qA95JBgz3VK6OqDaXmcEelbdOsxIf8RS3KVPAuyFk9Vvp1d
DCqLY46gpp2lQZPhuJeQAtccOIU4ui3rhA6LNEBAkWKxtFbzhrpXTyJE3oyKBz6p
HFtot19RZ6IDPQg1hWhKCBJ3C+6zFmyG8B3OCizYmTeGg0Bwkc3pjGVObThwla2r
1A+DUuQeHR+YoctE1xW6Zl6J70uIau43NVBgA3TtUEhKfZDf1NsarfKvhpQjLtNv
r2Qjja0JzG6SshB7i6B/TlhWhh6KwNeQT0qgxTG1ITALMJir09QfJdcPcI33CJ3N
GUtHi/gupfER78DfrYMzW9BVWI5pR/bRMh5ORM5puKIBav03GV6psaWMAw5oy1Oy
Q10uhshuY4uNxM8mIpC8mOmIcSPc/zgXTgBSx35LHjOhnpLo4rhrLndkChTQoqwV
1okGofsicciJRc5sbQNryed5WAQnJF+VeP/DINiWA2FPeDQr71RHHA6+mxQk+ZWK
qPIwzeMm+S4I3taFb9DExhGc29eF7YyGrDzNGh1w0E3VTJml/08QyIR7Sh13Uc94
3sIbt02zZvS/cYW+jpSmn59KJObXfXZCRQhADYlw95s4wwsi9AS/TdG8Q18HAAE/
14jIeCaBAAiB6Zxc34Z0Qbl9XQfUU2KWwshQqn1EjQcfr2RzGLqroBOFmtnZzAMV
Kvo7YWvxDXmNiB55zoA2vJuwrL89Ff68j6WaQwxO8jV1XsC1hJT57wsnTBtaFcRs
Jwo7HwWwJE420jGtMkqgFGGMBeTV1BTGuFae2ejGtlZUtT33WRfcPh1BTtrUDRA2
+fOE0zWR+Zl3Ykg2vQx1PKZG6caVbbtDjuHJPa4J4/C4IoEKg/opvElq6ulS+HuH
eVSN+9o46ud9V9BRoZ85uBFwxdnWbgWdEQJMGfydQjryNWo1qqqPhFbCYA0ONyoW
SGRv4cB6Asd/KZl1r6kkANVrYIHvMfyztQ9Onf7gw/t+UI7AO/yoH63Y421cV3Jf
RTOUHOTqHJwitCQ+S7nNYIT15oUBu/fSeypA2p+aR7sC542RTXpHEChK+DYDm2VN
SyLWRZ0jTpDWK0r/n8lvvO7hh6eJebwVRLcLUMa0PFzSfCYQG9fSBjHVGQjTqyNf
mu8IZXmdQcCnajJNRcPWTXTCJUFPg1LY8Wt2wxHm7Kw8/AERrYssASbutHFCjYcg
I81TmPEQAqSUplUXmMVTUCIyXuvn+55350i3xadwavUZALBf4FXpziYCtLOtFvZ9
+7rhrjHfr5sLN5NHOY5ipRh30EYL1Z5OQkf49PV/zCA=
`protect END_PROTECTED
