`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s2E3ATqg0erp4N8qBYUVL/UIyWbvdllvXcE5ZE4r5Reir1+oHwB6XZNW8GefyQIS
4rPbW9ubXFkUt3LBgunjyyZwkv+JLj3NXhuCdDg1bA8fJVGx0fsDodbwUpzKEOnh
dxHdvRdhmgzyRDafRXbHfklqhIbi2laLPGUc+A3o9Bk6hzYOhIYTMyk1XL4n44Om
3HgT3owWdIpFr3/x08seK7p1WbkvlMVfKw/qBsUFZCrqs6wluQWbhVZm53H95Prt
aOjAJjXH830Txq+HJDDMMqXGKUxV6z3GfKRfCreCbICtPZk/dXsY59mqPmbuoLY5
v3+n89r2XDRDwXBWHuFS5S7HrJfusZNj7N5ZIJeQfrN4geoSLFgoMVnYXnNm/SBy
RbYbPCc+q5Fbs3flGsIMWOQdIehEOnrCI2VhyxrF/oii5LdLd36Xy3VSgtbmXrKS
jalHoUJy4jBOutzGl9rk5g6b8n2eCaQJx130OMxE8qjMYaMGRsa+p24LbYc8CyYE
9KD5ZFSXeSjcNntEmwYcwDC5t32POb4z6u9msiUM5HhfhNa+YsWl9z4p9Q1JdNQH
K10dYL4pb7zEWgUWnGgy9jxIw041fo9oC5LVKskGv0/12sbh4lHhA3rLTuIF5W/R
iSnCDUhfm0pRCGL7DAOfylWFONXbh8W0PaPXth9EFyXn/AqgoFQ4WyR6wRGxMv2z
Wld0KPg0UtH+ZJzJHchEuKYjJiTxqPQj7HgdyeHhELFR9V+aIUDqOyjscj2j5wbn
+nUfYq9Zw+2817AGmKyCA/qrZfDvKzLq6vKLjvhWcgi8bkNV9LBkkCTfzBZrcd2p
H/BGN36gdfMWEIKPzsCbvjHNPs24CV+fipVJPLqq/alZ6rA329wg3356DUax8grd
h7/CVJ+aniuXALHPnquBS7/bhTuIJeUSHQbsKQQZk/e2vzasiKFClmYWqJBoOxyu
SvsaP6tGjInTlrft80i5aWv27Zmq5Xhir0DiIaF4DkY0ECK46kujzpMLdDsMzfEa
NKKEEO9nhQXJM0GFhlDoWlq1WA+X0xeHy4+WqisnD081skXQwY5OAzOGump8ABhI
F/FQpobqzml5qzgjh6BelED310yA5LFv3jGwNW64AbQ9meFFhmY+/B1pKTlMntOo
OIKZQCTdvQcuUEMmWhdMBv5DztlWrtTfWCimzEzX1UkEyV9fcUZLApIS+5ygks8A
x2VF/Yzcy4APDfL/Ds5NU9GlqhT8+StziEL+Pu4pYYsUeKbJtQF+D/rIkDSwAaCp
eGND84Hx71xXEzI4pKfBZn+ZyS2dRTdIKlz9Soot/0qyJE1xjYYC8fEGjvexBLhE
YDLJoEtR1RPaCWyaZXcNJQTJKIxJxRZ89YWuwJVx8PsoPLdzF11u98Q3xI5FSq/x
VLFW5J3lM0AKg+dTYQdr+d3BdH1bIlhbW3cidFFD/eneChofwG42pw5RLH+q7W3k
CZpUGj6Vol5fxO/yjyLsGff5Kwd6X/M3/qERm7bRWyA3CiDC0uXy02OB+clHhXKp
hdKI+ciYyblN+BXlE0l2G9us6XThkx8vz96rM4cRMls=
`protect END_PROTECTED
