`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B20dDacmWYu+AarzjKmeilUMiZdmbLxhA5ZyGKFxZTfjDg+iNbuw/MPvthjC0NWr
hIO8oStHrctXaSvwn4j2hc9SHBcIyTFs5Q4urhqlpLoHxoanp6FN6SS2WQLV6vWM
6rNR8ob7jU7jJRF/4d3NxStWIcHyWF+efRPtU6sqUUn2rRJouAXjg6QkBEkzKxKe
Yku+AaOZWDffTvFrnNvcU324DNMpameJjpBS/NE7oS15/uPKUUYPP0s9njdXlbNq
ZpG8opH/NU6cVKKFyBSw9ynvYy6B1FnpXetzHGXPI6ZSle22PRsEp3WyEYPUkBKm
vdntOet9uthb6NOGU0JvU/Ez3+CqVwFStq1xMrBGIG8GGwue2H8oiazn4oL1bWsQ
YOW77S9tVxkR+7GWg7OzmicHkYIeMN4ZtlQ5/P3nVZa7ho6xFN2bh79UCGTCrpn+
pGk3E0FLFOjTFyl1NSEDlaJmeu0R4fsB2/oAdf1Ao002Iks0xswhQoLDqy/GYZoh
/fKc9gYkvvJbhaCwv6nJxZCXILdmVLEBbZywDlJTFnU/jYyLCRJdPid3hckuVuEL
nDHCFEwd4TnXFard7rqu7T8n0WjakbkT88ifwh1Gr54rHqYO1u3hxtgka0JFVcUV
3X/tzMbb8KeGrIzvUd70MhGMkbrfBwRoJeOhxcigMOL2ZukSlSZxbwTxFO7yMHC6
Sz8YdHb4ePadRxn0zZSO9i21U3PBBIg1c/xF9o3tKVRxk/PN0gICuN43S2jn7U2E
l794LcjN84f4GpF2XjeRqA==
`protect END_PROTECTED
