`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+7041mFcWQq/YGaZUtV36TOGX02wccnei3qbKzZlknnzD8BmmaZno/hnsGPpqDui
vJSIz9Hmkec/jgQrUC+xnwhvL6x6KivaSu+EuyfWQ9TlvaplOIuXK4kILMeMlcSj
oiRxPi4EWE1RFyjYy6H+Sk8hIHy503fZ7bx7cfv6EuMRyA3B+s0QeOxXUnAijda6
JBcdyJMNT0RodG48pcususUomPXUvaFlW8WlknZXrd3khupGxmy8w8UNYTHzqrkN
zw2SQebA77L1lOd/BVZmTUMURX6GCraxjc2ypJoyz/0p9aA2ReSOwdJWt4MZkkrV
D+BFMwmJPoD2D+26ldMmzSiTK6xe3UBjDPvsjgbqzGLf0/9iGpIwvixu6qsxUZQH
3jQldGkfDkpP8OrAmwm+vmYLAEd0feeeUyPfJcIQRU4xr8FpGakBqFan2NYaGWX1
rHwQZKtwbQC8lU1z0uFDc8tQU9aKkmjDORMB/6cju0b0nNkPd0ZHvcwnYgfHx1Ab
JFLPx5A6g8GPfXL3IyDyDoQLe6ikm8a+973gzNOaIzmFISK+p1otnAotDI9vHYe8
phFf9VyTvuIDnesoIvXK4MakCCd2dTBaB3oFYJ4PH+PZzsIYO9A70PBJe8m7ML5M
0HYksMXfUyfv2DEQ6BiJvX0mJiBWdkQWF3B+BM1tHopVptJ4tR8XHn/tGilfF+px
qOXVZmY5nEAkvME8TtgxGRa+2xsMJpPGACj2+hBFWLNgaZ1C2TCfay2mavrWupZ4
R/73uKfItxajZkFzH7j1Co4y8SssvDcpRtStIJ6rVlftq/N74OOzLpuzIK2nCY4b
UaB4EvbAeryz8k7TonJtnVBd7XmhVahl1N9P2f4XY6ZYAXpptl3LZWdEfI3IIJx7
Nj594eMAVy+rJyoxGotHAU83X0WWdMQbgTe8OsE9IQdWWSC/db3h6yhXlztJw3Tr
brTNbk4uOOF3roj9XYKPuBD+FsqXqBu4FXYf6bIJeZapGb8WJlysHenx1fmRzF4z
lgJF9z5C4Vj6Ql58Bd46/DiRLYtNPtgZBUglwXcVX8Dm93+1FUI7xuuKChxQ1+v1
wVBSlQPow2HIlD4fxsCjk7KPA5Q/mpXJ8k0cmndVtOuvBW3qAAaLsNxWgmLq44eQ
hxDbgTrdkg+Vt+WEnB2dHOepWHwIYuoZirMgGruZ9s8tHcR2SuGgaZXBKCOPf7xK
PYzPBcHuXqXp+OJHNat9/AEq/1wvmeF9hYGPYBGURn9U7RU+lsJjTqEhzIdLiat3
KIoKhhbFNdTn+FrnFykCqVMARTYLO4i45xz5JAidofVimdf5vKVWN2KE+B4O2mJ5
S7wLCYuhRYKitKtQBLfxAUCXfR6Fe8kmgETnrcm4LmE=
`protect END_PROTECTED
