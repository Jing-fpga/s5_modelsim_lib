`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2b0nPRLzVxsKRreu3iBgW4eKRt+uOlbqmsIL5rk9B1bl0U89UO0w7KRjSfjBiVBB
YdAoWKWsm4qKBnNLn1O+iGgIY1ZpGHiZAPhoP6L4L8qR1px7dJZnukPEulKaAyRw
HMcvYpywFCzav1yCL0D866fyluMU7cHBR0XiVv5QoIq+2VssvHY9Njcww/hEP7Zw
ZjJ7KCroqhxY8NOy2hO+myuLwWU1SqcjEwJmw3JCvEH9Gb+DKOFOuEBzXm0zPi2J
rH+0+JNILQls2LFX8PizAHop3B9Tfw/xJyBE5TznJ+6yVXeF+ST1UFN1C3CQggul
Xpg1Y7An7C0D4CljYR8iS/oHJHvYoXDCjp5HOM4azGuGHFlyd3xKbQXHu74S2CHn
up7PZy73MFlVGsTbJiWyrxpfhw+M0EHyWvDlNDaxzas0iaKnQgwgt7EGnM3/LT+H
7rFDmNqfT4mWRyR8GSu+ChrY0gT3YeYUeubzYqIiQRIwaMGfZ0sko/UC38mm+24P
vuHVTpfZnsvjnpYDYHrjXB1yyBLK3Ij3fBOrzAudiCLkoL1mx+SGlVhdnNuQe/bX
wGBwYdFw0x9A+g9/KFXmt4kF7h8M1fXaD7YwAkFJPAM4WVGWrY3x44jpdGFfeZ9S
PjeUV07KyC3+QJaIuaZv3OtWCJcr/Q8jPonfNzbh/0g7T8HpqrWjrxLLW/kg7/RI
IhyHbacO1rwyHrwLTutdF6Tz+PTMF+fqaB6Rxgvdw+Y/pp0kQIl06Ca0q3/38YWu
sXgkKhYNiOFnGrmukbV3tRSyLhU2INrgYWQc1kgKqR5dzhDN8yRPdNxJaDqQ6Ucm
xi42r4sY4RfGlybhTBhjXonpDPqMunAgqa9fuY2fCVDFlZwn998UV67a7QanLv/s
QCYI20CkE+YGjv+d2BvLghGqB9bDMZdYVAJefFsZSBzQj5/ntXxEtqT6EZE8THiv
QA7wQxKV37Zb+YLdajRiMoCxYOg8VpdsfsvhfN/i8w8nVDapKAcPEyxkpx3gPMJQ
xnTYhkX8ny+fFdWRYp7S8wGQVZsykPdk7zikGAPt0BzFpGpfqT3ZDIjHjzj/fnD3
W53E1Yn6BNT9vrrU9Xo/2NzOsRWsWVtGxHC47tRqGN/wwfbTWE7P44houUpXpXP9
O48EiT33Xl57YT7xit4y2nPxJuwEsKSHT53DqRN7cjWBeoc3ngXjVRf9GV2+iKTv
UdhyHCXf8oL0TGYbAnz/pydy5xhvWeS5uNZ/sFqGROsRczx9nQkLPZzWO8zRX65Y
r+npkM3RtA0LeOo367UZ+cRx4EnsMZXSDwao8OvhoyC2Oav7rNMk93TOUxjtaXW5
TYaCgmG3BBqBzbEoaiMj005zdl2dehL8wxE3R1zkPruNY2194C31FLmYQVigZT3r
C7IAjNwkCi6kOWqpCc0AzLWmidjEMIToH18udGnP8Mbm5Wq0tMRTdn4SSbuNQIxD
D8o0zuux1NITI0TW+qHiMV2ETfD+yX1dcrdLpTJOkyJfPIMU2oQRUL0eliCaVbo5
bOBGczM13zhdlfLx4mpswWgFdV/Zt02GfpI86ODpxlnZQS9JC0qsqu0qJ2yMgOHW
t2dexllyjoD6GmKpYsUGElk+d1KSxpXSFT6Lb8L4tLb2LRvDxZbiuwarzu7HXFkl
kCs6lz+/3Prf6PLepUo481/oKzQ0lnrNshv+bQjblu6eIrkzEgs0Veq+bhLqAegD
fMU2XUUq67TEBB3w81obX88GC4QhqzqVeyOwOmSahbfw+ukXlXQPK+JOLE3dhKuD
6fz8DjA4vXk89vGquyvzw2wZyOfXLqE4ccazI17SHbE9rOlIN8uToiEbGMCg/S7U
V22Ff06gN1J5c9vY4hWMPw41MUAhEcODJE4EzveDNcEyYm2hxpt7KlO5c9YzYf7H
tBe9DeC4JwuYssEsebW1pp49bbD5eflkiXDX4BpHgz+Nk5gYGCjnSKtuBLzjXYF2
73/4pDfK8Jvn4MNjKDVt/jvX0/f3GNnEGdb33CGhql6Q87sXP/5tCz6YB7Arc/9c
MQA9NAS/silOmznEgvwMgFdqdtliLIsZwZGBrJhHnyzYwZ3r9N4LuPKN3kK9NDCM
g8Unu3XbwP0LSEM9jFSHJ29PE5FeeDvJEXW9frazTWlvuXpsgQ5GwUKy2cpZxxfk
4ueyXs+e2YogXbpzLvqC9guqwmRoX/iz1va0K/A25441mNQCzS6qCDu8ZKp6S3M1
3ijtoG96tpoRQWAY40/xZRpLWpShEiUP1K/3psJQnASiHnUbjCqe3F938EPZUxwu
NlL7cXFNcrridzsbUvB9zSnzx/kreQy6EGFJpSlPzcQfaKRJM9x0Pk9KhgTyUIKb
9aK0zaHWx9KHy7VTQm57Syy/Jrqvw0mAEDVVcS8Pqy+dU4vYiT0LhYa3YhHHltpP
z/eY82JSw0/2vGOTqqZm4/w2DtnbJvlNgSj9m6YX9nsdjkRnv5HohntLmMm5YAgD
LIx+fpFLVde0sogT6Aw+fza/RJ5S6pKO2ZsCq1wB4SEhIHKsn/YPI/hU2ketwopd
ZV/Wzl/0m8l/OkxRa0Z12AR6PZOO8uKGZsejD2k5UhWPOjOss3RgAoVwk2KW9vj7
Kt+6IetNGtSn5QB7Avi77EQWdhgGEJuRTwBqcCFLDBRqe/SBrC59plqlUn2MZKU7
GQiEaAM3+rrKZt7P5yQeudGHHweWOUSo2QZwxqnjGYiwAhLd0Xq+k/4jyIezYcKU
mVrO5piAndd+x+vSo2UsDZoQHCdHwfBAL5Zzh+XKSXC2dXng0nF6e6jIJrxzLOWh
/AIWED6h3v993m204Jg3YMSvHiSLRZZJ2OD2OgRqvsA1y6XNqvDLEsZ7+sVzvnBt
yeMCbuJVNwuKZ1RWOpQv0MSMV+atHukR3Dmfhcm1/rnIHeNwa80pMKTB/hKhEXN7
ijnZrb7ABAmIiN8g7WLppHdO9Qr0mgXTpzjhaqwQKQrSCUibpJTktCWLNiw1EwkT
Xh0pKZ6lgoOEaKvhAYyvOf4xN1v5ua5smjeg+s3u9JH7ySUvtLDevKjcQPMvuSnI
ZsCFinmrLlHwZatmYAosy27L53uYJOVUGcyWBQVRUPJ8hoRfX9/APEB8+Dl2JroO
b6wrXi8RffX6fBq+O5+R6iT0iYQBtCHPFf4yJOZmNRh2ehWKNZBrmepuo0VY5Osd
YTvG/T4XMXKCR66/8cRY1xjkiJ9otDe1ecNnhrSVupY=
`protect END_PROTECTED
