library verilog;
use verilog.vl_types.all;
entity stratixv_hssi_pipe_gen1_2 is
    generic(
        rpre_emph_a_val : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rpre_emph_d_val : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rxdetect_bypass : string  := "dis_rxdetect_bypass";
        pipe_byte_de_serializer_en: string  := "dont_care_bds";
        rvod_sel_settings: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        elec_idle_delay_val: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        elecidle_delay  : string  := "elec_idle_delay";
        rvod_sel_c_val  : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        avmm_group_channel_index: integer := 0;
        sup_mode        : string  := "user_mode";
        rvod_sel_a_val  : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        error_replace_pad: string  := "replace_edb";
        ind_error_reporting: string  := "dis_ind_error_reporting";
        phy_status_delay: string  := "phystatus_delay";
        user_base_address: integer := 0;
        rvod_sel_b_val  : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        phystatus_delay_val: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        rvod_sel_d_val  : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        use_default_base_address: string  := "true";
        phystatus_rst_toggle: string  := "dis_phystatus_rst_toggle";
        ctrl_plane_bonding_consumption: string  := "individual";
        txswing         : string  := "dis_txswing";
        rx_pipe_enable  : string  := "dis_pipe_rx";
        prot_mode       : string  := "pipe_g1";
        rpre_emph_c_val : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rvod_sel_e_val  : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rpre_emph_settings: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hip_mode        : string  := "dis_hip";
        tx_pipe_enable  : string  := "dis_pipe_tx";
        rpre_emph_e_val : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rpre_emph_b_val : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        silicon_rev     : string  := "reve"
    );
    port(
        avmmaddress     : in     vl_logic_vector(10 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        blockselect     : out    vl_logic_vector(0 downto 0);
        currentcoeff    : out    vl_logic_vector(17 downto 0);
        pcieswitch      : in     vl_logic_vector(0 downto 0);
        phystatus       : out    vl_logic_vector(0 downto 0);
        piperxclk       : in     vl_logic_vector(0 downto 0);
        pipetxclk       : in     vl_logic_vector(0 downto 0);
        polinvrx        : in     vl_logic_vector(0 downto 0);
        polinvrxint     : out    vl_logic_vector(0 downto 0);
        powerdown       : in     vl_logic_vector(1 downto 0);
        powerstatetransitiondone: in     vl_logic_vector(0 downto 0);
        powerstatetransitiondoneena: in     vl_logic_vector(0 downto 0);
        refclkb         : in     vl_logic_vector(0 downto 0);
        refclkbreset    : in     vl_logic_vector(0 downto 0);
        revloopback     : in     vl_logic_vector(0 downto 0);
        revloopbk       : out    vl_logic_vector(0 downto 0);
        revloopbkpcsgen3: in     vl_logic_vector(0 downto 0);
        rxd             : in     vl_logic_vector(63 downto 0);
        rxdch           : out    vl_logic_vector(63 downto 0);
        rxdetectvalid   : in     vl_logic_vector(0 downto 0);
        rxelecidle      : out    vl_logic_vector(0 downto 0);
        rxelectricalidle: in     vl_logic_vector(0 downto 0);
        rxelectricalidleout: out    vl_logic_vector(0 downto 0);
        rxelectricalidlepcsgen3: in     vl_logic_vector(0 downto 0);
        rxfound         : in     vl_logic_vector(0 downto 0);
        rxpipereset     : in     vl_logic_vector(0 downto 0);
        rxpolarity      : in     vl_logic_vector(0 downto 0);
        rxpolaritypcsgen3: in     vl_logic_vector(0 downto 0);
        rxstatus        : out    vl_logic_vector(2 downto 0);
        rxvalid         : out    vl_logic_vector(0 downto 0);
        sigdetni        : in     vl_logic_vector(0 downto 0);
        speedchange     : in     vl_logic_vector(0 downto 0);
        speedchangechnldown: in     vl_logic_vector(0 downto 0);
        speedchangechnlup: in     vl_logic_vector(0 downto 0);
        speedchangeout  : out    vl_logic_vector(0 downto 0);
        txd             : out    vl_logic_vector(43 downto 0);
        txdch           : in     vl_logic_vector(43 downto 0);
        txdeemph        : in     vl_logic_vector(0 downto 0);
        txdetectrx      : out    vl_logic_vector(0 downto 0);
        txdetectrxloopback: in     vl_logic_vector(0 downto 0);
        txelecidlecomp  : in     vl_logic_vector(0 downto 0);
        txelecidlein    : in     vl_logic_vector(0 downto 0);
        txelecidleout   : out    vl_logic_vector(0 downto 0);
        txmargin        : in     vl_logic_vector(2 downto 0);
        txpipereset     : in     vl_logic_vector(0 downto 0);
        txswingport     : in     vl_logic_vector(0 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of rpre_emph_a_val : constant is 1;
    attribute mti_svvh_generic_type of rpre_emph_d_val : constant is 1;
    attribute mti_svvh_generic_type of rxdetect_bypass : constant is 1;
    attribute mti_svvh_generic_type of pipe_byte_de_serializer_en : constant is 1;
    attribute mti_svvh_generic_type of rvod_sel_settings : constant is 1;
    attribute mti_svvh_generic_type of elec_idle_delay_val : constant is 1;
    attribute mti_svvh_generic_type of elecidle_delay : constant is 1;
    attribute mti_svvh_generic_type of rvod_sel_c_val : constant is 1;
    attribute mti_svvh_generic_type of avmm_group_channel_index : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of rvod_sel_a_val : constant is 1;
    attribute mti_svvh_generic_type of error_replace_pad : constant is 1;
    attribute mti_svvh_generic_type of ind_error_reporting : constant is 1;
    attribute mti_svvh_generic_type of phy_status_delay : constant is 1;
    attribute mti_svvh_generic_type of user_base_address : constant is 1;
    attribute mti_svvh_generic_type of rvod_sel_b_val : constant is 1;
    attribute mti_svvh_generic_type of phystatus_delay_val : constant is 1;
    attribute mti_svvh_generic_type of rvod_sel_d_val : constant is 1;
    attribute mti_svvh_generic_type of use_default_base_address : constant is 1;
    attribute mti_svvh_generic_type of phystatus_rst_toggle : constant is 1;
    attribute mti_svvh_generic_type of ctrl_plane_bonding_consumption : constant is 1;
    attribute mti_svvh_generic_type of txswing : constant is 1;
    attribute mti_svvh_generic_type of rx_pipe_enable : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of rpre_emph_c_val : constant is 1;
    attribute mti_svvh_generic_type of rvod_sel_e_val : constant is 1;
    attribute mti_svvh_generic_type of rpre_emph_settings : constant is 1;
    attribute mti_svvh_generic_type of hip_mode : constant is 1;
    attribute mti_svvh_generic_type of tx_pipe_enable : constant is 1;
    attribute mti_svvh_generic_type of rpre_emph_e_val : constant is 1;
    attribute mti_svvh_generic_type of rpre_emph_b_val : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
end stratixv_hssi_pipe_gen1_2;
