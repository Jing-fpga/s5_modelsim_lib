`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3JgW216HKPX2dQe8YHJpvFg1ppdGL+NMyk1VUhrHToAmUWZnv0AeydYCYZ0KeCDP
4eS6eh/oljNAKwp2XMWtrAP38QFXWWsFMn+82DLyKK5mbOeM2QPzTo9h0Jk30pWt
YhywM8NzVC/yZsbM6nKchE9NGAiQqE6I4F4cHtdelD6u/gHfOShHIoUmewk2o590
EIRpqP32OzThs9tN7miVaCPCK1eUKfG78tU6+Bz2iwljE5W7oLRjh7YHVJwYWBUk
0Aycn1jwkacM2qgiecJPc4Nr7gymJ+tLS9Rd2kwSL2g27s6EIbyXEeeFIca/5zcw
lnvW4qqGV7koWgrV45VUfpFDlpD18c8I7HNDSnxsTEOZKeuPdbymVk6uAksOjPnK
hSpIKDGTpgEz7QscWzPJTHY0+9+geJxq5oavC5UQwhcdEWArws7wIsSOdfuxaqBW
9I3OA4z4u8bypZdUHfwaqlR8MnlxAfagTKTZn0YqkU0=
`protect END_PROTECTED
