`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XILoMpS7+rx0XteL37dWEe5yK59B8wgYCy2V/6mNklD9VkCOGSQ5XcyDBJvSaFaS
KT4AyCctkiEDy1SJFZPA5QrJAbWYtcAccTU/lauMePJh0oT7dFV0SmB1VUrYSbwc
7sWmVyrcZp0gQzWeUtJueVo/nGaPOuKBVa0QKt/QtAO9p/PxLU7whZIglELHA0FR
2Uxo/nZ2S0rhWYr+g1ptIbczTnhII1lq8VhKZAsuDM0gD4Of5a1hygKrOeiUjsKq
XaGuwgRDHAATo8bvdtCs4xtMM04aIik336vm41hhfESncOeasU3y/JqdCBoNwmnL
IOpqlFLE40BXBDHRfWw+5dt/zAxR1XxTzHRdKxuieCmWAEYUU4Aq3U5ds7kIRX3l
CuZxDZBZgaOVhuAEThkxjoa4b6uoGWSw/CaFwhrYarlppSK+BQ7Xm44VJ4nLH3Qu
3bB5304DKHriC3pNiS+e9rSU05i4Bsdx6251mK71inHGUe2tSKzPZVn4Pv+fSaWg
scTp3N2hqmk/LNXPCkEEq/MOCMPPU9xtoHUuXvqir5PNEzu93bxv8kBiBvCKgf0N
WlwLOa+vRpDL0RXH5Ek62RvB27wUuuxXf1ujuGp2AFDyEjbCjb7eaBpFDOvnOmCR
mY4lUYRREiBkmQ+MmpCspo4pivf+bSTMgeu16BZpea8BBOljXxIuG5kQNpey/ZEE
8VdyRafXePby+L7tri0+ECTm8t1MNjSaVlun/NCZLo2H4Mr3Pcyi+pJQKDpgekCc
aOkpZj9HIgLbLWdqlmdnCMUAyZBGW1jFgdvlQ4vvs+6fl81sdm11g8x1ZWj/ugf0
YCbTSPPC5grGWQI6ztgEdyilBCinwxCAcrO/pkqrRXeCiWok1qBWCM6CY0CSQ9+U
ZWKD7z2J2gHJkNfT1OrDdJ2yB8X13wXTF1PCZfIlIGjbyN1Bjukmqs5pVsQSBTao
h8VKywRhS1h1NiI3P7LTuF2BBoTBIy04LIIZpXU+HH3eejfeObrV4e93DMydxoHs
FU9KMX/Qo5EVbHe1nxgPcbCGT1ajOO/6vu+eL3pCiuJCdaIkEZvAdiPswmnqlum6
ffzF3fBLNcuUzA5pl6xL/8FHkXUXclWHXkVlAU6NpuNu9fvraKI0cEpPWnnoJ0me
wuGlgWBwV0znX8cWTWBSKKhhW9o/tvVFeINGzba9SPaUngRJPJDJX4kLe0k7p5V2
/VqajGVOvzVZ9sTFKEbQ0RYr9jPXS/h1Pe/ZM+yjprOhzkP1LbLa3Kxxl+29ZgOK
JP8lmQL75XoXGybq4ahomXFqD6gB9iW6Sba2FKzIueaUwvABCEMuK58JTo4H+Dsd
ytb2ukONJvegwr7YUp+d+K/ne/+sQ8nElOKbp/0kDh9qxuOnXm22+wLfi4Wy5ZLN
KSNTmEtrE+CMeOgfR8154Mccq1N+HuN75ZDMjVfKutvGHM667A6xVItH0xZxLgXs
7prEk2xKo3bCT62JSNa5PPU/8lm8m19ZGpHdmX/ULzgL62Z4vpmBdo9ue0t6Vlx8
3tJxLFdE/Ar1cO9DYHOtkMKpb+lLJf3Jpl3M+JQBMLwSshIIVjqzJPHQJyV+eaYP
lKCy4QKOznE8uVnSDlelV53LqCMTXH39Cpo1QrdkC5c8IAlnjAajT1AICbLdhDm/
pdTZ8DAQSNsuURlzMmLbL4haXLz1R82Q/DvkroqG8OL96CRZ/ugi01UkEkEmg7YI
`protect END_PROTECTED
