`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
26zTV62MdXbWHtEGTjM/6rZkegu7QpExy86Lgzv8u0UaZ+yFkXX3OGFwzmJ+JjPs
SYfkXHKGPsl5OQ+pOrsoRUa1VpntW3qXJrx9O2oQGfYis76ejJFiFtZV+FR03Uf/
Rzp9A78bJPJLjMeKUPgq9XQamAUK6q6Bjr/d7XIcaQsOpo0BiBRlNMM87C3CJayL
+CAb0BueDUBY3w1D8j2C2LjitAE1e6lSveOeLVQ3cx0rBCeiBWUeqCLSENxezT0o
Q6ZMqyi2Zhs5FWsRkKN3JOXOOczqD1FwaTaPLWaNPdgGUox8aib10xmUIU4Fr0Q7
bLv+A87+WLXwVCXo0vo+S53YpRagDV33BylCm6EbT3yJIRsQVf56oKLby20OZkaS
DnKU3my5yq6yzy87HTuJ+NndZk3COeKsupJ/OxPnfe4tRekoLYbJc+efiKFMJ+XB
AhGaQhHWGh+GWh9LEVBJ+uVe/y4koFbs7jyesowfpvvYYHwhVhtkRfxZkoOCRFC1
HBHtx0JKJeSBBg1mwCdcJxBuHtDBkcjqbyYWIS84ZHv+AmbH3alLeAHdKzkpU994
WqMmWrjYKEjAXtjltbc7V6/jaUZZHOI2/AM4YCs9xmIYLs21AzfAsGdenZnAv+2H
nTcJw6XJ5pQIPZ3gflgQyb5gDWHYk/O0Qf+vDeiRAxQTXNBaS2A+CtHQ0NbIFaCZ
sx2h5p+TcToWC2AifDfcKq9v6tSRy5vwzfR/kqYFGYXT2mjWEah/Pi3Qv/qMonxP
y2Kb7/pHfjmpNcICI1psJNeJEd3rmfcapyElIB/s67w/sgp3nJy/pDvDgK3DcWB0
o3rXehgLgjoXV3WPuKs5oOohDfxmm4l7d+7G4P3T3dOItHfSwpsSNDv+b9SUPlgI
GUGfm4ng61rMkRFOdYP2VV3b8wyg5rSw1QdbWLksshT7OarHsBsZIwFWP7bdAk2B
btM7nIDOgEptxmiLK5eX3X3vRv8Zpi/tyyGp9NoAEl6o9TLVOuYHD8Up8O/pmS/4
NhFU+q4nNsv0DWvuXbRgplnoeD+9Pv6TjHvMqOOTzn3Usnfm+ZyS3zpzQbv/XfcN
rXaULoz8bc7Axg540NEFiiSQVK2Z1qD2NFxw+XPcvB2jr4ctJxTtvfaOnyz76ME2
jzGSB0JmlAAo7+FFvweLkYmg0bTN2M062l3XNiIgEL6NuD3EmmhOdkYKF9pHwLGk
qHUB2Ss1XyeqZo8AeGz2EMJWktxL/QLMV29UIm+mKYPEumg8VX9b/t+9fIDU+h+4
1q7ZK3ZjgNotsxKcHB3OgrL1kNX/qJM35vnyM8viphfLwDyyHCZYzA/Kw6Sy+F2k
9y0HUoWyFZKZJWsSBX6FCaPhilLxabDagdS4KR9hElgB33e0UqHC9nzyzsGUaq82
vNYDIz0ILdn7kXi8Vu8iBSPqBvKAxpdCKGjFysW1J+Xbbv3vzhi1TyJLI4sFHtZa
8BVzwHbg6H3hE9Xf6M8gkI6G3AmmleP0lRktxA2EuMnyOqfLYUH/0+R9psD9wQ+8
fv7R7asY+IescCdFQv68e4+7aPTlqStdQ8r+xA3fpmDMBvRjXOU9VOlCYYUfqD8d
8qmZeFWbsiv/SvsnHIyKonsAeoD8fseONTKNXxcvBPUkzuYFQJFNegrT6uSXRB2y
YpS4qLTd33jZUY9a6Q8JOSyoH7yMPbpzhaE9zKDfudC5Tho0/3Hlml03ikFceuVI
g8Vocta4qw7BD1XUTt3LPaf7rLN4CjClZfgpDjglahGDcF9kMh6cfRJuzn/diG1+
fkIUUbDM+Z7MpaPOS/PbdhJg2VD9jT7vRxW9gLVPhtwFW5dVJx/XnXTRoEDSHpzl
TXZtlWAkICWr4fY1wH6XiwaLyKJW3SM42aRhLbOU0dY9bZy67zyTY2AydpRa3oXq
HpoAMSsMwX6lxYGyCorBO5O+lY0Ri1ejUl0P6VytVVtvC4h5jq7QJtxMAHzOclcp
0yl/8jhkyPQ/vzfRBioxi25nPVY3qSj4/we+XPfBg0oFv/2TtLdwk6PoMwvAQ24l
h6bqlhUQmV/STPvfuyHMZYtUEVExhp3jDCJ1guixtP6XkJKE8EI3MEjsR9NmXQUU
n4LHPT3GesS392H0g/qnxHOS5cqiRfIpPbIQWllmuHbKSvowyOlaQO1nD76D23LK
23UiMGYILEFzDvzmrpOwUi6iD73hVMx1Ya5ygeQqhA1a8NzUOvfp+9OV44dcBkfr
WJi4N2q8oRJf39nwH5H+Zch8UZ+aMlSxQSaAC6FXVzPsWfWc2+HRSfljeHd4jJSJ
BVKah3vSBgpCumPEq9M/GSWk2tE6U0OwY0mXpO73+HDMjPp6MlDzg2EC0fd8KkRY
UcaIeZZIh9/xouawh59HiGSAiUiPAApabhwUQuswZO/JpRE3MMI9X/B6Tdwwbjdi
wAPPTVLrRyf8ZE2T9kfyQqngA06q5ytcuyh6kUm12DcnhiD3E74h2sgL6uPeGZoz
dZ7vgWPp9zXmOlyECpJeAvnqlBOXc1iRM8bC+IDsgei5tUCN9grYmDXqwHfZ2erj
iKVJpBMXKZCvqY/4Ym+9kL1D1I2LMKP8PZgbc7JvAZn4up9z7UMfPRIwy/Cf9O2S
tBZfi0Tli1FLQiZV6Vi1QqcWpM0UIQnzhwH+jFYAKE6tgC3cSqK5dYXxX5ZetYCl
xGXcpygUbLkfKR/PO14suxW4L8hKP8rFC1XcmYbOb05DqWO9CjVnkNeaVzx8MXD1
cOLaaORRB2In8R8B6PLbjkGvvNg/l191kowN7Z249w2vBOFa122ijNPeMpE5/vTA
718gfShYGQ9lmAiUJlQAgpdWTyY752gnngnSSNCW8Geo1QhcPzepV7nXsra+v6D6
n9ozb9LUcXgZrcI5POM3LzKMJBk3BPpa0f4AIavTFQropYaP6nbHJ/ClPXqaZBrM
2T8G+5Mdocq3ad+JuhXZTSqqtA0NrCt5d8hlesVjgmWmz3aX6UkhN3Lk8qKfGwSZ
F0OB5QDQnD11Fq5NAnhjgjpBEsUOZZxXsSH3CbLFYqei2zwdaYfC80ywuWf8UCiC
lf+yw59wM3CCC4L8lHtXhWz/Em70ogwENOl2BHqBFnRfP9xbZSMu8CXmlo3qT0De
Q/AKb7eOu0J8A7Bp0IsUVXgVFaAwoe2umvb/U/joaQaex4JkBEKbwgM52dUDqhpX
S9GR/G0fbLGK8BR4B3KZktUbimuESshSEiCtu4JeF3skbSMTzZF6V+B1E6vh5ZXe
9HKNxT6UHO5V0SK2A2+RPVbyme8JgTCWHtHk7H6t3oHFOMRLh9oOmKvAbKihNSWV
AcMlFCMXjmYiZfK1Er3GxtX0x+Txu17Ki05IR/PFMLxciaQhvoZdPKPRRANys4m/
fz26L5QdbhXTs8VL8C6jnxN/jcK+g7tzbNLJUwUjDVfL+Or83ld7yu2H1csOAQZK
b5GhdjH4wIqSpRLpBpnrAxaCWQ1yRIKWdbFNcFlcyogVZAQjvLUIPOO0OC+xvYW7
ZB/dwaz+XLGPOqNG8Wqe91ojJTR+dM1DdAiXBqGWfQqRfpsnNnbx/BEBoDOUE1oT
l8/XmTreHnDI6BV7XfxN8NFzKUFvFMrYFzAkBSo7YTgH2OQrLxhhtzJOBrufAR3D
xb69S9ItOI7pkdoPo/G0b/DSFMA+xV2JONbnxPXpaBkePzySm4dbyqZsNrm1OTaP
iLhx3fN8n1y3lYxCEIIDSayF1PJPNVyYWCct6pqu6L6LaJj1hbWKhMv+sfiITVWT
FkKWak8B0cE3VsCvCe9e9o8wf4b/0q1HnPzlVZRZ51n1mjPJUICkxxMwgogDGyza
sUgv3Qho/1kSbQvMplBquV7ylM8iC2WGGU8lsu78gL8c/I45Cl4UAwmaGZw6GQuq
GJ7spSfBqnWYI2TgDu7xTdf98pbceimpyM7OMYPEKOhQ+3SPaAzfBEobRIliPxix
gbegW+Nh/iA/FVF9kKuDD4hQCNCfRqGtvE6ztquN7SK5g4+aQOwmRLmnL+x1mfM3
4+i27VAhyWrTnY3jhkv+WqWrEEL2b19hEZV7LpCVrLQK5lP1s5EtMNrxk3sdxfEM
ZOklBBhIXWFpYJD2vPwwvi9aGQeuYJqEXuK6la5PnDojzAHus4E88Jss2cPV8HPC
sLhrF9nwLgKwGHaY25vxHawh3eOCmz8YkKh/ABM+DhHYIqc0rz8TeNHNun4b1f8I
tS7ZVOY/Bi6/xH2XxkUUMyL/5wfoT+9SH8Hzhl35lKPvVVITLIwapW+lE7YPhbMp
9GtZyy85Vw54/X40m1i3sweCCzxcYDNGpDiFgHz+gwb5hFtOUICkT3b6YlBwQS4M
98b8OxBnoHQDxqhQzsxKi9MoeN2h7bk3R4HGOGwIgOJj8sTtUdmLA7puvswjWY8G
30m4n9/hWd6rWORmAkewe/smrslRZ7D6Ivh+EXOSv0lxUM9+g6RBqha7lU/EY0sa
CSWXVhlxfZUFvrUResP+Me3VG/uc8SSYhOWJ7CkEpUgRR0we3gFWJ/6Qx9lGiuYz
cqiMR8O8bH7PpKZYS6P2WCtl3/OQr538ZrUmtdu8G4E0gg409tFrv/o9ExKCD8AO
AS1dLUC3FkvMA9aGJ0DjP9YZo4QpPslqFZIu/GDyMrSdUwusnRPOwguZjVV3LOwl
EcMATzVs3z7IgsevchR0rj/N+KxvQwlWnXdPDZ6JmYsLmgoVIJsJiHWyweO2i55/
Q3u+Ed3X+WPzfgPh9E2GVq9QpaOPlGIxW5pLy8GQhFvib8NFt5YDsSgKa+QVZEQx
/v2tvORje//qMvQYgsmY/ln9AsI8VdNL4aHEzTvlw2p8crM1pN8cY18CqPwXRPNr
GpVnWKPLp5LBWUwqT9hTpQDlp0cD8OEQtpEB2OL4AJ+C3UzFokP/1q8Az113eG6Q
79iIDGBU9EMV6NrasdMMst78cucEqfbpKau8ScTRLJROHO/36KfzbLkra4El1Gf4
mi0SRMDlbPTW+L7pVjeAOSzpoMcdE5ZcPJPxkkxmOz2W28agTH3SVTWYN+N6SylV
HmNeFagwkBrpiTl0wNTj3UOerVneBn9OcbMUZhlOZsB1BVVtdu8Y8SMRIEjannqX
TW+3iwzpZZbbpHyCYhKZ+QP568XrFQNrD7VF3q1WA8228x0E0OyvcQXhuwTo4gQg
QjWphlQqANSinq6A6FYpds6XSt1dlw38zUUt1JwWZqRfM1+b1hpL/RQLv7IVlpvr
vWt0kkmeYMAgTj9P0WZTqkqvhF9HBl1YROdUrrPcG+WSUvH22gJM3051GNaZ2AaR
afr+djhLSgSANuKmUxiTHm6oh9yqzp6JKzWCNf+9dlu/yZd1E8BDjmwWPNaxb5fY
zHHh8e6ODkIfXlF6sdIfySJtbgpK7q31geKKea9IX08OtJ8VlebiKuPVjuJ7m4Vp
YC5hGwccPTCwaVpehl1UHjNcPk7+MCR7N4lZHiMEtO31pMyiOeITkqyXDSqgUQCl
IpOQN+aeSUH9EEG85P+V/JMQoGxRmoBnDvmTjcC3+u3WoQiGn+rWQa79FpJpbGNQ
go321h+M9vm4Xp0FxX/Zk8c7/08TP6k9A1OumviqNnIW8TEb8H0FiPX4cNKGrzpW
WGi8cflo4ypA+V9Zc05CMIDh+B71XEAei+LMTn1LhLuo4fqegj9EnTF6eIyKrYE/
ayJoHVNsi4Pd9j/6bl7fMx2UWSlw//RMnCWpygLlDJ8h5Z/Eu3GVLhspSBMv1sh+
RgyV/HCXoODYpTzi0tcPps0aO31bjiSGGQ9d1Ee1OE79Mm19gcq003wbYwwuH2ci
4H4ktnDzxaKMXTJi7oaHRP3pkCrm1vUT0drmlvSU4B03NKfzWLw+IjSVSAjdsLF5
RFj85abWIuujmyg1U8X2M3MJcHuMZilyjU+pvN+wKhLzKPGGik+YWSnJY31vAvk3
/Ld+lzt9tXj04LeTNUhLqqzgjgI6KGNjQsUBXXwyBUqhJ4zIPxvI+sKkk2m5jnEA
nqyQftUaWLYg8Ki+SD9FjOLXNqTNfuH2TTvToPRhzl4osau/F1L5WT9xXKYFkpM4
hyAUu+YkpYhS+g1+v1bvLPOoezsRyXHgqeBUfrZxjR/o1HHg9Yw9gkGJqpOEvNc6
XYTsFq3m+izRKuheUgx0j5M4XX4+nFtbqYXN0/+B4beyN5qmT0EUwGFyeZ5WEq3p
5diOVtZmsMC2ZMqZ/h/Mk1I6a4XkqTZ4bzAwFWSmgBjg7g3dfpP5FklHwojso99n
ZJ/RjEbzVFNOfSFUUYJQ7u5MXmbwU57vImoEdSdjgv1ZNwQciLDG39Q3dceXwxJ6
ZgMRnjpwA8oXgiNoFvQGGeO0oRn7aOqGmfXsWmtGLvtuMqHT4DuDhVUO3tqLmKfU
+NutG/VZMyFCjsVorxr0puNStAQXGCJneqLvgT/GXGvNKzhfnVQdK3DtE9bU29O4
RJXp4WT/BZLNctO9hGangxD/u9i4AaBnRY+9tcG1Hi593YisGKUUd6n1SwhBcEvg
3OPVgdpUx4/2lNM0cUuLsXxZswG9Cl6NwJUSLjmJvJMGC++U40rlwJcxTdfqgvkI
F8fH9Jsm63smrr1gvrNvLhww1w2nOx93pacds2t7hg7R8TtektEXgimT/GR+WUEs
LsrBJn/0w5yfi53ol2g9FGOeelet/HxPf7xvRJlwk/SozkU5HTkao56tLP1PBDKI
5wA2yxpMK34lNIwqmgCZaB9xX403csjnQDMex4Fs0TXqYordLlzP+ejjsaPFrxqp
Il4kKEWfzp60I3RzDrYxtY2N7/hLWGGpuYEcSGIzD2ACEGlo0YmOw8+FlPGV0pLS
E1PmQRw3uZE7WERClpzgCjyoMNHiaVj76vVIknFKYxrQs/RB3wz8pGNS4WaezZlO
+HRutEk2JEedUnud7EdaXbPSWm0EPTIc4cTjzp+f1LfRjI3Rj4qW3kJ2XAKbSBOz
96kuwR4vTP5N1uupzbx00kDXz/bmojRCxcOPcYVfYre3gv+12GA3uURmr8N7U5+2
Bw7rwMfDeHv7sbR2XlhVV2wd8NeLlV6OVsUkiPSCK/feacTscfWhttViZSZDr8ME
cJRSVm8aidJ5ccKgGAlDq9u0y58w5AtOaCTNeph7e2l+nJm9ErHWaKo/99q1T4+S
os04WrKtNy8CeAvY/ryT/zHQ6Qz2/oHXLo+Ry3tBC6LlLAsdjaAb5G1tjt7tv0C8
/TLzbECawysHrrvexCson8Y3RlNb/ZFBiB6sWLivpTkxA7S3OkUvh+krfq9eUpuw
yL1wzFOZYq2qcREWEzlP4tDD+4fWgZbJuXGKwSBg4gkAfhAWuzPd4wrFKpAZKDDH
29c5Z6kR7VKZUPbL2e5oiaIAOGBhMQ4TrP28ulGm1cn7LAHp9wPBF03bVBU2Db3/
RI8pH7nQBbEL+wD3JuJBoDorXINnJsDslr18L399Qtli9kUiRc/bEz6XOkMUE83w
qJ76vhZpqJa3Y2HgEsBg9XMaIgrI/6cDpmlfD/ngrqqpGnnuFJRQaCJZgyGwkGcd
Fgzzy+UaWRGkP6VtWXs2sG1XqK8G4Hkn08K7D+s9F5eufPd8TuICCrdAKujj6k2/
sv2DgOdxadrFFFr3Ge00Jr/6oa+ff1nPcRIxlCLdOU1Jz63cN8vi2OWzybOhqtjm
4FbXVNw/8PRTjTzQ3/PbBlTvcZGKGFaHbLKLJJ7PbC1djcWAUbcgExVVXXKqkdzT
03BqTbl8Vc+bncZz30oEk5lGu9063B2Q4YR8xk7x8ar3eNnVkLSWsKWUaeIH+TWF
L4s7vSgDcqyLz324Q4v0pbY0EdqlI6z8p6dnGnYqFkO1a8aK/Iir9c6kjWKSpecK
og2tLxW1US/rdVsomrJETMhn7/88XMOy4UXZGzQtvreb+ljzXCHRfTdS4rigjwtN
MhjKUuco1CqaMPwni6bsjGeLeOik0ugy6zbbBUbuPlRUFhs/Z2h9pkguvSAvRuBc
INaGgKog/Fcl5STawAMvXRWhKVfuSZAqz4Ov3y9E330/Oq+fDK5cvXrfm2cwa+Df
gDH4/OaYx5BJSs17/eYNseDFAVgAbOF+rMewKPu+qRtTobO6a6zL4rocEXYR6FJf
mNoxUs5oZfaPPR4DsSgtiGy/wJ6sF5xY87UDqyn6yrzMDyOKHSPqp7u0Si6q2g4W
eO14PFuQbijY7BhyM/j9X2z1myYIQslt1t/HdU8Kvz43876iCtu92yYFuyrqIyHL
i0Pv18uGQAGvC9raKU5o2miZUEhSZeLdUZPFUEqpJ5CW+Z8EFnYX8HU31brvmsuI
jNf/a8m1/SuAydX1ONrYBubTNWQACqE2ATGocOlrTaVHlymgKJtUSv/EHr+/+SZ/
20Ifi96oi1FKGhYYP1qEKybhDXy+N/TyemKIooHA0z3xWI9Ta7GvmADsckv40LWM
AwqZBChXlogy3LNrHnmYWGsvlNxr73CNl45AlVOJcMpS/k+Bpgt+2ZcBBQcG/UFj
bgkJ0YGceXxLYMoKWgLa6dKyOupA9gBc5fWEhQlLyov0NB7v5GWs/0aIfyXtD70Z
4yjSuf7gB/ZoPsb6riLAfnGs3ePJY7Aiq5k6VS3ZAkvvGV1fILsfJYyHoEIBgd4T
`protect END_PROTECTED
