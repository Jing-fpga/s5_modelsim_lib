library verilog;
use verilog.vl_types.all;
entity stratixv_hssi_10g_rx_pcs is
    generic(
        enable_debug_info: string  := "false";
        stretch_en      : string  := "stretch_en";
        rxfifo_empty    : integer := 0;
        rx_sm_pipeln    : string  := "rx_sm_pipeln_dis";
        bit_reverse     : string  := "bit_reverse_dis";
        rx_testbus_sel  : string  := "crc32_chk_testbus1";
        rx_signal_ok_sel: string  := "synchronized_ver";
        force_align     : string  := "force_align_dis";
        rx_scrm_width   : string  := "bit64";
        lpbk_mode       : string  := "lpbk_dis";
        ber_xus_timer_window_user: vl_logic_vector(0 to 20) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        frmgen_scrm_word: string  := "0010100000000000000000000000000000000000000000000000000000000000";
        blksync_bypass  : string  := "blksync_bypass_dis";
        rx_true_b2b     : string  := "b2b";
        wrfifo_clken    : string  := "wrfifo_clk_dis";
        gb_rx_idwidth   : string  := "width_32";
        descrm_clken    : string  := "descrm_clk_dis";
        ber_xus_timer_window: string  := "xus_timer_window_10g";
        frmgen_diag_word: string  := "0000000000000000000000000000000000000000000000000000000000000000";
        rx_sm_hiber     : string  := "rx_sm_hiber_en";
        frmsync_flag_type: string  := "all_framing_words";
        blksync_pipeln  : string  := "blksync_pipeln_dis";
        rx_polarity_inv : string  := "invert_disable";
        prbs_clken      : string  := "prbs_clk_dis";
        ber_clken       : string  := "ber_clk_dis";
        rand_clken      : string  := "rand_clk_dis";
        rxfifo_mode     : string  := "phase_comp";
        rx_dfx_lpbk     : string  := "dfx_lpbk_dis";
        rxfifo_pfull    : integer := 23;
        gb_sel_mode     : string  := "internal";
        bitslip_wait_cnt_user: integer := 1;
        blksync_bitslip_type: string  := "bitslip_comb";
        ber_bit_err_total_cnt: string  := "bit_err_total_cnt_10g";
        align_del       : string  := "align_del_en";
        test_bus_mode   : string  := "tx";
        sup_mode        : string  := "user_mode";
        dispchk_rd_level_user: vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        dis_signal_ok   : string  := "dis_signal_ok_dis";
        frmsync_clken   : string  := "frmsync_clk_dis";
        use_default_base_address: string  := "true";
        frmgen_sync_word: string  := "0111100011110110011110001111011001111000111101100111100011110110";
        iqtxrx_clkout_sel: string  := "iq_rx_clk_out";
        frmsync_pipeln  : string  := "frmsync_pipeln_dis";
        descrm_mode     : string  := "async";
        rxfifo_full     : integer := 31;
        fast_path       : string  := "fast_path_dis";
        dispchk_bypass  : string  := "dispchk_bypass_dis";
        rx_prbs_mask    : string  := "prbsmask128";
        rxfifo_pempty   : integer := 7;
        master_clk_sel  : string  := "master_rx_pma_clk";
        frmsync_enum_sync: string  := "enum_sync_default";
        crcchk_clken    : string  := "crcchk_clk_dis";
        blksync_bitslip_wait_cnt: string  := "bitslip_wait_cnt_min";
        skip_ctrl       : string  := "skip_ctrl_default";
        gbexp_clken     : string  := "gbexp_clk_dis";
        dispchk_rd_level: string  := "dispchk_rd_level_min";
        frmsync_bypass  : string  := "frmsync_bypass_dis";
        blksync_bitslip_wait_type: string  := "bitslip_match";
        rx_sh_location  : string  := "lsb";
        frmsync_knum_sync: string  := "knum_sync_default";
        dec64b66b_clken : string  := "dec64b66b_clk_dis";
        user_base_address: integer := 0;
        descrm_bypass   : string  := "descrm_bypass_en";
        frmgen_skip_word: string  := "0001111000011110000111100001111000011110000111100001111000011110";
        frmsync_mfrm_length: string  := "frmsync_mfrm_length_min";
        blksync_clken   : string  := "blksync_clk_dis";
        crcchk_bypass   : string  := "crcchk_bypass_dis";
        frmsync_mfrm_length_user: integer := 2048;
        rdfifo_clken    : string  := "rdfifo_clk_dis";
        crcchk_inv      : string  := "crcchk_inv_dis";
        blksync_knum_sh_cnt_prelock: string  := "knum_sh_cnt_prelock_10g";
        blksync_knum_sh_cnt_postlock: string  := "knum_sh_cnt_postlock_10g";
        dispchk_clken   : string  := "dispchk_clk_dis";
        dispchk_pipeln  : string  := "dispchk_pipeln_dis";
        crcflag_pipeln  : string  := "crcflag_pipeln_dis";
        avmm_group_channel_index: integer := 0;
        gb_rx_odwidth   : string  := "width_66";
        stretch_num_stages: string  := "zero_stage";
        control_del     : string  := "control_del_all";
        blksync_enum_invalid_sh_cnt: string  := "enum_invalid_sh_cnt_10g";
        dec_64b66b_rxsm_bypass: string  := "dec_64b66b_rxsm_bypass_dis";
        channel_number  : integer := 0;
        crcchk_init_user: string  := "11111111111111111111111111111111";
        rd_clk_sel      : string  := "rd_rx_pma_clk";
        frmsync_enum_scrm: string  := "enum_scrm_default";
        crcchk_pipeln   : string  := "crcchk_pipeln_dis";
        test_mode       : string  := "test_off";
        prot_mode       : string  := "disable_mode";
        crcchk_init     : string  := "crcchk_init_user_setting";
        rx_fifo_write_ctrl: string  := "blklock_stops";
        bitslip_mode    : string  := "bitslip_dis";
        rx_sm_bypass    : string  := "rx_sm_bypass_dis";
        silicon_rev     : string  := "reve";
        stretch_type    : string  := "stretch_auto";
        full_flag_type  : string  := "full_wr_side";
        ctrl_bit_reverse: string  := "ctrl_bit_reverse_dis";
        empty_flag_type : string  := "empty_rd_side";
        fifo_stop_wr    : string  := "n_wr_full";
        blksync_bitslip_wait_cnt_user: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        pfull_flag_type : string  := "pfull_wr_side";
        pempty_flag_type: string  := "pempty_rd_side";
        data_bit_reverse: string  := "data_bit_reverse_dis";
        fifo_stop_rd    : string  := "n_rd_empty"
    );
    port(
        avmmaddress     : in     vl_logic_vector(10 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        blockselect     : out    vl_logic_vector(0 downto 0);
        dfxlpbkcontrolin: in     vl_logic_vector(9 downto 0);
        dfxlpbkdatain   : in     vl_logic_vector(63 downto 0);
        dfxlpbkdatavalidin: in     vl_logic_vector(0 downto 0);
        hardresetn      : in     vl_logic_vector(0 downto 0);
        lpbkdatain      : in     vl_logic_vector(79 downto 0);
        pmaclkdiv33txorrx: in     vl_logic_vector(0 downto 0);
        refclkdig       : in     vl_logic_vector(0 downto 0);
        rxalignclr      : in     vl_logic_vector(0 downto 0);
        rxalignen       : in     vl_logic_vector(0 downto 0);
        rxalignval      : out    vl_logic_vector(0 downto 0);
        rxbitslip       : in     vl_logic_vector(0 downto 0);
        rxblocklock     : out    vl_logic_vector(0 downto 0);
        rxclkiqout      : out    vl_logic_vector(0 downto 0);
        rxclkout        : out    vl_logic_vector(0 downto 0);
        rxclrbercount   : in     vl_logic_vector(0 downto 0);
        rxclrerrorblockcount: in     vl_logic_vector(0 downto 0);
        rxcontrol       : out    vl_logic_vector(9 downto 0);
        rxcrc32error    : out    vl_logic_vector(0 downto 0);
        rxdata          : out    vl_logic_vector(63 downto 0);
        rxdatavalid     : out    vl_logic_vector(0 downto 0);
        rxdiagnosticerror: out    vl_logic_vector(0 downto 0);
        rxdiagnosticstatus: out    vl_logic_vector(1 downto 0);
        rxdisparityclr  : in     vl_logic_vector(0 downto 0);
        rxfifodel       : out    vl_logic_vector(0 downto 0);
        rxfifoempty     : out    vl_logic_vector(0 downto 0);
        rxfifofull      : out    vl_logic_vector(0 downto 0);
        rxfifoinsert    : out    vl_logic_vector(0 downto 0);
        rxfifopartialempty: out    vl_logic_vector(0 downto 0);
        rxfifopartialfull: out    vl_logic_vector(0 downto 0);
        rxframelock     : out    vl_logic_vector(0 downto 0);
        rxhighber       : out    vl_logic_vector(0 downto 0);
        rxmetaframeerror: out    vl_logic_vector(0 downto 0);
        rxpayloadinserted: out    vl_logic_vector(0 downto 0);
        rxpldclk        : in     vl_logic_vector(0 downto 0);
        rxpldrstn       : in     vl_logic_vector(0 downto 0);
        rxpmaclk        : in     vl_logic_vector(0 downto 0);
        rxpmadata       : in     vl_logic_vector(79 downto 0);
        rxpmadatavalid  : in     vl_logic_vector(0 downto 0);
        rxprbsdone      : out    vl_logic_vector(0 downto 0);
        rxprbserr       : out    vl_logic_vector(0 downto 0);
        rxprbserrorclr  : in     vl_logic_vector(0 downto 0);
        rxrden          : in     vl_logic_vector(0 downto 0);
        rxrdnegsts      : out    vl_logic_vector(0 downto 0);
        rxrdpossts      : out    vl_logic_vector(0 downto 0);
        rxrxframe       : out    vl_logic_vector(0 downto 0);
        rxscramblererror: out    vl_logic_vector(0 downto 0);
        rxskipinserted  : out    vl_logic_vector(0 downto 0);
        rxskipworderror : out    vl_logic_vector(0 downto 0);
        rxsyncheadererror: out    vl_logic_vector(0 downto 0);
        rxsyncworderror : out    vl_logic_vector(0 downto 0);
        rxtestdata      : out    vl_logic_vector(19 downto 0);
        syncdatain      : out    vl_logic_vector(0 downto 0);
        txpmaclk        : in     vl_logic_vector(0 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of stretch_en : constant is 1;
    attribute mti_svvh_generic_type of rxfifo_empty : constant is 1;
    attribute mti_svvh_generic_type of rx_sm_pipeln : constant is 1;
    attribute mti_svvh_generic_type of bit_reverse : constant is 1;
    attribute mti_svvh_generic_type of rx_testbus_sel : constant is 1;
    attribute mti_svvh_generic_type of rx_signal_ok_sel : constant is 1;
    attribute mti_svvh_generic_type of force_align : constant is 1;
    attribute mti_svvh_generic_type of rx_scrm_width : constant is 1;
    attribute mti_svvh_generic_type of lpbk_mode : constant is 1;
    attribute mti_svvh_generic_type of ber_xus_timer_window_user : constant is 1;
    attribute mti_svvh_generic_type of frmgen_scrm_word : constant is 1;
    attribute mti_svvh_generic_type of blksync_bypass : constant is 1;
    attribute mti_svvh_generic_type of rx_true_b2b : constant is 1;
    attribute mti_svvh_generic_type of wrfifo_clken : constant is 1;
    attribute mti_svvh_generic_type of gb_rx_idwidth : constant is 1;
    attribute mti_svvh_generic_type of descrm_clken : constant is 1;
    attribute mti_svvh_generic_type of ber_xus_timer_window : constant is 1;
    attribute mti_svvh_generic_type of frmgen_diag_word : constant is 1;
    attribute mti_svvh_generic_type of rx_sm_hiber : constant is 1;
    attribute mti_svvh_generic_type of frmsync_flag_type : constant is 1;
    attribute mti_svvh_generic_type of blksync_pipeln : constant is 1;
    attribute mti_svvh_generic_type of rx_polarity_inv : constant is 1;
    attribute mti_svvh_generic_type of prbs_clken : constant is 1;
    attribute mti_svvh_generic_type of ber_clken : constant is 1;
    attribute mti_svvh_generic_type of rand_clken : constant is 1;
    attribute mti_svvh_generic_type of rxfifo_mode : constant is 1;
    attribute mti_svvh_generic_type of rx_dfx_lpbk : constant is 1;
    attribute mti_svvh_generic_type of rxfifo_pfull : constant is 1;
    attribute mti_svvh_generic_type of gb_sel_mode : constant is 1;
    attribute mti_svvh_generic_type of bitslip_wait_cnt_user : constant is 1;
    attribute mti_svvh_generic_type of blksync_bitslip_type : constant is 1;
    attribute mti_svvh_generic_type of ber_bit_err_total_cnt : constant is 1;
    attribute mti_svvh_generic_type of align_del : constant is 1;
    attribute mti_svvh_generic_type of test_bus_mode : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of dispchk_rd_level_user : constant is 1;
    attribute mti_svvh_generic_type of dis_signal_ok : constant is 1;
    attribute mti_svvh_generic_type of frmsync_clken : constant is 1;
    attribute mti_svvh_generic_type of use_default_base_address : constant is 1;
    attribute mti_svvh_generic_type of frmgen_sync_word : constant is 1;
    attribute mti_svvh_generic_type of iqtxrx_clkout_sel : constant is 1;
    attribute mti_svvh_generic_type of frmsync_pipeln : constant is 1;
    attribute mti_svvh_generic_type of descrm_mode : constant is 1;
    attribute mti_svvh_generic_type of rxfifo_full : constant is 1;
    attribute mti_svvh_generic_type of fast_path : constant is 1;
    attribute mti_svvh_generic_type of dispchk_bypass : constant is 1;
    attribute mti_svvh_generic_type of rx_prbs_mask : constant is 1;
    attribute mti_svvh_generic_type of rxfifo_pempty : constant is 1;
    attribute mti_svvh_generic_type of master_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of frmsync_enum_sync : constant is 1;
    attribute mti_svvh_generic_type of crcchk_clken : constant is 1;
    attribute mti_svvh_generic_type of blksync_bitslip_wait_cnt : constant is 1;
    attribute mti_svvh_generic_type of skip_ctrl : constant is 1;
    attribute mti_svvh_generic_type of gbexp_clken : constant is 1;
    attribute mti_svvh_generic_type of dispchk_rd_level : constant is 1;
    attribute mti_svvh_generic_type of frmsync_bypass : constant is 1;
    attribute mti_svvh_generic_type of blksync_bitslip_wait_type : constant is 1;
    attribute mti_svvh_generic_type of rx_sh_location : constant is 1;
    attribute mti_svvh_generic_type of frmsync_knum_sync : constant is 1;
    attribute mti_svvh_generic_type of dec64b66b_clken : constant is 1;
    attribute mti_svvh_generic_type of user_base_address : constant is 1;
    attribute mti_svvh_generic_type of descrm_bypass : constant is 1;
    attribute mti_svvh_generic_type of frmgen_skip_word : constant is 1;
    attribute mti_svvh_generic_type of frmsync_mfrm_length : constant is 1;
    attribute mti_svvh_generic_type of blksync_clken : constant is 1;
    attribute mti_svvh_generic_type of crcchk_bypass : constant is 1;
    attribute mti_svvh_generic_type of frmsync_mfrm_length_user : constant is 1;
    attribute mti_svvh_generic_type of rdfifo_clken : constant is 1;
    attribute mti_svvh_generic_type of crcchk_inv : constant is 1;
    attribute mti_svvh_generic_type of blksync_knum_sh_cnt_prelock : constant is 1;
    attribute mti_svvh_generic_type of blksync_knum_sh_cnt_postlock : constant is 1;
    attribute mti_svvh_generic_type of dispchk_clken : constant is 1;
    attribute mti_svvh_generic_type of dispchk_pipeln : constant is 1;
    attribute mti_svvh_generic_type of crcflag_pipeln : constant is 1;
    attribute mti_svvh_generic_type of avmm_group_channel_index : constant is 1;
    attribute mti_svvh_generic_type of gb_rx_odwidth : constant is 1;
    attribute mti_svvh_generic_type of stretch_num_stages : constant is 1;
    attribute mti_svvh_generic_type of control_del : constant is 1;
    attribute mti_svvh_generic_type of blksync_enum_invalid_sh_cnt : constant is 1;
    attribute mti_svvh_generic_type of dec_64b66b_rxsm_bypass : constant is 1;
    attribute mti_svvh_generic_type of channel_number : constant is 1;
    attribute mti_svvh_generic_type of crcchk_init_user : constant is 1;
    attribute mti_svvh_generic_type of rd_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of frmsync_enum_scrm : constant is 1;
    attribute mti_svvh_generic_type of crcchk_pipeln : constant is 1;
    attribute mti_svvh_generic_type of test_mode : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of crcchk_init : constant is 1;
    attribute mti_svvh_generic_type of rx_fifo_write_ctrl : constant is 1;
    attribute mti_svvh_generic_type of bitslip_mode : constant is 1;
    attribute mti_svvh_generic_type of rx_sm_bypass : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of stretch_type : constant is 1;
    attribute mti_svvh_generic_type of full_flag_type : constant is 1;
    attribute mti_svvh_generic_type of ctrl_bit_reverse : constant is 1;
    attribute mti_svvh_generic_type of empty_flag_type : constant is 1;
    attribute mti_svvh_generic_type of fifo_stop_wr : constant is 1;
    attribute mti_svvh_generic_type of blksync_bitslip_wait_cnt_user : constant is 1;
    attribute mti_svvh_generic_type of pfull_flag_type : constant is 1;
    attribute mti_svvh_generic_type of pempty_flag_type : constant is 1;
    attribute mti_svvh_generic_type of data_bit_reverse : constant is 1;
    attribute mti_svvh_generic_type of fifo_stop_rd : constant is 1;
end stratixv_hssi_10g_rx_pcs;
