`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EsqEXO8EF59N9qt+8lLQolVBcfd9LmF3Wrlxb+4YJlDjhSMMpX+3culnlq6F8Ymx
p6dnBHus1j39z2KelnFI2EIZDUDraBet4XfJs9NyqDPsVX/QxnYHHSam61P3b7hM
B3Qnqz+HKwa65uJttXcToUGNmAwrybnMozttDd+rjCQmLWoBPy7mrEnY+pyhPGYp
9ytpvZglYqa4iUOXLG+mBxjf+cCspOE6UBh39fCZi1cYOr+5rdF6ken1VwMlCjQn
3IKY8VnhIuI/092CYZ81ZgMkFu0ULYeJ2JmDTDY6zVRJxn32zOaDzIdrzSLiAec6
ETOcDJmWIalyblWk/RpFmJKcEQcCSTaL8POtah4fGAXOc+d9+/7v/lp6e1967kp+
bnOSp6U4Eaj6VuAKED7U5QrvPa9TprsT8BerUrhSe7dqATAjMygtmuY0+ggghf5n
sVQyYFk+ejBbWjvQFWyNg7QtADjeX7Z2aWTH/gMFxdGErSL3TF/iWyCeMEnHVQ1r
VLC6DRmaWGSWk7//IFxkBhH3v1cJzptFmy2jPNs0JkdeCvtwtH0yYoYiJPlwijRi
0ibHXOqPPNHUKevSme5Kreo5AQofSzvLcAG3XMIbSD0io+Xl8WUVn+3AzE6VSOKP
LcR11z7OqzqjtLvmrP8+wtkVi6pC1dF9Z2dVCpcOgIyQ26sJE3TI1RAro2em02I0
84RlEDh5AempBjpOFwboD3/amO5R8yv086zf8Ao4pgQ04QKMBKlGDr939jVcKFqC
3vtkBZo79xQwIhIBeh9zdr11Sbto6aHh0bCD2zzikNbBetNcAME8N8v4oogFQQ1b
2Xpedz7BNxTjP60R4NEnGsNakwldA3re6pK2PLo3p7aCkFNPYFa5zgYnFOakuTHN
4m5DfbN3yxyKFAToIHIk3Tkh1lzXXRbJo6TzOWFka39RdRMcpZKvHdxoMfHjUXxh
gE03fwru+DFNkSbzNtUeti1RsVyfD8J3qWFwizsLCiYywdlTyJJV7v3lHx1NWCM9
/ZsHPPbCWu5ZeGD8Hca/QgU2tPpb0Apj72pVnEV8Q5U0VVXA+S5BuAE/XB/Y42eZ
1zsofH/TX8potSHLZoCjujzHQx2BdT95Q5EyiuH2LFhxSJ4k4cb2lzaMm5etOuX3
22Ns2wjS/9YBzkJHuCyHXj4/2mhDZgaQtB/8XKb2gkS2xM6XGflHSLUQMOTggn1d
g4l1+q2rDKL/GuhthZsUbYwRWu4v93RGjh+xJeB4SYm991N8saS0epFDO5AQmw+S
O3r47CvcI2G8GLropZT2taHlbUT0fEfWUYfLB6ZEiIWKTKkT4rjf6ZU5/nNEYY82
AUgwRinQ70hZGsz2L6cBWmf697qWKoTOB781LHVuUp8AdcvsckHXpUrPWZi65cJy
BcDLNnVW4R8yU8A5oTmesKPP9zbrufWxTJhM8Xn3EUfrc5hklaqfTh6uCqR8f5rY
8KaEsoCGqVboCXlDEImJwQ5IRA6yb/vWm1h34325snueedSBygblAXrPl76W/wjm
oYTM8zqJieScPiCrZvFXPA1yYZmvjlFMPfReeDESp/S5gUYEZgeOF6/5Hhryv5Xc
wHuwbLOGhNz4kDmC+8v9Gfvhw2yk45fxUn/k7KsIUDBkYjGSqsJAswPUK7NG6E8z
2fJqkOsKbpbYTlBK/3Va0z8ligr/FeifBVmq8tu/pT/gSuZRErU7543RdjYkGqjV
Hb7JiRXOq3Dg/KWv1r4ir4xTnS397YxJ/Q4UsclNTkg+4pP0J4Y7uzbMf/je20yh
CWXnFR3Og1cbfQcL/bbrM3JsxFxNj/PfrI3L1EW9BaLNrMtZlpzTEz6Thsy57XRu
oqCVlljj3rUbWb8PrfhSG9dPIr+aJ44bh9qLMjLLTaTMHCYzGaBvbK8kpq3CFRC7
4pxVPuGiazM1RFkTtGvb5Jiar9QhfdXTi607ii9YbpsFv9W5vLzUc0gTH7t4fS8j
V8zBlOVKVuC3nHOnQiYhb/4KhnxwOBt8m/P76+I87m+y/1GZZRoAcYbR7Bph/I3Q
UureMmx67VjWMsNguy4iE47lnK5eZIwLYtJhOpZ8siCQ5xZd93TEPRPATC99Z5Vl
KCgmXkQvAXO2lU/aYBz/aQc8LNZh/pspZTG27EBFU13Igo5BooRjRE1aj3ZtDbTP
SmkUoW6wODztKmN173yLsUGHXqg71vfA2UJ1WlIRsmVKeJhbZwC1RQqw3ATLT3nL
kdQqI/8y5SfEuJJSSk+QrfFhL6iccGPpGMAHw8fOuqfOPHOjr11GCimi5DgIOozh
Te7jzIZqC94RWJ8vTGth7kTbVSDWYTaPwA+FUmUyNHb/0oZ9xvBhCln/3G/knlY7
Cpjeozkhb3j+uy4eOocWD7KZW4KSpJ679o47BLRAqeZu9oqkxBHV8K297e3Bjgk1
JBjcU4g/35IqoBz+U5LDL20QI0GGSi+F6LW9cygt25zW4FMMu8B5g8Y6QNrfU9mQ
gmohR2keQPd7a0hlNl7jU4IkpEh4hW/HhjBA1lEcHG6T+4fCOqcthQjUmEp4aQVz
vpjgXYfzk/aJGPuw2MFfB8uz1TbIH1F/lIsTbb9ShOgFANYPQuHmKEjKfxkdm7b+
JM5R/6g0tz+0k4UI+xjG7y4+SiHqfrijJfqRHHtz4pkMrQ+VMuKpS8t3yZvngaXS
cHNNl5HVyHHwz3Bo3G7sBRFD1lTMTnpA4GvF18Hf0Uv1L+MyKN228saGFyf7cci+
fxcaeE14IF0w6ka4wtuJkV0ui7JVTmEYSjwZth7PF2uwqHTmgaRykhlhVwm2aqXx
CAR0RlMF5iemOtZxp88KVH7/91PIAWDEGKmmGgqtBv6PmW1x8HjP3vxYwDpNHz7a
PoHnJuUw0f0uVNUYWod4w2WFnhsGaXZx9OGbOp2lKonGisvakqNUK8tZP+2KSPNn
AXIgvr8tK7fME3ZS2iD4VlwJeoAgTNP5UxAne94wBxyCb06toCMEj+rSJ2q58+5S
hyvFuiB2vmhZVOr5zPb6KZoIwHRyGkgSWdFeUpI0ArtxOggNK/UPUzSZ4cKww0A3
iA1GZJ/LLb+4jRpT//aXTmMgGeL5swXKozdCFp0u4dqRj1SPG3wl01fglE5pLvsP
QSrfarDCdpXgvcBy8zQk3gIt5R5rGpaU5VG12egeAHEpncqR/MaE12K89rtJRd4v
KqgDJlWZe+fn3CUj96r6IVIckoSCJ7yKjEzXq8RJTRd9cOaMhQDQePcrEaWmXXlt
ISp+COtfmgVyJwALm25NXP28p1tx9F/c0d80cIOH97Xxn62l59Pc98qLRPefkbjh
+yeqJC6tjEuew8bM0eXDJUeSMdf2psxdEfypU8tioE/kVpvaweSvzhYr1g606HVk
37SXIz9pnmDnDpX3Evd+/nzn53mhsiEmk24fiMQrnkvWvVAM6Fw+O2aLT6xfMBr+
`protect END_PROTECTED
