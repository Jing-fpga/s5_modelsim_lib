`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TUJbuICJhUnJRm0QUX9qtj80dM6V3hGT3juFAPvktufq3xnBh0ixrh2opXYOxdhg
ZWomh4DPwzgZcJkHCVY5bb9FYP9qLWpE5O4+LqYn5KJH3zRPFofSu3XeRcmwi1LD
k4oYgnJUZ5+b4DhxjFtar+khvkrGG14FSLVpTZcsMZV4ehdaOFaFxAt0py5e4NgT
PUIOQIyBaTa72jFDDcah4XyUuWYu2Eka78gc4xbTdv4VZNTaIqJzJ3svPvwE4H3B
OzG/lx0OGgn4brxVSpEuNEUfHcdQTAEglxdMJ3PgoIp7XYybnjnRj6au2XXBLBJl
Oo66OrrG3M7wymMyZVG8+Z2gbuChkIFu8QSZWQK6d2pyVThBHDmZzhbkDx+HcHRT
8FL1u3ts1Kz34FIzDcbX/qd4SjlffyZ74skNMl5NTVZ403xWLluqncy2Rzwzz3SQ
prLKf2fhl7hO4fyAETEDTGXNotFwwlHWtNDwEKeVEgXSUMdBoYhwnZxfqHUd72i9
VRG5nEcht6UGYdwzWBo/U7TNKNgYrWA9bg8xEhUL5wcaapLTVVD/Kj27kns9QSmO
sbW13VODoV8/Blqi4dywEZ2FWg5t6Njm9kG6MGs4BFWlUi4aV4YzIJ3liRkrm/AV
KLEMsudEeCnXgK8JxRSwhJWlH0uusQnczqgRz40AvxMBs8Ovd1fT2dAajjPBC6vM
XYyFpyyjQImOrRXfifkzSA==
`protect END_PROTECTED
