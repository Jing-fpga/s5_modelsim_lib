`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6tUGa7NSRqjM9C9fRN8RP6j3m8FNPh14RmaY6JuX5tXC6esHzqH2mtDrFSut8SVo
d7twRy09qHYig4vz4D6y5PsNhegHzak74RR54iofti+neeBDKFH4i7NCMZk9w551
Zd4GvOBfz9RvMUw3BX3OGnMcX7faI3M7h4wYb29QUmcE4AymprgFW3u9T2jbQQrO
HRf27Up5oSJzJfsjAZ+Qo5axo09IVL6JKDk4eApucFD69Bhj/85475hVO2wvSJPX
8JcMAMymTZ2BBjkkUhtc7/mlUmEmxyzvuLh6QKILCx74gNOgN17mEqXgs9/ycoAh
OW6tbcyHYbizL27zZyzOFnUgyJf9l41QD/DlxMQd1Di9U5lBN5H0ICQEsABFjarK
BNh0WsEPsBP5OCouHRAPja+/vNejpESfLsF87XQqW5bTp3P5JNIdIK4mAEQkyX4v
kbyvEdkAoTIHvXCrj7tCdukyusO3tTyyBdwzi8GwKVWXfPO42+QRYhL2LSm1VWVe
tGMPtjj2fR+eSVo+HXg008xeqwtbhbGlmGf/61bOsGmfP0KWGdfjLm7Kt0ZtPX3c
z/+I8WW4wtSvysrBICdsYNxmDNGv7NVGQMyAuezM4qUOJdpbHsqu9K0PdLlGX8hZ
T2HU/0s/zRST2CZW3Rvk7n6sNbkeJHea3Oad3FJxYrxJC4T/mNHULpLKMczyEbgA
GT8ZLF4zCcv5BvcNzXkSQWXw3mDhhWaa3e/TabxC8usK/CVfMYHzXgPLKuxIsmGF
+EHadi+PXEi9jhD91qy1Ssl0yvQouBoLjk9rrEzECN3lUwK7xvYTPmjISMd9a0ak
aVYPeGZFAgws3GzkyVREpFFEP4mYFp0V89yR1LaKddp/c42qKrIUZNNUqODGfb+p
dXQ6OYT+rrj8AQkLYfQu1ivC/8IporpYNlh33SossiEQbypmj9iIeVAoaI0MXgwo
6el3FvPPz2D+hoaTJLIoFeFR/+G8fuwWfKpI0pQanRsYexkKX8RQBZMPzQWjHv3F
uRpI9VaEk0e6X2CsW5ZiJduTK2tddSxzFjnQdBB6Co+exxIGYgiBiKXlIVxDz39a
L5xBN238QKMn5A/bjH4DlOIBXnbMFZrCE2tL0MxV/4m9ukIyEchVpIyV5Bh+NRCv
GCbPpg9JTGB+i4aGGbv5L/+ut7XGyRk/RuEJ656iHaDqwHWAT9n/7MI+mAn/Ud80
4bEEezKIHVX1z61C8cDMhXYbm1jbjH7OgRbecn5KDOyuEoqlLPxU19kNJ5ilXgZl
N0Y+azIpn1Zfdl31Q1erCb8kx9PtIw0erYFuBy3laYOnqvmg3CFzlNo1xdHO6E1K
VD1ldc2UERVudFCA7chw7POLMrsGKAuXjzUkdiRmtIba2tmPHTT2hvP72X4SZRLr
9YPyuBHjxX16pU7VlWNorpVzAJTlyHJaEbYXH0LIT8OFXtR20Wki1MDlURtFSp8G
w+4GV34V/jRTVAU9AA9kfw==
`protect END_PROTECTED
