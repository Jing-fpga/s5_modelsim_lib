`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5wIzgqoRga2jVIu2Y4EvbpezNSmoXJ4qkFsbdsCZaSKEFD9R3A5SMI88kP/Or3rE
MPXDiGcN4sTD3rGQx91oZshko41bjkZ9fCIGRszN0aoiBo4mWCIxkwMjHkd4KqjV
TjO3AeVoK7jRPs3HZ79VUVBTZlxB2HhfTb0KqxWIalesaW9RBjcBmVCepjBFx95+
11GhjUsE1Vo3EC+2AfV5W37PrlQWrNHyd9U1ihXRKhG0jHSBtik+qVc02YV8rITs
pZZcWioDpIZngiZj3u0cMPFq71WsdykwEtEHaMR7Ax5GGsa+Ayk1VdXyYgiVrV4n
XY2tc8pVJw4VUcGjkweQEQRdzZikF31Uow2wTftIKPXAXhvCsSxRqq4zEEekFqfn
BJyZADSDALQXl4F9qvAg8F9Qsb9Rsr12W9AvcW1PgPb6OM6vk1yQLqsZwYXGJ3jM
n7p+d0HwjlJeLA6UuHdNVqGn9V8UZU5OsVgBOYxlpvEyK5O2ZVgd3iIiyzvsqyhq
u3tHrvdp+WieBRlh714e6hZoMI/yBB75K1kLjDiTEFnQFxcWWDyosJL9ZMzsRRYQ
/ZW07myviKJuoA2cKFLhrgQIAan9dpxg/S5eIYyuDt4rlDCgUsfBX3ga4UfSSWUi
WMYYvwQXgNSLGC6j6sKQvdug2jleTXZvyOed7lMxVxOup6KFNtOIASPfYPBCFaU0
cqOTtLInwN/DMKh/D/vBf6fFKb7gMJ7f0ru+pArZ1Z/hshqu2EECouyw/WN/ufj4
/0jUMoTwrFHfaBR3cww/I23/kwW2BJ0BUTz8sX+85O2bJd17Uc/Oxv0qfLonQcJV
4GUMHOke9DMwy+kzKL0WvoUodj1twppC5F8b3n8Mo6s7gZ/zU/+xueMQ63Yzjqgh
BEA2WEsceatZj0aDimq5DKWUYkIP5bnCcszNpY8A+zyyGxbxZucT5Zs+kurHrPRM
L+mheTpzBlDVZ4OlSwS4dMQusk+/d4FssnpUyu5+b4VwNpgjRs/oO0jdtzKIL6oO
TYEhCOFQTQUaeJXcH+wmMRTw8cRuYsDef9b1YcPtiAU1IWg3K/U1ruiol5AaTdNB
5Csk/3uQBpLfWvq1OyzAGQ+dVPewfew9B8t/ccDanu4pdsgjVIirc/I1SEpDO9iJ
G+aunTCPWqcPSNvoKg6PvLHJHiCUwSVwOSOOpARUbcWJksIvvASU/WM+KkhyGfqM
UXhFzSBVMLs3OlgsteazN3Xjxi7G/+cLQFX176oQNWLp78AybLoX2ld9B0xufHt0
YLYrGR5JNYyqo0zC7D1wokXO3itPwb5LDz1UjLGWqKBbOooslJi/z2dDfthelN3I
G946aBqI7Lht8sx7jx8jGNXpWvLin2auC/nOx547FGTfzHmYXDAvBB4ocI39VzBt
MdOzmv5PkagFy44gVDabAZhyO7SqacjqPAwjd7PO+DFxT2XvY+BCXG+GRTTfRvVn
8IYRtz2IBc8vJ1k8q+zd455pO+XNv68IiuyDApxJvJO8nyaL9EhqSAgoAENDjk+x
HuSKhNdYqQvKRJ94S19lxuHB/nJInN3nqic1polvYa1QGH7tR/sRvNFd9NSg++WL
v2MdGhDjIt1ptwJS+8zRPrH7fa1ASDHouo5Z4fUvOFA7+i2GMOH/lgZQt5s3tz9c
48Cv63qxjNgJ70QlkjMPU6fBf+AjBODrnfZnSGKrjv8qVB7tJF1peEu+EM6nvW+E
Vhl42H9iN41XkGhbLiYL7olH8WNxKeqmJOJ9wEph1/oHaW67AIJjy6SyO+QYClcR
3hnDMHZVXzd3SrNfwKThKAggOFu5JPacRCVN37OYaZvV49m2nMPtw3l/92v8+bCJ
j6NgpqkUUmXKWvtdNS9DoEDa2IwApTs3ht6jLi3zSXHJUwQCCSYbCw7ZSoF4+1tu
apzgjZZd3vpQCU27aW9f6saHIqtTtiYIZvNrJ81QHAod7cEmiqSBQy72RaTpU8SN
wl5CYCA9yC7bb63z/cKi8WTPYOZ651S9wf4nsofzixDCi+v0/942nbBUN9ilANh7
zOJbKtXc9tqstYCcTs96cga5kj2VOxzgQt0FcBIwdIxdwhRZg/WgqSqZQ++TssJ4
d8rfniCQewQQMw+AZo7mKox9hvtqn/h6Y99eNiNk8gIdcLzUIIl4yv/0+ep7zqhj
LxFVdCK16kZQA5QB2C9wpJPbnSQiZ/2KKk6rjJ7U+GNtPPPhJFqomDXCcjeAD3jn
2nuR5h0SrmipEJD60LlQZWMtunmWcx0FMbpITX2tZ0UQF/avHUl9DN8QoGQwa/P1
qkIoUZkjVeGvxiXs4U7hJFgiXfg/T0vzLyyM85Smz0WCN71gT6Vkh7ezUc/gNRUN
UahNqV1RBqQ2Dnl6uzaPsIGFNZCyD20vIAl83Q5JZ4j1D40I/8WrXvO03DxANCYd
7xuayaht8V44Z/upfh1nAJrnYCRsSzl9GVkNDXXhB4M3CTkNskxuqpDpJNnXNbv/
mj1HhZN6S855MRNDCLsnzwtbZuTbbXriANG+mSH+Ply7VqBN6lo76K88LmPZOm3+
Z+dFP3Sv7T1UfZUz8HQRLLdcKPetN1P2fuC5L93k9UWuDVd/DHoYzenG69rtLG3X
rSkh+i2mMvTuaAHcOLHFWodT++bryWMm9S1eZiIX7o1elJC4Ch6enFXnkO8bDnTV
lGBPSO5M52dl56jqeOqopZXl67hXyHRnD5vcozrEgAjgrRwBe7Pxx629fO3t0PoJ
ulNvsYdUB3Oe9E7ujnJf48mQP5RsEqzXRVxXj84TkX/1WV41qLIOSkRXsuEUXnLU
RSz5Jl1TAUzqj49Ws1El1E1fOBA0d8WRci3bF0BNi8G0LXptRyEGuKxro1bi+5Td
ASe7KstvbH2cHby6MbED/DHL4VBMfG6WmaI8tUsYzCDiOp6JnsyXffbznSa1rEiK
uzj2NNXNonzdDEFkOcg9/SLWVjRhnaATCnUNdsi12RMYI/YewP0gvLQuc2OleECy
XeIOBYjRAg0ATd94qX1V7A88nIP6+P4jWDJfkOxHe0ZCLkSNUEbxwXjMuGmntCN0
8ZnZ5avGhXJWwc7V3emexsQrmj0jKRqzK3UoHoOJqQ7HJ6LxGR810XVdI/p0VRZq
JEhzLDva/GCZrtJxJZ7WzX0CTiLw1JwuKObJl5YnbCtmG06dP6xgWv5ae/y+yX2L
aykj9VzRhwOIYxyB0M9Lv/QEfwYr2H0FYrcbAC6eIC5avhbkhF7YufRQtHQLSlkB
8+gb9flmVvR3k0NITkf5rJp2aajrY/AVsPRWNadMYeYutm6bkEQqMzkI54CFNYza
ak6+VJRpWMlVxcSmhJNQVRXDLZ+fogF/KSCC8MyoVD4Hzkysb2pxOCmkstUtAsPw
C4Gyxy9btV8nmckOP7ZllcR/Mz3c0tI1UQ3yyLF7eiJ6qLp8taiMlZDXJ9z1qj5W
NKFT84zZTpBqwa9C6uv4TTYhOZ/9HarMqU99ncLYUEhsbunmjfR1iYj9gHMT8RX+
GVdc0OApDiWmBSuYIN7pbdkxLzblFjPgfJxoFkb9N9mEtsQqyUman1kjmdqgM2/S
3yLC7Myp3DcXlVmSac7Q/I8zN75vgQD+Qz+Eyzw4VMBklZKFPIuDWHbv8kx5CEJW
GcPcDWiarKGJZmeFwXkgwEtowboj+ZwiENnFpPBCKgDM/unA7ohv9tDRhrrcXXk4
s32svS10DgeCwywNpQlI2y2mg8YdcUgd7mZSBfKgSPVwidbe6VDdoVDIeR0f7RBD
msyE3BzsegXlzTtjFuEj9ZCtek+Y14u45eAWhg0yvL9YqX3uunRXM62Ftm5/PE81
C00p1ZWQ3InQyn/lWxNt+xx+yub7R9tz3m2z0T95gtLiJeB+uYXLf8bCqojXBPNA
aSqcTHQYlll3sD0laff/9BZ927ZmgMNDakijlZ9l0rYXE4OJ7MQDbWYIVzIyM/mT
kScRyofzN8gjUkjdqDvdHn50//wRuiz0DixjwPwfomZDdIaXPe3N5cOnzo63lInb
T/84gdlQSUh/cRXNMQq0/rnrDQhm+HUuUUbR642A3aaCDhlO+8kwf3gNAmRQHZEp
8SE6FHWx+fQKNqo8SFAwpO9E80/tyOv5HXlMmgEK8KNk5flvDRiUM+rtcj3E0sV5
Cm6IOs2Z8iyVfdh2PiyrekItaW8il0SBotMHsqOeJCRNAtOVdMn544TpxN7CRh9w
unaCUwFaw/vklduO25cMe9lAfvpVrUjoJg7rvom9sb8a4vgo5TDWcHS40bXf9AX9
w/tkjZDRy81MS+pN1Qqt8XCKuzqu7nvSWWXlLVTInCg2R+AlY5d5E/pFOtfwX9Nn
/HrVTQMb6EduSxFoB1f1T/ppVkNx3+FG5R6+kPZR9skYt+5ycV07OZtqUZTamRzG
nRhPsGcVkyUOOfg0R09LTr34yswYU1cITNPl5LSJNPP1H4PPaeW4W+zoGoHiycu6
3h5Aqz+i6XcoCBF58SpWOSJSIsDcutMwszjnXc/x4PgDALyHp4Q2M2pCWc+uLdFq
yKoD5ikyXmihLuIWqr2bzyUk9HkmlZ3r4E9oNukx7A46AjGnvv7GO856a4YFFl4C
5NJePgewm6ntmWzfBhm3gVnGY3F3gHoYNFkD6oVjcVDYCkyx7RZgVFlEAgU3eIn/
ppSzBkW/A6zyamkc5fJ/UVRbJXITuXPD2LLh1TBXf4V7yRap51J3dAlnLrQ+SP1w
jrETj9mHArHWrPyubcJkVOS75UQMKFVrIUsR7XfL6UzaNqikrxStKJUmy7HH2dL5
VhkU1ilE/MB0luQKwQ9H+yhaI6ie+uRX75J86Lsqep1065lMRf86JfptGb/BpvSM
0TX2OEaVdP5jjKOhXWsfpDl2KdsfIR6zqG/72HTi5nlmtVBiqDwFNyzKk+MNDGsn
LQ+tV8dA9aYw/epUAETz/RO1/kejwq6dKVpoQHMfLCqDU/8XTmD4lbggasiOlKg6
9P4RZeY2VjQ+dEG6H12U9bfA6Cg6XIqquUKxXvbzvd2xG/Qm2D5zIVFleywTRJKf
+q8S8paZygCudGpWXCOEXAiTu8RsNVjfrNbRd3S8BIenBswZ/7wRdYQb+vNk+CPR
NFgtjiZoWw+SQ5k+Gzdahibi+M0SlNn1EGjRXxutq7hj2M2XV6m3YkgVd/iUyH33
DLB+4ZW45aD/4PvBMkU4VMThTGHCdiU5hqvIyu0aHKgkwlZ4ONL7JvfpXVb6Blce
z7ihNNxxPcbC7z49dTEZqfl725HGVZs2rG/aYDTaCC2PkizDVfSXBd/GZqRLIk1g
szsFmBhnZJEwDtUcZCEJUbcvT/lnrCwAOV33wWMKk6AQ+BVtqUSE8WMcnyDx6wns
ooSGW5djB6q1bU9GAh7s2QK/FauQKv1L/weCn3lZI4/nqdA/AijtGUdUtCYRSmwv
ijrJD5GLgDYkyH1AHpHeZhH6WfQXKMIjOQGNHOQqXITmUcLgjv/kCRswCFZfnHlP
TaFTI/Cd2/2IWtU3FhMZ8w9u2LeiKpTQwC3iRzR9wYY05of7y/ZPXCUGGqejTZcw
PyTovwCIYS4EqGSxoSfSGdQ3R9LnAynxcmlrt9m7RLpEBhXNW45NC/lzO9qR/4gw
hq0JxSaiW1gsn+B8PRL1LHb0zMkgWTqYVggXkVHk41Ll8K0j2EUkNJ8SYIRloqKn
K0axnXIBOMuuTm8UQSYDTV8R88Wu5RQKYMsv5ua2UXwUk3eBwFJoKnNYz3ljtWWO
eHVA07HWZBcyQos76V8DXPIolPiEFf32ovN9J5hfZZk5tuMgGlRWRmuM47tJkn1M
71j0lnXXbKTv/kFy5q4BKIQiLp/5Fd+CHNb9H90jfsiK8zH6HIKC5imRzWzPung8
/c4ObB0C9tfoogt+fE3aiMX41OEi1eoYla/qM1b9t2H3T7oWPqQ7ckw3aaRUPFec
NRfXTvUFpjXYxp/sPU7/sIiWpcZwnUDsyeTc0gVjH+XFL4haUuIeUFoezZBzcZb4
hODSF6n937tdX48V+hIwC3lw4ltBDq7Y81ZhV36EGJb8+7l9P1l3CvrBlBUw9MF9
Qle2d4kbcFbV0RYE/9HiF7pX/J2RZ8LfWuZ7p1G8Q3/2xem6y/lECPq8DvZ9aqlI
NW2LGmreNgmgkqzgzx6rXXTzDtlhGE3rm+6frsBK1aLvM6/vsixdIW592Imo66w2
ldKiTbpfXQwvmb52bxQWF7awNxRORAiwXuqzCYsXm3LFLncRH/voDeRvzQywq5pz
7MCcoBd07k5Z1nihmVHjXE2Q/drgAXNQgyaosVzBKb1prOeIMXbpe8uuJVVpYh9I
acxwyttbY/zVrX2/E2ER8hS57V1s6xbcc5RusLAfotypNtZ235al0191/i3D9jYf
QYO41mJKrwKfwfd82HjeKJ8QZ70o+fRYgiRrObcFGBkOG/SD8dxAw+ufsxvCmVxt
bgR/9EfR8c0z1Mu8nCfOCWrsQc6YDVYRinxRP7OU83ioPjGOmjmbHyIm1FjAVlUi
oKJAIBoirMkzYjsb877g84yjm1s2wVoJjryeOKZzU3Gg6sjG6kOzBOxK8E6qk8PL
etAHC33hcRZPnzOlY4e1b6Bdsx14AlRbrjvMmFKP2bpUmP8M2+juHa4A6fnWSGLH
`protect END_PROTECTED
