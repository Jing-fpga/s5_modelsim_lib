`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8mIkwVAh9p/d8h1qKwf9dGgH1SzOlMcQnC4AZo1HIR68P4VeR9FUMlsKfo61c19i
MLPYEcGCcLE4H4PDU8MK/0fjwiOXQfMGoDBydN8ST+ZC/BYu/5HeCKrUsliGWB8u
HDTUHekV5bBFRaWfM/ycAtdGEbHB0e06XDU5nsqxV583fRhGrAD5wVEq6kpOyPpk
X/zaapgI0tg+AmDei2Tvyn9BfjmEg5f87FM0NbM8sLZ/XFGfGH/UqrGertuFZmzA
GUg0Y/2LYEq44TBf7dLsRpcgxWMDOHoynn2x9poiPVHdY62FH6u1LiY1bDmt5zgW
rEEPi5Y6EfQibSPLNO3bB+P3e6S6J3EpmzfqkU/r+2sAz0+WEhwJP455Bk4haRzZ
inuAeQ2w5rL6t2MTiAy+Y3PhcjVNQuo7MueRhankxQ4OtNZkaPr5S6Z7w2A2vqn9
E9T0K0fRSUA25dx4KTTa0iW6pjpkpdtwp6RZ1HGomfvomGaQJaSWgSjGTNVAk/oR
ZOsBkYU4C+WcrlgX83hbw0Cb48IrSFQbcdNP5p8hNJHYaBTTKJ14d06coWG8B+0r
cfZo942sBJDc4C2USAw9V9XqS70ZZ0xihV0b8m2kkc2LBPub5RSBNaFMsx2Ojobf
Nimt828RQHoCUZtvFN+ld6r7Jws0mc5L/UoG9DhWGpr71vFdAo0RRC21WJK5azQn
UPTNVV+mnPIeIMfGyJbfeJtLG7EcJbiLgM2p7w97OtlHv2Rq1xSLE7f6PfRLm8IJ
y0u2tGD5d5y95ZD27gTNAfjnR9pT6XcvvSD1uZHBh1fXscPQdVmWsmj5lS7HICv8
gwyNjp6Yoo770BN5eq1ifVJcahH4l9/27FHWm7sIKLpMHw+bU8OMtE7hRbnz7gXK
iGEIb26SC9hWv2X1100ekP5c/xJOGikLonP1nDMDWNibgRpGXzjfP90nknYKd5/k
kcPmGt1EaiRd1dVEobfuM3nVgckO7HDUf6FaJuc5nk/SuQ9jfyYOLl8XOlI/04kK
QKVFGuUadiPDbO/sFnW8iOnGyqKeFZnZg4AhROyDwOM1jV4UaSi0DK0PNC6fFwxG
IP8GsL6gor5kgqcYy8WBNvRdm8j7dGd4P0y/CxUeWLsbf2tR/Buc+CKr45EBQVyf
PLgCfr+nNRnRbbvwrj1fgTLNH/fmWQj3f7FxcaLWBlT5+6WVEx8zQIxq1YfNNbXK
DKPQeBoeUv0o5XmVzXJps9ZXpDpgbpJsukBoVMgc7vmANwLxLCcjwcShm0Qwgb6U
69y5YSJSGC3DP5xKkQe4s/wkdVBj4zc7OyyHvbxFbH1GdxP7bjV2k8VCEBYELA3J
7W2TaVQ+O034u8EH/1oEGXokEK/6gW92OMTaCeX/EZzTcjIwSrTuptKiqW2WBri3
FnEprvm4wyvVbUl8TtN6rMyjrKmegYFJGzDvfO7WqcelzYmlV6XNVjCC0iyhK935
`protect END_PROTECTED
