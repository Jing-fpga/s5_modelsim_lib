`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rXKC9Mj8LBv2q/xfCkIn01gQTUtqKF8KPV9FaWN4PdrrG5gxeGrSBZQg7Clph3MF
klUaH6sVCcNawGv+ATOTS1FO3YE1pd3l6B0bGP8qCsOPtnOL/qYjaLXXSXZ+2gyn
nMnrSVbMFxpfdlZlvPGp+ZbH+UUX12cuP6O+5Q6FjiGpRXjpiH2P0tDrxRqtiU/W
V0VHTWD16MKoJ4DvSg9Sr5VaLbUK15ewiUsVXDpUxTwEiFOSGqelOk4Fw6SgYfvD
+cSMA3h7QdvDbFnUB9F4oIi/3LFEmKHvJV8VcKzdD2DFf8vDM3s+fVDJVh3xSDuh
q2CVUg+JfhD5QBtECtzISCEM3u5u6E1v5ArPmTzFQ/upNd5uHx8lUnLkm7eEbDKY
E0QhlUC4OjCLXn6IVsShmDNojJ2VQnfBZRc9Yg0Ohj7hoIAPpOJP5exNqeeNNCZZ
AKoJQSth1DwJGZLcMKT282UOl4r5RhHgXjqg8Z7IBzVT5iMiPT7GTQjRnYxqV1N9
ASZQvfOQe0Bj6DYD8eDxituhB73+xiQhAsQ0/RsbllktJc0Ksea8VCVc1Kxsizuo
qtJO5HOfzGJjvE/jHg3IXzvq4cXdaLqV8mCbP0E1rZa1QIGGPu75aTp+c4HTIhPO
4plG23JC/oqP9Pnrkli54jCR8I+r6NEBZhENCs1pKerNhi2boQ6QMIlKyyRErVJj
gMmHIE/YI0fv1fxB31tE2cM0TFYzt2lc66Cq9boPyNc2AR+G4qrmcNcJpqNgX8Bb
xqGxTjk3++I1LlVB4wWFLD5FyrM0libV0er+c8kg5TAE8X7eWWTgKThqyjl5YsHe
dhP2HqQEazVcAbpIVpLbMetdJDDtu8zp5tMouOKKuwg5ei3sWsYymNgmfFZ09rrl
1zo/mCLy78T4aDK+2qdeqCGs0vVnvJF7HqedEFxsHFhAzJLvPdED9swpKoeU2Ppz
RX0PkWS+ft2ZNxLIDErDDIgfBX626KC7l5lzX6KOyBixz+SHDE4ivgsqWlr1EZ8G
mZ6QHm5QUUHdsUoDOMS+fbyOn78+AybKgVkuRCWwV3dzTDLpA0pFU29gBMCFA3dV
tW5PtX4KFHVYqRe6Q2QWtw7Rw6Tf7u9UW8JYUKQJh7wkXzGv9131KusjmdBrmiqg
vkJWxORbJlHdeGGJktRzLj0xO1nT4np/yvAa3qFvDyJ98SyUXVziK70RqXUnBCqV
+FfajnK6w4Q9gPH1b5gm1T1PdpQEpV0DMnLSO72p69G3Vloz4uAnrOwINqCNEvuT
oqsgXNp94qHDl6uEpn0l25w0dR1vybhW+Sd4Hbae09mzyt05Wye5VMp7nXPT2Uet
1JjCTkRYVC6GY6LGO6EXkCFYH+QgJYk1/G7JfTKlbB88Z6WTxlQlw/NUaG4nfzVG
u1OTWiDTxAVnKaqcumevaYUCE74DwcmdkWFvUNo1M+Gkluzd28gOS4NO3s8iDRNB
JQexS5dFxgr9Gg6TON0xrOvrlB8wnPfHnrRIdA6Db1b4R5qXfYMf5BJHjzW/9iED
zUrXQvWkodSlxZohUZgz0vGyaiVgQC9PpJDBOrffSYydDgQcgZHv/GWCqtjSgIda
KRoQ/8Q5k8+nAAXH3U4GK7jlNa2nZz65+bEro8D/SXvYy2IqESww9xwNVI9Cu2zt
bPGwsg5DI1rXLZEo3bZ/IgSPBXYIfM6+E1a9qwhEj/NpQFE/kmHOu8qbApa3e6oK
JP4SU+gOg6CiUSkLGykqoVQKeWV6rzcwaPF50cSpzCTmACbo8ZyZwRoiNa8gpmh/
MgMjjgGI+ehn8lP04MnxrXIHrYt1v4amSw6xdjyudEZlrF4U4y9YP6rcz4bgIZ1C
QK/b5rxKTSV/dN4MpEmpiU8DwgmEqe2DuWDG/HByAh1qEWwkSx98A7FbO/0XE3TI
PCrq34QJ/LcGgfY/xx04+UKSoAdKnBm+XW7QKFwjwTaBxyigimcfHCx9QIEjQeST
q6tMbxg4WuxGQ6lq3Fywtc2DvcSvr3uakih6FPCVlcoVfkJA+41mZ4USvqbAliK2
JS2URSE8p/eVG/dIPeA+tLey7bH/Y+RN4NifSDZyVkWfkPbZUG+bVO2Jmue4plwf
ttwxA3UhCecwx76eAMoxDwJW/eY9ETY5hNSLDX44I6cydi1qQZu/9bGSqGnxCR+B
P2OxJkf9uQ9hsarRWSJ4IgwMBpnJ9puvX0dry4ydWtW3xmydHX8xW2OXu4dahWGj
vDabm7IH5+ANFQPTP1XaVti2SMx6Zkyk4XSM3uQYWB4njzziiEnCn7AxsJy8RQz8
21KE30hqCERgnXbjeAS5NE/eenpEIEbGb8m5Q0Q8enF3uqwSQkJvL+RAJSpbj6nG
qTu05KbpU/0IVXc7GRPjQAAgH76eC6q4BUEBah9NlRdmGvnz92dTnl/Cv1b7ovEp
Jj/Vk3yleEN8+FsqZleVKUqq1IXwyF6ALZ9msiJdrg0cFxXfHcsQazHWZp3S0bBx
+1Bue7ijug9GCZcfgXUL15VeJHpUR2kV7b/KJwCtTSkQ+t5M5rdCPr1g+5f+guLM
nVfx7lrjeyuh9h/OfSqSnz5SCv5erJDo4mWDFD7zX1mtsYigHdX+Q4ayLgmVE6ec
ZvJYfH0aCtFpe5o5OS3+AVBz7cEKBgPzWZYXYhM7ktqtW2+KqoPars9jQXyGc1Sc
M5bgyivK7FToXpimJBL60pPatQnKvXfII2BiBATTXhqYpHyE7AdIFNEIFJAgC8+o
xXIn9HRSrX7BU3nPVA7DrIsuL1JLsmukvbjWaa4zoiEblOHv0N2Cptd3Ut80DxfV
cZvxi771nOc7jD9vMgAhZMfaTg+Sucdb4CdqQs+9sTrwYw+dVEHBaRTxUZSJpMuB
S/2+wAP/6Wj3TIujESZa+tpJ3SNQs/6M5BqbwOHQ5e/phhhQgiyUILwgdI/dTkdi
3kzy0N06zfLlWb7ctm25OQc8M/i7CosCncu++2xMysuyxp6nNzS+yWLb/0L1/QzK
b7JymLCMO6QT32+oxAvycxk9egj47IS9Wq5/nJKeF9+sRc3AAs7PstIKaAT+oiK8
/XUdrBMm88sz2D60j0STwYzQ62fv0Yoem4NgnOPKdTpQSd4RmRRbi0o/odGaIDQt
YIwh5DpoeqQmMcJk9khFjvDex8p2hPh3WBeTcKufTk9HOEJRSTkm6+BaZ5Yit7Cn
qQid+0adU+qNOx4CRRi7EDFw3G9wPiskPmZ7ID2n2YRMNSIjy2VkxOa3HpldWegW
+xpSvdjikmiJieXCHhE36vlWxlthCyPpqPdB2Sw65rxnXhpWovPPGMLQAmBdUBK4
gAlhSWhn4eWIrCFagehV6Cn9SixaZezj1rmehDh7/Iq+a+X7szJpDYFs9Ind7Uy0
xSPb483vs+/ikYZhtJigapmRSVzGVKS7ztxyQyC9hScWl1eRvQHmp6Q23xFXPcJ0
p+j8S9eSpODtrMLTmFhTSHpjpU6AuJ+mompHwl0PHQeJ1bK5v0+119aDhOschb7G
Kxa31XGW9M2NPcS8OiLR/jvnOtvhLVjGiEnMgSVuPd+9NwVv32EVPQJYrWA/nGuQ
6zEOuMoyMLiXsP28tuf3AYdVSZgZ0Af8hJ8xddrmrZqx1PI2cE2mQcaMWbLoZLCS
0cVh98IT85EIbZ6bj0T5D9M81BOfQs1Eb48gkABO5MVA9e8Xm1rEECZStNHFsNNt
X5mga2PbdY84d89M4frkclq4XLrTtowK0KO6G3tVMWpNXwaaOruZbfrUx613ypDD
HBc9/A+fW3Fh1yV7/P2zE3sweafPqw8OX1IYIc5OzVx2NCga83oFETXCC6omeap0
UNortwPGuSt3f6+lUnq15wIfhFwV9fVS+kuEewHH21m8aphioQUl/5+1uyeFZjRm
8Tv0EmjixnhRdIXmvsJ9dp33lEIPpvhmwjP5OWDNd192k6gHNX5aj6qUXGxTMaVG
i/CcxmEB0fvuJD6ZUS5hiCBvY/VQqRkRcpJrXnyBFOCOvkS2tv38aPz8199rHh26
8e8CyUFC6XzC/5T3Kha6eUvxRv+knFg5DLMB++rri8iewMvJs2w98fKMpv3BF6Vi
cstKvZCIEODGSqqP5KFNI4CLvML5k7FW/4GTANxnEiJjJ+8fGtRNL9K5O/YDbbO0
c5dJXwAaXEFx99P3nudatonJ5J4eoS34tMZE4TEpomRObsNtlo/n6tO6q5QqN4zX
+XemerkppiBQ+9JEzj7fUP/dctDrKCa+vU7keXjHAFMQF2vx8mFis0OXyIxnZoKy
M24rFb4NFeITpa3clE9mrLXosqvlPjtQTsRQ7i6LiRnV+eZOhUFXGqcXm1FTn2CB
11A+cXIaF6iMCqcPd9gqYD8hNmBiHpCTkVQJs53CeNPB6A1eb4Qh0gL2JQ/yoB6X
SJehS2JYg+HUhEFc4MNjfPsmmJueaT056dqbVU1PD/M=
`protect END_PROTECTED
