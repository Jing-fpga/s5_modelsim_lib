`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Ezt8svvVD5ZWPAtmvR7gZBPlV2s6PsQ/oJuvXCzTgj2yGLUSNC//EfKjOHk8Pko
hpzknGvX3bdigz3dQ6tLJJ/XgTduB+00rxYOZqVtKPMnVh5k8XN40Y7l4yKzQLo4
NyM3tH9hnXqPRLyXPKA2sakbjEiSyKq5X04w3KtoREQNZQL4VfGwoVBrl0rWF0dK
o4wg1wRKKgXoBDRd3FR9RWFNUQztnDKV6Qo7JV7844g8hu5xvn9mRTGgprMKqYyB
15R/NgXlVEL0i6250tsJkC5YbJczbOLh8aZ2A0juTZj954Hduj9a51pW3Q1HyCRe
NVtdWA4FXBKaZ7uafUag5Zk7Vwgjwa3/NL+/juez1okqEYHjAv+pHSDwlhdpAy+C
g2Z97tIyzbBcT+7yMtXewMC+IkSjIBpcOfyn6Cm0jlU7hFXv69q6A4Y/iTVorI7I
tmODF+x59QerYFgKP56eV7kHg8bGqrcaliEPhHbr2+XyJszQIBVf9yQ2iGBwcZzW
wZZx1XWeq1uBdM3c8j3m1R+GdlV8wJTJxhUahHvo+kVdL4bXLsNCwYtbae+XaSDu
8Kx/Q4F29H/qrd6utscfotakIRg0GZX7461sNpD3cZUrMR7Pm8MIGYFVgc3NzOae
U+96TSK7p1EM0Loxv2B6jabiq9Ev5mBY8Zrv7TAd21Kt/tBEAlx34+3EhKYGqM39
KV33BYL7YndlGZOK5cZyE9Py2Oc4ChCtCiguD3Izhv++YjJ953yKbgX6AWji0HDZ
d3P1QyltMijKN0UQpdbVbDQ6C+bUQYi/1Ssx5uKk/sLTxLEqrhiKRAA7QqOKYATW
1UpIn5tUY4NApIvIrvVmXa7RTITx56KJIbvULiI8PhHNJUYtIdRXuD7wYS3S1hcn
dZrUB65iXAZV+KQTLf4ru/gpo4/k4y0ijC/GZIruXqgHSdxM9DUphhye2dVR+Run
jlAbYvNqLm3NbdtJmsI6VsSrIOZNOtcclT5wIMjhPd0fTbWqZHiDi4NGJ7w4cKvi
cJQEqmkcNpi5nmDrY3Poev6IYE3guu6kS6DjS82MrBVOSqUl4yl29YnDQ4ibKWe2
jERpoiAVaL+QqlSt/3ekqPwXY6SDIQy7/IFktgi8wUGmwvRWlSTmqPIBwCz+pBYS
5WriHWgCaM2iPIuXsGc7xya/3hzTSWwTEuQs20iMXJSdHrONfspp+6UoJHfkBAvE
/Bn9m3ko5hRBWIjBAC1fCKJnHJ2QIHifZGdMeLF+AfQf9ePF+9ndJT1i6vQjz7Ob
r4e8r8mPK9kgaxFlx8qyNe5ZVzz92gEJGoAj4Lfsxt5RBRBGofmiOpZeA37miHgv
F0p7fj+/lNexqqvaAz7lbu85uGFfNS6+eBxwl5S7big=
`protect END_PROTECTED
