`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvrN0/7OZbyATpSGrJ1Yvn9MVzv8as1MQTbabSXe4Qduxd7QeeTiHnZe04EwrnqS
pej06zN2W6K6NJ+xzKaH9jVPnpAAYFq4SX6I6QBRYuI8VZ7kO7UvszKP6ICnY3M6
F58QuNbA+a0PGvBkqBxooAfbCFqVWSrtzHab2eVhWLpyIERedDy+xAjnPehQ3/6z
W0p5CNLwkVDuLrYOVxWyDbu+GsIXHs99izbRd7oS/RqA9IZYzkEqpDYw1zYn4RrB
oDYXig7rBy+jdPC99ji5wtkgeT8dRboX6eVF319dynip5gXSaRWUzXSxPnV13k9J
4tcfwOLVvK95BOG0bmcHoxnfqzXIQ2yrtnLXhXyPEoEpUjNaR1j0Ys+dAr/68eGe
XYGWFBmTxkxsFqUAm+sxsgr3z1FkO42RPWMKHVaNyLGi3xz8hl491B1kRZ8gWWVD
6LpMxwCrwk8Atm9mYNkMEgjXsj0aIY8Nkgwn63IyJe35mt9tG90FZgsGiTq5KLhM
2CQeMmnEXgzUaN18tQyRDyQYULHJfQDIbk5uoTGVsYriz+R8cgE7kgqMCMUUhOhr
q0tweVywt3LlYtEi32QeJTRaSPDy7OWNpveuDryNiZap7lEgJO4+zQ0fFLXwkGbo
0kAIDZ1JR5y9t3tM7aeURxcu7JNDindIUfUbOc/OAh4a/PgirX8ssWabXRMYVIFS
HKGpCg7XQprhq4C+lh8Hk2/MQO/yJcntC2PxRansowUrfK1U9qbuAs+PNuuZSGPs
ivgqIgfAWHms7vBUNKYj3vdjA0yvI8tAXORZGHpi2QTR/ih4JHELUsXGJIkgajue
D1ugEWE9DiKumzlqO62fEmwyQS8zcnj/LVGzOjdGkSLcqHMX0r/wefMni6uqSV3y
b5ZwLFMzWTCbjY4tGSUB30aLTREvwGQT6ugPflZ+fE59cVvmMG2WFUXPGlENePfh
+Ft+DT7p5V3ABjMd/bxM6IR9QdPEut9zvDa30vBFcrVoD/L3MHJ6YcXXMGFVp0KW
pJvEMuYuRoCxnFAssS64kBL+K1e6lVGStGtHOWJnQV1FIq7QMeeeOPsumSrXWvtn
6MIinoCGjwcPY6vS2NUzEcQ8GyA/+ge681rGBSBZgByOk7YYqHwtUlavG80mhl/M
tq7znklFbxabfJWxk83t9Czrn8UMCTrMgojhMCHHmJJuSq7Y/VG/YM2Bs7hwOcG1
wyWeq8OAzbjFmnrFY3rg7gYiAGgRQya6uMq3ssSRzS3nAvTFEBu/rzqHqO4RGX1z
usAbOaCx/AYVSiuZvR765hGNDaTI8B2UMeyK1CW01hy5OBMxyrsvbmq7N7NnNtQc
t3Jkws2KdKhpdt5r/oAu1SAGRDOXLeXo57RcFQRpEeNug7kM6wpoQpI2Dt54gCcH
4gsu1kgzteu0oknMcKh58hrx1NNQxv/f1DqGqDrhsYqVyRyIsJzQKND2ZwVQXycJ
qa8qy+iBkgDC586ZTdDoJoYZ63pLi5kCRaLVDe6tlagyXfimsWYP6JeOrJhl+eCK
1I0v7vkcCzyCDfAyJ/ZgmWQlJiH3sfGzuvDBgZdhWiZFEWcZAgl/mVAiDodBqiYX
S43573GWX2wBRRuAJYNNUGM4B7Z7gcNW4ySoBKkJdMjNTCwQTdrgc9J5/YxMfv3j
xfb6KCwWO7HNncOUA3G5iyjhZ8+D38sIdhb/H+s49NJh1BcE5fiouUjDfkokUV9h
lepr3pcGeMCKRgW2fGX4xh8u/ikmunTq3E0hcTbgF/LCqG4B6ZFNPwEU8WVXn+QK
2N9dIyER7c8HZoeJImfy6J1ODFziy3QDSvEN/ijBiu1le70lzysCjTyL5WpdcBuK
NEiCtG7wJS2pdP7uyQ1DJ4FZ6L/DoDtETlx7G0WO+OdJAWjgfxSpeoKmiqSHinOx
NHC5PskB+m7iBaau+L6Jv+6WJ5xuYMVa84xuzzipQ5SJWV15Ktv2ubkBNaR+W4xp
DnbbIWEpTjKUzWfAZGZabDX48YuuuQmCIlOrcvO72qB0VzQ1vZzBjnABXsMLrrFG
AREG/Y6RsDubw1u6u0XbAAPBkbAT1FKWiE03hyaERMnzGrgHyt9qfz9tFHmoBTxj
YYrIpZOvVwKYRjSzjHd+dVSRCeUJJL4eEO/yzUeiYZdbjknKByG/nXft6s0hjWyA
/01KdNcP1z82fJOfXYsR8MXDkaxN8gKFONUYQ2yz6qAts93P86rc5i9NRfa4LvpY
STJ8SF5Iz8a1NvSwAASf3qhMdmLXJxnXOW4+KdHgcqdzeTjbpmrmED6h+oqZhbZK
sQrHLmw9f35ie/jx5+1E5+q4VsxLEYjpWQ2tdRxevfVDRf1KSEGBc4EMG8QSUFO1
4MNe/fZ04/UHRbqL7/Tuv8MuBqz2Qq6kd8Eyjh4W+QYLOfWpkaaNrsg6IZswHGoa
6CywXBSiT3lsp/lAEbWEaFOtL/n95kmFg33+dEXKug47lAMqvN2RalBktu5F94Vc
AD/qfq7PlREZOaSx/2ofBy5/d9k4aSpt6gdp/tmWq7CgVNkL8FeY9MvUyYeM9m1Z
qyFTTqPDFJ1RUjFdqg0VUoWZTkTeVO1d6l/Xs6Yv/85QAMDo8CC8ZIsCTbY7hqJ8
YIVng2ITY/onJY0XlCcwXrCEAdK34FuU0SCDUDgKw7UsxCu7/hzzJ+oHsvysLpx6
VcCyZz7ciLXpie6dCZz9wwjv19NgHNqMSiyn0WrB0Q3rVMFPvKDpKdqL8QWgdkvi
gDnk/royC5Z8aEOUcwRJYb56YwYR4w8O5SndUSiXma65FCYjTHfKk+vVVWUNSs+J
W8bGg15u9+5tyrFjLl89JOodBQr7WFX/SxL6t61b6mS4F7RTgn7N1/3wqgjqOD40
LLvyVrAdTz1kViqNcw10FwxNctnXkKP1xebGptTrOZKr7W+PdBHjqkuXt6+fvXjK
0NrBKiePKmY2PQIIciA/D8upCJvO8zGhAf1xOkKK6CIGok50AYpBUQKrE1iyE+fj
Bal+CEZDpsGifVc0y4BBqhJlbubidNkdRuowLYD+x4p74lECVv7xJa1JmgXuxaH4
+xaSkdtCc6d8kMUGnFYHLTON9hOOkElFf6FbdSOpqMZydV45dH9EmIUj8sA4A8Fj
BTXJ8tuRgr9dxXhFgGWMwfMrY8QOFzAk97x5ruP3c/USVYqOeEY0qC9+TjpxioX7
lo2v4Rf9aTiGwnwoa//aIJHfHIGmpa0DVdsd0Nu+XqmDhoiPXfex2tkDdD+PoOcW
PJfAUKcsqDcG+rEO6gH1x+Nvcp4PelJZ3ECAcuDhITsoaFnK47tuFX4nsZmd17wc
aQSCHuxKL9ZAzWpu6n3V/LTGWyKFlr5Aurc8vnUb6+UhnZ1kCJJWcCW+EyXqz14A
o4dbAZH9XrkpkVvdbLla2RLMqsjQKk9CgNxITnYLTy1ejx55qtMJ60kdupNS2mOg
Z7JgtZjDoLTGgqzn74PgycjVcYw4yWYLcIYbOCJHCnMl+D4U6gRbYpwxtKnQR+Wt
d61dqUaEOOPCv9dWnDj1zaXnUKIatrch3EgX0WU5tvll0P/Q6ndvo6sBnWJnlNLh
A9hwaY+oTDAWRuPsI1sy/uBA0RGu1Nvl2ails5cYkOAOH76vgyikHJHpq7c8l9zo
HoxeUy92qkSPT/wcM5JEGeQCIzCpDJNvXgRklDnjQ6/d8xJEalIrvr3rfJOXMWGi
L4Pcr5bWsa8hjS55EQh+72dHHP+KK4NZnAeev2/Lij0f0XWwFKmsg17e1UxdvBOD
Qz5mp1h7NwmeRRBveyrzUdQIUeYJ3HOAR6aaTOegIF6eQBIgmTbccTdLA7V/Zx1d
1LtiKRZCqFr+09BADjGJ0uGhEY5edM/yM4Tp6LvnrlM7PT4NZ/4HGeHtxZFpGca6
WM+HSJque2amQr/WPptDhwNh89or4kzm7xDv3DLmpXnTyxdniov18Gky2YrCRhGn
MWQO1jdBc1a25NmW0EP7Ib7KO6veB3qxG3tQYxcZxVckrUWh/mhE4gPPtWZZcxiW
XMcUyZuwTepn+54KZCA5H7XtzHt5hoipFFp21T4cP6AKtLNQ0aKHlDdv48Sn39rx
ZchuDJpp3PQ6Fi7Le1qXVt/xvAHXgYDHLdhJbEsdP9PR6MVYt7Ogcptlflm+vu9a
2+xFNpz4VgZUWnYp3nGorqGdzLfOYI65YAbzItkBxS+IJHfPp/Y/zQndkrwTwwzQ
n/OYhKIuFNzgoQXSYtSghCvQOVo23J15OapkU+j5cNRt2az9MCAjDsUO9awo76Ex
yoeXRymdEa7Fkjwz8QGoOlEHZMn0kRgy/tGUN4Sqzp0MCp+69VpnmcevzKAFKmUD
Jl17RCCSjrlfI6zBaE/QxzEqv9oucJK0T2pd5yxQKRNFqfALPJFNIYFWSOLJqTOi
dg8FaM94T0E5SlFX+zcMxpCXiMhPLIh53P5ocK5N6Z+6kJ3pR26axpx1CtHVy6Qi
ThQLVOPGoIRkoZvUr/Sk3Aiv8wsjX+WMVg9bru1/lgvGHji31MfgHvkn4MGa2D9R
C/Cn3sYztMGW5e7nhuvzZLd+mddAKd3y5bh65IunRBfwoEjbdYwavy8mW73m7g6O
wBCaGOk1lmOkMrYvQ/Ayqafh+9yS+czC2ZFa0MwwAWNGptdYOiC7rlnBMm+kaIrn
DmSDT/BbAfFD7yZg/3QqTOLd4cpNCyREC8Kizm57SSjYPbbMbwkFWt1/YSzx7qZi
HLf/sW6/eDgccWxRRcDnjhfZG6ctKXS2tnVY9B4XMr3+hppEhGJkm6ftS3bk317V
oUp1LmfpfFfR4FbhGWjQRQ==
`protect END_PROTECTED
