`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ITt/H6i2lKklIe8pOr/oWUqagF2mUxP8jVGXNF6nKrYqI/kEFGzG6aR+NwYKnGPY
qKrii8uZHXO+ILbDqvp4P0eAO+xTA3sKF+mKilUcwNu5TlHWW87pnHVgqugH7Upa
/h1cs8qhg6hX0SmTfC1u7LdHqq94ZHnwwbydMEh5rSGGzsMIAiwdU2anRWpOKlWy
edM+N7k1aD7E1ZkpfxAyXXDsACQLhfETTdMF5+slLuL+6o/lwQhKfzboW+6Nw5HQ
kuvw6oAn3Ya1GiX09GYvSMqbveW/VU64DiznagF9eRCJ3EUUEWNBy+sx7FZ3KsmW
FO6l5Mgun5i2ZQ8+opgjITtXPXlBAg0JMzkUGaEe7iXFtXSoZYoKy8ezNimCccOx
xgtx5xHckq+38Tf6yZSxigFKskp56Dg85sDnq6HTLzdnMI7S4xGq+NqWbf44TonB
sofIpOmpblqQBTdBrW90Lb2O8X/z3OLJI87XFY4c4d4=
`protect END_PROTECTED
