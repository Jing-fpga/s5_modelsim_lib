`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PYW8fG9B/XCuZIDKQ4ZkO8uM1KkoFapzlwZ8dAiURNjAIFo3rUSeMBXCj73BT/ON
IkVJdtkn7YzDQKxmBcYcmbz7HvU2LkaBzlSvosvlf/EvN33XDvdZ6dFVjtufAD3g
2g0fGYPvQvQVq1v0gQDzbT6E2jCi9OIOpawMQhKhCZE4V73ZDEA2FkkEkJs9JgnW
fL0kOknqLYmQVUzDN6NwjyKbvVSfc2bgu95Rdo8KgRpWtYb5GxlcL6/LLrZ/Ehfg
z+6n7fCYXuvatrkpi/AqlNBe5IrrCWugARSSkEDfUcma+bJdAfvZ5K6Y3EDNDwys
jxUIXTCibMlAxxkE5IMtTJtpGEFB37KEVQDZQyd7IPoWNhiljUa4XL+7kUW3E3DX
X37wa8WyStURxPVnjqONS1EZFzWKRqtPypmiPZqIXngJTv6LoYIWElCg2YSKSuIq
8tosBRkRDY6EUuXfFzmETmfkTV41QPZsdUCVaDBwsNomeJBDEBvBQkqtMFt2gc81
+81v3Kl5iSysNEjRCJHX0hsO6zIR3vLYDppAI2hBtii5EmAMQX2Uu0BeV6q9kvUi
Q42qn7WfUVGrnPONeI5cKI4V96HQIvvBl7L4Zk1GIHH0mDyCtv+mSEySrCPp5Qwo
ahrlQpFy1DMt5Fu1iSJ1FvsjPfR9+sPEuYrLp7dK+dNGbvF5UOuOFm20dx8e4RtI
nlWwe1fnYHk6AOT1+ql5g/tqgL8I15fuEzz3TSaLTWozvrbxSs4sQ0cNoIgszGdS
cW4tPpr+A6DM8+DJ07b8V3NWXtZ4mkiUk5sTd6DrjZCNfy/osWnYA1lTh7HsRWU8
ptlNj6mDqHk1yUBTj8WX0gRaWlN+AkUKSxxZFYgUH6N6U2JYLBbb90dbkjk3IIcX
i0Nlbjf+3x5wPDeYXtAuePSX1I5nkoJlkDMNX2XwdoAzW1eUTk9JZsLx0mk1UJOs
h0iT0/iVib9eXYCdVujHx6mx7mjQ1+d2YpCInY3Yi5eVlyX4UBuxxlvf+2hWIv+2
4rjo/5Jnc0qL/9L/RKtILJhUrmBbZPo5oafs1odyXTT7L4ZB9naPzB5PN1Z4TDvW
EP4EKHIQ0Hyel84Or+mOIiHcFLEU/lObxdAnNHtYDuRVeDF2spYF5AFTl/unoitN
a+zmQ1qwW04OP6QzE8B2YSS9x1AeM8KjZaK+NjZ4GuuEnvIK7exmdyflVrLDReeA
cXxNTLlE0t++/tl/1WV550Kx40qheN/7y7dk9zdZ6TlzJhz6HbBnXFEbS4zEibnf
VQSIZkmgVrR+C1/O3GSzEBEioOFp8kD+IhEaCxnBZiMHsxTF4B4oXGIIj0kG0SXS
YCLU96D/7loJ1DvHFmV5WQQiFJwRSMg/2isxIiZn6RJxnVuZf8KKMTerLK+UcSQj
X7uYks9LSsgyWRZGjP8Kiw==
`protect END_PROTECTED
