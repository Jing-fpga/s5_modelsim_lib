library verilog;
use verilog.vl_types.all;
entity stratixv_dqs_config is
    generic(
        lpm_type        : string  := "stratixv_dqs_config";
        dca_calibration_block_input_select: string  := "0";
        use_pvt_compensation: string  := "false"
    );
    port(
        datain          : in     vl_logic;
        clk             : in     vl_logic;
        ena             : in     vl_logic;
        update          : in     vl_logic;
        dftin           : in     vl_logic_vector(20 downto 0);
        delayctrlin     : in     vl_logic_vector(6 downto 0);
        coremultirankdelayctrlin: in     vl_logic_vector(7 downto 0);
        corerankselectreadin: in     vl_logic;
        rankclkin       : in     vl_logic;
        rankselectread  : in     vl_logic;
        rankselectwrite : in     vl_logic;
        coremultirankdelayctrlout: out    vl_logic_vector(7 downto 0);
        rankselectreadout: out    vl_logic;
        calibrationdone : in     vl_logic;
        postamblepowerdown: out    vl_logic;
        postamblezeropowerdown: out    vl_logic;
        dqsbusoutdelaysetting: out    vl_logic_vector(5 downto 0);
        dqsbusoutdelaysetting2: out    vl_logic_vector(5 downto 0);
        dqsinputphasesetting: out    vl_logic_vector(1 downto 0);
        dqsoutputphasesetting: out    vl_logic_vector(1 downto 0);
        dqoutputphasesetting: out    vl_logic_vector(1 downto 0);
        dutycycledelaysetting: out    vl_logic_vector(3 downto 0);
        resyncinputphasesetting: out    vl_logic_vector(1 downto 0);
        enaoctcycledelaysetting: out    vl_logic_vector(2 downto 0);
        enainputcycledelaysetting: out    vl_logic;
        enaoutputcycledelaysetting: out    vl_logic_vector(2 downto 0);
        dqsenabledelaysetting: out    vl_logic_vector(7 downto 0);
        octdelaysetting1: out    vl_logic_vector(5 downto 0);
        octdelaysetting2: out    vl_logic_vector(5 downto 0);
        enadqsenablephasetransferreg: out    vl_logic;
        enaoctphasetransferreg: out    vl_logic;
        enaoutputphasetransferreg: out    vl_logic;
        enainputphasetransferreg: out    vl_logic;
        enadqscycledelaysetting: out    vl_logic_vector(2 downto 0);
        enadqsphasetransferreg: out    vl_logic;
        resyncinputphaseinvert: out    vl_logic;
        dqoutputphaseinvert: out    vl_logic;
        dqsoutputphaseinvert: out    vl_logic;
        dataout         : out    vl_logic;
        resyncinputzerophaseinvert: out    vl_logic;
        dqs2xoutputphasesetting: out    vl_logic_vector(1 downto 0);
        dqs2xoutputphaseinvert: out    vl_logic;
        ck2xoutputphasesetting: out    vl_logic_vector(1 downto 0);
        ck2xoutputphaseinvert: out    vl_logic;
        dq2xoutputphasesetting: out    vl_logic_vector(1 downto 0);
        dq2xoutputphaseinvert: out    vl_logic;
        postamblephasesetting: out    vl_logic_vector(1 downto 0);
        postamblephaseinvert: out    vl_logic;
        dividerphaseinvert: out    vl_logic;
        addrphasesetting: out    vl_logic_vector(1 downto 0);
        addrphaseinvert : out    vl_logic;
        dqoutputzerophasesetting: out    vl_logic_vector(1 downto 0);
        postamblezerophasesetting: out    vl_logic_vector(1 downto 0);
        dividerioehratephaseinvert: out    vl_logic;
        dqsdisablendelaysetting: out    vl_logic_vector(7 downto 0);
        addrpowerdown   : out    vl_logic;
        dqsoutputpowerdown: out    vl_logic;
        dqoutputpowerdown: out    vl_logic;
        resyncinputpowerdown: out    vl_logic;
        dqs2xoutputpowerdown: out    vl_logic;
        ck2xoutputpowerdown: out    vl_logic;
        dq2xoutputpowerdown: out    vl_logic;
        dftout          : out    vl_logic_vector(6 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of lpm_type : constant is 1;
    attribute mti_svvh_generic_type of dca_calibration_block_input_select : constant is 1;
    attribute mti_svvh_generic_type of use_pvt_compensation : constant is 1;
end stratixv_dqs_config;
