`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RMnUtQIX+g03U1dbhPzfTHQkTb/9OyayHcTDuGv7QcOtz+zz1dYOjaK7EVxnHhPe
mQ7LS2qApEb7ssWBElg1ZpNvUy29yTMw/+nQ2VvO7I3d1ej7IspH4cp6n8N6fkIl
MORYlP4/MJb2dGSm71XjetKF68+qNbrulcqDqp7BFx0D2iiypaLU8KmGIqBIGU2B
E39mE1yQYesvC81vsCTwNxMkUqp1QiwwDSD2fbj3kljhRpjCNNcKEKlaKBiKoiHF
aUBUSgndsCRtswl4rNeCGTBcKKTDU7iY79iajHj7+yREje9CTi20s6qARj+wPzCy
YRBalH7DTrQOVMl+gHSSe0v14iWYmeWmSLBQt7t8ArBpkg1b+pemt6mF6Jw0YUZ6
iIM41EC6A5PFQD1N5YkGqT5nvM35PsPFL436gacMo64mdi5jf4StL3jpiVt3j/LR
vr6rZikZ6+1JqVA8+1rqyaSxm8V8yEoeKtZLRqCWgwpZk3wLp7jdY6SA4eJdTLbW
XKIxzRyrfoLvW8mkI95I6NvNUWA/Iux69yEor+sbMATlQ6qngtouWSpFSft5iL6R
Oy3+yi6hD+lX3TXxRxDyroo0AwChP5EnFXnl1PkSAdWAii9MPgj/sp0sTLPTERhn
SNrAXgjHoz7gppwRKvf+F786bkM2UpIVcye7t05qjBJwjONb8tP7Aqj/7DYAgYYF
dRdszOA+sZHt4u9g7LmgM1ajpksOvxXg6jy2tuunN+pFijEZE5fXjBubWilbf2yh
`protect END_PROTECTED
