`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jRYFIkJ1p32fTCxinKepbTqzdwbn/Z0LTmEws3cvBk4iMBb7GN05PZZnlIlBOAeQ
gsAvcUeWf69fKk31X9cD6o/bfhPSS7rVfejTTuDLc4sH5q3t7f3qrvSb3GRf0wJ/
J4ROwwah6X7c6lU/gnIzYDwYa6T/GUrHE+NFMjLXNCGpd8ltDehE9wM3EGHK1fTv
HtkKuvslJK8EF9mIZnn3bZ8tYrBX/KM/3FoKjY+KnVEmn8zKoxvpvsO5Q2+24rnj
W34iIeNX/4/mx2azYO4NKA8inDCI7WEvdQWZlTpyQkVGAeeuW62cpmCJ8dg6cDxI
9QoIdGG5eaKsyHoHmPh/YL2MMF+kI2YlXnNgGlueoECYJxFnAcoR9IxzNnnWK3je
k4AX2D1zfHT16gHjp99HcdR0Dnu2CQ2R7b74AEvqRVm8ArxUyf5vaRMOIMERJ83k
EJR1cRH78UU44AhkxvjubGNIF8+c2pzidx1zlJv3w/txy53WjOrUJfaJucTfnm4C
JzY5TUEp9m1/jfi71nFCsq1i+FMG/w8SQz9T8cAqde9K2nod7CEvvk5+biztvI/b
sU9QRB+Wl2zpXQCP4O/NDdQ7vEpF+FuewO/9LWS863SwsJ4MPxp3k3Akv/vkMjBR
3b7hn2Wvr91fRp1vVcHDHdZzbHlUb5Nqz0rO+iDyYVUB2yGwORRFOq1m3rqcbUrT
USq5lsV8n0hASEhCrBHkwef3o8QShGuQZf3W13bM6pf/cHuhBsI/Q2Fp0spkYkrg
OgT8jsJuZWY92jOyCPeW2AnHqxHRKBXX3p9S/W2vjQf3zGdmTK7Mefytn6PtRage
9LZ6LUa4jXjjHyGEsJIX7vD8qHSXfsaoaaLXAdirZ2+CRPQEgImSUE50aYSj8gY7
sfcNaqbCnL0fRiq/xoh4RAtG0itu2Kh6Q1jeBkuZGQm84oceAJ0g4zBl1t5rSTWZ
j8ttMBeV3zSaDQVVoL1ZmZ2g1k2KXOIJYEYa4lg/eJn4S2wDI8LGkCGDhwT0Vpwm
SMvLRabM3Wtvyq1EZmGnN2emLNO8/CzKivekP+DqoFxk6vwggCdSDhMPJjo3DUIK
ms+Me9gPecUSHIeRLAqd0aA+/LnSnZzsKSwfcRus6JM4KiUSFAFQhLDbMwyXG+qL
42DUMDFqEt3g30H/tfo07qXz7XDZM/WgIs2dG3Fc6gYppRziXtzJpAL5GfgKfCz5
+Pi5Fi0QSHUXFJqdDHbKcQ8OK0tVjAeRNZtT8kdlAqBMMDqrmQX/yw2yf9OtGVxw
zebxhY2tSPwoNY2RQi4yU6uzj1cr/Vh032HdEu6v/ysZgnV0/HLH/eeK6w7m4rjM
eC8Ui9TsFhCORw8XKaIaTPYPXCUfHZ0uVZrvmdxH23zzHWVY9k5CpKDut6cUzlUC
L/jf3CPSt0JYXIFF5aX8sXuE/0ltLcbhO86v++xVWZmdPAXoufNoGEHPliVHOS1z
wpA05CSL3g3iV50gGc6N1V1cDYBi7vJAZK0GhTyhfRK8nyA+U5atfTU/3qPmeuT4
wQ98sCVZLdh1buhgbuTqUx88JvavghOd+gwMsPSLjWLZZg5kL6gAE9siRwuPDMIk
RDOLGNN5aL/SSEgFwO6Bty0cp9vXppfJpJPiuulgDsniaSxuTXTJfncghdJ1PlYO
cVxyTLabUVnEXjae5LUIsyXFDLliyxBUrlNukS/bUOCOI8t75CwB2vS4PJ94MgjP
2ZhJVJkolF2gUGV5UEwCYrgBRvJWW2AJKNRbaHkC8m2SUF8MHd/0WBUsjRh10IhR
OY+1kCLNkXuKxbpC9j3WwIVsvpnuivzHTbKaTRIg2Ohz+zabhTN7J7+bl4cKn5hN
TPPztnpc1jGcMWLF+QX1D9heCicIr+UFgHf+SvHy2i7RieEsXAUwN+aZ1TJqhsXf
1/5zprw4ti1/gdoB9Mm4mLFYyOMQ85gOIeA44aTh6oHWjcVcmtkGNi6dsAHobbzO
99+L7joTdTKkD3DqJ3bKLtqmfbYj4VKTmEWIvJE6L33TEVp9vono+uQ4/jfc1PLc
8uJ5Mqr7+DvbYFF5FPIwMeLO33yEs0rHVyBYngj12GgDevfEAQNSd9JRO037jPOn
A7XlyG5uHRq9GjpBHymRZCLFdh5lnlRtd4Y4YqY+/tMQEUAB1wqsahOK+7pg76+6
/iRAbfoeVpotr6baqNq+YYrQOT/o+kwk3kxnOQRfX+qcKqN898IPrKP3PytLNaOQ
n3XzrKcczFMsTtV7a0HlIVU8Xt4tS1gSNB1oT0pBTtUQDEK2JH+OOfas4uTVXEcM
+FzjdUSw5IiA6w/p9Khzrjwh4ayC6B+nyLIKGk9pagmtap76s1RkNqwRigB+gbKd
gcXCn9tiUVxQfTU9lkwu78Irve+7oDNp2oMyUUIq7XSQL8VC+yEfre/O1yxmdh3R
xEnDCqoG8i+NcxDGVf1vxSNCpHXGvu4CKAFUBOaLuZXTjr9Hd88GeHRLApSApl1S
ZxPAxHO78gY5JIarSfuX4CxiyObk2AKGCM08MFTRQ/zLm9cPUq3xFy+0cLexSJM2
/0/He3aQMdJbEkrABOFLFr7n2pDZ03xRR3Byj/61dT8v8TxjDv4SKw3X/O2M3SBM
7rhLM+rfMeq0mtg5DZy7lDgEPOw+pKJYb9tjd84VzelElYkC87moSUbs+YEqEbYT
4eNtiykQFGcEJivXswDHQ3MBvsoT5FOFfCGlsltnY0ppOCvaZqIiMvPFIGTQ0vrn
kaliScRaFNPk3uDuyywktEw+s7/m8X144FoH4xTUlA2ovipF0kuky0wA/rRdTSJ6
cRsp1Wo1p9weYhWbuJ8t5FaqNx3iA8+A+l55FNU1RZ3V9jnTu65Gsv+JmHrQB2zj
61msh/LKDjfKAW+GesejcUjgXdp07Fi2TehCVW+rjNyaBFOBen8BdQYsNw2kOrtt
5TEhMRM73IeC/YiV/snAmUxSq5FEq5KBfsIUmFSolP+HShtCX2dlzLcfes2QwQQF
L/wZUnSKfPEgBKCYlyvfZdIvsa5YxhdcZ8WURmRbv59klvhrUKO+3+gfJhC5PQqm
lzhDEoB2zQVLxetIHZurxb7HKHyBZkhCtYuf/8nKU+Qy4WpjXmKLptwOPRMVDoqP
awnNtSq5fZUVSOoJOA4tO6BHl0H17Zsod32WzMiffYy6N4ywwd78QOqtM0fteHWt
pK1mcasSlN3rQN49bhSixYosGjAbuumssJ0RPPZbmz6uaYBBBIVdlxA60u0+dvwi
XJZ+cyg0jE9ZuKf9VKQUaC+B2Wig/Jsrvw4D1VJkhkeqDA+wbmqrDBWCwPkXb8pG
lyKVYe+1Bjc7BayE1Qj7TEtOdb2WWLOrKP3E1Ugjy5Gv8e5+nxbTYelJF04J8Qnz
iW8d2JZ+sdgzIOP10Pr39rPKJ+NEJ9iqJCe+7HV07z0QFmPiYccYYFrAVqyb2A+Z
/FQcYt9voUSoHFv/c9u1wroFLxv/Khco7wsvhmMt0U3Hqa002Vgze0QtkFZlF72K
djfp+hzxhruRKiAk5fdvvGzAdnjTeurH24cugP5rOM92QAm4tTjcjuGOJmDs0FLw
NBtGg6iSijEqSALS0YgajD6IrzVmcBl3PRAaArdK+pvpjevGKf11Phwtv/J/JHBN
VJyjqyyK5mCnkVqMEHDnwTh5dPP1CQDt6Ch7ee34pA53zPtF6mm2uTSIr+TUy+uM
bcKffRm1lr0ds9ftzIJogJpZrvCgELW6hdZA7Zl7idpDw2YtSwItoDdNShwM058C
KBP/uNLRpOwzJSOjVPDfSLTaQ37pwg6guxxWg6aEjPxqPCNhHZeTfv4JqyUyPkvc
AJt5G+oObOrdz+i8/A0ELaQpiF1C/1XG6JjFw1XzHXMGZmpOGQcxg3+gIggYZpEj
qdZulpPJQJyD9hc0oP/1y/mhZkl396Xda9OKui9e4rPAVDfoBZZSelibVnr4LvMV
Ifc3Z/BegviPxApTYq0aIZJPawsp2xDheD+6nG0NJxWpluTucdIo+pulh+4rReVj
bA5iji7hgT2U4Ipe6Xj+BO0XZscqSspsMEk32fddXQF/lEEPg+/PPgeQtRUkPOm4
bRCJaLWdBcWS1UVJzm+v1xCLaaLbSf9oz7x3Y/9HquePYBwQSJ+nknP2wCieFIbe
9QVE75wHfLJkGcZ7+jC21iVPvyb8Dx6el2w7ul8v0sbYIiQBqi2ISfNa7i3r9SEi
1EqzcSyhFNDuLyDnsgJcQ4hY+dFLJDNvDzK2Y/lTqutwEZ1rEgo0J29iLrzGbouO
z/GUUIAVwyT8r9H1UpgYids1V5szhR6gJA3zk+verYpyEJ4m2s3T5wnu97fMjoWv
azA1vCEZHRBksEVS0eavBbTYQni+ZHAa7Bbece2UYvpT8NUmuzWa4rkheiXJE5u0
lkJDklFUVKASoO+fITeXHqRcPM/Ov6rBt+RfkiyL5FqDpvnPj7+Nf47DX2vyHcNw
oZj2xFA8QbEgcRu+6OZVP043Fi5NTixupIEzQL9OF7xbLHyNGJXk68k9mN5WcKVj
8yrfNuw70I2tgMgd42bqkLzviF+eI/D0tJc2BE17LXeIbJmQt5Fs/smB97kM+b5o
9VkN/6+89ZR33CvZua4aVYdI3nWj4II7ckoC6G1ACbZHcTpdBPloSDUWyAi/tto8
eNJfSs+wUiuPakpuNrmWA90RhPuvR01M75P4FwRtHb+Eb3Dx8vb0itQNQCfByPgL
mC1HezO3g+lJYUZSNaIh5A==
`protect END_PROTECTED
