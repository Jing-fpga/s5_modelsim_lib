`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xseqzW87PSpKuYx9IEKeLAVDT2KdpXW5+0VtVGv0rDDDxouHRcy9yB1LbB7mDy5J
KlHYzxD9X5tUh+X3qZ8A2hi6IrL4R4g2sSTCar+acct8Sp+Znv6eYJAmJzpvszT4
h28NT22Z5KjNsSHYoP5TPp0skPZRQWtUk9hLXFE9Vbp8SPhPBvUWP3XAdU7Xh7/G
QiI6B3AxT56G8qqmd4PWbRwFnVMO0oqyQi7NZ4b2Z3Pw35YKdGqGLXuJUryDnjDb
Ziow636UdmMlDAJ62m+pvzLGG4wlzViZOYd7jwdEZFV87pPz06ViQp/NAf/69HFS
7UlgEEdVRdOuw5SoQbp6zGJrEO6sLX9pXQP6NTXuPTG4HxynB/U9O3S8QmWNXPlg
`protect END_PROTECTED
