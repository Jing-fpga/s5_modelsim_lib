`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
75UP8nyjI1PRb0+VHho/bHEdu6+Db2ZPTh1Z3+F5KAvXis43OuYxRgkxskVEsnPI
Si52ZkSA+LjFAJKn08/qI1Q+ibYQBl3rg++arZ1nJfxAW73mNqb0M4ZQ6I/SgnPL
lx5+lO6/qG/fGvdBCrdVPRXOi1UuRBbxD8tjnzFDHQIf9GalHhvn269oed5PalEO
R3Bj8295C0H9XM/oRhvS0lrhGUTils+h6GfRM6f9cibkg0Bfq7KHchT2NaLL1ujT
riEV6AiASP3mEVDjLvhjlSfB1GkPsUeTmxh8MGJhq7IOvHY+1sdG7qb5P9Ypowhw
nsVu+mB1ftwvvOa01r3at7J2fHPZh/Im3pWAbcr3vwZFLnOIh8A5IieeMZtKHaUU
yBj8DeaUF0IQ9/pjpwDf1lFUVu/P8s3Xqte/ZnEbAvekgAp6L2hjWZdBTcuK3rtL
xJqLDhiVPj29cX9DHl8QZoeab+X8cGPFuw1GtQEpWUf+ejtmXheN9/XnkdEiZMXo
dOU5RRM77zyxfGPB3cBm6bUQcZrF5W6Q8Ub7p/RnJky2IM2ubPeVYTWaiT/8MF7I
`protect END_PROTECTED
