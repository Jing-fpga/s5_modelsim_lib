`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q1IyL2tK8FvsZuqAib2i9tjcMb9mLQ2DwWeQk3I0rVxZW/AhxD1A6SKu7pojKUai
aTrX0iEXSM4IQX/IFhQiNLViF/VrFHeFbo0zae0Y0QedqhnJ/hyOyhIp0EZQBALd
Bc10XIJyXLbsJht5/cAAQZRisCfqnBIovzmfe5jceM0gSX7YRK+Rp1hzbIMBLphi
tZWZai+gf4VCmrKKre3bMbWjnBODDsdI7etwAuoUdCCsr8YRePM6GqiSEOHE1FnA
c0nCZcxEiSFstBw6K0GrYBTY2HWK6WWoRAa9Tx12SZe/9J4Y2CDGGh21sAw3XBV+
/HPAFWVnQ7HFj8IUcl8929PdbwalpNOkFe5tBZ/pqjudOcXp5f3i8sQZOpHwN/TI
HZYK48VcsMpEy4u2rEGPCuKl9FdX+PkQg/LI7ehtgpd1e+9wTbwDK9cDSxF8btwk
JCddZdKQbyPEv217DB4UmVysn9ObvJfM+xBJZWhJEn8/PVH4jp+VrlvRcTksJknz
/BTpbt4nJdRtPsAOmhdacxtAmCQYCsBWNx/x+h8E13TvPTU4zYCRXLpU5O8I5LkK
CKdaZV6z4Oh6BX6SO2N0fFeNmE9Wu+8mbdcJ5AVpE4hb6OrYOSJJgH+gGOz5J4yk
/bXosbMs/vvkq0B5fqp45tgd81T5FKnEiyeUBCz5jwctL52CZH+TpPC+D2Ckw+5U
/xMHnUvLCFjB4YtfezK2S3jfcHJHFbAFYt+vRch5DlBKZqrDoD9wVYSd6bTAcdJf
YqYOynJhPhVOHVEILbOm95LvBNzEJBGpa1HXXci2xNRtzUlAUrih/tlx0X/Vm9pF
k5Kkfoos92zk1/Qf/C7Sh9GaCbzInv1TDCExK5Ehje3v3bGF3bRLw4uRObw3/JYP
qUKjPOalIgDEjrnz8xPXyJl2hQ/okWvTM9DdyQF2AvEVVJW3bFHSJThmyVMYu7Dl
bGKTL7FjV8UxikVFKOhL74WnO0h1TGx0RH1rMVOLHIHUbX0xRlmxj8p9EPciMiqJ
swnwYma4gdJjd2td2pY/Qf48z6Nvgm82ROydSccO7Qlm8I/Tm3jMuGS56mfKklWQ
JgsbAjRTIS7sJFKGa0o05GkN3ZwenRNZy+R4+cecFTw=
`protect END_PROTECTED
