`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D9cGg013NPWVi4qzCDfjtqU3VPCJuXanLcQyjRH8EJMDJlPsDRcXMQcyfmNO5YtF
eZ5zmeTvQJ2NZ9JSWNpmwq57nTCZVjBreeBfJCeXDA35UVgeDBiacapkcj0JI+ye
mY6NADY+JKWcFgiHOTtZzTZnxaXy2u6vj+9e0frlfptMIe0iPBl7NL/fX07r5Kc/
FDEhtHK20eGNONwSPJtWJMCVP38A8+fk3ClT1+zRlQeDbRA0Kebn8Sx2BEBG96eB
s9rmtmfvx6HJCUvW7GlY8Nb9IuDFy7ds/lc5foB4lzCY3ChRdRBYA9WWJ5QPann0
wLSkdumbdjyQewgz7zVVGXR/zt9muLr9fEq30IbzGH1KyUd0HAlBKXTztodro1do
owfwXMWhu6/zVr11Mv8aqPXntqyZbq3ftcekvinKOQ73B9xt8hYQcark8B79VxU1
ks2TkN+0rlC0EWlF/bWQILFcj+N7V2tu1v2sWh4LCd7siCzZTPGA5Ms0+LHezHbT
Yh060QPtQQVvnAmQQKaZ0JTWUdIRa+++D3fnBbMMUCarVQixu86dMdxsqzoQkQtV
b7Bv1WAnLwjtS8IMb4M8puD5exoE3iVD/HzVinH414JG4UC4NEzqX7xrXg33MflN
JZNdREwtZ0XUejtnDVPfNU2arbzgF5kHJGeakPSsBkrwQ9qJr8oRPasttmIY0uk8
bTFVhVZNjYcOEYeGhS09QjlDFt9ZgWe58HuAHye8IgeqBvEGPn2+hOsB4b42gzNR
ctqByIelVhy3HGqhzVv+TDBqRusdKtIiaqoMoThSn/6A7OSlTLhtSgDBafRBSfdk
c+C7r2POBze9mH+dz25HAZcgZ7k+icsqLBf8pOkR+KmZ4rlWNEajL8NuaBUI8c1m
cNzIMWPUPPkSHlwy/TPeRv8VjV4KHPdCG9+ZE87A50/XdkaWyVNDGySNqp/WjYsG
ezF/O8yMLn+kknTiKVjfGTKuITnV6z8iMWDkfW7quar3kIBhecTF3LNAt8Im0vnT
kIrVUF+nvXgfxCHamo0Qk9dJMcVqPmdrcsFi8CxDoswUK4xy/WhTPai+47k7qiKh
XbPwjQ47ZJaGsD2QiYJHDJiqbSr7ZFkec7qXCZBSmR2NMXUdxD5hBf4zi+7sVauS
GRJj3CBVeYoFPIi0IznQ4EhCwsd5WL2GIhandAbUQH8/yQzhNEyxMz22eiXNhcRn
Lbd4lsaS8vOTmsye34uT++u8wQ5ndbtI6nQrbNMwKC8/Ezom1DEh8k8iecKIG0J/
Wk83WSIKOb54JDzRaBwt0GGJYjIdm+kq2tZx/Juxg+xtD2/Dypd5YW+bMg8bYlpy
7Y3dRnfuqxymz6e/5IYM4PDTlBHtHnjiyO3rEvR2MpmkbFs5juRlLUOEYCaAwADC
GHs1DJ28U89w5I19T3tCxIodas1ZVgZ2J1kCqv5qv+NdQSD0fkDLdZZo+9YExSnw
++dV8/ChL3DNZ1gRqMDoGTuLyqXpXYsmf5Yd6y8M0wsKHUa8HsCsyO226OnV7lfU
iR9zcuYJMv8lKX39iGe96rK0u747qOHTaRuc7+zwX83qwa6TypCu7S3OWGrpXqkl
3nIrucsCCqGevWuIu8zOmAL1giEjRUg6wuDp7VknD8LI+dTjiUZoQAKW/w2y+yvp
5cvlXOB8QZ083GM0vPb/SshRHR2AcQwblz35QZZI7nX9mCeeuvy9X0XUtrmpAgcb
AVCb0Cu338gCfYmTth+GSQn4k69RWQNuHLyCzRQ3uBEZCjMHWacFC3UGyKdhSbHq
BfPGrKKOWJ2ptzMQ0cSj8A3HrrZ4v3CgOzws/qcY70fPfa1QF+/CPkfR4eyUt49Z
UPbxwJbCtdky7xQvrP9uQKu0G1duUHt27QScGVVgs/Z2Nnt+xggT73RUnmGNKZcM
7JjlJGqDhyKFUKdj7GU1dOh4PpH1a27fT1Md4azXg73giSd8biP2AhIExKomxp6l
z7X+4M0luAyI+b1Vi6hGDT9RPfOKE2dYD+lKW9RKumMgokhz2ZounvoHvtknxZxg
qwNDLbgao7sGzYJpJ4D3BI2Ap5FFHbiBO3+J4mHWc41wMMjgtbBdVPaNlmSo3/q/
aP6mJhVnnVe0CWYdk9YifPfWiErb0KFyNiixMoGeRI113gSFBC1Qydp9470Izxlf
GHXSNBQH9U1fSH0OpVb+X3S9bf+Z1dti626apMKpzvjt3+rOzaYMRukiio/kBBZ1
EfWhiAposoBIo+WTSX2O37v0KCj5lxrqqP1qxP7TM7XI4Bw7PncztaLQ4BWTOk8p
`protect END_PROTECTED
