`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
141+ovgU41rKfVKa7wXbknmEMkOtFFSFMgdNImwx8NuEl8mfGXpEoA5RIekKxDRK
0no6fwF2qA3QsT4SZlE1MRXVSrq2MKm3ZkT2Sp0ApSBVRUxpUDuQqiw1ERuzcFIt
WA1BmNTcw+UpUCKT61dOjzzjBjoHb26KPhw1L08Q0q+XjS7T5eRNszm/qTtFjz6s
oIchyxPgn67EdUq/fjicNm334QagrmcLOmvsnUVkR3syNEMSJQ+OjPD9I5otEmha
/GXfa8GiXqK4o+62sKn7P08wGwWfEJUnGvKE6+XTOUNAkMbactk2ww5H9B7H4rwT
6chPi8qyeyDyry87ZkMAHY0N1igYIN5oiIoJnIzRz2HhwPW0UpsOqVzThSu9SorP
aI86EJZA74VJYxlw0bxX3tR5ptO/9QmPuMfhf+w2qxFpAHbh9Ag0SlnYrpzHzudx
ZeXFgbzlTALEDBR5CqOHyaIZiZ+J2QEbKhfMSYHaZGsEuhvy49cOHQOIbS8uona9
3PoFhVSg2N2PuEwZaCrQQbE5gnZHjaw1FdvwqDxFZsoh8onuh5jaMdbg4Kf6IdVS
omgh+pro56r3KqCjcGi8ev2rYyYfFLKfq/cS/7yClnmaJbotjnMSIsf6e9MWxw64
F2MlUHddmWzQ5KD5oMYe0e+yOAXjBUlsORvEbhKHHQ2XkK6ninnsbze3hx9VNo+K
xH9UnvQ3N3aAXQ0rfCWaAYct4YeWFVymerY1MfBsPRs7wzz1ZHNm0Xql/8GXPX8M
oBmyRLE0Oejiac0P0p/TCW8VcRxSIXDKs3CrNSJFUonrQ3laV+g0kPj+2T+qhS4G
JwLiDsdbe06TV0vBgGqofMTI0qASN0GrrU9nCtxI8KtOcTJDfQO/ynzD1aRXZg7+
F2WOVJ/j7+ErXDvgaXfFN+LN7AgJZnyuKTgFDvDtgdMKnwjVtKYym9y1hB2SfoIf
mftlL3HPGQjDdsErzEEn8w1hq1sWPlmsH14QFHoIzcYLfWueSuLlZrQh71FS8EKr
51aP+JGD/q0EHYNximyz1F5G74Ix/KPvcPDRZMv7DnlWG5VPr7cI+YnMsDBi5oUO
hnzCkC5RGhpzGWWPKC5YHcKkdVhYNfmR8MVMpLNY57Wgw6T6XAESMBMgEIzj61uN
YKAULqmqv4/JrLuFurHgtBDKJFN9ZQIr2+6BtKzw898oN2IlcLuBiotWnglKXaLZ
VhKPefrgvTdU7oAyHCWp48uD9kodkColepWCZlBiktDr4STX876tKCBRhh/DfFoC
VvMEU3R2Ah4nPkB/Gn3Sr74l+4+shJ5g4KDQR95wT7/GJNjwk74VarqpYVZtyed4
UD+9HwuV88DPesQAmTeKs7D7cRgtavvPQdbdyb0tZpq2q4V/cuDwYBYGti9zLQl6
YGWtPpoNbLpgfw9ZQOyfj2Np9D/yX3RzEK6ZMgieXlLG5bFNgRxzvvP0XTsS5HiS
M9pVftQC2cotXACgciUdePcNsbOJAdrnC5YxQqRxX8aVwbNPlCqorYSJ/Y+Ky5Iy
+1M8IrXwXf2HzCxRcNd1PyFM9+u9ncZ4J1J1oldWjJUlgXeoINgrkYa/iYUPsE+z
6Zi4i5HWfqyOCYO6LmYvn5c1cassQa1N1ONLtK1iIMPiJW3afSeO6EeIhN8vrnAZ
jfxw3ph4ypzNtew4QZTAD5VMQLQTzc3CsO8saDZJrDbkMOKAccoiwqrgXHVp1J9h
qiNr0clrXz2nUkIG1e0kBFJ/Ps6tU60YXaBn9WS6L5Sb68qQIt4cDDgIRuGPbXTy
2PGJdLy8ZjVUu/6RLAQ39EpsH9MnmAdfKZCJgWumUeDGHpG9++jcDSLoeAMLsuc4
CvR8L25HwGBpFoB8KfahTnmf8ZDfX7MvPV/mMTfqhVFyI5Ib++awUtd0drzdnhu0
y9bkvgmmQIn3eW71M3LhU2OIcVSNORdSIBjjkLHHezwjSN5dMOR1ARxQthjNgf2U
7eAn3Uxap2GPYsRJb7oxCR/ubt2JiihBxj608DYv6uk5XGRcBeskfKmOdrUwaAQz
GiCCHrfkiDmtsY/8GgYWQynCP8Uu2e7UKCcqNvaysWI0JJnxkNukjda4JKVcZC9i
uN8qX7MrYyGaFTu3KuBv7e3dHmwkrpQ+wX28pcwDil7jYBJGIdUCv1RXqn0mjB25
da+wOAZ6JpB17yqDgGQo7GSDDPG3LhqElESrT+o1QdYt+ifgDqFZQk15eQWdfC28
jIzc8X9tBCeD6mCw79Jdmarc/Nr3WScD/+FIq3THN/npLgKcQzLfmTPWtEFMSo5R
S3DdpPT5kRumwMtNLGU3mFHBvD4rCU2eGbUUarqs5L4szVm7oUv7hETQyNoyTBLm
Me5nqcXCvWuLzn4VqN881bsMIlyQGnWnTp1QnbT14dLdkZeBoxLBRUDg0a3b6dFa
9x58AI8+E4GYeox6W9rC8o1FhnL08choJu87jo7BpKxHrzd6ZBbk86U1HmRSv09D
zRIoE86uOfsK5C7PI0TMHwl/UPaZYmcHLkHAZck5Tv3o/5a4mbLa1VzLmoe4C+GS
DFBcJn4pwzXY2GZTyYVYj2ksZz4123YONOjcWpr3W25i07RlE9lV4lGHywuSkmQW
jQqfATX7yToNqt9w0OKrsWUkBKrixAyi0v2E6l5SZRkpMlEgyu9SUTAcZqUsePLs
nCjXtsD0wZPxeCPYALVrNpWoap3K5jFgoP790sBMfRlQ230e/Faypj11PTuORtaH
tJPblsxuRuKx42ra1KfdaHrTmiNwhQXlflWPxVP9clf4VgcJzq5VBK1D405fEiEz
ahwV7JoCOfPxU8x1ktNaOerZbj7lzsG2c0YafnLZpkLDHVAJ3LwalbFYzmtbncNz
uMqYK58c4u1H15lAhCb/TpSzag8LRgci83Tjek1ZNf4IwJ/HPv37fY9yodnlUpMz
7KYXEAtZjxaHoFpwZGCmzL0NyNgg5S6PXo/xGhZar160bRkgE5XkGnqdjRTaSbvq
Y6eGZsydjHSzwhfmdrl41E+FsazCFoe3t+mbdYeJUAhUdkMe1MRWTOinrXtEzjsp
vRJamF3LBYLI3tM/nDjPPjPsJ028nNIGYZG/xBxUdvOP0tQIzXWuO1v3maikvymq
vX27Z0K5t3VGcOJdkzfSbKzTakk/u0tOEBdEAR22kghc3QGq6tPI0wbfgDeFqx9j
0q74ELW0fuyxqrV4ydOlhy8IaIWE67pW9VnSFbyaoLOGR3Oq6wZPc4eE7hu69uvq
2WjUvLxtGVCJDBCjJaMVMuG+Ig0ohrwm9seUqX7oGowRIwB4dwz1zd4QwynDiDeb
GwTo5UTAfjk3md7TAopvSIwz57XYgxzr3PBmtVOLVCq2tuwyG5vd8d7EB9MXWq3c
l8Bkfm4AGm4wDWuOkEX47hcJA9RlM3NL1R/l2zb/jlx7qaw/z13rfHkByRuu/Z9V
5+AyodvywYRH0e5bou4lN3tz9fEe4JLD8mas8Pha06xDD7mZAF6uisbyFCXsaPtH
nnqSqhVohEdg5Z/EWQ9IdpaeuMnUhKuz6lGMAsBOYj0+YpX/BlZeCW0q4+SW6WME
WEUN+qurMybmWtAxC/44XaynTZWHZH7dJZ8GaLkBaEa0MsUT1yaO7DNkTGG7b5OC
AZYqA+juiqUyTItKk3Snh0ajSxa1V419wSJwDIBdjhLi4gbxU/cqDZNb7ofsdLV+
E0ngh7OU3JZZ+VeV7xF7FoQUx/DCEq/GdjadZQ0lIEgGCCMYfXU0uIOZCvZXxLmc
eFDrjXQscPkZUY103bw65Aa2rgIQgCravOjN6IpiloEZ40eDvwVTusXHsBSZ2GQ6
GE28FL9FXZiypFNK9JdcoOnPZxqhoxllm3gh68bnVcxPSm/X9QaxT80hs4FjzLSg
MqOB96tOsPC/EAegMAOvG9mdRgN4Mt0UM4h2BRIj+AKrSB46+zzmT4LX9xE6FWS/
Z31ag54S4kdAwux6/RRNvA2cNYkSYIGc3uf4KpvAKQk7M5xi6Pngp+DdNPPqJ30y
V3qz62PR0gh9nMB9WdYiIWzB+h93i2JlpFh0Q4LkYKbe5yBX4+Ka0SyyDPFey/u4
RU9FV2ar+QiSALyfo08tfvQw25pScFfDuLmdtK6beYl7+32QNxlvk8QWALirgFrB
xlIJgSU/kh2i6eDRuzInmiYrZkdaJjjHba3QAi6JYetlSqlb6VXwXbvLQK+RVxt3
/6xaIxR7Vk910cvzSlxjY3QhSz4w3yr+//qNllI8l/ghr+ISzn9cP1pL+SRhwvjS
wBl38eZ3nlHK9O59FNTGD6tdfVN6tYwqB5ntxpNANwxwiBqZNE9yg1sdSNF3Rlmw
tdYwgWKsIpCFKJ8jtvPqP1uSMp3EPx4CuTOhzvEym5C+Y6DA1ms3bIRar9RvSaag
6pmzgojqNVMw0SKGZE8TOSNWhKrK0hn/NZBz9HgxlVU5ctptyz30ZuxvWMx9pQAa
epyHBguYANgGOTVY+9z9WVQzzuUTbNclM3/O9Nln3ZA5lcyH/ZY1Sj/ZFM2BOVNX
EqLpTktbvyQOdtbYmCGOGTjxwkyr6XffC7p5FYKJ7RyQI5NZeafw2J1mWLAKUt6X
JcVaTTyMKLg50tVOTcd8q6sok9gMNcwq/eizD67+2oq+7kWwQQ5YHdYSI/npO0ta
qWveYxKQYMUkhzDDIGdYjnpaypTP4fPiadPxKuoZ5dfusLp6QmjhEpEZmajBSrUY
0iEoB230WP4OWslrKWw+OyNiyySYK/BEQSRCKMf3UA2dRZt5AjgLGAsqX+v/n58t
i16d17i/TnuV7CZFrCsOB+AjQuqYeBumYNdTnV4IhceLi4oBS4wK2Hei+HUPLDNp
HjuQ3FbXzk9aWe/mrhndjjOUOlOjZ41iLaioUHo0vYX5+hXJGrKlQE/5b/utfRpl
Asuzm1B16Yccckkpp7B9QKIN2TTSBU+6uYDSswBKhnlxo24MGAkMUZxR03zH7mxu
X49FoMBMFn63SzPWOav+oVP5aDQuDQJ8wvlm+45zkFdxlWfvqGRJFMCaHtOPfgjm
xyttnRd8yRefTJ9JxE54av7PWLM2heRqgDGcOcbFsA5SC7Fpes84J8xbf+Ngby5N
TMvRq/v06m+BP9LpAvcmE27RJJGl6pYB66Ah8zrSNq7Zfmk3+rxqwJiORHEOvLFc
4jFRnxtISF7d0hyS7oXup4T2CzWpE3yu+cSqJpbZGKCwalH79l2RerxLANsQNYdy
VdYHkqkxSPQdLSTO73jmt1Fo7+mxxywgjAJRfTcvSeVuI5ONGtq0Lnse6BuTj6z4
cL6+dnuywsV1B/rDnciTddChd5bFyOqfTUspXl98B2SvYGI/C5RKB2lqKtJjxapb
CSohVD9Ik8VEswlMNCFU7BQ9u6ByTLljXFEAwF344ORAYNLiv0NZ+gIwlIkEV+lh
o1URv4cAS8TJRPJbGU4xBzK1qBAXNbFYQbc8gB6hNDtb7jIdiMb11WHjscsA3BHd
1n0p88LU+4KLwyOMOcDIQonvGTSmlDmomIWbohc0QJ3k6Zmanwb1lEGQtAEkhWNt
leYK01TAG8IhSV6xWGBCTI20R0OQNYORRWlbylHVnvJsKqeBCrIXue5xoZ75aiWq
7rTOCEXqumcaaKUxVKLKue6CRUT+MY8AdxmWn8sfjfe2LUI5w8/c+KxJlDLkOWYs
csm+Ak8K19H+tGL2NmRHVccsfVoxJOSXU36ITDgV0e8gElrSvGsh8fGRfSpGb/qe
IR2e/gYREghTckNYj0HM7vaMr6Fh3TbryO2cfMxdB8kRPRFktFu3SL4RpwKSYXbM
cgyEdfHJP3iki5htHGb5QY/39zUcu0bdAwr2HKPA0ErUgykQ4aIii7bg3rGjtezN
h7ykqMPsruHr0bgvcefQvjOKKx1c7YxBnjt2Q+DZ1b/fm6tEnvPULzhFuCsG8xFk
Yjh/47k2lxBUVeEOzSvBVxAT0bHT4Wzucndvp4QZ2k1mJ8MTb6YG1FEPR/cxMoQ2
CFK4YGtgWmYkSmsKP640dwrYG5GhMRJToDZb/jxvzSErUCyipCDZzU5MZEbOBJNT
Q9P7vu9kJ+liOX41DiDkkcgUAZdYTCkVCWhNELrdQRtbdBtuErih6Wp3GfUN+w1l
lqKvazaF2e0+GM1PhjiyCJekImJptgiUrhwL1wFLiMVKEr6i6dZ1p9vw2J5g9oWf
j5Q/wyl7Eb4bWEfRVACaxvfrTSuZ7M4gXNCdICoBgpMfEwv9TXb1yc6HTp21PKt7
leUWr8PvePWNf0IMunPRpl4Bc5JzwN4im48yBAAbN/4mX7dLPZ858yLHqJkhvnrb
sUBHTpUsArT7SyLTqIOcD6+7onUQ3UTUJHgJ7DViQoYF/BZO88isdtkaqg93rweQ
V0YAFtqMCH+o3UmsLV0WDBb8dyklNkKGPIrGcqhq+v6P53mmhs8s+ocEsiNQ9b7v
WwU/y2b877g6yBPueh607CqU3WGnFw3H1tlk8PH+NEKjDD1fJwPZEj6ptk497NhH
26tIQYa0hJw8Qx/MCv5ZmhpW2VIJW/8Z72uaOuGLDmIeD6zjBj/EdohLCM/lKCKy
J01Bz0HL+baMNPggkpLTeJxrvizsgKokvJfYM6qNWF2Tb/DUMtgvz926yzBcfc1B
1wnfgAQpvBVSiLcZcwX7blMYhfbk51hk87BV34iP00X5zPGW7Bq1ENVOMsu84c0T
E77+mpeoDMlXEZ/sz7Ncvvu8ku7yNPnw7Z27NayYwd4E8nZEkRVrwBkPuru1q2FI
nrUkvtmde1WOvv+sEWAP98dAmNPQx3/GD3lKOR8ZTEHOrm5XJI5F3hBxapj2ff+o
9UJbZanZ074QWMDh/jdeV2cdvmErPaL6xvNCIpelzs9+uTxfLuQrP5bhUR6qluPy
dfwWB1sPtvbxlv0xi7iI/6/w1SZHc3oKz7VtyWq7Zy78qMZgd+gfPqpX5OnSXjL1
sYu6V/3zpG5Qm4GRjf9iCJFJXOSBSOHuMtYAI+GSSt3G66bXQ+VPAMzPDgyH9kc6
gX/fclUdG5gieZVOhchMqcZfSkcYvNXeNTRolPFBrvfJfX0K5lTJV2/x2q0ZUQOA
0M//uqY9RD0IgMo4Nr7gWo/4emUJiXRCTSXTuQzywbw9M0njpRKgFyq1sFLAIdm6
LXgnctCyaFM8R9QzsFpub1Yc9jtB+ZrliN2psrjNK3IQWGe0Qn4fg8lfArnFvTF3
02h6uyJd+0P3NH0rpzZR+QhmLy+3awYmorAJt5RR2UoMzLH3iGLKLQvfsjyDYlXp
pCCB6IKBNpQ/VZiLN7f5T4nFA2ydWUoob8LDpdnv3GLfDCZaw9tcC2fVMCZzkUTJ
as+61dsJr4BoNWxXTsZ4CKTq5Impg3vy1uV/xPm0tLJ6t+cug0zjGLciVo0tznMq
bKjUP1k9tS8i418y6q4H1OlcX6ulEQCopCXPNuv8rFQzp8z6LqesZbvCGTpf3OPy
CN2Pbgv/BxvAPPsjOotMnsqpNGe2ItuOY7bR4vEhzptIKsG5Q2NtuhcPTbT9G+p1
mAD1fd6AIVQiFxNBtE2J9kNJfnja4tXx/bIThe2vOb8wgH2ANz9j3QhcNh/wD+fu
njrIXH/UxQPzKVGTj10dpyLIbqk4P5O68DzeUoDLMjOzhFYJFTGHDQycviBZJKgS
PPS/CNwQ+f5pFI3i89pYMzQCYa6J8j8Sb9wFPyYc7zpMeRRlwTvviZ0njH5pjMbu
eD48Dg7c+eZ6HXwnioJjsfCo50Gjo7cEQ0U3DzpoTOeSmc3RxuJjO7jz39C4zlr+
ABE+QEdivFTE35PsMLxXRMtf8UHXdhdeFf0mPMfKJFZ7/LspWVaTxPL+Jf3p8aA4
cFwaWAFdJxGjgHy1V8UwqgpkolAS9O6ss6jDDYiJwTal+Zag2z5/vqGje5RVR8sj
y4ucVDymfzjNIea2zkn+oM6/wbKOQhHIc4EQypy01PZz42EozAAQW9EOOoVmh5Sh
VnNJ2xYvQ58awjPa0g6vIljaaK2VpXey3+Oyu/uVJ2qyiqKgIFDS9D7Qg+RwgyQ2
lWt0Mahsa5UTM75scekVyTVAUJUnaUbYlsok90tXH3Da89FnoKolRqT+4U73RVii
FpU3UHh/woTVoaHLmde9pdHsPUetuxBQ+YoB1pGAM5/BGVgCapm67F1zI75Xw0Lg
/7NnaLrITbhNO0lMNBOtY6dOCZY8GFn3hG6TL+hUxw38LJiWS6pwzy9spheLxSQZ
IwQTZfNhni8XPGXB3Yfnpl1xMJw06s4S3wxyyuXeZHBEH5am/jZDXELZfeMTLhwR
d/10+RnnL/TYp7tsVWfMoUdEOEQ7FqlbLY8Vp0y/CUSYREexX92W92nqqYjy8YFU
i+0egNAsGpz1Z3QcBCzroynI55hXVqK0p/aPpJrLbG2EMSD/nC0l92mu+JY8cHNE
zTiUXwKgejESU28vtfwN3WN/UOJ+XsxMARfTL0wuZMLAuOIgnr0aYjsXtk9xz4DC
Yw37+IzxBopQ5ryuztD03OCzGJk2KiJP/LeWHof/NyWzrJYs5IK5W8/wWBExE7w3
bieq3bbyU38hdWAbtALID/sHJidoEQxGGF6DTFr8xTSVtp/aYbeyaz5jErv3HEVU
cba4W0elaEWbz6pooGlIrhki6HP1HAOAJ/LRwgsZudCt4ziJY/mCmpHau4926Q2Z
tXfyAm2qLQv33D8aho0IJjAqFLviXgn6/j+HIoohcRawHBZSim4UNh1tjQn0IDq9
q7Zg14oIHY6TKFvho5uVA2AqzGTN5m7vfQOjv9rSr41UdMTt6gpAFqqTwEXev9Zf
33fp4RbNCXAfkpfgE8Ax8xs//2lgLpzXXpfsoIHbBKWqw1iN9nNk/TUFIe4va4ib
j0lw875l2gq3XY/ymOmbTX68fpYTmli7LL0vsf8yzCTWinEgXZIMRDOenWHO89eT
hcGuH4G5hq1ifDmvOEG26COqYLFn0lW3scgFmYcIld8Tl2DzmoBbMqvlX5uVMwN5
MZT6ATB5uw/dd1db3HR5OUB11cP4SBh/YqDHWqOnFaoIWCQAhYOsU2KdEkv7x4+q
onR8v4F/cQtCgHL43yytPvvDjxtabJ/VAz83ZJClNh+hu4oyAL3zghjfNYFIg4Li
qBEDnaTzH8GsRflXXnKHhp1azMQGmFR3n1WNADfWRPmwq08JfDafTWwcjF9tcK4z
4AbeXxn7kMshGT3LJr8dhxI9vVUynODDGoWSYmG+4mN9aN/Gw3wwkWYAcjmvuViW
jsd8Kib1K1rHfBSVx9DO7i1tqldpbB5lsLdJGhrI8A9B1Y/9XLInTZGv1XSqlDeM
NmWbReL4SoYF4VwgUqyYa+afJjenjmh2XA9zGjfCO68LMDUBrocfs5lt865CUxHa
F/F1Py0nz68iklJRs3dwFlFnnPVpr6ARjrZQvbsGrGl6oxQCg8w6der0BsO1eDWo
aWBA9BTITLzbon9XeuXo5JhF5frrRJYeEDnIySK8aSXcW+zhw/OjVm5PbWrp8i8R
Nw7MRjB+rEE0ivRbUkiaQ3IPfpJOBe459Y7G295er4pQXJTRmx+uBDzlasbwGA54
Qwbu23vEKIeQ+a3Uj89bxe/rdfNtYwAjVniwr6gzHnvFgumGsH2woMDDGpDg9b7C
ns9lKsBjiR8IO2mY9fUzYlXD459YbFPhCKnidlVbJSxkhXal7xHkgD4c/9523xOq
sF6sKwnJT7qR3onmgSXEmAXk1S2gpVN+YTRV9voWApo7y3H8RA6J3ugm5MEBBUC8
HXldoOay9vWsiPIxK1UH+gypkop/1q80ui/n+HeY0APjsWwCeny7xE3IN9a8nQgO
aZVDmzESXxnucOBcRPYeq1rIH9JCU2WMMtXMLNte0t4+yDJblAi+FPcsMDlzwlur
2N5qwQnW3SM5spTaoKymOpqlZ5LCe84s3SzBpxSBf7MIFswrq/DXDzdJpqdajGcB
kS6qjGnAd5Uv+PUVnNxJDJkALxoIH9pCT3HP23Zi4QxO2J7n9Ih+XEvXXypnLbZA
4sHMZTcTXPFY0hJmiy4+1TFKz+v7fIEYDsb740Mz5LxbWeM4PrdYip5dGnJCihnZ
/aCxJF4SEaVFqAalkMXIO2ouNlB9YgzRONZQiCCrFJuL2R8kvssBIXreVdtWrdv6
5JpPJqOkUnxsiuwR2JsDt+QNI/Tu76LHSzSaxWyeIWmOFYGsQ9E2dAIdX1RjYDIj
RBcyvwFPk7CmABWJsIVJhPMsmi1iJ73p1d9SW/iidqNDBmDLIRmY3gUru5gi0TEJ
eE9zujjFtzkIdxxoC6NoxkOUU1sxLGRDDVh6WqFOgAlRODKEO6A1WWllLvIIkMCi
w3Q937/3WV21PkbKPQ7bZOanKyf2hRwxHYTZ8POXIlyE65qXwHEB/vZKryXZ7WrB
YioIkg+5uyKj4tVgIPqCxNhOPKM1hLGvqQb627Ypruvg1/+tRsrAgwSQerdqBK35
7ZgorCmHPhbAGXM9VpCrOXFMGYuQvrkxBu9ErFGCzBE6Ea/OGYxzxYpREMDhdfH7
G+KoETX5/rMiigJ/sNVcdzoh5+xQET+hdSeR46Ntzt+RMvd/qUeTc5VYmK1Y63FI
xRhVQBG+pFXj4tPToCpHzi1QHhDgHUNej0IiHzWMhJZ66yh2QnjQRrbI6iL6jGtS
KjTAqE69ap4HEPCF4Gi5fOn0EJhR1xZU85SaGdjnzo52a5pP7X1hXiNbKjKHu4gJ
2uk3axGhw8W89AOtPYbi40J+SI7yPnQeKTbUDprWboYNq52DHM5LxqifAtfbDcQ1
4qv4e+S+cLerCEDjf/XS9TRghTu9VlN35wIWXPSxW2zl83JXXztE60tL7tzTqmIx
hvvg6f9ws3JExAUJtWyulgKjB14odZ2aFixvg/16/3j6f+pWhLCEDRI7MEuYClCd
w69s/ysAaF4dKrdlXFYJg7oS+OnA85gzscbIj5awV4RGnnDuEs5guEg3gwUE2VUq
4bHQ/9XEbUOpy6ipGKhWHwjMFlfzoW+/m+8lOZYzDqxjwI2Q3PoRn8516a02JNUA
8v31WjZZy4Zf2r29pR9wX62egxaABFNBAaW/NA0xYAtD/kyBIcDjoKfDqcu2elYp
7GT2vz8he+BHOQCcF27hVJQMelFkgDTeQ3mkwWJq9jiElnZ6h5b5LC5p9PboEGp0
hmQQ3tCz8aqHzwyuzsf9vS6hgGAhhYcsVWsVinr+ulFV14nEg0O9/WaqxcLXzKE7
5R1QHEiEd1iTuXLG9YNQAAutxH0brqLep2nA/Q7Q/7YABvqnq8OBraWBc5KN9m2G
ezMz20OmwnA52f9qKINKEjvbHSRzEkQ24CKFXSsFieBbwD3xK5+u3dvZusGIBGMO
6TLn4hw8cF14MYWE0NtjLvz8ywf/ZRVy/CSugxeALQS6ZI34YuMRENOv7KH4uZqA
2w3NWMSUR5cBf0ElGbYDRiZdbm1SbVKKWm86ui3vwCX0kYL0k/hvTkoYDoQD57Ok
SO/mjOh80h3DPT3RH50s0zMNAkxT1D6W/r1zbHpdxVfcqFYVD7e1FlloCQ86CXFr
pjMeJuqidwouM79pqfLnN6o0y+7aKcdA5yjsaLstyIlsFHvCT1KWBidm/NJbnZ4p
FO9XAUdPr01f60gQoaPE1SfFzXlXwKR65z4Bu1l8FNcUCrUne0UR3m1DbL/Uz3Jm
+DqjhHD57jO5O6RT4MDrBEgR0CHy5PWK2TP+/m7r6sZzIxVgZ/IeErFt8i6JMoGx
QGbOFjtxHiKs2hpFrrNzs8f2jqbPkKYAX5qYByD1vRPqUInPkuReM64qxo7OCwt/
jMoGq60jyvGcBYGSbNiD2dDTg3BtADIJHPEydecCvw0dNoI5MzcmFNEl1RvvnIqe
hF+0fkXqTQYIb9fHwA323+tp+hK8wqJMA9ksWPWOz94cB12+4BIMt4RJewsFo9jI
VwmfyerRrQaBQHXc7K6lhrAtAVDif8LgcJA3LZNs8ztHZkUuqraIdl+pYiZ/OK6G
jyF6iCi6X6ecDKigg9DvLkkz+tgTn51W2o8RZgIY5qcBo0krVYlFKURD/Ems3NLr
vRanGYw75fy2vtppsQBEN5JaJugrKbIAfWIjItHBrDyew7x71EEpftVsuH2nGxct
TpFCAFupLjESUIKiw8xoKzBnQkKcVAmWu64QMAd4bElGq063IAeFAr1HQ5JTy8By
ovPLRrZHZe0Dv6qmbORV4fS1VFtGFEuWNOgoJhbwrSoIr3fGKbcGah/MkBZeZ+w9
Aljebta/CnNbxktWjda5Uk857hGNr3DSXGerZNkrqqGls1LjhLxKaeYnl7EBvAkT
hAjzDW9oyHDhALU3AJ8m0tOs3zdFcwerVMXfNHVTKHxKMQFWlYc5QiSEj7J19uNE
NcmZrrUMyfVjVdocLN88mQvNW9a6VQ5rWkNlFkS1nVLPtjPRbNT6W1dCCydRpPDX
HeV4RBkLTWKkFJEdU86Q6jRvirFRJ/kGV+ohREkAXZh07cXZbzWjX9C8Y+8JlHLn
9IQmO3HSpIyguwooA9f6bYebX638Z1EGSSBTme4B68qZQyQwpkNnVAOxGyLqKlm0
qJ6zh39EgAwxHyOq9Le+HewiW8nGNIkY3DPG40HrNqgCIktzHv6DTCGqCwxcnpF1
CqAq3NKEIy5u3h8run0jT3H9BGY/ZFfiBnOYtTo9AP15QGKbZP/YCWODOQDlN+5Q
ygsjSiQIQkmhHPd3YJMXak6+DXQDRETXo97LxT5QzZy8zHYOg53g7pvSbl/jOx7y
u9bsFqyMCWWvQnIOlgTPBLpiZ/m3+GlD8uaAQEVT0i78RcrvqQoyzXgQS6IFVcYd
p/g6KuZGrZg/c9rD5/dzODb+I2y3wD1iP3M1lWfrjbEqXagvt8M212HilCFJK6B0
8ZVW+ZBtSseMaNaKLW/BD0OWJDQnSbFQSmNYr4G4kOikbm6ey8ubJ2vWhd0Qk+Ji
ZX6SSYfY/dFq6iMcFwgZ6XlDwnFNTeg6S/4/39Sx1A3F4EAanV3M49nlJHcuKFGK
sk1wnguWKqOI195ydW7kEMMNnalUkqlTk1kdvFkxCBZtoE1eRJ3vwoDZMKKVU+oX
/d9KjpxXNO7aEInvkTRhn7CD3rDEjEtzm8SK9eP9CpfseQhDwV8cD7sxeviR9E6p
/i5+X/RYHvi5/hVdOIfBF6y0nvyZVaCwLzOZv4qKw78+HlR3M11AdXZ5agIO+enM
90UtvtdzpFxMi3czpkhJsk1JskLx0NPktIeBtK09xNMSmfJLIIpjvMCI1O3Ll4z0
nzwALssE2KGmp0Orl1TJkUIzq5ikrlsFsCgPWJH5MMH+8DX0a/1n5xNn+MpJjLVT
B3Akp5T3qiV6nkw7p/UUxwFudFp7HLZUcLzZTXVEiqEafkBSBeHDdi2dTU7GCzKw
1uZsrR8AdVMY28bq5aMX2CGDLfcKxKMSqSyv12xY7DmrxmMvx4Qenm+bhJQiqHpE
jyBcI0CGhhvWKTefonDHykNFOhx7RQ8Y6z6YilfIF37VKWu6Gj0RPlZC2mwRz+Eu
WqXIuwjU46/5Aeh2T/tAnZqti9oDnl33OXcDQQkSjN/SzgesDEaeGWL+fAx5hTcy
vSdv9nF0xMCT8jHeJxHuBbFYxNP3wayoZTXUFlEb4GIy8SST1bAbN+S2jVdGWuyw
MJgPQCyTBG/JO/KEOTZh+M9DcGmTdPO0aC/mT4qKRmuAqc37MMmRReArGIfZkPy0
xF6aZ2Uy32NGLjQkFdIilL4ZATEVRhCD9Z2bEXJmznt27FHumMA1ufGcF4vSsGdw
ZtEwM0gC2HAXXz+xlhQszfzzJxCsmYDXqgjmvi3N4RB4QLEMOG5g7441/+LfcAWt
H8SS6IRmxmpakddtFOD368xP+zZ1KxVx28mjQERPuuRudd9Zf5vdH89nw1buNRPt
aof5qeOi2TV2WbM9zj2OkrnNbVRrcdhTxMqKU1OzimSfKXX0e66wjlYDLw0OV60t
s+0KILin4pJaYQJ+3gs+G6sFK/4tTcJopPajRB/lV1ICBPyzWZ0hsG6OC+yykyJ1
oRE5gmsTyi1Ckmu005TsUvN1HGlW39fqEoyd3QO5/EkZtZztj0SdAahoNy8G8gHG
AN5CGBWa487eEm+Gq94VUqEblyE5nRkFVh9isGaQYLxx2mKLIh6FM7OjXMhW+9+X
qoiVuk638r/MB25TxPcRq/6Y9LUxj8fGLvsZ6A4d+ufT3QSgmmVXxb+lY9j0IJme
ZGjKdGisJ6hUaRyu9L2JD9+ZTlYXlOAlv9aomj4aFOK1Vm/hKKs6gJcXUAKyyptU
hUP7p/5kydBCbeSZ/QpeBssjdtG/7s1JmBbXEFn9tesshd8rXwqMkSqrFQqfqHA7
XmVccFLvB6xIW6MoTmgEu4M/4r7dq/iWS5faypCWKPdinSCzNfiWPSbyo2OiJh3C
6BZZ56LnPw0KYF0Jj5NXRtr7KG6P52cSNoChrmjr5MOfStuvbriD9DrAt70Qy+Dw
Jc7YoUnTTg0Ueukt8n5bEDYItvlfcgyImwV+M+Ebh0byWdASTgR+rUQil7sIjuNE
aQzKAA4i8E7/Z9TWphM6/OYA2gKTrVaP95f3eSdxTlTRnlzVSfX2G+N19gP4j7hA
0SzhbAmzIen36ut6Deym90q32dS/DWSmem5t0faSRWLiUeLR6kv7HW3iRsXx6AJU
aZ3QB64j2x0Ug41Bu/A/RZueNnpwkl9nC54m0rNQSCbEYDhU9lncu1GfrDTrjS2E
t75a/hKeRJTlWo2EL3cwqDWSdnM1PyULfAzlwMER6X5+Rl9zMxvPZyKXrlk4/sqd
Wv8tmzELYICJu6y+TDKWwiH7ffUz6zhu2c2xqukmVC8gi3pnD4o0Yf63G49oFnJG
JyTFIaMuc1q4FHV3eel//9ybUZ/BS0Ezrghhe19CI7mu+5MmbvYOQo69I/D783+5
RqxD6I35joN9ogLO6o/ajGN2Ec28qUo/wnZ7MeW4vZkJluOBxwvYL0gW7e4J46BB
h3dsOJMGVMGlC+x7clZhMpVSaorZt1csB/eLVJ+P/QmhRtnuiThEYMcEcpVVxRpl
3FZVOqkWv+0hTas2DPgWFZHCnom6YxGOe2rapnCtCtpxRhtTj8r0vUoaKeobWbcJ
uQwez8N/UW/FR8BvCi4Ahrx1cV7EoOPfDZvcPUpYD6Uiu165AsMe62KCtxv0RlNZ
RNuNbjWc8YxvGUB3j1yi3aVdHMVviiIGl5AzeQX4cyERO9dZpVIkRIiHWs6D+Hv7
J/U7XsMewRCSxQ2/0U5aizqKJUbuwsEP47oc9mpd1PAe4GqPiatks8NYuchkZDqk
giN9c3hBPEB8Wj1qy+enNexHs2z/iuF9rJCHZY1mf+n3eQNOX6pUv1bHhwNpKIWH
07CtSfMCrRbl8d5RmdL1OsjgI/YSh8XXDrMP9NV70++EEY1zTfUEvcabDEhmSP7+
efNfCxo4GRMsxLdyJ1xNTou/NoHweMO4UlJIqXZUte7p2Sa2ukv52BskDwwSNbX2
3YC3/qDAKul5yii194nZFOwHEf9yu/iplcrmOn0mMQmUTVAOBJNUNRLDwLlWtMTI
Urg/UXMkHZwVvCSOLuAS9YI0OyR3bm7pa9Ed7o3htBlWGHGmGA0Rh51OTrsZBUUe
bNsmbMsG2qurvX8AV35rkO1n5f8KAoX2WOD8bRXpLZOpQgwFw5wyVkaHKiiHmL1X
zJLhunnRcg/t+fUg6UlFrvPIB48uDRji5H7GCu+vMy8GN+0p0IVHTB/r8/BQDgl1
NSJKMp82pGniBz4SyY3WBd6JApSSqFkZZ73QHSZVFiJam9l2HbMCB0rg9T0waOpf
bRTFq9NSNvgDCFhWfFADkGdrcB+42OG5oKWln4a+8rH+T9/N+YoOi9rHUMWOMIwF
/+NMP46zT0P/o/1FSqCxS5rvOWGlavfSOHK8aKEgm/hIbP0WRFeBl79CKhS7OBU8
yha3pcMC6XZxehUoxAOsUQt9Om2ygyR8pq5FqJvT+/Pg7N2PldIZTN1RjVwgT6VU
pgvv8nPFAXaL40mKuOLMil7/7fJt/C3NydYJtUnWJ3TTf2s6WhACTT4A9CnFOfVL
uWp27pRwctXsZmUjMIJY1EbOPaO4ke0Shpncfhc11uEQiz9T/btVet0uFwSckWmN
7swUqxsW99C/yPs5hTHOPe1kg+aUP1uRI4e70pzooSwL/0xzWqatNPj8+msaYtdn
OlLc+LMkypcjQnccY5Zr7/VfJfkcxpXFrj2CG1jVXo5U2Qpz3lrZ3MP5Ws3NLGn6
Vc2BU8jYkLAKrr/YisMvOpwwbUzSlwCzueRUIl0YRtoV7/v1oJUPLz7ae/nvkDBe
eZx0MNd+yblkvmLEA2RIAq8ZLaIJWauz9FwZtbfa5xI+LRG6Ky+Xaa3gkEmttpMT
47vdMXzRS0Zu7rhk4awJvB4SvM3EU4JteVSIFKZjJYDHmNxzQ3RJIG5O24a4pkGi
CXVI9DYHFIO//E2IWC0oNWuYtfEHK3t+NLSoN4x8PCq621ahtCZZKWgtm+EQZqts
vqXe7BmHkPEQ9NdDlyV/C37yFyKB5z/DngCelRrwUPGBEJctWq7j1P5Rl48dK8Ie
feIEGc08ybcZ7P4Fb0TKvlX5QQ32U7zLlHvQryY06TbJqFX1yyXho2txcdiflMT5
+J/ql/t+asr1Qg2hNLDO1BLzJRzuLpiHsxYbwyToskt2xr8YE1ttNL2DaOlo+BUe
qcCr/p/eHL6CxMaSXj7imA7blolpBnwqm/L5jEWI0ir9jDkBlGw+9jTb0k4fK/jN
ADlFQ+SHxhQhGGE2SXDkIXGxHI4IEHzdS6HRN5P2uUIJp0hM3R+CTiB4364kQZb/
6sBl5Y/Rnjp4XozZmxNYES3x2kcUZRi+Jz9tPGQriwnWANb3CempRKJeNRxyCNsq
O0pFDgRGG/OW2DEP/Ot4Wx0Bpx89FQXqaLBtZL9Bh+GpvMbc6+7u6HzGFklMqLRr
KMOhEnnTSXEgYNsS/iHccO6Mty8X6qznzCMdt3pnriij24wR4PlZd8wiQ1s99rCY
KB0qX5e2nWHyFFAFk3x1PqoPYKaHd3XWQhb/zJUHZwL2rgCNJg3fvi2tKYJQ6dNE
ZO//fhU3KQg96O9ZQuvFJenX6hq5FvVUnWixlLJRE16XTYE/fs8SVKitt5M2+Mdc
hnHemF3IyGkzyRZ2f6MIPAcCp0rZ69oioQDF6ZcUh5taHf50Vm1iBYyJ7+/1kvZJ
lnVFc1sDZ+2h+0/nh9T94ozsZS6TU5HnIS+u8zo8sQjRAiQ+3Bm5OBTHV5t0538o
mf9Ms+IaGMqKxqu4S6QXcfQxogHfSftOi3S2617b7ZpLE8QqeBTHV/FkJgxozmgm
4ovkpKmixgndpWum46zXtpj25uayz3pFFTnK2q2hGyVs2rLBZ/WtSzadAtBizBKi
UZxCz5/+hRARk8T45kOGotscNxlXC+Sqg610qt37GcMuMddLN5QJZrhuwWs96fn7
YhcG7sGZNeA2WMqr7eGkTlKjTbHL4rOpuz7SpKJfbST5e0NKLLtQMEHis3eLNqyY
T9dHSbMimPUobT5cYmBv5rlxo4G9xlljgyhjXDOxA8ZHYkMT+BmFjammFG4kjAwx
78IC3ry1HowdWqT6vcMAEnUvyPOD0//SCZ6fQ9YviCzgLs1DkT2GhJRJoxXhjpEJ
JWodaTzJBqny8OS/m/+QluyCAAJXOf2BHNZA9pFGRz7TR3CDDJ4kIJ1mMgexVN42
4g1MvPWog3xyvllarg8WuqE+ZOxlM9OdWTyhX5xpPxZQwHndTwXf7E0Z3gy1lj8l
oM0BLfY6bnAkWcPnPJKvHr23TRkoEtfxAqU34R4+9vBfPg9zU1wErZhtuH5hZp6J
gF9d+o9fM2mYKT4naFsrimiYILkTCooOpyMtESZ8ACbALKFYkBoW0xCGEiJW8L8b
o90pK7w9iQHKv1LX64y68vhawahOLw7uo1GQVbRHRkdtPtkajyzhG36mJgp/iLth
jrthW4MxAaIqBzjOPpvu6guV6GZY1z1Z/zZ/wxQacV1quDE/W8EIc0ht8C3E9Cll
ScT1clanpNiYGYUyytNkVmfYwQm33wbFFJkVjoUs/9CWHuBoDjM1MAcdODrTX3aV
GG7qNYU3BTAcO2JCAlrysDVvcbtVUSZwLrk+nWbxEWWOOyl18IH4cGInKmLLZN4J
oyAliQwSIv1ZrDu2kSnRIM//H8tqVBHbRvCf8CegdLjkrMeSKQuwsYR+t+UltAAR
tkGupywDZEhrgEqfcfmZxY3+dsjjAA2gKiEoJ/h3Aw8AV4qgu2WzhMPFKH3VZxZp
tjZWJFI/qhqGPVd6svp2mgl0XvQxQx638Iz/38u8mNMcA47ipuKAdMNpLu12xK8b
xRvx1xmFUzeSQ9CBniH/o3CfT3RZLTZ/W6bgxcxecIBc1tZcFdV71MZBTyRCYJPt
XCbysYu/dMB0r6YhnXjqx4OhD2kVtAYUapzAoOf/BTFlHF5IhFBIBEuqUmXwkleR
6BBzHVVhAEgfAHlBVNFUoh4+xL45TQPFXfj0QRDb+alTKCK2+6pxmsLj/63Ydxty
Iib3hWu/faRen2GIX78huJT2syxE49YP89pkujnIrdFPRgYqcG7NqvmIJb5AmWZr
vlOXvfzga1PnGznKskRZW/I4A5bG8FuyPurR/UYsADrBGdWYRC0NgOxGGETmq/yN
OnH/kW4juCRTgowGMLnJFDPB++g0fEkStja3B3s/cb+wICwqp7o922EmK/+Ffq8u
XvtDkQ2KvRVWStD5yvfGkKFTI0jrzhxrtEW3P90Mur1LeUZZqJADUNM5tRV76Nqz
eplvpZLStgh4jpJSzjW4qCXDJsS/cvmOKSgU1neKIz11F2PgMAcV3eldltVrERhE
YidZooIl0UcVApC07EHTlUzNrbTstbsC3f1jTIL3xgxayAMDgqF0eHHA3ARAOm7r
Xr/N6fKPvwSWT/XZ6lC1WsD5f1+KX4QfV4wP2t4DX5z68B4jdutsh7pIDGQwUubB
2ZXhvVfzgy/ZMYmjpeyKYm/57JIHlWAUFyGP+JpH4r7GYLHZNLqd1QjMQhnoy1m9
Uq1hHl4cgDfPInNb3tbaPFI58OOI32xwobJ4Xb32hjps1z9grBSYYpX5HZcxxLLc
rCejGGW5vDqAyX12pJyMVhu7jHib57Nwmm2rH1y5Q9vTr1AuSBaFKH3C+1FNz3cE
bOcD/FgxV0gyo+k/0BMee4RGr+7TfNoSvr7c7seyqTSDxmrAbQTn3s1rAxbFEK1H
zsd0vI5wPP/LjmV1w99bfeRAJXuNQGXvXOHlTM6smKDOhQdqzuE6VAjSMt+CZwtr
8MMi/G0WRUzjSDsRk8YApCdhNLeV8oHy02BfaHvhq+HHmt83mACpy2oZlIF8qhUG
Lv2+4/r4twpGWyjYeqC9LxRI2QSM7k05O6IPKnKi1XfmHHFOGFOuHSscpIbumMS2
vA+XMIabawk03FhKHgF2WYgmKS7Q+W9iQIN0oOxLaFciIRDj5IYlK/IlMw5tAe3o
XCTrlNdTl1xTBnzJW3PaZIWnFYAZBNNJxLdaCRjE+YiU4qUvgMOvaouNR+1r76u0
dxYjccNKughXioZMjjaJV7TkjG9WrsHv1Ze5eSN5gvQgkbVhVf5cH+7NGwfWuzN3
6I5WHehJGRIofD2rON3hV2NTA17xfOQ4EizqoiexNEQO5DQgCRPP9WY8GQNmbAYH
Z6Sp9Ql9nXlY+K6ezTU9UpcdCjST4H8JBQg/IYXWnZpH2n6bW3AH59b3jheTj9V7
OKf1b3vC4+PY6M1wivtbWvxEPsjRKtOdBipH0DR+UrRG8OO2vFyrNms0MHqhbtIe
DGj6Hj+JmWrg/P77qryz1r3DOQW4wkXpiW33xfAMqazYpR6TsuMTNo8O92UIuKja
LIYvd5/gC5qg32Vd/GEBcgvwaPwW2w+FQduAXmi0FYjEe4q002DJCWkcPdCR5+9d
hqylmwW6fVA3JyKsTeFPjNgSx5lddHviGSota5JuR4xPfywnZSqIgdtRIpQvU2Nv
qkTopDxmb4l4MO4yRiE8e0QWYj7sxPel9fZW8ESuH3sr9TaLeLilLEM5WUbs/Jf8
kGjYzRi1gz8HNz9ePkqNIMEP+L3bNRd+AmtTeluFoHPxdtuN06Jnu2yKFznBoey1
lvXOTvHFTXnSiJaDS+/mkax2c02kZjnDGPCqbYrFuWHklcADUX3/nYqpvuB97csp
oYi1Tb1Wo0uRJUNGEjx5yA1u6syXynjWtWFgLHAomMlotc0nd/qDYZMvsM3kLXwp
7AC+NaRbSi6sCouaunErR+EMwa88ZClOR7otKMd5dlNsn6l1hKvem0rwo5mHOwJU
cKndkE0M1GOxJsNQc9ACF4DFviMuOK55SyAn33djLL+oDb+vwODWIgBDqYkMvxdH
nFZB1Nz4IKcNqkXxwk/z/ebbewFNDEowyxQR73NiyrA7+m5X4k/zZepHLlWxLZkL
+ZPq+Zyx4T4JlIFpdQWa8PLk7A8dxw8Q7SEkn3KQiohWzVolI5GQflMQHPNe72CH
XdNO8/NAaTppBQ37jLtmSxMq73452w1pqtLJtsXhbXKfmuaj2staMY79ZnnG1JoY
ovCTKhAu4JyzP6ySfdLcJ5pIhFt/yrtQoCnS1BdgLTYd62elpXwxUgbLavKyx+0h
23LO3JTG9PC853AAJrz4Y+eNjuL9eZ5eF9GBNFCArBAD6g9dWKU2ie6B3rzqthv1
BEWDqdj+s6FvSlsKKvkxLFzsY8t54qtZrEQK+k5WVR5+K23GaUMUqxpEHpwMvNLC
603yRYN/nlKZVwsAlmXlfFslmAUfD4BrywfoLLjlIz0buMXpaTLfgiRnYHL+sup2
kCDW4CcC0onI1mrZgVi1ZF57LEtGwCer8WRlmH2gtvfU3y4yzpMhddXfGc+0qhAZ
7qbZWjUV8Z6mJHOl/pfl87lREzZPolxchh6reXmd9cZAb/wY4kS8yTrhs04Itip1
/Iu/lxkje4Cgh29/5PolPeSu5cz+/DdndbuvaxN5fbZK0eyG4x8wKw4e7JvRYsfw
xrzkSEaUOs+ggxSyl4dGUwkygYSnE5+goXSOLCB1iF/53M++ey1gbWnzmuGLAa6j
4ebSfwRJ/ZQcdSnNi+wK1ePEiyOH86yH5ZH5QI6AL1j9F/naS5rKklWV3+4ZsZ4d
SoJdhNSE0uLzof+Vahl9BGP+Ce6+rUIvCEkdiaF/AhbhhsEqmvwD0/cOWlGmo2Wl
JAwVUA/uTG/nNsJfHbzw1UP4eMxQcepBCB6tXNuohpR8duM3pF79+L8mgvQZ8KTL
P52AcVXxP/RDhfD641AjorNIV11GZYpNGU3YLLxL45/t9gfLBt6rJ7Ud/B8L8wrP
7hLpueZt1zfEm+BTA+tVzAhKuCG71Xcu6aU/WHl6XwLgG+BwHFyNq2X04gJsmBp5
Xp0pwPTVYrMuMERXXDNPvllXqS2tKF/Zhux0FsmM9MrzT14AHwu2OuumafapotEm
XjBOrbCmGgPsa/kIw1+rfyC3Z94Kdc7N7IpiuyvQ6lkNhr79Oieg2mYshPZ4xAD3
b8MJ716BgDUC5TiVYHFr+C445y0nY/Err18n1Am3iKDmGwzQC3e9MR4e/p2QjkZB
7Lx/CeiTqh07gS0YKqi2+DxVZNmffaHN/hj+h8NNJTuFtFvTXkU139Hl2t4hi3cv
hNqf3+HqD9RpAWs1zCeJ3OPSLHxQya95YsvAH5PWx7NrO4alPvMMbb4SpnzIm4MH
OOKdpjtARVtyze3zQ5nL4aBvzA2IUS+JCpC064JDSL7TyEKH6n4YGIoldfL4hZWj
Cki06o4VytkWX/i0eYTaIcAjArNXvM9acMBdCaCXtqnFTY9cjTp8+nqD1rMc4I1E
S/Rg/PBcMdq7fOQJbBy3Qd4/f1qS1M/BltQN2qagmZ0iPyCbBSTcr/SIGBZ0TKmt
xihD9PChWvqFMxbHwbgHshSC4jNvidS7Pr+re8QtFV4/ip/cLVGWg70b7PjcllWl
4xcO1Dif20e5U96sw+Zi+VBO0s+KYno28BoZjDHcs2UY0ZKR/dSTLNHOW9z3wVd0
gZ/Jxkvfk8MPwQvBTVKXqnA3FRhkrUHq4GkRDl7hEP3TwxOjBxv9j0r/71n9kLWA
kOnKHkeCDQZ9em7un0PA8oiU6p+m63tJ+hJ79zRGlaYayJyN0josf1I1+RJ9Imae
QEKiDk+3ov+PzJ63lt20jCBLoIx/maBnhgraLcsgeqnSv0og8bCodqzinLtJeZqq
NtVad8Yos5V0XcEHBZANiDSaBYHqMkGhBG7KIoC6+VnvxlzPDjFc6IAlnkGUYIpy
DNnYcO/3kNLsj38+Zz1HmEoqPac+pGN6fTpicevnuSN+EKLIEQCQoWNX6NvTc52H
1Ua7da7htTMqXWLABj+Avt3luenh+pc3XPp1fpOcrAwNbiJcA6ukeU6zl569jreY
yalXO3IkqkYQN5b3EitrdpzJmUIkpl+5hWTGbth4SgvkngpFQDMjM2tJGcnOdP6f
ZoruOjRJd3zRQ7er9MWAAWnjFdViq81wbajf89MtX06MeQfdJOl7utdlTKcjTdfa
YN7qVpNGNoVeXBYGSocVU4e+AGEJ+T1YRqqOgT32gtjCkCZOFGE7/pxmIPSkyozb
qAf435w7UWcgSa8sEEqLaxpg/V3nqNvIkKM/lSvLrUeFD9lEnu3aUvJyKPSOmYgl
GENLOUPeW0rio/uLvPbm3NpOGRrVrkTdrxesY7hj/lWhg2u61M4DLJ5vLscqbpJT
75nVDUFDEXvLiA9DrNL/DWCgT897YaR+dKbjHPQLNmrmMZn17c1e1nWj3nKjaAid
WrMzWlMFimda7bWLwtOz07Q2tm2vlForJcM21pGRnuYW0gXf9+BRDUZCtuRgWp1w
SRaFYJa+9HbBO77IDuPaSyMWd1gXsMztgBzA+oy9qwM/uUhkMrHBCMZseWMiCCbq
sy9OZl1MVKpsonuELftKR5WZtgKwscmm5j4CMxnP6SJ1h9HvEs6qJbjEb8y3/2/D
FGbWJa19U3TbS+s8STItfN7drRtG0xpTRR3XjXAXpdxa7e2Vo90d/52BrsvW/mMQ
n37h+Sd9J1U0t7LR/7slcI4kG6h4k3Zkcqo3KOQHvCpVFTAlKdxx7W+e9Y7ojLJk
nJD9z1rTjrTj9wmszFxbtW8N96KIHWaCfVGxCMqsmW7uQkDQ3RdNOuBHKqh29xSK
uUy1Xk3+X8sReVFRKL1h5kdXZ5wpJndKfE4SjmU+yzDJqJgIzXmuqOP5jFqBRC4e
BtBKEgAEzHjaajnLwF765rHgw00H2IcbakO/syCGSLVDm755NpzRbF341KFKgKMa
Xd4DWevaQwEeuMw7etse+EcyDN9w2NXL1h1IBMWJdW5KdQpeE2mZxiF6HJlxsh2+
rqHO6vqscWmASlEcGLzHuIA5cgfXr1ORL2eIU66s152jsXVvF7NeMOTyFq4UUUIJ
ligIiSQ7ZW8LQ5QTMrMBLJVO0xZ/u9qkIVmeyU2HYi8B06jDqz8xlAvKqHjb5mhR
l/j7W1LrY8+lEl5rS4wmUeK3rT64ACS6PXRtMddP2gbbz9cV1Q2QLG1LR3Q4vbYz
2Cd/TuHgxBNNBcfybUFhlYhNaDLVRlnN4otc77lHdAhOb9ASjkTsoVao5uAW5XMo
eZWKXjlvgzRwqm6EvssS9V+sNNEYzyvfpbYSwb1uHYnQld3UhPTpVEBNG7MABA76
VB5K+2PI47KNbGs3AkPCEsyEOwwTd0jOSwY9IgSMBIeLzq1f6MNlOZy1huPtkOWO
bJCj7j/DNNcFACUe7xyFJmpNkIReWL3BKL7XBVAXHCENL2Qb/K4lZQFxDTp7IRT2
/ttfkABuKcYk8Edw/bydLTxx1YH1vqmVsryvR1bKPlEchzyiq5axDDc0n2sLdOOv
Y09x3c/B99Lo/2RS7DWVKzdGFIZiNzUc4bUJU0mhrDUm9eElt4AlRww/y6sZ+QLR
s9wzSxtiVoGgvwxZ1pr3hKEPi32fOdG/Bc2Sy5h4qosxgUFTxequb+Oay1RbCyIk
BKOFQf4qCPNWVckIxREJlDCPv5MD8Dl+JZUSXyYie///TueJN1GZ5L7jMPcXRgei
gpCmsVlE0aak5ZHeYSwdV2bZnyxxnhM7TnQlpSfJfRbVLi5KqPpTdnwHzibltoPb
IFW1nIbYyeQtCtH5rf4/B4Q5fDoZy4VnEYOwFA4Rb2l2+oYy1qhLKtFd7DSc7PQk
9hwKowcXEmnWFPLuA+CWLXzEFUgOEVvQllk6ZHF4AxGQwE/iptlsGjHYtuuglqvF
Am88Q0d3t16QCitGB3JfOPxuCnOlIEQjG8MdhM0t3PWXTOdxLLCq33qF9zqilZEb
VSh7yy+dlNDr7Q6cdaiQo6JvT+SGVRODhRa8BmiZq3ion+egV/LdPeSEFZyOpyVr
CsnPSCbk8WKOCSSVkHQQEHPPpG6IoxhkEWCJ+vgV72CZRCi7kD0WX3ykf+sVVZ0j
hWm7pwEcg3bqHp5+S2HU67XQ7oOuCQomz/CutRbuu9y+BCHBTqeKpz23/mFyQAC9
jc+ZJBzMhXJunbF0yslEkbowYFsC7x6mSORQrJuUuth0ixikBKerTqYZ0GVpu83W
HLGDUr9cAOdSeTnhKINbznungluIlb9VuCIQ/jxy2OqFG9YOglTSyhTdssfzLscE
7GNPaBVUBZVkvQn4Jf1hQhj4lFsfrAjoziFmZUMnApnUDvQ0TMLHhZ43rq9Jogg9
S2ZfTfOtMTu3K17ocD726I3r4KiQcbZzmVGUNCyyRGEw+iVIp57NtMTxnIPJqIU3
jOo/eKY9JgNmT6wZwhwuDp0IEiRj7KjINlPOgfUST8JOAJtmDQS8ONYCHtj28RkK
9v5Mb6M9muiGAJ14+goYtC3Cs9/sAw/7ZB4AwQAZKui9v0iqCgQ3/5FZzZXZjmkp
ZUthJWObdx25X7FImsYNV2I0+EBwcRhO90TFVfhOo9RTMJjC7KbjJHOFO/ywV+0K
SIOFYfmfpyfGLN6ZgfJ721F7Foi4xDvfo631Zm8z6dwDQu4FKvlT4ENf4NvSFBnc
RCOliDcqD/k+wGYm+4uNBY9YD03wC6iL77FRxPFHng8EfyZPRmVDAFGpHHgGypyb
mOqIS1fsCM5R+JukJW/SJkAULX+zL+Du28E8kOsFHowR3IIIceoZWdCMusBA6kdr
uTD19Ez3cnS0+k/Cmk99i4vG9L2S4oYL/gi9GkwA+Dto1T0uK6WwDy61JGSTh40D
7I9nAaUgDdxN99AXPdHi5l3RgRvnhZkRcAc7fLMoc+Iuw7/inF45amU1zFIP8RXe
dYRVbEF/b6bqWk/I2Yl/1p1h8Vu+use8CLD551Z2IWM9s71R21tVNTtg9Q4GvIgp
qzyncrZjts08EfngKDji/q4+xSNMVS5CzZhCSz/3s3+eRY/SbomG37TzuDVIQPwt
83E5x7gCSb7jrwaKzb4rCIb+ZOxnokpfxiMMH20RtwNky2vQeFmdIBOxeLul9SSe
Kn2kCE7a04x87cqNzHUw22XdX0hXt33j9OeGiLS9HFqsy1BDhOTW28qOocTKEz7D
N1TdVMqoBQ3uUgP2SDJvkJbWTuqSblJdG1nagJCY4xPi/GlnJAjbwhmzivEEkRjY
mUSZLHh8A2dMMsy26UWgxt/PHwFn6FR7fbBB6h9n8MAIc+bI3pFwkz8WbwEHrTT+
AiCs43o7BhdtJsmOvjznfhR6Tr/moG6YZGTi8QZY4mxSxVQsvntl74oF2QNtio2m
br9sWoG0Ve/Bp91y13ymMyw9gJ9A93RUHQBaEzcs2ZEUYv18TShAkDDDzFAMrkG6
v0LoVbyWzZ7whuWsA0QwKGdaCwaPmlDPXLRHyC5ERN7PjFZsl8yZ6wGhXRsSkVVy
YIt22NsTCarOKA3CuCkuYaESGhYBpStDPT0YEczUXVaHm5OROeNC2d2E01MoueKT
aIq1Xi8tOh5KWkpQ2vZJDbQicvEPEQ9oNPCViPHVTU6NSACTYPSZIT5iX+E7dczT
yLgXPMxWSMd5xpcmv2jynhA5E7aOqvS0b6YwA/Ddr/HXbpMa8tiUcrw2ilJEA7VV
SN04nYvQ8mlNDKcgjHIxAvRfM+wLMB1g6yiAaUWMyjCe0Ckqir5W3BMh56ICO/OO
s9dgJuEjJU72Kwnv0M1YjrFQP1s+ayNr97MF+H2lifzLNiCBt/AaDyaFPytXwruS
Zqli5K5CZf7diHldG27L37MrfcdAXATMSwDDo2KM0MqQ3yxedhaM0XQ7BH3AYOSL
fIa11AFimoiRB37zrNZ04je2TdvPTrseDWxi3xndTVWpQtJPkoCeD01dDRJatgl5
yQYhGOh/Z16Gz4amaRivW/s6vNeK+Y9r12qS2BftcbLIeCzWIQSqvpQPr8Ke9f72
abcHGi+c4dy2TZkuCQmW04T26p3F1a6+iJnonSSJXMM+EvFNEN0iRxt0ih6u16EG
WPM11q0qsoctXanbep5RcLxYOTHtcuIqWr/Vh8Afc6XOlGDASTX0NBerlMA+0ufn
ivZsvFcrRN7xxxIJukAIBqMHwlzo1dqoREdKnWtNx5qmSP7v/c+QQzz5SQg3jwD7
aO9SjJXOE+mMhU9Q2k1fyYn2JbtfETDrFtuZ0vYBm+jOIYovdNghN/a4YLZL+yRa
82H7XKVzz8cvOSmoXcvpk3AtWGNsjFpG0WmYLzaP4FyU2TtTf2/DwrCGmfFvxSVV
7YZBlN4kVz/C/F619Xwxwqw4CSXxktW4HWjVn/6CBruTKzqfAoT/er1WU1dHTBSP
dolSO4GIUvjGJgrp7q4ttT/MtdiKYuuWmkgtIC3weWm/p22dwTQjlHno1n4nKUjk
/56V7PzUnY0llOlzJlL6T6QaOROMdt5eLcFkcF1TC2qU7W72ZtFsixAY4vbGvpji
TjgvxSLy/hcTBCvXbxWxlnDrzSy9qC/kAPefJqa8woBHUdR2vmdjJQ/BM2jXzPo0
RlfFZF2yisgfCTF5OFA6etg+Dt+BG4FPUjXNCs0d1+fAnGvggZVtJb2PS+t7r7SP
0B+OxLLgJfn8iBJYhQLg2iiGc9E8rlYJvwSo2rO6ZFW9+KtJ1zW2BDvMBn3YMIG2
7b2BgKTQyaG1dlQuiDZu6vYbSsW88wBzS8rCz1MhBXVK2e7whO4Hs10dRNgOqBqP
svuDIhl2MSC25h/0kYyNjOY0cqf1DI+tMuWttx+WHGJV/+SYFSvezLXWiF2QLT5Y
czmG8gvJFYxGrQBCxJS1wD2r/sGSGekvQdYew0jnMh7CDhddjoiMoFay3JNaBFEy
ENHJGawNGDglJd3FBqtDKipKYyZj9JWWj1gpTXIAHki6aWXCzmHi+FnZGteRbM6o
qTuAgAIL5FuXVTRJDTEcZBVNCy9g1c9lE7tppRzzV6lH1gRFvADfASIpLtr7Ksyn
Sre+1Z764IG8o/azKg8UEA06nLEFBDayYDaYwSEQ65qBtcFerSq2V2f+eFhKGkK5
57w1Tfpr7sRPabzBKIGIPpOhEK+8rd+1Kl3ZMe+iBZ0AbovjffYY51FYlpoZucGI
nfRVzjG4Ji30sJkCFy3LsB9fVjcUaTCViSJrsF1VbkxtQimOLWJ2eG4boWHuLinI
lQveXsoul5AZceA30Gu/5ie/xYiMSOTpvnPEQDT5Rrzx6qMZvbHyRFvuBJNobRw8
WxY0zZODquujFSFy5Enij9xLhY855RPo3fGw6kaLFZXpSrtxNK4d/h0id20QzImB
Wmfqo3GdYmd3CFbTmnUNeXkSboa/IcTtOtTzPgkbLj8G9vr+GTT193EZmYLHATg6
oVPsmwrs/enW8rnv4LCQ1Cck62VF0deT0WAgloV5Bhsbu+9dHtYWARk37G2ce2J2
8h2XiSxvskSjja0XuU+XXdHpjekAsRsw4tgA+7h1Nj9GVYJHzrL/LlFtQlUb/vDd
IGd06a+dcX/bxxu2QKimkuLQfJSf51k/b+3IRl6GodydOFuz90YM2RLRcI/UF8iX
x2PwL9xOTBaZzuOhCzcYsKT3FD3iyydlQFzeqUIx7G74OLxB6O8xMO7dR4fNFnrB
8boLgXtwOQMY40SZhQS7zq8Quei+/7xoldraVB5rqeJvr9ouovtqV4ZSeJe5hzYq
IRGG5FvKnkyjicrXmwRCC7eXELlZn5MuVfjonhl8fk8eNt58jmpg270kJRwbj/FA
OdXB+R/Ebjoi0wDhyB5cDVivxEFMYjI6XalzHb5rTqR7h+qVlI5Nl1vZSBSeBJAy
A4rIdqIHuia/FUGWGfVMcfRhjsCP2Rhg710pYa6I6PoDecmlBuDztySMTZgb+V+w
rvlIf1TwxIFvCH1rWM6HPUMgepZ6/UcyEP9GoAT+OH3dETHCzX4UcyXfrazxdN3S
k3euEUBAcNEIOqTyiCzxEVG2YPbEh4uEke+MV7Af2Lz/tykluaHbPE24BNZ5nmO2
ZV0YPeuawVs+jmyMKG5t2+omRFqFfS5J1ghCIqICg9LPKuK82ovWRk+Gaup1fMWt
Gt8bFMYyd0eZwsTQOnHSrmsCNqSLItWVT8xarp7B5Q3BqRXxt4EfF67aSClcUsPl
59WNV52zhCSC6U4osv7NC9eqENv1K0jEHF8vk4/beGAMF+4K5NtZ/1ZL464Zp+k3
qmdHDNYQLttlN1WJkUVl7aVDlbzBzqW+tWaelqmHvz3dQ5o3DYDvcV+NSr0hpDUA
Wl6sFXws6/SG8rrJTwsbLdiuuFuYe9lG4tMvE4hk0ePoi3nEcms9d1AwS1b0hbvV
OmV8cxiJObPVwjUUhPSmAu/QVAK0kk4Wn7miADmT4Q42zRZXp1GCnhGb5Od7NS1T
CTsygCHtayd1D/xCOzmqrt4ZzA2VBj2yRBFyl90ahDC2ImtfeZSFq7gkPOS8yhPP
z6gj8XaXkf/LVd5/U8m8V4XMTHpSnzdfdGMbL0Dcj2oImiK7bVeI8/UH7Y4/um8p
r9TopDaDCX23XPCGIIb5ZYuyRRZXhJJlR2/G5AzUNmTuXx/IUM/qnvQBdz15tj4a
8imIzEZsrHkXeLBYrcv5hvt0/u0gW9fDH15NThwLm46M9OCIC9EGN3gKrvJ86rnN
8uPbdG1BZVF3HdWzBgeOmMfwwI7vfOWFtdDXYOv6JE9yQgZaTM6dBXB2CQSjzyRy
igpLK9DdVBnTlceE3zplcZEVfR9mKbM9cUDo8aTaMp/9aTjYz4ihcpaPGdhCwel7
zDK2MksIXs464n0jJHPgIqBk8+TpErjDDTP3JOCm+JndhN0XrmYcma4+d2GMwcBt
//8hizUvpY3g8/8+fVrSDGbrOfcVKqVhslGy37Kr/ZxBdfac+1P+gvAxajLrOBE1
tiCBtopp0Pc3CldlEiwknsynu3HCKmFgbca8Expn8agYmuCrgUc46BQ5KL1qGG0U
cv0u+otWAlucEo8nvbvjgPDL+F3x8dOY6YaXynfD3T5PhegY7QTDcR3bGASHDq13
tL2EG23fxVbLw1ZoHpeHJJsGW0WghsNH/09voUq2c8xtA3fmnwXBp0nsuE+5l3Fv
PpEI/XkClcmoClSA+mZcw8mJQzkTpYcIO060CSLJYYrkIDLWLfSxrt6KkNNrEr21
Ol9SJp3ja/QlhcaUILWFEMRArKyBOEhzBt9K657bbyvEEpSsUJwM2NVN6VhSJgG9
av9RACUeJzOThxRaH2ti3jeb0HyIFWX/+A5Wbn/P5ETWzvCyewz1Uh13FEhidHk+
RFJF+17yxgzdP9NFw6yg3tkKqhkQi1lXyjcP/CO7aT/4eMPXO0PL13E3xigEJ1OA
YrUgm16MUtrp1JLw4sX2igY3gyuv410DkGS2q9ayexVA3bMMA4QNZCSqiIKl36CK
vabeB/EkTAF8TiRDa7+x5PVfRRupzKB8zfA7quOahqWf3++AQoryeuarDYvYtFO7
Q3chZJVCW1Sl1ypSUTmoRJMfBpAHaJuzKkKWwQEYSiXOHOqpEqctF7zPqfFo/RPv
D50pnzhMwFn+cPJA4TWiwB9v/Fy8Ua5BOfQGPFT5RaVGuPPKV0+cM6sUaZvUjyRP
ZtJJJ4MpZInN12ryCV/XOx7maTl4NU7doOL6Jy9ZC1ObTDMGjR9uyeLS3ANx3rxs
jQH9Miz1J7/ccAK4cEtNtnuJljuqTzAh7+cSZwj21S4L9Bp6nSont9i/ioQn5HSk
1s82upcfzQ85AMBiIlOtnuhQJL1fHXvwTWhwv1jUoKN1fPuVl2hTV5cSe5+swciD
ItRFwPl2CAQdf/frdoevd2vdOwhMJRKrkYEmRyOv3v5m//hQ/Xu5eKgATn/z0u0o
s59+Oj63UskM9PJEOduimpZi0157xYIVnu209X0cVTyybh2rndbc4iTO+UbeqwnI
cWDIwJbWIEk41K42XcQm0zkMocmJ0ZUs/QdRkS2l/uYOSEwcPAMNEzLQycaPQ7LN
vPYJtyT6q4dEfzSIywxzPfl2nmx6ybf7RA5/Ss//AS6YbarsO3eXjFMYYNQvZhdT
Jtmf/aCL/8EZCgg7pWknbf8JDKjkmpSp73r+YirFFRpUtQTxzOBBBVvTnFloeN11
kmHH+26Z/wjxgJu2u6iP66KQQguZvSiEiAZwb5H2jDY+Cj87kf6kRsDec5Xn/wxj
RH7jnVXwsdKUIz7TuZTkA2AM5vSwiYA39xeQwlS5qeaN5fe1LDmMsfXOmYWClFQh
N5m/Mh3f6yz8DqA9m6/Gxfsk+RIzBYNW5qwcGZXhu1uQ+ljtEFgZZGWVWz+9uXog
aKpXyl6zxUDM0WJuzUhNIMs5IASAvWAiezy/24OFOmU3pmrtgCPYxw11N5cmpgxT
ROEL90TrJWl9N6zBun17Gugj/TEoMrBGhY9513pgqEBV8qFvfkdCsjxYC3eWHOv/
mpXmwV1EBDbAE6LfKGvficzgWh7L6kYqhu0UFZeuuXqEWOXkahDiv3M+q8HluA3c
yWzKUkz0tb9fe0QyVb1cZAB0tfy63CqsA7pBHt/vex17SOKx4qxG0r5HFsYyxLx5
4iFK7d5QF9y/f+G9eVErmcB1GXvhUsoYSqADpYVGcsKYJretd9YpIPVnvVkqKXgG
Ryb/KnzCgyPfPd24A4KhpnQobwuY16oZGJj2WVvyHHuIkdj0TMvr75u2rPKZWG2a
N20k8ACEwkNKzqi/oe/2WWDcWlfFX4bSwF0+NgDua7QMI8/Vlj7uWiYL9sBUzBkX
NyDqjF6t9A4HbQwn4Ieix/JH4NhjG32itznMwyAkDXO60R/9PBsRFbB/fYPt1gCI
2NBwb14vmtSSUjLAFJfsl7R/S2fXJNJ8UBpdC2BRSJMFlKREd3PDYN+7tXUVfrb/
kj4gyg23q/IgVi9hrV81C8AF9mwmGuI3fj6UuIy+HuEMSFhUYPvaZBB8TdMTc5Co
4l8gU5Jd/+S5kV9rTf4UN7l0RO7Gv79xuf4UP4SUQ6d0NiHGyrL8VAUl6VlNovF8
it+E7ARP08X9L25dTuiMwCS6QUIPv+TITQHl3zrs1qzzMFzxM4pWyU4xvXc64kLD
SvlpnhAj9FSLLkylzduQ4NPYrOd6G2uJxqAJvptbtt2KHhyJdPdJ7WOBHeqm0JRg
8aBCpmY+7ks3BgY+olpj3wjfTrGxUu/9TeAB4KhlN3QeOSnNb7UgAX+e10JrFlBJ
Pnv9oLr8ilX3gZ53Cmf3dETKT7fFtxYCZWxC7V3axabZcXvgks9eemiGtCXY0OQJ
m2gqceY3G2OSwh7rTl2wTUA7bJGbZ1or8j6pLTJsSIUzHPVP9pmGOdjIR1MctNwL
79twYJKBwA9M1nwuLlPcwIJrB7rlgQBZe7xjq4DOapEtbQWBvHsQEQNwdiDBIxwq
+w2Lw9TYI3wY9PqXbf/Yv3txrx6DuXKzbMH/4ZVD4ltf4Xh3bKoqJ7BiyZOZ8Uqf
XQ0S+Wp1QozQZKCi2fj+ePAxl3CwrY7wVCEnKhVWNyzRBaA1UuGb/zHf7k+CHJco
T6oU4fumUAZzgTrgirgzaH3ZU079S/s3ot4yC9JHyMbX0mclzPLy0W4oknODwakC
UljB01PYwZqFZEPgGZ4ZKP+W8e+gMhRxaLhCjtSjiE8Wp5peOfwoCW9fiMvZ8913
3Kf6167YIHLHNDnlASgw4lryVZpTLzgAI0Z5NeIBXCOLjIy4lnYRn3NtImT7RhVK
bBfypYzZGcNPIkCOGRg1OyWdqiz2eTi0BCT2FWvhZ1qSy0lItgevAMrFwu126Lbg
AXZmf0afA2khPII4OaLMiQetc9a3sXPT4SW5CzQut8IbMxKkTew2DciKt6USKH5N
EkRm9vykXjNlUuN5RgQfljL/rzgR6UdvGCm+xFt8+21rDl1Qn6/ja7GpxVB+nB/v
kkyWsknYFgXFpRcmk1UdtKqbl77P/lBzcWPgKbz0EyVKZjUaPOz4xZ8nrEA8D5Ai
p5eLZzuNK1NgyvpFvZC71bxP4hbSeVzOmbdQMtteAEEA29QENSr4Zn3vzsAO1b2n
u7NAmMHsHhktc9ypOjxZblGB7ZGn7LdGXkQQZb4MHz3bK2HBYSD9/wo17ZaeXaAS
oIziPDFmXiHUwHCwk95iUnfGxolWiXmWpzPpSpP1ov0bag9ONbI1u+MO/SqIRFDA
f7mma3lLsVoM6AnmLbQPPaNDrn6MDYXYVHnpEoC32UXuzC6oEAk+gyjJKQJdEd5F
2TBq22md3JuI/VbkY+0LLJgMdyZIeTciMJ2h/eH2B7vTCoF0YacP86/Psu6WdrFg
CbRxFuh5KXDEnobYqy6j6Eoaooj+teLq3njDgJXekvSzZmcUcH1I8kGHzDEY7Z2B
53oboSZzZlS7Cfg8HwZtlyAWT2NJSxl5PlwLbrss0hZiY3THD65mJtuNAdh0iUhB
slYbdK4Rlbq+mr4QXkxJEaPDQMJRAuO9WojWsvsPORhJ00UhJso/3CVTCfuokc5g
EmuFDt6KJP4JOgQG2CHFmIuGZ9/vdPDll0yrYs3b8IU9fbBNtKTqJMJjO6yX69f1
NBnI6Ct0T+HnmEEDl9K1DxvhAdq5g93ktLHJaYFtt3EnmETlFto+G2XV6CFATJ25
xWryPNBHDisaZKNTYoJdkyC9OfhJSNFFNJJosz79CD2/uECQomcvKQ/des2bLVzy
lWV/OMLQiLzz9kpqHxTmpNXAGotE9mbTBrcfs0X2WzQIHmuLere+OaItrHtudzvw
PBKR7HkO2VaPB6/WYkvvzNOO1ESIDw+Pw2dRf2HwcIENC3Xxb/+SDLpgJsfIXLSS
uvGFYPZNv3MqZE2ikgoZOR2Rs4+DZlqGPX1ywh7EYE5DjmG0jbQrAvv3ymhkO1UP
IPR/oU+wgtspTs/gxCILQw4gf4i4oH5I2334XOCVq8tAnlIPsBhJJenjpRoz45pW
4Fg+y7VtkEOqSygf1CMccHsWq0uHIEGIj5MrqJecv7MdU2NA3G9QJfU+XaTjibYb
qIANtaK4rNYbJr2aH7BI2YLWNuJTnZITrtz6xdLP1munpXeNByTgkrVIuQoF5619
6UA7skDVYWYT86/3KONldQRGHNmGb1DNLGMECi/Y5QQd9DZl5gU8NiVWfZoyRfKM
EyNZXPCem8nHNomZhM++zGXCo2vfGP+ETJeG+gxPm7k8MoweHX5QTWrekwdER1vT
4LJIZzunawiI3nvBPbhkTWsVm53qu3lo1f9c0GhjdQlB9qb2NJ37EI7951Sq6xdC
7SdXnVUL1d01/N6Q+VeYPY01WU8F30fXQeEm+T7k8wVnYKIC7y8OldW6GkMkNyor
s/VGWEHCD0IPY+RpGglit+Togv7K/mW8oR+EYw4zERD34nD8q+jM3udIA4IU57CM
a5b7pldiIzINWvn5gQj9FW/rxbsRhSeS3Mi3RZhS3DW56dpxejn7Zz6kxrRIMX9n
ZHB7xw/LSTym7HMgtf6pxX2Ik8J2pzUnS0i3SkNpyG6Esr48sc3w+Kq0ko2yl7N/
xOtoObP/OQY6yWjIoQeg02grZ1AGeP7yoiv5fuDR/+Sq69uLL7qw/6/lBLHaBYzN
WssRTJxXHHpkRikVwOy3j+4tqQUpmOYsWuE8JZNc8Dz8DIr7WTQSZwXnbgVavBPA
J5mUVPfOdOy5C5r5nvy+lsBnArKwy7SZ3VWXvqfgJtI7FyRmdea8tx0xGU60/cdj
TDRSCvP/3zTu7El1lh2qArWUw10TdpwD5VAxbFuN8naF1qPR9rNgiSBoWYWQcge3
JVKP8w5IRfw+hFghvR/wy+st5eNzJ7ocuCCuOq0jpTJGw/ND4lbN1xkAb/JO72H4
SgcNLstM3PpkqWu6DnkM73EoSVtgcHvE2Vg3cUQ7ZZjTGqeUj0NfjugxV3JBjcVC
FytGgR6Odbcz5v1RG2jY0CAdkd2tRSYtltFBu+IVILEmLj0k/J4PosDVluni03wt
8dTuEkvV3T08fP0RMNV4xfkaic4gIEnoIgtN7rs1mkOSb8sVsqcJb8bYNgsPh9hV
5kNNOMAwYDE8qjqAFJD9/vaRRWcfo+W64lmvNAYdrf0xEsndHJsBzbsz14pQNwsh
JpdUVR00JwRy16KkZSXgGa//lIUOEaEhSA8qdErCK1kwWRoNX4DNZ94qAjBkBt2M
IoZG9UgqHyJM9wPoa+7wf8wPkJq+2ZAgutRNYHNO98K+p/zF3SYTgsJsJfUYwRN4
7YWTnUjJlsJF748T80qX7IBnHgYylI2ycdeGQwLDqnVvb7TCAFwE4D/jcshykqrF
nwd2HJIjNs0BrSvJbW9VebQv5JzMgFWPSXG2KC/QbAbuSw9rtYEHVhujYUxs23yy
A1rkSX9uTSt3zWTbCZMdsBO7cUukoAa9ScIPXHLAvn8DYKl15dPjsZUQiATwFr3j
NvBp+s4Lh4Hs6/Dqe8FeZf/k9d8Xqp0NhG438vmXCsxGlB2XD//SxhKkRQwWv7p3
tjL7059qq52b0aDeB8CvPNY+K2sXsQeYa8PqRN/ixTnTZJOcdG9mFBRgh7SHzC3F
ECZFU0qTo6gPvtTzkX4agax31/rlFmME2AZMX+GIVv8AKH86UXhaZCXhWwSwjqmc
D8X94GMbamE6b2EsCVu1uyN9qaQnxpLpRJCAmAcEssarW/JIS+B93CKraFVBUzWj
z8n155el4L5TA1oMqpT3t+Pm9/DkKQDLmnquOFp0SlZu3zFajSIXxpcNHDMElHIB
kU4zZCE+eNbqNPY1usGprYKtrDsucMzhCC91jrvm0VsLC17kzrh+On5R4qzL28cA
0TZeUGO1b6W93ou3sTf2Tz5u4W+8a1iY6p0A1qvYL58ESfv3QzJgXTBL/r7oI27L
WA0tIkNj09wKZa8WJH6UQxSuWTj2KK2w9QJAvLiNaddZMwoKxTF7v1aE2jIk0Mju
bdl8MnhP20Y6StIUqNLfT4uZa7G/X/bz3YVMzBvR0AEfRrq1V3Ms+IZUfMwxvxVK
reWmZypd6C2OH7A4hFw9O6alQgzLBca41+8IouUfnFfw6mR9Kr56tkM30ANIfsCR
/gB1n0+IHIanniqWPj6qHeyF2mIbWZEiAohDRXjNfZx4vQD9DzK7cB8cjrv7sk4b
OgBpUsDLv503oQLHaNH3+8bXn3xJC98WhOgwEaO+UOo/e4qtiZczIJbV9ja4Sg2Z
DKDQDiVHNDv+qAGwSzm8Ey24+fvuAA2gn7N9SN77WDYx15wr2C3+6yIKuJYzBgqJ
cVtbf5iwjWCdkH0gN/kunCboOVrNcxT1dCpmlJF1u1z0STcZ7uSzT4O0SYfujErj
+nAjK0/U21kXqpT5CHpf78GzSYYlNpQsyoqgdozLfmO9iSjFvkklguGoKTJe9Bc1
TfqddfCQRdDktSanqFtXh3qrtRet2UaPeuckSizfF50fNWZNn0vD8DnZ5VbrR9pR
Wmx5cgL7tgOuCEa2KXD1T6HoTcccyT7f6/A4RRppLSyBC3dLAx4JlCLc8qSq9/Ic
2fRm8rvGIP2e2ltnBfBEUU3nGUSLFsdLfWy6qav8TV+9VryHzTFJpaxv1uQcCLDz
gf0U70r5nCRD5EMgUedr2malzYSVIcO0+WVS6Ec+N2X/6PasyXtBcioA6DZLkyAj
p4TbooAJJkkjFMVeDXmKyiaWWc0SfGq+65zgBUV7B6bQ70gSQZlyE7IWKbXYAfi2
/cvmlCvkUlpbEA4AdTZCG99gyyY9/f/t3zye5QI5V0Hadt0MGVw/anLZnwFLPOZd
fsddZN94uNL27P/0v/qVFPROteu77QaoHP2k3xnXdOf3mY6iRHVhBgeG7c8ZpbmZ
+CkwyBlfSU0jcC3uOFae0IjkfNX5zQPx1Vx5KRDdSFTZbSPtUA9sLJmJMwutpDqS
8eWtHku/QFdg3Et9/ixUe3MjZupz3itdfxgh4Oy2EmEQs95vbQEs9cn+P/Jv+nJS
eajA6wNgoJhI6sIiwnNr4YJsIFE+mv38EsA1shdoD9Q9gU81/HnG2XLuTs4s+hBN
gXM6x/Cu3AHvExV23fjwJ20i1KWNLVkvqqxWJbiTaWU+mK5HByZ9G0ypiXZNOrPj
1xPmNSZwo9vvFucTKqc8g1p5A91E0om14yXW5ymKogQ1zoO4uXJXZowHvx3AgVH2
qjGiRdDN3OtJXGXtZTpvyVWImoYlHzBvGQ27ZJg1UVLp4Tp/t/wGlfAxj0/9KjSX
0CArfHWYyz3kvAP601cyKjX8rg1OMrqvWpGO3VKKMKbx8gzdCpehltumjmh4ndNu
tFFe5ZmSLifP1i69/dRg5XosVddWjkjzB9ny6sHMm9H8BLh//FCPJrja3fM84/y3
jaZMlB8uPMF/hEXCr4gF3sAtahyAySWIw4NNCjqlLUBpOfoZjjcTryVvYooTv9ME
jEVzoB4F7bloBJqqztET/uPrli7Z8nfuFXg5ngB1J8LQl7YVZtF0mNlwhCJ7sGJa
2G1Q2uxMGH7RFsrvrevF1Q8fTANLqZEQEiU1dmCWGW6nfXtuid8392wClNCgTu9D
0bXZVBVtOhOQAAj9anRWT2qWyFSnoVebIyNyVrTcDxVP4kPNaUTBhTxxcWJPQePM
pcFoEFpCZi4PI0TjZ4ilh6oA6K6WhS02MZWgVMo2oU6sWzPoPq6oQyyqcB3BFNH3
9Z8BZ+5NbisSY/lvnxVa1VQ0Bl2dQLresd/Z4lky84dlAiYpaXCFVaDJ3QlMIlVl
o6BD9+V93MtCcjIPFycPWLFP4/TMUfK07Nkj+f2k2cfQXprm23Hjz5pfv10ZCBf2
bftgsPyyARsJQFlOi+POcSjBdv49qks/z6JkVrNWMIJB2OUhpnVxV/6KdGE8niDw
dejUXm37D47UgO+1rxuRbjY09q/hnUpY3VQUBIFf5rTafPbhu5Y7Z/5o6wdZxxwa
2j7ps8zxWsfidYtLWUsUpN/HkTa0oSkRm/szi+vvtn8NMH4hWa5ZswTEnxwJkPI2
tcG6WI9WPKGuB+2bNov2pnVwKfm9ngml+vBEukinKOsQuO033Zh30y1z4pUNjmMv
gseuHbIofAGC0Rl8ezZt5aqPu0WTTIVjRiqDGPP3xH4s2Gef12smHWMKVSL+BbUB
zxdcaLXDC7ZKEcx0/0R0natVxfnvTo9Wfux+4JVlBcwoP0Y0swPF5v4bo2HJa0FW
idAV5ifsyRzzw58YFeAlsg8/smtnMCLTBpqYg42uK8FuNiOEc4YBTg73OqN4qoLU
e/CqC67ZRzuUG788y8L1GYCvQdjrGsyyLuTsVaJAheDqQ0qTTb0LX8dRcycRqwur
npmRJVyozayzybzUvFgK4mugpWRIvxXZjy6w4zELNIJAbyZICEgqHASObqfEgEK4
kjybGWM1uw+aikmXb32fUfHFsWY6PPJlHz5lx5Gs95cHyg0l9OG8g0TkULBP7frm
azjhcP9H/AGQjlbBFoNr74jxCA/yj6BI9yN8URzPtKzuCmZ+FND6gjxQ5IG8wOKA
yKBe+w/BVgwlQ01IuHmpcOLz4Hyww/zHj8LEg1J/zZ07qvpFLop3uh5XHD419Muu
1rexFg85RBTCAVX0KvIrA4NoREAHXv63rJdUt14By44UReZiCzXE/FwHYDiZl02g
7GBMrfrYRQdGjktBNhZHG22f8pMqIW7VkxT1bvqgILqZt4RyeEAe5BJT6xtJnTVn
GPPAj8MaoLHGAIY3CFyJmm8q8EPn70bFqijDoNbuL4e/vbFR9+yEI92/ChuiyK+7
+JdFi3IP4esahYvDmN7AGOXk3R9H8mJQYzrZeZ0puwC2QP/Oe5uZx3CwGMk93lB1
D6vOWb8x/XNl7F57MzDozL5r1VgccdB2i/F2kmGAqDtQ51PE2va53XYQpIqFhqLl
sLgxfwF3EmgGtHDha4KE8RhPBmzrO1g1RGGBgi0WGa06RrS8S/IqDMvefRC+V6BQ
rCsw5NounF0OHBJ0Oh2On91M8HFV4IyE5HKR4Z9/V+p4GXhLLAs04f+2ZbXljEyU
5dHbrjKUL3WdV5gj/C5we3LiBXDH7daBp8Imo7MSoUNayT8R8JmASHzO1ZQgdqbJ
8GvY5oqhzyB2W/sEEYOBL1skt9j0q4G6kVfgmjHlHKFg5XdhJMH0c8XAN+C1pgdI
/rLAnVS5hx3RLpuGX2XGr4cqO8bKH5bsLmqmEG/2oL/nRF4eO2YIauE+tHalZl7V
eKvRGkPdZKvpRgP3iy3v2BqSL1jD4Y+BLeSpgsrXypwuF4H2iA/I/dx1eGbMT++i
GIBq9TrG5oFr+onCJQnAyEXAAM5jO3Wupv2WDfYlIVAj4GWtssbpGJN+LNdVDMzz
5IXBU7q9iCcAB1bESqeZWpfGZqEbd7+KCynvrPuUD3gKNufnK8uHyVqjs1MgLJ/w
YkDzMm+u5QTkn4Rn0H93M3Bygm8HqK5udnnBH0D4kVsztvj/A1q1XXyq9jYJmhxE
JKUCyl54HPZ2ZEZ+N7AIOpjpfPwzqI/DhQTJ8kItA78JRj6mVD1bAegNdlV4uHsE
BAjZDGf28cch4a7UqqsWhiDiX+cgHEo+eLKbLWgp2tJ5AR26mamZ0dlRVBlMMkk0
RKoOqBNTICQcIF8DQg1m95SfJCkvLtRbH1RDT5cMOu1k57ZKbM/jmlbh4eXFdwtB
/XsO/eZtRvwTlhZ4p1AeokPsXWZKtGZtZ9YD8FbTdNyOnbyCmVBQW+phtt9HyY0L
BQ1HWadSCqN+KVPAvkWYSA/XUf4SyOsHQu063alLxzHZuqC76utNB3pdDXtDZWMY
iCWnFdVTfUFvNHOYyGa2k4ThEgYqZ+CGIsjlPxzVH2MGuoTy/qylhnV73R/o/bbG
qWGNahi5dLjKuAatlvDDYwvLMNtYZb20RZOusa8seKXMVtRfajEAzCmN8+BFgbU5
oxls8Ubku/EnuLnx5oppV96tK4wYEIanFG2RLbUPX7TaAtn4b2vgJfvAuYacMXwx
dTkNWy5V4ZrZd4IW82H5OKY4iAGwGoy/0RQs6XpkOmEGmGqSF2FNcs6QQPENzsHe
O8KZR8f7agVSg49fVj/3ee3zfRPbhonG6lxwONhfYTwH05nFiFvKJCAS97g/H+4I
h1W7gHJJaOLj2vVF+vtQJe8EQUTjL1D9qbVr2FgHhnARiuOLG1B0BSr4UWSR4H+G
RCwrrzIbwU7Z5wQG5OZnaud7o4rm8+3YrhIe+c3p2w2pp6RksA76Hw6VNDgxFTpH
Y8rzJM5FXvs63UZpBGhgBQ/p5AgAMemgPyMv27LNUt7dlT9r9mAO/HhnZV+OfwH/
Ev4ytp/E66D/VtUkfmK+MgRkZiQDRvlsuLmz/cgk2wBWAVCZ/gdS0ozKdbKBGlz1
K87PGmM199JR+X7hVHTsA/LHlceMFq3DO0kA7VcP9XwNJCK0Az2/vuN/3xIs6+HY
HevkpxWbGzHLN+KgmQaQJ/Blp5EdF/LnKFNrbwEd7j1zGd70zFGavzIZ2vW6Qu05
PaeNtDN94qmmzz5AfggJkO1SiE65nXSrLg435awxIz2c5Fhl41krkLCdJ8nZxalu
NpwN0n+5EfJm9AGjQNDWMzkpXNynzxD5fkS5VS9wEUqF1Ele0wUyn8NOgCnBSDeh
Cd29axMDGMmk2I3CtWrT9fWNkpfmQ6O3EGzn4lSFxSfVSFQqH4z9QeNYt6u7oz0y
tWbQ+qetrijqVpsqQfDzU9JHw8ERgE0Bxjj6k2dpM2VHJLw+4gAExEDjuN2zBEhr
OXXmfK5eyObaBEBdjE8r1vHXHhEZzTC2y+eX3S98yGdBqlXQbHfcOlQiZDJqQojc
l1WikShuDKaNqe66OI6G64Ul9tk7VLUrNllv9GKwdo5e7OHAu9lY/dzvjGiQwh1M
OBI6wVYInSofLw1oygQxQUYhXm3hm9vsM3hEPtOFP7mFVay0U2+I7yYGM2he9Ip0
KapGhIyvZKl904c5IzChb+ngw7gd1OyiStVpxn6UzFWwm8Q/EAp17/lfsSr/Wt/6
g25zoT+ciRYSZtNgJTF5xA+QAPhF34QwdRo+NR1y66MxS9F0fYFyN5u/i5Vamqq2
SkLj9TfZU7/uA7nq/28n4LRgP1U8icThYOZaAAAgliu7fYhLK4c+F3ibI11/uPy+
jRysXovlcksxkzLFmaTVVOdRDvltGOZMpS6ejM6dz4dVbCRUw3beybBShm3Dbc7o
KY76baD10Fw+Ml/XIu37qLESW9PMcgDwwi+GULyH4qnWZouBAh2i9aizwqR9dnDA
ZbbxEiHeHpCyVEChgLqruQc2j2Y5OAyjKIMA3OJGlJqR18HNSFnOcaABKQHHs7ft
sIYaTqa7klB4OeiF0+skZZHheblOPUHYT9Fj1JLS+a1WFBKx5i44R50TY50MJSFo
KUXxuY0c+n8am3HmKJvKJG3HbOvD27lnSGXG/vSzihBLP/9KsJAudNF9JmxqCVXK
rfP0YGwqBdzHD7oz1MkHHPJuIRcwydBunSDyu6ZFMsk9/CurI/0GKkfejmQj5P1j
8O+RAGFLDzNX6bo5HmsLj4yghqlDzXnDbKoFXzMRxEITREXLQAtSwbt0I5P8skMp
i64MsXbg0ZPTTgfVBpofL+V+UOVp14tZhEakyBAUs21PiUP2RJVgyqL/X6YYd1SP
AtqAqWDhJGzlVKJzVsl8jAw0298h55Zsknqtak5xIj7D7ZlqqE1kgeZZ6kX9dmH4
m7MXZUmnPxsASMLH6NvvR8DxXNPuTPgpPtyT0fMNeGtCs3S6D3CebwuXamPKsaFL
GKqqC3sK4mSU8+EymcVyLK3cNvwqhgmqJo22SZ8X9Lc0p/kpX+9o1TSgcAh//luL
wgPbf1A9CxEcfv96zuFaCd6E2+bg9+PvJR/3R4142C0X8tcy+51ssk1/t4lBQZEf
ntT4NnPZLlM2ZMbhiWyLJvyq1JIICysf1J1dSZ91jCYWwCxaOxpXIp4BxkTGCN7l
8j/XWZUXU38/0KXoELORxUFloKPswESW0wywTb2czsUhiRu9tE8chk87OPc5H1Pq
vtHB4eLMpB5WsdTQj+26GPlAt2uuH4RMgOH4QhoNR0AD7GXG/yZt4HYDgvbOiPdF
Z36lc2iwFHaUOjIDlLh9uOI0KXpOCBpQXV3XxCkEZpqnMZvnD2PH+tQ6+HyjktkG
pH1YC9WLd41VJV6ADTPhN5lCRrynqyFINO0WD7eYe6/MxQsxmaoSMwkfKmfyGyiS
HwPNBE0qC/EqqyFh4ke4C08yXBkm880bR7dfu66J0KGL+UDds+MuRzPSikAKVaJR
6Zyzy6CFnoAsyI1yeicfsdxdVcxCWYSkLEGrMTRcgEaiiMfZAQ7/pEjqLlnIPR5+
7svEtk7WTZ6yakmNDB9pJT7hUVMTNlkn1AklcjBZLIHHo16KVCW+pht/u4sdowo8
7Wjc2/W61KdQb0FCLzXfsFy8X5WTEEdcAfMMExFOsQONJvq3oz/2DMVMKaal3lF0
0rQllCF2k4ZeIjR41F1u4mWl7gF4plVyeVHxq1Z14WUbSUBScPc17kQox5ev6/VH
NRe9Trl3JkL/RR0bEaJhh2aaAd6o/esZ0rXJvKtzHKJJZA2AAjr+ulOrwwDs9qse
PCXWg9DrB21jCO6WzlO+07gtcG/itCxAqylAvA9JmSzJ1od4GwYI7QK07mnZuZvx
t1vjaPiwKwYJ7AQQ61U6DNvcyq0Sn6wWEaRECD5Xq7XHwHIRdPjKDTZcTCJiX87L
mqPa+/sGPogVatuID0awoDFnbSFJ9ZcmECcMkScnUmEYOIsHxkM7yqwVBdd6sBXj
C22Yvito5PybqsV1pYagQV2+Zk066ky0wlUjEDRs3zHhQ5OJdb43Xbl0SGgp3GkK
ZH7nRZyV7LPywe02fPtivy6vnFCX33Fkq74eQNDK3v/VSx7u1FW/o1R5UwvfmsED
r62aU36ioWCp3iSlGs6sp7k7iHl9yvVyG709NCRke+nUULTixkmWDXDW9vs/oWyA
bNyiItr0ybwc44L+TAfHUjG/OlzW18lMFxKeIiWBIcswu87D48EHNriTbLjnd66s
4MFO2VCGAun/zlSXIIwb4Yn8qShDtu+7NbWoHSVhT5RgKpFAozNyarfxDOdDkRgA
MKWwAGXVpC78grwDZYNnaR3Y7j/MB7Po016G8bQReZElwMrsV5vvbrIwW5CUYi2W
9R69mc0c+bI+IGIGlksR3UVg7nAVF2oxeY3PY1sUUz6ElD4TxlDUdSUfIZUn21wK
tRTAnSp16eqxdFfGmrRVjqCDWs/ITx5jdW+m0NfMcWLotLx6b51xJyKToj0LhPhY
GXKNgA4IQpGRFw2+l7KeprAqdZEd8UwymqFZlNmLOOX11esHuCywoMkFY37/+y+G
w/ZRAykytvqRODEA1//kRv4dcMyVDjqC5r3ttsdURyK2/bHlwuKCLhyjqMOBt96Y
cY5l2ObyZd+3CefzoVBHKxBhogYwpOEK1KSlETy75bPcQQgC9GP3MaV2/o3lbbTN
po4WbedaFC7MxtHkPjNLx6TGbwMIJ3zJNqB0eWxt6Rtc1nxrCs40/UWjm48R/BcZ
sw9sq9sVUWzDvqoLQetVPtbL/ETK5FwlRvrQpThRnouX35sB8A3lh6pjcNFb5mBT
GVLEEkDSlNWfVdgqD7PuwoLhYypdvVnbRJp2Jc74VFSwLO3lXlFmMW1BF+OFVas9
A418sNvZYkORCTOMadM72XsgwWQOR4V4Hg4sAKwtFaLZON4PhfXP8qjh5LvOR5vs
5FHCUYfTJRO7OBoc0/Fe2IY3EDaPnxI83lgEbkv4RRBM1csHwDKuuq/+G8BOHytd
6tQOxzzlcqE5y9xbSZt0VoCWCEunoMLkrzB5HJWeTDfuQuYtiEfeeAJe9L6/FGT1
rUalxR3Gn1zJevvFKOSoNdx3m8If7T4U4JrCkNTt5zTS95k496nzbS9/NI8lhvcD
DhkdbYqX46eYi2kxQeJg9IJ8n4wHDPJDdB1IZMoH0QN9y7CpGnpwxlSodcWjiXNM
/VYJoDfXFt4v+EKdmyXknkmXLQNDgd0k3a13IgX/+e3NGd9WW/dMfXcVuivzCpPx
CXh/0gYkOnS+EMUqpRdUEOVFCR+h55cxYb5PysLCieceC4xoEyvpd0cR+WCc8bNh
cyLcuXOUhTXsaMdqpqf81ZTZf7gg5T8BW3/MC8HATm+CxpDlZSjWo1440hlLCm7G
jEygp8c/6duEmX1XH70GuuFKSQImP0MObHLsBSFnFUBq9vOMf5e8mg+6J3OTWoKn
CI/IIm868Nk9j/eV2NcMOEjHE3PKeWNv3UJYAe5087jVOy+hkvHk/zeKcEuAz30M
3uSlAvaurRhKm781dN11HMfBlebXfsKlooGYTH6+6X6Pzu0dO+4qi+k7Y1gIXfb0
EWpzSjuSnD3RVSyj4xcKUGQDCYWYMaMxTAfToSB+H06IIojBE9jAJUKZb3ZM+nBc
K3jLMJPF2btR1U2B14kl7bGbp8BzRtUiGeuu1nB5rkp+f7H06s1ZIvMUUevcrRmL
V5Nx6RDOwtLcZIbY9+WdX5LZtwf6lh5yiF0acBKgWdH/sHwS54zLEpDfTQETSEBQ
aVG9+ELf5kjlbTHxC4eiviwUt/mLGOVc8bZP2iU+6rI4wQ7vthxVS9azu6+wqNhi
w9gd68hKmTGc/FHArEk4+JbQQtwLPL8AYmWtv8rcYbNwJWIHVcQ1pThpBtESFNlk
47jwvHaqkh2uu22b9IqQM9THHHJowIbd8f7PKY0gPQni1RdNkuoes3u5mjwzNHzp
YVbBGTpgVuSHg39srXZDCX/lz3qvgiGRfq9QdrAUqrbJ8sen90vkNlJAsRMxt28I
OIk88hYpcu7KoN7NyqsXx3Q+FcXH+ll/xBWmJxhRzVCIT2qp2WR3ldwmwnW/z8S7
WZ/YxZpjsM+Chr7GO3qSdT8P2kbjzOd7fLVvMlIG8WZttZe9KZZP8hwgNcdyyWmT
80u+2AGuEaPVMxtGu9DFMTUjzqk8P3ph+yoiHoOSMcQUDBHo/NvLXFoRN7+nKs8x
YU8IPnDFdfsovvnlhO5iDbKpXko8w6qZOQF+qso8QZRLsOR/3cxcIZjP86DlmVRH
nCdPHhAriyx7x0VEMkGbMDIctSNAeMM+a3HRxQYZj3owBzbceqiDIk01VDdf07CT
rSE7TlEscHqUh3fx5vkAeJDFE7Q0HJnCR13Ak9K/TmwMcnQf2bMiSGgpKdl57oK1
Ibvu372PukJjeggCMPZskqmgb+a+zNScdUdcnAQZI39hwX8lwUSkPnuJhDYTCBi8
w8jvuM6yUcXH+HnLSDzPY9KC58h7tI5sPvKU7S9v8pTv37l1qn4Vtx5MWRr4PDEy
DqG9/LFeDwZvLsFCgkULPc8GH5QaPFKWXTH35QmIM3RapG8yTB8eMQzbYNV7vR6K
EE/6OFeVyVLzVJBZqe0wuvxxXgCwEsFnmeMsWCbLKKN3NqHUxKSbtkl8uvG/Uhb8
q95x9thUqKUnp68PRbs8Iv6YFTxOwqtmSksVm89/J0xAP9aBnN/8tRaoX0xnf9y+
BqAV+yVRWVDBcAWyG8cGJP9BSkK5WdB7vin8jqUvlFHtFvEeqmqeCKFManp+GC1O
IlnMcDg9j6XJ97PQXLsh1Jd1hS2DSk5OIdjQyWgtpyM4KzQr1X5aCoKdXwndFwoT
dH2EQSm5c8rMaE/PZHrXjyQ0ywae+GgPHyPNaayB80RyeRsfqC9FMuua7zdnd1LG
B584PMvtnstc0LdFICUY/x1WzvcnQrtCfRh6yGPaDiBGCqFQ+a3qBR8Vw77oDPUE
nAUhA/1XLk1R+UOlD2f/REZQixX6+XsEdMysKt+yDLd3+Lt7jzQaqR9JNNlc9LP0
8oLAtPloety9uOfOO45r2UjFuA0WfX5rsw7619mxD4Bmuk10GqA1Fz9tz2wL3BAC
nZ1RJ9cC/JTKuKEXf1I2MzjfhPJ7dW1fK2fDioCi7KZ7IiFO54/9J8Z9G/ACnUAN
NbjgklszWS7sutUVc0DTV8nz34pme5aMSlX6q/dnDglwvz8nhgOLMwJ+40HlTi+5
XAp6oNWz9W0JjLyJ8SgmvwZB206K+GvY8iug/a0ioa18/p4NWGiN+BD4dwc6qCyt
8njhIj4LwCa+W51rzFW0z12AkZkSgSKiBDbMu0e+hTNBblxoaeiLJZjxe4Ec5CMf
RK70T79fyy7iExZUEjEISopePc6NxpdIkUFqWuUX1GbXbEe4I31qafFS/Olndc6y
kO0uha8kuXPACy/Wcvk6CpXfVLo+0mL+Q4+3BbxLjS7C/3gXQkYM4Ie0iyMXyq6e
1xbfl7tvlGdqv0GL7NjrrxX8vyqSncN5o73KgNuBmQI+tnG7ktMBbM32E0A2sVeW
Bm3QVGH/eT3PM5BBrDlkGL7R8dq7NByUfhfwC3zC//NAmSqfysRmH9Lsm7hkX0X3
QInnzuOUY5MiNE/JDu1OJHBOq3x7p1efEc1bRa6aETmxGHSINnVB/+/uCbFvUZ+C
LpWG5xooBw/eBjLUnzD7FlqGbk61PAxgOby4iYwrP4NwjCQ1l6xk7M/PsjenWQqD
K/4JwVNuNOFY7MXqJ3eZNjo4KN2tqnlMkS9swY8y6rw8bOBeH9RKGLXSaCAnOPnE
jDB3WFyiKze31EDwgYHdV3Max9LUQhWJK84yd4MmugDV5b25x9FPI2crt1+7au2t
79GNkdhZs8TnuTVxsCev/g1SQW+CKCx34u2/RltBa9ffpHLQ6BzJ8TkmBdxQJnA2
7U33mL5+02qKwi3Yc9IAmOpiZ0Vx4QTxdJXvhO7Ln7dQDzhaqH8FdP2ta8jAyy3v
qHRFg6pJ6+wXLahT0un5SVY8DFy/JMpDm876nJk8Dowa3rcpNMAWLamhkm4TGIqZ
hafdU9A3hTCJT6lY8Sd5i+PJ+46ZIVWZvlD/i5KS0eVX78oyHJJNTFV+Wraz1UYv
I4HcikuOUmxNHtfmNhr67nqCTqS7uD3+0+93zrSyj2CNlDYq1wQZRhaLWFe2iSKI
zD4nxS1fNzJmDn4e13a0CR2I0ioEQ6z7MEqbnfaUMGn7bQR1IGjUGXUjywOui/jn
ZlgO6dG9s6MNWRr9GMCFS4SENq8UQZna8LsGtUhQFp9ZkuVz7TehHpYBm/OQ1aRQ
hqgLVPPzM2HnnQ9EECmnPto7HuRYcDDqVZpDsLL4V/WcSloj0TvVZduY7nX9XSNu
tRUSzqZM8CHGOAh0285aJr0auveAtmdwzvQ3OEwQ1f1u+EIPcNRuS/jUGrQJuq0q
OOVrKyap9MNiHurv1eHZ/x9ETM4uCVs3xnrtpT/FeCAefRD6zcCS15Y1yD9K3ILG
/AsHzVLXxaQ7GA7mgLuKgfeOx3XIl81BmRNNtwjkrDgB5qgBEZfcNEClN8mxaN00
3pZv5Mp3j0f8jYHU8FYK/jgYr4vb3I9qa9VTGDZA8r1rnp6W7MTlxGqSrz88k2Qp
5Y0Gs4LF7XEEzADXgICzVpjC46xy/qkjOV11XE4qH+K7R6pQfG/HPloNOjWuARaQ
8/XqIl4cvZzJqfdffjEAszBV/DegacD7ZnGg/39FfV2KZcnm5uVcl7Iof0dJi2F3
oUGNjE1FhSAb6JsxyDWNsLiquVNf0eVrZCpX5znxSg0z3eNSVHYb2mnrkN8KGZdP
ZEheua6k1lBBwyRL+d2PBWDtxi6o+EL+lAYXHKgJqWFjo3dg/iF1ED+sFKKp8oGp
Y8DE0Ei3l0X1x924UylgPvS2HvSD9m5PjpTK+CFYVRa0r+l8AI9JVG8RS+Zu9L60
oFg+BJu6jCA2dICvfxA80mDIPunt1ItCbOmWAJ64BX7eN6uN+2zE95F43lts2XwU
RtNm4pphVtz+b4q+T/RZOMq+EplDBdByYKu12Ux6Fj/RP/xuPVGuVPpeNCF7JWtF
lz4VVMSb0eVw9nKTlWg0+6v5hDYgFSGB9JPpjLOVdJLkqPSgx0kyNGIur+IW5lLO
7MvZCk3oOTqkJAzsVYguX5sBPR5JSG4MWOIgQDaADECvyesb/IPLTETGzmz46qgn
9wJAl7P9Z64AI61qRzCqGu2KDcZNYqIwgiMWj2CFGJTa4gkE2hVn4Uf2Flxwk7NG
fBfCTrsTBhWiV2hQ52DOaeVlPQbJt+wtgmk8+vaK0EReh5L14eoZo/ZqFrX15bpm
ib+NPhwl0nua5xY54owHoehq0f5hwmXeyQHgXXLnEcASMXGJkrIwwIkivZd/ZXN0
ntDmg7OLTqR+1BEFyY1ysaCYwx6EK23KbYII4dzNCUterdhaMx6AXm/rG2D2mwEp
Tex5He3SKeJbSbv+2HzUJqT3B1rBYNqJfrL6dt5BPgBE4HDsjnUWdKvTdQGsodaZ
g025meZyiCdPOX2uC0ibPLCZ4T41TqkTYIpALe4+3Fl8mxP+CENXTZ1NQ0fXWjAD
pFNLmTjnm+H+Rri9083R75DBo9KEJbipTHo+25i/4m3Sa0KEKZb4toLUlrhXBfWt
UjwhNYeRx3xT3Coln+XerinFwzmSfsWBl79q9IlziPpaj78CKaO5rsVomVzhkpCf
avxxoq0q0zB72KHZ7GXrAgPWF9a9RDWFFFFQWci57QuISog8RAaVC4YXi4AGAZNJ
oaE3i1gF47TPZV+0CN1U6APvvfX2c3yXGqnW0lqbsX87Xq3dBkqBvwjpAj/DxJRd
T9kPQSuUM3tTWb7EGkqjRT/DgnIlD8UvlTPV1kdL+SP0LWq4r4pF1rTEQknaUvfq
8Bx/r0tFTu9m2lJ2tFmqv+yoyv1aQNC0mBeGUDxqdJIj1+3u12E99z0vvRZK+1My
2+FdKeOEmiT5ta40+AW68TuFAbzgDi1Ui/f81zamivrP6Ite6AlAO6nnwpvy/tkX
NGOEfoPHJYFlG1c3h1ntwnIHB0ZxUsABTGvJSr97Dp1ibMC0nLcfgQKmBPFrXqnI
BOKGlPLbBEg9mt9Vmw5ItWvtQRydwcu9u8wAbyzYOg5g15PiqNCxTwBHNTNjCoZq
yDAU7CSPzJyyiBT7RH0yQeamGO3tyhbsfVmpkRc/Ub+rT17AU0kF0nm1SfpJuMH/
616/xVUMe1UUAyjdnHl62rgsFfyAihFkJOnYUKx1gAe8sxm4NJQW8FuewnPbMs8c
fAsOtLoFCuZsNQ9xl7XSm/2dG8nFEjiRZOiNhJld/jl86qa6ggExw+xroia1KMGN
kDrUNpVtfzmpXNz7O3FG+/pFhdG+9ojYo0HY58tg8CDiS5Ba/k4F4Y5KYeDOc7Vj
sdnT8kNUXRLZWNllFb4aMl1JP6HpMgjNb8XUIoRkynYwEuRS3+ahMTLRogqM+Fhe
U8OPo1fMYO2H12wfejJJoK8y0WMMVqKMa74pSUFmbj0UP6UlEgdZxkTX8l7y9hMF
v2BG3VbEGMTmk0nT8iTwB4qB9aFSSr0bhuMVUB9CZqGa+63rPKztPnbABoq8aQly
Emcof4bYCTXt5sIidnB3ArJamuLETBr6lTJEW7iat9r5E4cTXChmFxVivtekMZJ5
z/Rz38QRZL25j1eJzjZSp7k3AvK0vSOtEldZo3WwoGIxH2Nvp4jq6i2Y7bjPRE6d
fDYo4EKgYT94IABt+LiyF+Zcd8jL7wyXxjD7wV3QYy/fPW0eTJaAe6ysB3g6EDxI
J4FBAKj6e+Lf5WeMAwHu2jLHF8GKOgNv5rciMaa0Fswzt2sbn4Eu2/Sig0eSo4+2
gdx0KcIwhwsZx9IBoldoDbpdn1s117oPidzEnflfNnNDVdUJZobikYC9ro3MmMCM
hMBQeY9Zd4DvPZWM/hMnpatoj2iBIoIoa8yKNMifjWqF3IrWzlmm21iz7jN8U/Lz
FXRfYFVPHqKkr7x1ui0jV/4gkuiseW2vU1QK4Qta2zRvhgyGAjdR0NHno+E075jU
CV38l9pr4G+QADC8eaTlXeUR2zmr/QjUZGwDnsUvHorzGAXwvKew1gKs75wkbGEZ
7TQLAtrTtkhuLNvqqOa6gLrRGZye08CEDrVDG/Y/OxgZTxLoHU+KgQa+zGxH6E+D
W5Ly3vNHimNtjZrzyg5fET8NiLUlakKHfaKEHhaWxSKSXG1C8+6FKGTsVuKTmzar
bL3vuPIoHAf4W2K1FRJiI0EMwVm6a8tFC0H4ZiYfCk9EU+Js1EQFDQBy1m0+E6Ge
iHslpQua4+XUHpsFJapdwoeVPvaqvmYzN+128kX/BTulYpISmTBp8mFpHpHXatXM
xvR0xQTFeyk+ZC2qeQRIpF2drt0Yo4ICfmkhfyTVio7N7cXvJjfXmXRkUW4+3egF
O0/EojKmhYVoVg22yawWDV35B1D0cpliYzUXruyRTjW/wcNkzTFziFR1Vwo9MVC3
gmZol169AgN4lwAd0M+KTJX0LDvybNQ0GemseaKTRewt4/HKOd3sAkt/baJwLGNt
IVK4DAadZ/VgTaxzUuAbTpM8N3pVaWy4kc0xgZGmhD8kQ0SiRDIfy5zn2vvB4cpN
fcJPkbDz68qm789JCoO1+NV98xGxRi9HL5SEamSMi/0qMd6h6tmbTgruvDTW23L1
TYGgr0RiyC1PJ06G6zCMhOUBC3wYm5WYp4kMtE0GFQJg7eYmFbRJCKF8+/vnB2SR
ghBB9jV+YJakl0EjttHNBEzNh0ySnZoPFYD8JoHviIhuPqUMRLiJmULdNfN+n60M
ao/hWibp/f4SqhZEAFNsS3nmAeVV3yz2z85iaIbps8LBIJQGbP+QlVKB6OFPIQwM
9W0znMcibcp51DX/8vQ1phIJMS4Px7KHalQRgzjy6/xEHnNPOLH8TLBpaac09fiF
zLepS/MavU73EjgzkgG9n5/rE6Toh4UVs46xvDCkbzo4aiIorhuY77RXZGh0X53A
6laJByyvq3GX8tYhIXDyfXemEfiL6bZ1ZHr/DZODyBc/Vy5a57bZcsuu5ztMbG/1
wvzidy6WqfxWFbBTttN2GJ4USJ3EEiR4Yk0D1nrOOpCTkN2zbsfSsOvc4ocS8YCY
/yHcppR3MDOpJTy2pa9pEg+wFIk6Hzh03qw4Gl0vf0fWkc/Pm6dtP5Emi3+StjJ4
ZLMO5JlLFvjQSTry63NVDIUe52Fm6g5PLtG9pPxcbj105mHadVnXSLxD0/kifNA+
OwYyAZ2A9BthSaMkYJcen20lrUbBaC2fYw1zvRwtUi35jF0o9UNjEl8ZnlL5+ua+
KtwObSuxMpujHfPr5q8XZj5Mhd2B3ME1HwYb9ZB8IM3lPWPCJ9UqQV2whFaQYdLx
8vBj25ni8gyPI/S8QZ26fLJ5RdhT9nwytJx9aDs6lti6m8PI9dND1Y4r9WkYzbsH
0gcRdB31sZYbsr//4dpoFdyVYANFskaNW2yhjDIzHLDXJ4IkDvTZgMgnorXIw/qE
zKyQLVOeu/KPRk/6MNnq51iafxvVqJ4k6gh7YKdMxzrCZ6v08w96af6fQYUKd3TO
CZBfnYrMRnp2p3GQDWNAvV6WSpmRK8bC6VHKW0+1aaMIzfSrtxnj3Ic5IVlJzwvZ
HebG6CmPV9sHrWBtuMtUI6Tx6AS18zsuiT/h5mpMt5Tl3wxNq3hOB5Rxv2StCjrR
fe6eOLASb2+dQJhDGNMjIPC8UuR0emmjv6bUoBXyvH32lS0D4TfYaooiPeNJkH/y
fFCZsUk0nnF5fUUikjTvMBHKifQIMP1QRdPjqOd7lEcdld8aHjyaf3CKoU0H/vwP
YW2yh8tB8XK2CRIAmo/XkdUN/E0T/EfA/EaZ07VL8bs/egl1g07QRzoCbWEwBUSa
MDhQuc2kNzEfv7PsjMIYz/vgsXjmGGnTGCXtiS0KPLGT5DZYBeDyFIblhw+1Dr+i
OOggjjnIWdFmWs7QZV34WHczd6OEi9vcRCKfGLvdK2DdmlZ+rhfQnO1djjBial9W
+zQg6YBzRMasjDVGW6DP1jQNEHrCBtBx9qH0rTmrBrKOVHF73pswRM5fx1qN+8td
Tv/L0RhU7dMNccoqbbEFpafPLG1sJShCrURl7nePdcBDBoR2MSJp0H2B+mmouva8
a6R5OwP7gfDHSj3sKrt7yVuZpjJ0Pm/bXJ3ljKgAjlmh6dsd73TEV/uZQaUcQ452
/hkIl0sfXUunkesFEIvqpVrVzTT8W98vIXsode1W8732SVczOJDfKKy5/ylOk8RD
ldvK+PctjsPbn2GLjm6uR0w6S/bBY3/rJu+WsHqJ6pwklieVhNn7AEj8wJPjHBWQ
XiWBxd2cHARFcXOdxHCRT9ge2IFzJrPgvCEYErdfqM8sAlCdmfiEhQ+/Z1p5iydM
7y5IMTo1pvgIj/8FAJWLPHLNjYySax6ANTjr3LlKC87eo5nlZ2L4W4nXtMLOdbCj
jChyWSzZPftpClkawuVpm8MBDxcK+GfJNpxevnpx2sctISoUnzBe4NHC0CI57zhm
h9I7POL96JB1b8EZabDkHjJs8eOUs6j2jO5GX2Mn875q9vj3j36EB+TBA2SoeUl9
FRZ6zexb8376yEcCmFCWj1uu5lR0FSL7N3FzmxImfhWEmfc281a7cxvJj8EuChuc
7aQqMgIPFd2J38v4hRlj1av8/gvWEyv+MbjyqzyRlakJWxNXS2Mkr1LvYHy+E4ua
+hEPWdNmi39SB1Mut9Hpg7LrZtoM/1h9Foebt7WjXmMlOSLuZ3jGbqDlMTGSYEPC
GS/iyal0EqBFKhCcTaS2CrrIx4xIxtFNChNuX7qnRFHRujMUgC3GS/R8mf5z1bQs
YLDawhsVDBwjXGUhadzPALbiYUrZSiT1DwP0tSnYGvcraqv9paUByQFRbUAARgVL
bpovmZVRUxLy3WXK9y/DvCLA4KL/XWhFL1eWIFW0mnHRojqoyGxcQkIB0Ds7d89g
1BmLRmfDxlkiow0XJGmdKJFc5KUK/LKsrt9VNlS/xQZwXUXCsQv2SDsHkxVxovIi
MrlyZapXlknebaKOKva1GiteR1wWczWR66MoM2EV3FKNyQl5wDQa4SLl/adNMDHJ
B1ZFO3UT0mzgSS7OYjL97xg/itVU19njSZ9CQssRucNFtOQRBrBVaCMJAeyL1p2L
SuSWjJPaF79u+TPbcarH58EcOjeYwgLlvjMnpZ9Ef9zfJtw5k1PDIMSLvJLaf4mD
lvho3jEtkGqRv/a8bVE4oeTTcxFlRET3jo9J2FE/sx38cAg6OKXE3VSyytg8PV9F
0uNeWPw5KF9IsImDEYq87qgN3soLS7SgEU/oHgxG/9SZxJfE0fxADnSQpYXTJ+Kb
bZWn/Yl0Ts8kkJzLHQB6u92CCQfjXeBPN5WVn2QmOnmD0bKRMUU16OnWBxVylhkF
A8sc0u6YG62M8M9CF1sBUX+63nCF9G1WbDA7botybyvKnAwM14IxWz3nwOHYmGVa
YIO7UiyJaUgLaJDvHAO0gEIUKZVuOA79K74XZoXr/hO9ebzs1nppNtnstK8yaHAY
lCgvLgMnNuN21UOOQ5vmaCDnFzSywP9I+25WOYkIRiy46jj+5nwOYGX9VvyQKWSF
UAvL3qYErzjrkJJwP6g5h5XH5JGNrFWnmttZb8Px/iWQD6C0VPbn9L987XBHglIs
3/6vzohbtESDXr867eCC2PKZ2LIN19DErS/kPmIvyB+bKlW7wGV//42zoKFuj/MZ
xGKpfD3Gna3wAjFz030s0EvPOyvxM/eLa1QIiGrw6x23d1rLotzFW99p5qmCnHZ7
aEltHkzD6rkAAGUmmIUstE12pn4YY4QG1Z3FVTaBjBD9TGwyYypXKHxDEm7/hoBi
alqDH89pRiqeH5vrfw6kxeKJiOEq7PXpFsvp8nmcWjPuXuwXdWdgrweE8fBJVRLm
lei60I+Pc7ChqgcinUSsqOT7LpfmBOTkEZkw50mNjAQnjqUCt11Z1ktaZv3qtV55
zII3vO2Vav18cJVWCDsSSihEORhdttv8ykYmli5mXGc9q5Lsidc06cwy5Vw2Y7z3
EAi6ilnpHFfL8bwhui2y/fOnO6kMMq8U7shjU9S3OGLa7Us+AlPGuyZa2fi81MsX
0FcbD4AeqfbQloPoe0zzD2Im+1OPAR95u8Lp86D3csWGqheQ1Vv2OpguVF7jCXh7
xmPU6FAXu2iGoYMFajCGAjVE2+7Ndw3pOnvRfV9aCDnkVBZyZHUaDM8YwoxiqUnE
664CSB/N8V9ukzxNXmScM/Mlmq9sALgZqrhW0yNL53pzFijsJue07EWeujaSR4gy
bf4W5XV07zUWwnOjQxrNm40UKLl5GgV/QB3bSRKOzIHHwq10vNOJzclHEytFelHc
2rlOUhTK2/4uthbj0AA0K+r2L3Ncy9LAOysaBxoHQEnd1hPRyWCCTSJOUv5i5ylB
1XDowmO8WjTGxSUq27vP+LUE7oPF3v/ywKfN8H45hfthuiuLWTEKkC1Al/a4Na9i
S8XALitTiYx1g9qEq/6vzvAgp3uuyy3CsjqWpJd+49reLJRY5SMuy1qS+++rWnAF
4v9r4d6s3ivfk9qaMrq6xKA5/qQi3TPC5mKbTyuZQ6mCv0z0bMwX84cPakfls8QR
rY/5mrAiOnSIR0ukysu9IbkYEjl6iAKPer4OgeAXA5ye77Xotl6Ry5mmWEVD7HX8
V/+GlNZE2p5zdE6YM7VSahJBOR1LF/n5ewXVBFK7ee/ceN6a4VvQYXOTYob3/mST
TOHLQ1ApPP3W7oFM5Y4Uu5SOZiRSoccqGQiZ5UQhKQb26FQDwHUt5+j/r+PsxAIu
fIJ72TC1PuaZl7BITCjZzSH7zFPIjSXkOSCsJtvCEFCJd5qw8GoNynQzESmdXld7
Hw0SnqGVeAdGpX65SpdNnQwRqd4iAf6auO0Y3EQZN2Bj83S23MCjNdpnmEjnFqIz
McwXea6tXJvjQvj4hq3HCiXwPqDYpds3ssV3YNj97nyicxT9pVtF5Eo/P12palzR
P0RZDzOhmeQzG8Si/YDPwE2HbeYZuT41Hfr+jkhejAvorKlXWO0s0cUTrSIt4IMR
ryRexNOKYghOuu0STKkyWO7xXysSUKENHg+IcaO7ZMGWxUHwfy7w5pjWUf7FbdgQ
H2XpE5NjSuw4qo+PoeuSyyDaulj/O+OYxdbvbqPnZsT749QaDrI1RGwEFFwrOlj2
/QPlj5T94ds7q2gT7VmJJ0GDZJPvqWSAWy6Iq5A0gIIIN04/QREQJdEFkxxmjSJX
deTAZiqUGpjs86ewIdyb2j1gpO2QFWEmjb6UT0srJRVJoVotbcqJsAkwkusvnti/
2KEK6rqbKohxR6zce6U04ee/25dhrRMA4wvFZFCBzJHSxKNmP6u1t37xOmdy4/Im
Z6KqLXM2GKkegwnz8u1tgoST1Iv67Qd8wW6vNRsuDp/Sz6MJKaCAbDX0pSKQzrTa
u9e3pDVlrKCqWEmXGbUjMURuiZnek14PiihNRSvT4b6Ex63kBjrT10HXab/YSaIO
DYl7YV7lLWB+m9b4qQt4zH0dckshVtOWPYJ6NAaNZsVTGkCnuMn96HgQRdPEk8oT
6KYONr0yYYTEG5rYHbEKTk5X8tXWkyv5C3fF9vWH2EgsxCv+sAUnqrYgfRrsEAaP
ajllVG4Gr1smGkw0DWmDVfhupznUW9k0xxqgWKSLrNPFQINNqkETODtvlL2kEmvQ
U+zkr8zQM05/XLYB8n9jdROLefUgZRrAR4IB3aB9O3EG80BwNZn11srZkWvtTuoL
Wn5Ib5ExDezavFsMVXxKPCooTQTvgvreTfj37NtO2FghQymJCNM+k4C3pcO2K3md
8XfC3AcskT7bsjgJEjxgSn3x0l6H+KhjcdGBkIGuI3mv/D/s2FJnzost7kRkcaph
sdqcfoCjZe4/Fr48T/w4n4d1jj0EjNnq0EXEAsfkOtLklIsVmWfRZBaM9JXCOn1z
p7tLop9mEKD1TdV/fWvhKXR0ACZUYUpjF5+10bo1AUZEO2V9xLMVbNs++yj5xG8a
MQd1ipmIR97E+rwwOV7YsF4Y4CYDwDTV4tygTVHqgTHB/ykCu79sR1h6WwJnJPxD
hKV5rcNtZYP0Z1ev7PNZFE9wAQtdrkDxGcHSZcTXSgnEzOeMIYHlHyJD5O1Q2BQW
dGL8zhG2gd6Y+qlHZnroF4qPBYgnM272Dp0JzCPC69uxAKh8SnvoKUbRc9+XpdWp
7WiUWfnX8eWze7T9Gy5Cf3bHkC5o4kMtmXyUj5NQ+V/c6c0QCgnx1y0aQR081VK6
0ew7UD7RE0PZKZpXcradFadjL24Wb9J6S53D5yOE264PgrHYV75S+fxst17WQaW5
Q/acAhx/gc6Gor+gxi2UOxWSMVjxCRkWq05sxRFrgMBvkFUrzd1dPLoY9k7sjmbx
pHYkAsvaqr6iNxxwFDp7GVR0Pm+9wGU3VDV4PAmWiQTDY3uz82mDuVsTZt5MWD/L
CAD9zfJ5W4jSGMuAa5C67WKezSTFL/2SHj0Vb4/ubL8bfMBe37rCXrbME8cclZXK
iZZr/okdKVqu3PGWJNG3Nq7wr9HPHigpUuRdWd9dwtHZvxpFGo/eiyaQkiduoq7n
RJQz5aOwyj+aViCkbUmtqgUf0AhHSx32+p+8fL0LJiiDvfVp/OifQVBRFHPhzLr4
PavTYI9GSSUL51XYfMF09rfsFKjSdQXq3cT8fdDQKT+53TDo/zYbuwujZTmJHYKR
T9WV1jINnBoGD2Hh59oienWDTceWvUWSRwmgpv9pmJT6rYmnypocFIEhsqZQNl4G
LM5yZIEswi9/sZpAsrkVaDv6UuaXgzoNmFgmJh1Z0w5oQCglNImLqAL6X6Yng19O
d2GMGR4N7sxUMt89bVcxnzUVVKHSRW5qAfy7hZwV9q+X65V9inivTh+3zHt6U1XW
j8gXaDmo0nE6ezjFspiUumpvIxzMlzVlQ4mnS4Bl7VPqisYxSwEGgiBn1Le1shCk
3XB8MDdOxJW/hsmDRJ9A/ojuwznl/vouBtHudNcd8iGCkPvlTqSh3hd/eTajBO9q
5fc8VjA3S98HmVXD4zgqFQPIR+3pvW39Gqyxk5I46VjJoeJlTGNZXMm4rAgCem+S
yz1F19g28XeYLpQnzA1pqs7nlvVL2gW9PsxAl2ECbYRiTjVT864hO/3oLC8EiDP0
Pj2g7TMlz8STvQpeVb0+SmfqzYhjSw4ToYohWg3dg4tWWQh3ISeS3fg/oFlMVhpn
f+FdQDuJoOKJ40WwoNNm3p3vY0wh5cNEda2xkrHJTEuK/XHqm5ezdQCJPTCJnX5S
Y71Nqq9oLRpB3+k0V0tOj43TyE9BhMOPZ2uCDPg8VOEON8qR4ywVCtwlYZmykqG7
Ii/Y6T9VgEHlxcP8KIBcvUz6ubedh6Xj+jNwzLkRelXYcJCd5hReednCY8L84Rgc
F3kTTz/kykiulxhwCTLjLSqKRnCL6cqM6aQ4a+NQ9vAmLMIwLef2QA1Crq/yakAl
X3ZsFo+f6auVvqQmhgFs33rl+RPmCozEm64h2ndaDbg9nr2Zs/I1vKgEHU67YsJL
DbkQaSIbM39Akmrznqqzqkw5d+7hdSQ0VKzFpxVl7RrRdow10U5rg1w2kn+Zkz7S
YWyXJTJtNG1WnL2n1UyWn1dJewnoHtS6eH3nOpUbAfTj5lOmNu9REVf4otquUYbq
CW+UjeC4VBMPy8hnwFi8LyZLENyxpIScLSIOr6s5c0+MwP1baE4l87hPJg4yC8pT
kZo00gUi4q8y/uor4zTstCL6acrhGmTucyrAnAcTjFrgPMyB+YSNlx5pUbgAGapq
NnnMTh/lg4EjlfOPsh2frAXl8XjetKCr3Xcvw8ZRkY3JuKscwYQOEXi6CxHy+PKP
XPHCuP4EOEofeZMdIXuNCn0ryrhWLcjSjucF1WYxjavdzrWbffoVacWWKlw413xT
AcKx/MwZb/BS4L1Qqc53bODEKKCSw2XOaOBH+wvUCI+KaSq/qcET0Bwx7INt8pIq
eOTx06s6fo/SqRc7sMNSJIlGkG3oGBVFpi3fDTOvOO7XeB52HTtt7FAmSSRXOt/9
A+4EE5vBm0/STFl90vv/B2ImiLx/jj5eovVckJHea44vQBqobHNoAZguLGPtD+H3
eXPdZyq018rMmzZ2qS/1Kj2B3eqtsjHKXmiw3c0pdzw+shjA8nQBHXp7AUsfHuco
HZTu3kLIsJYChkBWJw1pz8jgYVfWysTAtMH0r9fBMQl+PKMOgFJDL7UZI7qiRgiJ
BemQ8mwp4ipi8i+/Iw5d9uoGxn70zL4fn3ELKsFZPOhgCnMoHVQklbFdAhROM0g/
kxezfONPuuELDxH2fcx/nGmXUo1Z2J5MJ9AM70qFGr5okW27WJL/EGdB5G20/e7K
bctA89lsy+dy7oujLaOu7pdcNCzGZSTP4OCJrZa+Mhw8XXXM3r6+r5pllGwp/Nin
lzLr84vyxW1ho+LI/BawlREeUkvB3AP1LHKsn8wVOMNnB7QihAUW0yWINJMPPnbw
42qC/QLAb9sE8TBfl7xxNecJLz6+V4ECDatI+puqnUdgek4BdjFn4LXjNxfcu5cG
fWsdF43ipTGuggGQPb3xhpTMTsHP6Bs5d3gzb1tVxQ4Knlr+2mobaycmc1ZajlGd
5UoJeVBIsL2QLmjMRQZF8Y/sU4z/DK2HtRTKq6YeAVq6T0iV8MbaKI61+ZOnYZ1H
O24kkix2PIhuiIwjwokUIHIooHMih10q7eKhEfSZXnNqRymgQyNh7ApMArSFlR26
mas6b33fEOUW+Qv1na1fhHZ3yiN/Gnv1w+ORautiVD7LQjemOgFcVjPsfpeOnvaN
qHakI0GgyEC1E8Z+RDW7YqTXlEjBWbOe6KvCeFk8XaL6iH/emQOpGvBXi6PS6wbO
Yik9jUG/DIylDmYlKGD8tQXZ8A9eBk/RM8gIEJyYS7qBqv7sd9rE0DZs3kX0pUHo
XRdkEoDgKoXNFykgF+E2HuChyoMjkra1W7UcmrzLYBVD1VH6p9SGhuWNwMuC5xVt
bs+zSuWMHHY2lpfan9jXY/u9ViLdDZmFFGW6UPRTkeAZbtyDAG6eXu3y3zaA+/JO
im8cZBlOZCKZw0ValH5Kqv++w+yaNjxhpBe1f/BVQU/erw+VUoyi/i1AFa83BOwv
Vz8eieJ7AWENMmMq648p3CqhMRvuf7n7dcfe7i7FKMr1rMagD7O6BG7gdlgoT79e
SHUynKsAuKUKgnH88i9P6pFJKRkVQIjlsX8IuPyVyHGY7uO56Xry1j0piwGfuuPS
86wBvSheoZZ06hgtlGNGN2P7SeQwF09soFFJnOFsSndu2gQkafGIx6TJLuDZZXl5
Rz5ff/wEues/YRhDbTc9GdF2/OPQblvOlCSMjpL8iPO+NE1MB15tGLckMgMK9QCm
oe5CAHE4Ww17Z6gORxNr5Y9XvfNlOJllJ9k4d4SBiKphRWyjnYopfTyx6nhrrAh/
eqpQ4pUHDS3t6thK0yE0Kglk81OfxLYts7ZyqcZnaCyukvma0Sd9xwn55N597kxD
LUC9igIs1Q2Nj7gqvbJS3QhSh7/h0ECF+zHrOTSxMcdnFg/943aWXEukNy7LOZQ5
F5Eqb2H0VURKBlVi2GW72FKtcUF0gTgzpRVtiaZ1dup8ZPkfRSJvbBbtf7YFmDMB
D0eTlxdee69U+9FkBs2ptI/L6Ie4ZkhB3hJjr6VvuoWQHvj9qoUEs2MeFyv/0Xx5
DN8haYTaFsvGu37OUVuViIeCvnT+aTVKlMCkBbB3GsYQVxGwWKJ/5DZqL07qIOkL
BTVpOcRapFw4hY5uCWL73AK4oxZYbAyjdnlTrtMPPOrXov6yz12NCkSynnYRoV93
gqnhh3dWeQpP5OQIsM2n42Wk4yvEiPnsJhWqu1h+6FK1A0/1FyXXx5uCve2eM7Ed
lS35lJmV7KZJMLsBOge5gvDXsEbOIfj2Tc697lmNGIFR659z9HSIVwFpPoaTjeif
SYxR0OVXpebncy3UZeCy2wVDCHdwDIvdtLNmGROyxEfTYV/mYGiX+t0uXMVP3GiE
w8uuokbjO51R2nDNlZeqePBfPtI8D3Kc4/89JAZ546RGc8B6HrGr6o+YXYU/iJDu
r4OJY4oiWGGNwRtKlWAl+LH494zz1Xe30DZVYqg3le3bprFvlH40pmv6FyXupX+9
CuvQrqfrZDdm+zyxUuxbBOsXza3INizucmaGCddBon93ACjBq++vxVjk33Ma5lt/
Ws+qHbB99RL0rmd+msW6ba+HSp7TaBrZLix3mEdmHAUZ+3Pbh+PvjYcu4FY9Lya9
0B+Er+/HZoHwHSneK0thes5/MHXRTf//LmXxLeiFMHg/EkVAFiOtcmKlk5I2YfSV
o6wKCOqO4x21sgsXeNTXjNmuKWsxM60Om1d3Vt95PjV8J4tGdHMOBrltZZAdp+vu
wmjn0LKBMOaI29qiexCcOp9qXGV1Kxx8wNy6Cn2BCG1dV3bnuUxOdlP6AJ2CHFr4
RvL9RMfKawRkzLBvTi7RSXu54phAIc5EXyI4EvmJk98xYw4nGgoZVOseQYfciHWJ
W1af8kHnYPYhHltltaWVqaoEWTrT2aeofRO4lwqQIb6Ts4qdp3u/Xn39y38ovkxt
IGLgmuv6fsQvUtcBQzBBZAt2hM8b4FfoCOes43jEv2yZloVir4L5F+nkhtKLFxM9
4ptnoiDwCeaYgI+JzWyx+4reg6WRFmzJq4OzvEAcMMROqTa2ATsigW91YfYY359U
BYzwJHWfH+3VzZA82oFk9zJjnXPaZOv4NTKfOYvVM9JPLXAfyO5WNo6gnwYsvn6D
KmKbDEFrMOctSwY0cP1ApVJRGbpVEvPSbBP0M540URNDOicLRzU65VD4YPb4gtBO
R16QZv1JaRGXCu/K74ns5WO8J3FlylFJMCYnTz6N79hlxPRNDoDGBKhanyx9/qTh
yh/3NlMEKAOyyycWEj7ygK5sGLChZSaCk+KegML4GW/QqXK0vpS0QFwpk/Pv0ER8
Ign/1P0ww1gmwhHIkPGzGRmc4iBFMUhIMkrjeroQrazjVjUk/lO2iohoDz1iyDnb
aktoeV7ox5UL9j0QDwfhmLaFjiABU15gY2NFJS0vOY5vfy4PeJ6Xp3DAkVRwYUda
azpHMUWdDBriHqnHjpGYNUADZcQkdck5bsK4uPCACPQ20vVMjGlF9NsTzG1n25kF
H+zgWb7snC0Vn6o2akUXorqBAmzcJ1xd2hbf0aHrAt6nxKYNZrdXRvIB/T/QXHJt
pZCSdA9Kgh3qBzFc2jpyrAk5Rpyen3jlZ4Z0mDgNtexOSoM0COin3EW/n2tfDyWC
D04gVkm8aa8akcWJinsdwlnF3hyObTfnvSeRXvCH/veG08YYBD2j3imtXahZcq5T
a2rCwTC1KnFh5AGm4x3wQhY6J61CJMn4yT6XzO7D3F7I+XTH3fVZvTbe028IcP+M
Uag3IrwsfDQOIllRatkQpqC4lCLiDwNxYhyo31ZP+txbgW3xRTjZMfbtEF54Xtag
m+PUsP/fSs/G8PAhgltQ0/JpWCG2GERaD6eHXnq6RdJ+10IIuNcwhfUon5W4viDj
HZWa1rW+H3Lmo6O3RSjX5I5QTlE2POeqgNC2vQ+z6q5cPgRbcl94fTTHUM7PQhVM
z5BL6nuW5CYO5lXRwpdiPAGpt/FV3ZrllRb7yooP69/B+E947RmD1xo2YSwBY/Di
c9mUyF3s+EEs3cTy7dvmxitleLE9jq8aukzAEXNrml+yPItXf3u3rtYUhcoqo4eK
Hk9dUpzyBKdUivKW5mD3XJMJ7UrfQqYlIjn/NngKrBYM2wUdtaiTD0pyzXaZgJv7
Q3Wx1XsofdG4IMGrB/HxgfD77iUirDepTjWasPrCu9w1xftXdU7w3OthcuYyoGcN
qMsvDYk4w59QiIP0IbGr2jN9adAIw7zDHrBDZaDAg7V0kKII81SSXA31rIWBpOj8
pq23rU4Bg2axy111IWP98PRYVJeAaKw/Ob1yaceFhOFREtlKCrBt8laUC0ckDr8X
LQwA6oGLU9eu1Z9+TsQMi7cgISusdo/xAIAHD6ziHxL+AYzws7r99RcHmaUDZyXX
/kvnLD9Yz3mrRktynjrzw1SFWZ8RW49cnWNMj9iQ+4NI1XknIe/AqaxxJtL7NDfN
VylfnKnbJpSfyAEi2zyrGrL9GKJTuD4X7Lh0da6TVd8/T/X1VUs07LAtj+fg/5tQ
kvt8sJ5R8fP1f0dTcdJDWaUodEPD35Jx0NwqA341jVm0BSvmrKzmu0ohaKgfkQCx
MQdosM8SBgbrR+WmmOPUdJsMqhsllvyEnPja/qZBUPyWeUps2CVo6+ZZuKEnMTdG
Lk73qMgg5sdALnwMYCcdc+GmoaqJTTnzRi0OTOhg6fTzFhTbdMAux9PEOFJIVSYZ
swnWJ6TxXalJcnXOUuO397gPchwHaoTbO3Vsbyvh9h+E8cbm5KMs89BDcNpP8IEk
c6bwtPrk7XURi4Trt22V+OD/YQ8lkVyEzKqJPkrJ2GHdNIKLfrdr7R3p9FuNmCTF
c+6Sk4TQ/paY9op822S3ZjPrH9xYOJuCDLhwRTcxijjdRHkJTJ8jeoJY+6jKNyCb
iFU65olxEmaEIdt9E2sJlRkwF3hzfHDOk32D88nOrWT+rkHx/53SgaEmWQm+7VGV
qcZC+knxYJbEOS6R856n9SlxnYRi/uBLJXXtaxhihFXWfh0J+tVeVD2matdKF88W
6lWxnk1yAKNqeEFVChjYAyDr5LCrON44FTe7OKDt9i82QBOeJl33VlgtwlEwdLSp
zORv49H3OmtJg1hSQ4yivAm/7JrSP0HDsa+8Sb1x6qdMFfNitg8Ygc0fFhZIW/fI
LUVZOUeqYVvvZ/i9kOpwV+87bQ6epHiXgvXWydux9fHbvH9cLB/UyC7O4oh9gbaW
BBywf5rI2fAASP/0txTD9FUTmLoiMt91a/bbuePLatI18A4hdIgd4Ho1/bwpplEA
3vOzy5fLpsghoMmHOZrjQNKpSxUxXFn9vgx6xJcpAUyV/Nm2rKRGZLw/NykqkVcn
PcYFUCPIRXeRfayvDtyxLEmkISIR5dk5rlDcFbCQ20O2/iaph/Uf7S9qf86hDwyI
8zdMvemqzol7qSN+zHCSmUYaaHc6pZFiiWo45jWfvaszmIGP/cTDv6D+ipkk6f5Z
Q1t0nOOTCstQsW5AnGBOU6lWn7oWB+8Tayh8eaOcuPRzGTzfmJIm2vuHxtGyFXSX
mCf5UqgkIPSvn5nIgntnk0x5vLBxD1O2U26HLmm2kIDCM5cXuyAp9yrldGzufCeM
15fMrZm0GoZ3cJhezEuQWDNh9x8KXWepLuBxLu/lbcI9DP5R3r4qgpHoiVZkPydQ
CRq7i83nrenpki/0wtVHeHc6USpTc+LBiTBbiESw3+Qt2ghkC6kzrpiL42RtlC5S
Bg7us2En3Qd0E/EqReE7AHszbQnwmAHgQvb82ci6Us4uQmx7iEopSVN3xkPzcPKV
kWvBtxgaaCNeTEjQjvfvCsD9atUeh9+ZiGfJKKm1hM/kmQnlS88j69i6GQzRfSYb
1kms8TN4wTklrkVAPso/wde3hd7ohKtjkTABX5TqP4HBOgwHxARuJFQiJFqqUbB8
6D6DxIt1ZW35NoCFvwmdBMNuugVAGWek8mQrHzDSZtb8tdpw7yBH89uJqvdnwPBN
fBMtC/6gYzG53aA18ygCvelDJYBFNbSidzhiEx8BV9CLk/8qRO/TRaaJkF+Ixk+L
MFWnmI8y5I/7xkMVkPXimKwRSRrIRb/7LmRVZAQ5RbwxGtqHiXQve1tJ3b/7IoUI
YQelXxmxStzNSptEdZS5qLRYdFJUNUde8DEVe57LgKZYWm7LQjkHQfeh2v97okit
OJgVwsdS/OMcVF541R9xtj4IyJeYFnaIagp0F8QgV98VNJxH10BiV+9gUhA3xsDO
r+IPuTaFNpsk8rpyfsN4f8lYGN/CazsDiKlI9sFLkfESGPeRHeUPABF8jng8ex3N
uVBNr/rQNhH4maOnQOULGYo3CvSQvFjUimJGERg9AVQh5Gqm9IwTqXN5nrzpyTZi
kbNzquXsca+4bGUCE68q5T8N8Ro3lxdDlZaiKm3DrD6gayIYGuDH063uHQ63dQP9
cWJLpYy/1Qm8skCMpTPhMMpqzKKnGuYUCmBOiSWbzvbdUDuPI2NmBMtTp+mqIbYW
UB7Xb/9VKF1FU5sn84XCw7/KPMqdzQcUzYo7sHEUWgDmh3XZNZs8f1dhivWpWoIn
Gol5sqMHYGY/A+pqZWpPIJR6Fnfkkz8L/z5JEbWsB1jIUNcf1MimoR1wVxdVBuDM
TbnZFzQANb5EItvOcumf60J1aU+j83XaZvNd2TfVkvTAGUOW4OXG9FPlh5k4w+Ct
cD2vp7PwAemBHQziiW2Ob2bjVELGJI1vaRjNQKpFkhSpboFnynN4jKX4GB5NhdLU
x4UQ82AKuYIMDsHIi4q5Tu+ZEeuNPWdL2Rzr8VPIm1y19J4L0bwsmr+LFGIaX/1Y
THpQY5u2aWfOKL/O2dDbANvbsX14IqkyMwTq77lVNEGbDfo/FMT7Wc6nRYHiSIvi
3+ynFzR5bT0zFimCrAojaF0TOU5ndgfDB98mjC/C/PSE1YFgNsfxOYZ1tjBhAIX9
MKLpQbVSIHbbp1o2FyXn2cx2fuwdrl1O4406DAK+goUeYD+uao2m7QHhwaAtzIlI
n8jQHCcN3qfN1bTpnKCmkylp+MMlwIqjp27tTYStpHLkffPIZ/YGg48kif4uxdXZ
NRhg3hl+c6Nnbvc+2ajlwcLKQwiFoxzCqJryIQl2NqlH4KNY+4zzm8jndO8CUvsV
Fh+u0Y+RyEgP4xy92nRszKXrFm5mAYa1SVlIbcxLHtj0LtdyWA/UPpUXs0gjhsOx
MxKvUTlV76VJqEQJySm+bVt8NaSQy3NjbYVRhiY7AGkjZx7Z0DmfqACi3k5mnOGQ
TSdZpxGZjSGpi9obt6b6oNfBHZVWRws/Ohp5l/G/he4kdGFPio4ikGmplUxgp8cW
01h0gCnaFwHaUDyVTMFTCFy+EiqGuw+jnECjLbvpjWQPYIP5F4YVozr43IQyhNZ9
5gbAjSa/KvLR4IdWUDwWM3ANAlrOZfz+Eq+fi1sSwoOZEyvcNDod2Pdcsx0NLye6
tBd8zYxM22z8o0M72LABA5ohAsFVnu5BldlDixsLCSqLZFtWcljYVHoEXI+b6zRC
3rbxoWYNipq7htV3uaeicF88BbzWIBnqpkIVo2EjVpzBkG4f47jDOsy7E6KRxYlJ
mF2IQ2uBpVvy3dhyepw42mMnIFIIBiQObpEQl+nlBphKLWwj9dmTXrpK/68H3d4Z
w8lIjfO2rF4DFHlrDWjhr/RozPrUI6upmPji7O9tB6j4jfW3cP8E/ZwFuezNTDSR
7+4BT/pLVShVju6CoH3oOT6lIepHkyP4XpdpMtHCeq9eBKDdRjYpNJ4oypGIBLdT
8yb9tL/7cEpnvHDn4mHJhibWJY9wFD1hr+Hw8N/16d1ah4v0u5TqF05aIEvXanrB
NlHKZeZfMgwt1iHqftY6gqjRcp7G+yn2br1G4k4xF7TeaYI8l7Zp6xyBsA2+r9iy
r0iVX8iY0X4OQETVWj1lrEhFRNh5fZxe3EOXatxFSqZIei57VACBcutOSBXNJeXT
+tHqxQiWqw0S/cfdNpUnpKgdHfmWBth8GjKQ/O+po2k5VXnHutwahy6lYfwrKJnW
/UuhoIlHz2No99+Vi67T0NHeQV0OTxEGdDqomjfgw1w9u3sXiuCzYsQc16YjUPWq
gBDJbN6UUl9+9cNehoyx+MyTV5l89moEVZYqCmYn6DV+4XOGiCQHCVenfHRgHGP0
4i+Tb48qmabM+cqKaxazhbPCt0OnmuqJAfeafW38Jtco1mAH+Yx5P5FHVAEkaBm2
B2CS+0eX+eRDMEDgUED6SCFGM5fRbA/nTZeU43v8wIeQamjdGZ7qmFe4OxLdN0Sx
PcsrRJnbQ5JguXgUM04gyCsdhJQkt3p2RFfN6F2MjifyiACWKh6r0cE8aSyzdPDh
eNmCGx0Q7+y8+VBe4MNfv6EfD/oGnipbdC58A6URPv2nEjM2yda+YY5JHF8XKzi/
Qd+/SQI/rRUKiCa1SjzMyoSADsy8ZBVQk7kiLQbginRC5jOVlEf5T7Uftyk2wziU
vrkAusfp/fIi5cd6PTQIH80qf8fH52CTmBzmyJsLaHUTVSz7idL5VTCEkIKpaVSe
3ln+17fXYSnU0XMcBCJYtNZ4eHWbCTO5AMTdhCy9OdEDaHtuOUZOGv687emxVR0n
49cnePxQdfsEUQtrqChYgpf6kiayJUexN51hJTgMLQgsQhUFwnK3HaaHkww4iIbt
pZYS4mD0Ilqu30cBrSiEaZmz6fRuwpSUN0S14voKxbnfUvK0RIIhQ+l+Cw1zhX4F
vRPI1kaldYVO1GJ5G38kcCJ2oW1bOjsyz+VUkN8CVfsrjOxj2jV7P64jEkCETi+C
DOQKOhWDa0I1gIU2qPzh3feBs2xi+dpBTakzjW10lC+ZXt5AEPhtTzp0D/s3fKMC
gG2jlvcV2pSyaFLfRcQEbtw9Ipg7OXWyS39wUkWliQk9hvK6RfvGEU9zRHmjsTbG
bNAIgjq0Fx9mRoNz0flITG8hYrpBNmOvU193TJXYNQhtlzWh9hYDOdyCbppjLDRj
oi/rcaYL6I9O6IpdIJ/RY+uPVCmq++nJDqXVIjqXCx2QzEZtBy4MwcCQpgDw6S+2
0COH4ubxRxD5NFvOxExOZ4OIKb9Css0slwda407q9hdEsriaf8ZtiFHUpDS/m8uK
lZGEMMvkg0le529NEg8mx0wjVlGyzUWRNh75JszWHUgqhnRIASl0gbNXpeF10Uws
fUOmrmGDA/B90EaYIW3X8EGfzSS2ijv7EkcibLY+6B2r8maKjNyjO67Fa3MaOc/h
m9dPvuNbooro71aZ2VOcGbbOMa2T2kqL13/bgal+k2lC1eSPUJK2f6dKzLM2Tjx/
a6+maHIB4b/qmDgiBg1TaHqTy8DWTAIBiMSpl6iFvBY2AZmYyhJC5A1H0mfnavtD
650JIMHF3+kjwRYPRjSfg1wvDUNzI4ZsDAfEgVkWSr5iVzJ1I+oOtd/yuY/KFtMq
MGnjeMcqod7QHzhDxT/jQkhZcV24W519858JaRGqpBl1+m23v+NIxETZxB0Rzxtu
5l32SjfJfrr95CzRpb1aWwoT9IaVQy+CRrwzsdBlbvJm+tMewLP7IZp3RlbDDKcZ
1izL1e5fuW3Tkb2bXq9tHvTWBz2w4v1zX+0zE+UBMWqCcLrr0Zyf/lGFZf/WN9P/
p/lRjw53lU9JYcMDvrfPzJkaHozdEDXy1Yxw7dlwGYZOcFAIhOC72TJZfg6kxAUI
vF4f/ErW1h6RimXOjsV4pxhXk85/crZU2buj3SR3gXbfRwjaNVrEinG33fj0lxdV
pxjsYVIcXJ41V5CothlU603ftoIwSrIPqeO98XzEUytz+YVS091lunI0enXxbf5J
hEiG9RhcaL/Afe0+2iJSyM8q5O6neHpAJMDe6Ga7hb07uHjnC0at2hSMlh3Kipw9
DHsyXkUSn8RGZqGx2vcUaGJHAtSNL3eGSt6m01EaREq2LC9HhJ82WAX/aUcb6YNX
EKnFjQZPL2Cp/Fb8Y+2MV4/8kVVQE7NxcuGwqEFlaY3hKy0KIrmpx04ubJK4cR7u
IcAftPXQA//AACiSFn74GD1txjaecMmvTLaDd3ZhdANdc0l1pOuLaE0PvEk4rCNU
krTaweHSDrqiDc2+/tdOHfjN6zcGYRPcaTbtG0Do1knQ6mL8NdiTCGjqSUtSyEDN
wlh8dKFiPPHV7C1tr4GTrJzCAh7/kPixf4oqsWyJbfxLSeia69fs+GSwceiE4RxS
E5EkKEHrQ8ShMdiQIOKDirhiX1mwbGnb21PnIcPefdMzejaz0/+FaUEIJKIWPH+C
6oQLSmJjDfAeVGMdOOYyxCk2mQY4ypvTbL9AMhGXkusoCL+7pjtlMudRYhMSuT4e
u1r5B1iMsNoWsyiWcQgm08Jc4yNqWY8Ml5S0ICPUnarBAhHQPmK7oIk6bofbtee8
hh+Vq/BMGHBfOFDYuIL5wSoa+pKfdvYLAnQ99DpN6806yvmhlmMNSGxmB5mHvUPj
phYUDVykD6ltwt5OfX+BXct16gd5u5C5ccfxGWWx+ZfVsCmx4OWYhhr8dqzm3ibg
1uk4MTOm5w9n1p955t3BRyQiB/QIrQT7VOFHwIr1EaZ27iL8VOa4R+9B8yKsZLUo
Q2OI/hBEf4Vdau/cHLz7+iiuihRy3i1vVHVVJ2DK3Xedyah5XWBCImdvuXjbs33b
qJzblBQTQvJpa+5s1riV/WIL7yR7zbcdIHHKNSyN4LGgU4zY0EDRZCDSQ7mdNQ2L
UZTy+LMnMQ7m64F/WfszUrtdLk7yrNvO1XdwpvqVnFMAwK7VwIqyYUJUHEZs+mCU
1DWVTbFxnKxiO2293R2eP1WKn4DrJSmEyfKVQ8kOnCytbD3PamDteqGNSIrGU6bQ
0f3uihX54w2iT4AUAHGcE13dP8dHmtkFnTShIEi7sfv7trVQVsy9z0YRzvFe9oUv
K9NzZTFTzgADXqDcn9iafF20VAPg9Xk0AJaLZqDxJoBzxFQvGOLXfHg+kJG2nuRw
cShYucf4K3eYGtcaDvNN+duw8nQYvA0QT4MXlGVFPG+19Q25B/10hF8JnljRfYKl
zs8rSokna6Caq1jq+StYqgGlFNY6ahMTeHqZ21Vf1WH/ujbMsVNZkc3Ol96SSAR7
HPqgFCwLuGZITo9kbAlTck9wHILUu/5cXt0btHU5UycPif2+r4bSwaItTXATp2eP
Y05CJIVi5pM8u+ItIo++hbpv+VAp3LsYyAPx4hnmem0Xf7XAn3f2pY45i1nKSUP0
X8W1CvmVBoVTl44Y3Lcg5Q7QwqFZnIejviT4bptAB85DQhXpVChJHOPrK9n6yMn5
Hr9VOFaXQ2C33a+OLuZH1xwhBdUU8AbEsW1qoqzaard8mXhRbTWWj50WSc7/oVp6
zzvozbKj/Hb41H0waeTTssMuP7bQ8EAxxa/jfWF8/U+3fD8pvPToqItdpIIxDeXm
eEc8QINCOPpJevb9tDGSA6U6Tc0kMOfTyfUI5tSHS47IM71/G1lMWGsSv5laU9l/
5aUrHo/u2Zu0lb2d09Ojf60jBNyBK+SS51cn3SiFy0Dy1yXIZX4LfOo0oVZybhkz
+HZyZOSMHIgjh8GhtoHDaXEyVJEqQnLwvquXrGA9lwKbdDzo6P/aVxmQFg/y3Scw
VE7jop94+DR93EAyJc3i2FlHFYq4aGQQYFgcaGpkury9pD7h0sABY0KhDH6hiio+
ihPrzj57bwipzDOGOad/WzQLlVK8gE+yo3/1ey5BHMo5u5+/gRbntCZwEeXhziZ7
jHgKf9x3e7bEwKBsBbEW0g39JylVXpUfNnfma44cNbGa7zIP8JkoTXCynVVO924m
KrmrY10qHPVmC6fQYnFzsnFpSakj1PSvIpC0Z77YCCjo4LH2HZ548iq7SoUFKXKT
sh3/DKoXvqp/FW8rRB/J8A8euTjg/7crCNGASd1GKuA0iITHDuzCZR8JC1a08GN1
xygv1L5hiwY2PU2/NAiK+sfYV0zHlcq7KUIptr1Nrbt7wqeAIRyMhY4hrrcgZV5n
8dKG3lEpTs2RpRGQzXpXt4Bfr8mx3gp4mj19if0Oc9dsqhR45NEQExh5KEo02Voo
lE6p3M+tg8k2ySjsu79tvdzdkjlwOzVIyoRjbqx740t9Y9DbZPOxNUgt5VVsnQir
8LktlnBwa20iuU0AjgPJgoABFKih6XhR9gPPxgYINGDyOTiZNX7mlp+On/5sXM0b
Ep2Ky3L9ANZgaKRvnq6J2MFZEPnSDul2kgXY+DWNepLW/fbvhMRfPgPO+9odnEE7
2uenMaS3glzuNdZZL7HhODmuvdXbIeTyLRMjIMoog+O/3HyDn2UWhARYEkT7DsrB
BUped08WW/yr2D+HTUaS0At8st8az517P5vuTYhim9AtRUyrtOx2ZvVjMhP86ut1
yKyHMfc7Mf0UKnwGnNdKh71bPUyPCOPnvA8yEjet8VkeVgMlNo+PnA5M/Xzy5wqW
LT89tyrI1J3L6sJLIj+chvH0JWzMt+tXGTP1MgqAjKsFzeQ22mG+f6v6hW1YuIBM
GS5fjdlJA7zu7U5m3gOGHThQLA5pPwuwY0c+tBqx0EfHE6Nyhh6V1o67fxIrpDnn
IMS6LFnt8oB7c1HU/jMtrS8YX3AFzIR0KjjA9NoOqOTHUWZsaaws99IT8YlE9WL8
FDk9m2nPeZS4kI9H/Z5josBNThAEkTilGD4lk0SR0BzatRRV482T0moMN+SVA9xc
B/7261bQNRTchlNke2Bfa10J0+bn6mZ89UXQzfqqsvHiPMBrtRBCidwXwIOIZMH5
JvY93P6b69sho497lIbaV7DWmpBQYjn2c84zb50Gqh2pY8q2gA3bNyhtq43ltZsQ
Z0Eg9IlmAcBWQofJcUw0UObdO/iD2NJ+03ID+PMSBmxkE9h0EZisU/poKfZSQXkS
OubUjKMarxo3fLC+SRNwNmk28kvHU9vF7nWguxMBgeCn9NBg31ubIfZIKmliAaxk
yozgLGitOK7jyECawo0eA6NV3ddLVRzTUiF+BmnQQbXV2WFa3YYt6WiAjqW3wj5/
l1x9e06Ce/209hGnxQtDJL3N89hsCAxVILIfZNbZHOho3ido2HiD/8PS6y43Z2rA
sFpYl/r2gPQ9zw6fTAkgQ42WTf+UBC+B5tbVlq4KwW2fbXb1t8g7UY8tMHMDHfzH
wxtNqaIElZ9cCPbf+/nAWSsSYjwHdZSMPIoi0H0xjhY7wpVwla1VMUHoLU5H5Vjq
lrorpLsNj+2djMS/dJKDRhxg3jLTPQBaIngDci1/UMx0PquJrFi/IhJslJkACXL2
x7cm23JNqRwz5X5pt0eqtdtrGVRma9vZtF1y43+9H8q9Ti18FNmpncD2XRtC1JL2
3A147+XOOratG0/+sCOLc+adtUlAISnPJPIKqJyBAGSNETmCxUyHukIjiGBX4YCr
koNmm28UI4OEUm1eR+msJL8ldWG76Uf/V/z3/8lR0PBtVFbg2zkSHoerRsYDr3MA
DEoVZ/Ka9t0CB2NM6PKn4teRh6tnrrePj/X3vIOW/M+Y+fUbmAfB4LE/GWObl/qR
Q7wBD+RbJEyHg2G0oV9urwMER9Zn9Pc6mydSNxR8PYTpn3RiJcQD8OO6OH/KjkzJ
OXrkIq1l/HShk/a3W6xjMW0DXvvU08MyIsIPkTsCcupV61NyrEyb4q+TTBTcFLmv
8QjscP6CBErOPv8lPbRh65PvSOrdeqZC6rfpCDONzuwAvGSztwqefwe8vwsfRh99
KnBopuEC0y9UXG2x6xvYkrD/K6DJbrCjxVIqSLz6oqvXeZJ2a5KrR0j61J5hTqxe
H8UEZjU6mhsz7IuskOHWh/IAtXPziZKkzXlsB4vcPFhO1vyfnZW6Fuu0hRWov4Pt
r4dRnEptfP10JlYIsQyAyTEEP6Mpe4ALm4HVxqo4XRTzolFiCd17hXCMaMxdn3RK
lypIguu8yvYIEUmT1lkCKsYk+8fQHvXNma3rJ4wCjSieUHwMr7SmFvDUNshZiNZh
iVDpzDtYOHYTMN54jNGhuULycbShufjhNPB8/Mzx8MHPvwScjObKEuXqdi8IXhjf
Yg/p4rYRnN0G6M5GIq8PKhIjEITfzC7bp9zBsuL6tHj7TNSnYzupNgOCjbKMU2mt
bj8vf2uHGce9nnSocfKgXmnyptST5aS3Xs7Dums3sXKKpfGsymXiCGMDpJUw3orm
VJb2HTyB3716UwciIAZJb01mJzXvUw1/M/Y9BjXgUc9eSFXZkKT4Mytb2XIQhgue
thWvJkw+BOHCfqQKPvBT0TBxG2mDWikcL524LZhFVriNs+lqq5i9nvEG0zyi8OgB
MPZ3WfrWXizDloUac6PuZXM5WhJI8KlitV0Kd2cMFDwAyc1H00cuyqpS6itIRMPe
oGQYvfojUrFg/3R6Xf5BycaRq9sp2xH5bXmDZKgXFEPFgzZDD6TYNj3RELU9k5Q6
4g++he266nrJpcb0KXpd/BLZtJMagAKR4vRbGynroCFJnDlL1wUc8waJ9ho47HO9
Kff7BbjPZ3GkiWn8sA08IB8e1oVjehv0ag2wywKvdqse98XEPOrjtB9oFYHayDB8
r7dgaHMlSwxsfbr3XtC9AcKThLPalha/e2XtpKdW3eDQ1DujecjFUgu5LOUYP+sx
u0IKPC52AjzAwPyW6X1p56Ke5C7uT8yxsmRzXSTB/0UtRGYX83xAYspcpC92jrU3
LnAdqmnlaFekhR2Dg48HajR3CGCMBEVNXfIgmsntspVBY5kdWto0tJkE1dzjBwPF
8rH9wSFDFoTvJprrPkfD5fQOOHuVGcO2ruGqGSKzZTEfFLKuSzHtNRf094T4FMHL
0eAlJOIGcEAQtmpwwLOozz0MoQn11lIWeNWlIwqMXeQcDMrxy8Kv8iGAA1hcUIjN
9LNP9+Z2akHucy2JhjTlybwbOVmRw0HY93NIWmcBuAzqbDCC42sMW2jdMdM32zMd
HGuktE59RwAWkPwxD6qdSyHV7qaUMpfEac/g9T8pkZPwz2WNTmdOMlWVk4prZ9eR
sNKLDVtxe8hV7qQfBed2Hc0SCFwGFa+h4SbhMJCyJ45S2+b9fbcTUI40ClEoiM2R
ok8X09WdWtpUU9o1UyHzhejHOyilaGWyBF/kaKg6lQOIbbn2t2fLOTCOAp6v0HFI
LcBQTL9o1eHqWhoTW5ZrHM81QkbRZnCPXgo3cc6wTQRUs+AhnnHrYA75mM6itCTZ
kTZNZfkYnvLuUB69OLKWZlxSxh4TmG7cfdda/dzBTlz57GXvv5BqoRonz1qeygAO
UYDbCvu3BpGbRYi4NO1lyOkEa/a7y2ANC0ynkAHc5w2pnZCcjM1S99MPeuvvKXrF
C0W2ZTSSgmbAK9HaVfKDkgIgPMyV5qlcsdWZtJUYG50iSoQlD2V385mFmd3+ivLe
aYGCc+Y6ZNWdyCswPrZTFVSLpyT/t/o03s9b/IZz7mSlKXAIfsycQ5vHazo4+eu2
tRSoNH84klIKGY6LCmUqOk3xM/xp7HMf6cF35Ugtn6ztua187NQ/fJ/KryeoW+Xo
/YHwQRnRXgCtq9I/HPfyEw7tGffFuRQj1rZP1O1zqVb7KqW6Ozy3UkBGGqtAI/61
F/9M5uF+4Elo9ehM9o55M/SLUKkTLbOccQDOak0DusE1qkH8Dn0HIwKycacmQIi4
KZFfuv6W6mDDu9tCnW4pTUXWTSmjm/Dr3DpInAxTiPpmF1g01H9JJhEZwbVroMvY
gvvvi/foUF3CgHZjBloFwgZxGXUtf+xXPT55078c5iLESpmm+Ph3g4uz2p4fHaGm
ZjDNGQj6CwYY34CUx+uYQQH5ahLr04eeZLo+AY+TmCJWbqxzbEESsk5CeZuCIprJ
XCZFacO1dtTgnY56VCe8yqmo0CnLlBxJIg4GtN45R4ld9qcq7klVJ1ttlhSTmRqD
szS0GAOIoAO1Ke8ft4BEgNDL4VfQjQOuOj+xtzBobEg3ZzREOpP01Yc54roFlMat
7c0redBaLN8Wd1EmAi8Wo1TDG2LLl99wwhjZzc319YEP+JaTKZrOAMnI0L0ecfDy
dkN2KnAZEQzOEy1zyywcebS1vIzImcrNjA0eGOcZIJILVnEAqDzPeCJD0WzLH9/N
6hpBjVilogJ1bvmI3tgPYQvgAzw5DfnRDgg791O6PEZO7OqPM9veLLp8Kjr8NMJN
bnSDkmdF7QWOT06stxfio2Xg+2kmkVO0QRhfYuf5AySUjzPrTvNlasCrIdBsIn1M
L2uAIMGrNvvC5Y/zSoKPd9o9V5Y85UPW2P5hzdFdUlDI5SXdlY5GbaiH/D2r21Yf
5T6cHXiTSPaUvOz+oWEDAskNaHLqZ7hw4FDB1894zlfMhQciv8Wygx6DkXnUZ9dQ
sCoXacSw8CA1PEGpvo+RibLWcBzCFUHVzSZngS+d3ooLqM6yQN0fZlv+6fiSjQ9z
AFDmfzimgMfX4lFK57ZalBHui1B+Foy/BOBNdIHgAVAx7cIYrYtH0l/+TKA844tV
Fx27gZWox8zDtdWTPBT2FIICoCERU+enlkl+gvMd2zugICpZ3dbYM67dlkfYpCnZ
z3GvOJ6jxS2jNgmMzltyqzzcBS+GG0BjjYxceG8oqabGEZHTtV/e+bUSwevvvcFd
BoGK/BcYSXzeTnGZqXb9WIGLdGynr7Z8bUyzMT3OapU/WKdHB9/kgtvvU6axwhYg
dW8jO0CvGiUA8pBwFfr3W0w7T7OGaJ9qbh5LuKQMT4kQTy0vgDaxdUDaRsBpNiCJ
TgncTM7zxM2fOAWCpAfO/JsT72WlpVHpv6tLSf9ba0P2zgCN5RqVtzJI+m/fsWwu
4y+B5kFywXWlb1mrqHNDJG7Zl28CFquEz7BYIteSzNLFcfAyHqfjQ53sVE7DsBeB
+qBN61dv3kToKLRyXOv0VDWYnKAPzEmEVZcIgM150Xe6tJc4isFPGPT3y7005U3P
56Q6TwycB2RAL0iednLpdUwmvBw1aiJPHN5/b6kJa9yMaoOQd0442+NIfWALfJX7
JxkHzWZdKQft0jBYmrB49+4kMP5Q8u1cQ6rYJmsOuzbB+S4n7KYdsmU2m/ZKh7dv
Nios9HmklRL+/x0FxqUO4/BlY7WmRYXsgHZulgGWa5+mSQnfR/soqDp5q3kLcivB
8UFTL63NZdxxICmPJF4FF1KVrtUmUhM8eqDrhqIE6+jkWveyhBBex1JlG33YaCQS
tSrvw40QAkizothHXlpdhGmEVA34u25EGq1rUVgW/joXd0TdGFOHYeNJkH5RP9nr
i/skul0PrKWJ8fzHKGmeEEEJvJhIi5Y2nKuiEV9fE2DNgdZqrckoZaQ2ldHc9Amp
218oB729p5IU2LcgOrLRHgGdM6xcw0PEqyNYdUDEF2y6c9LZPO2FvNkiq+Jg9Gy+
alzO8nkf/7Sh5qKLZSXt24Fd0E/IOOvZsAHEEgu3thhkeIm4jf5ndxGcQyNGFXcF
qKmZXJh59xAq7IY5LXc/XvTwT8JWxWrjhVkhnJ3N6FHDhWmEaVmBaKUhgld+LcoS
Z1yybz098UmunCeEKroo8UUObHBd3zGCE+Z8g4LQyut0sQ3YDVcvXacpX4uAelT/
cXD54640NaeYrGsj9XTX3lugRmex+HYBGCnNwupddJlViWy/G1Gdhw0J0r6jxQxe
qNWxnCTeQ7shpssFbv2nALR43H0Vod2XAzRxlcDHjlE8GKoeeOwytA8H+1ukO0Se
Lqqvveqk55eoJUG6bVIgGw9qDwohSXHnNfisbh0jNhCef5WHyPgIdQdnfRalLBT9
nE0fPX4lpVs817I4Lvrgwq7wFkMyIpm6/dZuunIsvnKjwKhLVU4gJazXP8gowsHz
0d8r4gt3gAeJUaLiuTOmUyX++hNf3CZ66XZHVkpQ/4Tdf8p4aHw9DLJ6ovEsN5i0
LwcOclBDd0cwIbTG2rQC5npuqJ93MTX6ExW6PlvGQeRWvbsHoVEfckZDXM71qrca
ayAz4LnYF9z9uyA7LhU1CSgWLHCLtyBkoZq83NF9jckKNPijDv1j67pw5qB0FUHK
MOrjogMd78luENbdGmPA9RQDQJ7+fb2X+2V73Rw/5RQFTHegsHf2PhZCdyoSpiGP
xRW76jSVKgT1RSJfoyS7BN7jyj9xaFCKNpJD9QggaesvYvb2dnPb889iFaKeP7MN
IyaTuRXSoDTBQawo9hNureNhWQxGR+75+fhg4JJWiO5HAoCAqWBydnXwi1DMCv3w
LtkHmVI0mf5NTD+nDpEDBTn1hfagLQhFK4ytFF5Ewbsn8UdyWHPriCNrW0iedh0o
S6rgeRkVXzMCFvSh4w1optzC/dW1X2tqFtO64yUxRHK9ngxjtV1pQQAlkF/RNJR4
VtMnRWLjge7lT3EkpjYcrhTLfH5QzU0PpRN4sBpEUdVNcVtNmPjcxdrVgTPvAyIl
/UYXB3sju4XNJ626+qLFRR1Aft4iyQtatmT/sRmsGh2fiW3vEzFIcwbLEOCGX/k2
GBGY2lJ4zXOb/lM5YH1s+4jakoCm0UtTEIaSOKD3FCMuQ1REl0n31Gkk2DQj40An
9DM1IM0fOn5YtTynBoOyIRUzexhY8esXgVZPaWw7cW1/zb1yzZIfaWKMD721od9J
Y62WFP3PiK8+t+ip/zgeezRPNbMZQ/79qLFI77QH4ysk6DpP9RshUtv+h6VyARro
w219RQ1mJMy1HRpZSdNUJkE7CQpaFVqTFah3LA6/mcLLbnRl/NSoc8Y2mHMNub8x
IVrNt7Ndgc1/JDBrW2zIL/5QqBAL/eY4LlM2aLWotWMDRM5SXKChAPdSNDYNDK+N
4v1nK1OHMA2mf+b9xqfWWm2d+7hGi/9eYmnMK5VCG9O/JhgYlunbOLgbVTalGCAa
Rodvr9pWgny0yWggwydhxM5LbyFnbI9REPsyunhab9/SSwfG5lakI+NpGKesHG6l
OnbtvwjSYNFUhqHhyefvZVBvGTQg4sokXfac3Pszp7AC/V3pwq4QEnky9a0eAN0I
djHoVtntZGu3z24C/v8Bu5zb9OqkVEGzwaCOt3fVsC6kAwJu6MhIDceJekOVJhbX
ms4twRxiQC/3EjKKkH1wJCpKQqecAiZhE6C2rjMxe5sQTVZzg/FDu63jQHVw6XGL
Y3zC7eCk+fSDq4pp9rRkJE/k/+wzamP/hSUYQgM+Gm2OXapjTwa2sEAWbeAk613N
GAfqDWK1ApqBmcThtdGCJqcenEWzxfn57kv5KHPywULXgiHHWZ4iHfwmhVlQDD87
asV/rEWbpcWIPePq2PPM+uN1YBTwdcXMh1Mp311X+UvRn2NwzNMKw0uCIhVw9YeZ
RdzGn5clUaESM6Yae7bw6Nfr+Cno5UUkpxhGcqNxAXQNhnFVVhy4BvQmDWlwVKVt
u2gFJGf1HbUYLZwAKNBQ8VBtNd1y2Hj/esqp1AFOd6bsGuWsQ/tTJn4fMQTZqz3e
8TTIRNDZppjV1WHlkIv7OTgoSsgAAdnhnVYRNcgs5p0knhseN8/JyTRCeo5EHWX5
C00XAWNd04CTpruGzG33//Qnkg65kFOM6XMURlbVW2fO4AwyS2a1VaX0y/Wf7MDV
IK2JdTQqUBp2c1g6cnXQCZMUSMhwFQNid68MxUV14yMQwnJHirYEJWLpXTDrqC76
3ht6hyDPhHqTOgYpofljVt1UIterh4xMDL0Wn/mxiLR3HXAfg7Emg3kcLdPsTi5I
RYPG2xwka6kbmaOlPePhscXTqiSi8RmLgMXVtg/2Q+3rdGUcjHu05gXaffSkSIe3
U9sa0jwIvxgRkm8wWE9JHL3xva5wtNo2WYmq5JO4ozHDQSX27ENnxu/cuADy0lrV
bn8t8SS60vZKD+Rb7bmBZ6OTAHryMKHH/G/VNVHVcEmFfWCpraC9vFivMuffNCmS
5RqCJOy/7ereo1GfewmI4kDOprUxS9aQshr8RyG1FTfYKNRjioMrYYcmrWO5XZ9V
gseBdbWroladcufBsTLSq+ZwMGRu/EeT2wD5/eBOD64QW9HDFaJKhg3HywT1i1c5
XY33F+lut74InbUNUW8tKu1jB7bedLBiDOV00Wqjy61kANkt6UgCRBwBiPpyC0bk
5ZXVyPxZmQaI24NGqbXt9XCJ+njFRn1bUh5uLGegJbqH0ijyd+30zbP4Qv+rZcJk
mxMoS9gqHAi50Glv1q6Sz1WZSW6bc61svjTHpwFnWM5oiudjPROpc0b/6XuO6MX8
W6J056v+CRoKZKaEjczOL3C8aR4kdewYpKzm5/4QaCeaiXndwwkEkDBUqXv+i81R
BWM4VTa0J5bqiRQ1ArJx3BSa3pcSj6OAf5wz6Rs5kqeyn7SX91ZnMZddReqd2NID
qndiQy++U2gPM8FKej9d+FZUjLLtn9yVA3wBHbDGLHAg7DbRoEs5dZvNVB3IFtzd
P2Zq/b/3qQW+MLhu8IUQQ8JGkpZMKLKmfDqiJVo0SZ9U0SY5wWHk2tmZ+Uwy58JQ
sv6msg8B4CAze/gtZmPbCW4MGLwgnga0f2Xq1UXPIqei53KpOo8WmFEG59ozwqEh
42ZjfgzkJFZnZ7EvLnBAPNnOhpVbN3BFOmCCAxuOr0O1ObyTJHMG+Ea0Hu+qp65/
07GyIbWCvp6U86Qgg7w42RDI1oNf8gzJ6yiw7JUCnaAL5EWnL6AKzB/g+661KWdT
RZvo7vAcbIzjFHiqomJe86y4BHbXjalJIVI8AZf6JKeZXTxx6eB5V1Fd0SJzhuCN
NkdwRfexAeEiuA4LMC8AHCqYofiJSo21j/uOFY+7MzVN6jDXgH2uwn0G34KSlOad
etSioHL6EDcRppK2DraCkJg/MoLUx4VxCqvkCKLfvQTTiUJPe1ny/hEaU/FALP/W
xuUQfQ+2HZHm9gVmbam3Ue5fFD0g/PHqnloN9f4bAN8S9wRY7iW+xqkVdT7AbPh1
SgpeEZuZnBucLalwNvuPVxL3V2Zac2M6huaZaWhFwS+BVC7HdN+SVERgmFxbPYlZ
E2pQJCliOGP2/7kN6BdtLpfL3Gh7jiN1f36MYrjOj2bhBllrti0LRDs6UHopdaAF
UlLhU25Jk1FqcetLa1nSBwWNIdWyRG2mMHyg2nPUKZ1PrvjsSma4Ut5gvsZZq3yK
CqKgsRxQ3UB+ss53a7sYbZEhU5M8wcMM7ab1vDw1R3RoIfzR7bsnn5NPSuvMWTdR
pXBf4WFSG2LjymR9luZrm4WRNCtWZdieCp2IjAOz9SzZYnK/6jKRn4icWiMCUj4/
dV6p/0a1yU15HNNSxgSvmtzqZ9KRhrIDZoegaHra2nfmYOQlRayrDaSF4aulgvv7
5cJgvxMnZsZuevMV7+Bd8MN0pI5FWX8kyg7qJp6r2ZzulEElWrL+KJ557qw+y1nV
CRx6SDFU74/GFzzL4TxO6JW9yHh8klKhdiZMRXG1zUgLZh10Arq3rctbh4J11e7q
8JUeIr6R4S+vUsS1mI71+qMwrHDT/l7nCYrc9uwi4JFfailJKawHdFhMxUM0eYUK
1w8y5g8zaayoHr6bH6Q+Bd+2ueZiL67TL/CP+XhaxLMKpPt5qfslwUw1VCELviQJ
nmXpiMM5Llmm44Nyas39pT7oPjzpMJUg85NEfYGkDvdYq/yxS7P9FOcTTtMgF2nO
iCepXhyYbdtuF9yZMz5RHI4xVHOEXRggbQAGsf94trKq2HOhoOqggeUKs1rwNYPY
V/cl0aVdDiOgSmfpm6fbsJwtDGTVVZjHD2HY7yiYjaVeTppQL54G8/VFPWFH2gUe
wy2Gi4Lj87PsrHPwMz6OLMv94MzruPPEzImfae0rhYAgSN17Fe1S7XCA0/gEIjqm
QX/uu0p/h1vmS91H1I3UdNsU1PtRV6P01qCsEIZW0iEd2ZeGPtP4ivQDoOzlxr6v
g8+8veKiPHabOZ+BXghtLcbJWkbJMabf9SLQrxVd4HV/uywUnhxXZECBlETOFsYw
WQAjywr77+Gx+viQ6bsR20YHHgKwZBrXz1wdbkawsngNw2TUdG+rxlkOnHlQVjuq
YVQ5XPRMY4+WBE0S1cPOv94UKLMLyihR64/voIxW4aHVP19Zf3QdUxRNU94Km9up
qR3vN1ccQ4GN9oPoDffA5YalCW07M/2OQAaqw2+/qmu3V7KGo//y32lnAv0A7r7C
CBspKWCp7Gv6pY1b9E04CnV0IsYyak3mf6VSVF/Z/SeZHyFtl/RHcSExY9qPsfg0
mKcCo5sREEAonOpLoEbmVYbjz/1UxeCOuCn1jwpHkWXTypAxUXUFihisv0BrXda7
JCPmp53/cBoBbncgFYx4AF9H9h2yedY0S/sXMLbNUygdq72ema+1V6AOA0K82dfJ
pEZurw6PxvuTLxB84ohChGWvVnQfdGHMaQV3NLywolbTh5FGcdjaih9zCHJoxNA1
O+OzkvU9Urx1QOYDGWqoyLIB1nGSceHRNtjpRyudUUvG3OydfazTUnaN6ki3teK4
gS+0IeEghx/5ReXuuAFnHWOBWvXvVRZ6VH33zhV7VbVaGbnAMh7ICsikOo11n7f4
iPhOo9WKn8qdcxuEnXUCeiLaZOOtpuouQMFUVIVrw0iC+rSE8d6F0fGUl6B8gHZA
KZw8/rUdTfuqUe5c4LYgqmi7lCBHSxwHr17scwEvwYiJLBU6/PYK9WSUFdCuBYmi
ELLmwdSCE2EQ3GqLMo6/+5whPfMjhXkw3n3xDJzpGLxpog0KhAHN8w994STC2Gnj
IlLjcVsRcTWqkG3shb1zVp9l65Icx/Wb9dq/oQQ6iGPf171mzH+bwcu4DG6ZUxQD
bFMsBJY/8xX4/NSjLyJw4g9DjbORLmyHF4dsdoqP5q9wXWUsMX2viFCYClFQYctj
mrGdnyui0H0sXdv37zw5d0p7paXcaUhulAxLQ/C2cSC0dXWFn+w8lTfZOlQeh3Mk
bYxRuDPysl5W/9Pq2BEgCPHtK+oVZUym3ROSv61x/7sFE41ZaAPycBN/pgC40hRF
6yii9EIbM6g9cluDoVopwYdAHtDVVArlm9ts1zrI3WEPbMTktl0o7MMH3NSBmahG
d6FYV4bVapDdWtmR/h36y82tbhQiJLnZFEdyM8w6IevhYq/1hWND6xUadCyG8n0C
0b/UrfhW1zGYHi4wJ4C2EEILcgomiY7FyT83IZGJBysw1dh9BnRUqlXvVLhUrAFy
O4qBFiPXqMPaUoEPqgbuU5auvoSYPDQhfEG/L1jDMC21prtuFkBVgcJsOJLnjhv7
xlf+FAffyk0W/5TqkSK0HNBsXnD1SM7eaFZE8rwIz+q6XigW2pwwtcaOT+4UqwTR
YZitcJfGsXOUhQEkfOlUuMEtipBicJDJ421fmGW0dlfwO4BsOzbUXW5tFmnj/Ztw
R+5ka1mP9/7cADT4rvCF9camCcW0NGRoHyrXcueYL9+LvziSprAn4KgYULF4w77D
XnetxUA2hxKrCdYYPwAVDtiGbfy0MzyrHYbRgE/zRZaVelx05FHgC887LlhRdO/1
M+qQ0KLwTJC1sqHfz0fmQhVmL1bXrjukPyTYjZHyJELkvJ5tQwbz/rLyNbTMUgcP
O2yEPItX7UILlPI1natypYgK/WaKPPPjEhcg5bfKFOyIgLopd3zwL9WkfDePhaGO
ENJ0FgHP0vqT8VQ1ILKLG4xQ7JlpD987nTvbfVO6PAAHHHK9P5hZtGCBSanOsahw
jrViow9COLO6H4RItBs3GiNCTTp3Aq1OTTltWIupqvunvoifyug3J0Fhw/UniltW
YAkRuTw2cUL+iDhqWthjvEjIFqgb6h7hA+BMwIuPDTKDMyP02R6aJGbkOQV7R1Jm
8DY9Wet+v5CH6TXt2II/dKa4fvKPJ1cfUOYdWN551lpGlSXHPMM4iePLp3/BWsPH
Ntr9Iq6TTlEb3gtLBhtzxD86yfFJGkRmjd6Boks9j1pheKmh8OjR7bOSJuIuwUY+
uBJ1wu6qmBQLJyHIyLIn7aoedBQvR6ovgdnB5M1aOx4yLVWKDrrwLBl6YGD2QC7O
QZ6DNJBER8tf9Dqk5gWyWtC87PzBXRFp21+hR+PdKdvmuQYuoKn5GGSIpxkwY1dZ
q9QRcpC0wYOufZHe6ZrYE6SVcln+JAbLuluCePaMPZNnfT4I6C+KAQK1vKBdksaz
6HM8VLGrV0W3j7MKIvIikyPCLJo4ggpWnE5INTuCTtCvCkzZFLl95sqbFUxj7ueS
t0tVUJyeJdzlDfseNG9AKUQl58C+XEGqctruTtveGPQs2Bjaxdez3Ey9rVThEUKV
6e2uwGPue9xHN0mhDRMok5ygzaBDNik7+DzPcaFZCMmZJO4cHgf26G+YpEdkGCvz
pCKO9wPhrkGyiGpVR9GoWpVQk9ABUwXe/pTbNXeft118ueKIiFPMf/tc4QxMHO50
1IcsjB5g6eVbPzFGVeW18SY3W9NRYbBHsHtcrML1locGhtnbBj14WLZdnNdE1Wka
MMh9TQciVD+YrqfPDExmbAZFZsasb0sCTGuQfD0BAFNQ25hDNpiFKQWZHW3leqlh
ReF9zPvZdqaMiYjtMPTTShkvIeiXSq4nLZkhNi0mf/wfkPvL0ake3y7cEtRdsrMw
RkA6UhStm4u+XwqZxat6THuWbDABE+Hlk49jV6Q31cP2VgKcBUjmFkMm7qNarYil
GU5KyFR+nFtvlpCzDIzY2bEkn5ZaayhIgnWckDgJ9/MQ0/S+jhzTgBKwgLKXnBZV
KtenYySMD+LmFGZEw5Yzo1zt7xxvTTardtsQzZtZjgHGp7qWaV1OWmNcxVUpJHgm
4A+1qI95WKIJPGEfNNru4k88RFQvAftyeV6l9n6NRgXTroUGewhQxJa3dTBYR2iG
ux5xm/lpn2uSm6snlIOe/KzT3/EgypoZnkQrB6Mx6FuQsWDUOQrjj4R3Kdhz6rdC
K97Bva2RJ97HkL6/6Rf413oOAZ76OGTdqPa9+iG0ZARLAWkHLA74yp83pbqDt8f8
jxrIFLXPaZq8aSPIzPeRqsi9oPfUWoiT1udZmsPqVWGrWou2qStnZsIYw57seAv8
AEHoMXgrU4ih6Ry28k11Xo9TXq3afxVD+OoPbMViMJ50lPY0nfKyPaBayLkt+U8+
NDui+V7DLY2vhdNJFEQqSxQp1cho7Tr5u/ktUSI0zcTtuK6/LZ+drOpU4TwEUxUG
gc6FYCT2gIZiergwvBwHTlP/obnjI3Z6CtlReE9YtvKwZCBmLBqyk8dJZyykVBD6
bV2MahrVj0bVJv5w1fImycHjRjyvAwk2HUcOseSAe/LsKOsWkgZro9VX0NTzan/V
WI38RPiM6wXVnV99sitGplH6wpKuBIpC5qSNiJaPx9532QGbWgqycubyKghhj7DU
Z+MoqEpcu6ITb701J6XbRzyWq02pxxYjLFn0CYWn9361cjyzG8RX5SJH7zL2nTum
wjFpzx6W8gTQXfI7d3NBKWYJ5gd8+sCg/H8Ql45EguUu1ZaslBH4C37Ks07q7mMR
DHFt+1fllgOV42Jp9qp553dLThtMJ0H2t3rhoS1P7t3VpfgEKaJibza2VI/gJzUx
x2AIfuDmKDqlFK2V9tMeGkrIHVJW6PYjQ4RxpeA0pP3Ef2nT6e2JqxMy7nrxNBWe
7zClJl7IbhjWVC6EH+o70nyRTDlLHk1RRe7pcweT29vc3/OO9T+Ij8KnB2DV8Buz
8TWZ6V9mqzTIMH9BtqFpZ80KZgjVfDx22SspqcPthVfrrumY4QH7uNbPC+x+D0lr
f1gS8YYbDvIVDDYGgjWHN5aqharOOP5rF/KzpY6qXW+nk765hgqxovsN0MogpgrC
17fIJCCyqHla+4AhRzOgoA31qSItezt2w6Fz5XHNkFdf7y78fI0xi7zDafz3dt9T
yvlEO/Y9xD32XzdagapAhOR6GIDCpDooslyuFKisIp8A6YCybthZWmPDW7KmhuyC
UB0HBYi/+RkWgyQT+S8WFW05Axj7ZAURUmHZC93fp8oN0P219o78dWDoC9Ge+q3d
rCfo1hPGiu7jnzW32RhMftnnFVrqsWj9DDWIkMmTQzBuSRZ+qlWan6dNvGh7RR5n
OSEgfzhMinQxpN2vFfkR9D+ETcOuHstKTLKojgBWY36rKWNWltI8g+O7owJLdere
P2y8Ms+ayEVfQSzxNHvs+cs4033DH8ndKypErMnVwfsudxh0VKFVi6SrdlawuWbS
8//pGJaEmdiAaSNSRvFpcV7J/1/k25Mlka+6n3ymJk1XUs9UVO3WQLXXJV9KJX5v
d6l7s9k4Ybpj+Nf/v/QOoo9LeW3v9NEgyPSRFZhFbx88Q6j0M10wo0LeE34KvFSy
l/Xd/krF1ufJkacEhFRkd2P2sHKI4VSMQ38mdO/Xx3aMdg51bdbZtNJsyYIqsV4A
mo7s1wlsTCvpuMQPCX0TdHF9uy/xM4NPNcMBPz0syNEIs1xfF0QekxSt6bP4aHNK
qMbHN4zzcXg+T/Ypvohxii9BBIOwuUbSv2vGDaac/GFwTcX98AqlZ1xTGIz24BxG
AB8CoYd9rgQuAFGrRaZew1u/f+9Nv/V6VBN5QA4esF3/dJwM78gALmfo6EBUod1o
otiMnOBL3b9+AacKzmW4ECngfVyaRLGMRsqT5Zw205anC115xhX472mZmiD4ARO5
IJRuVEfP4GBqcbt4D88NSQN/Gz+UFsI1hAb4aEjt2vYECufvrSPAMiJlmt/0QCVP
/kCXkf8jvgyFEAXTSyIe5Wx/FvfdgZBOqV9ZWWnfCHFZOx970eDeJ1lKzP0CCY0p
ZMoIi2hF/7lEkTnHb75tenM+Cxljv32FPru2bBMHwmTp9qJy6pQgC/HBgDdr91Hz
EpDL2kuZPvilhpG1PPa6M4aF/llzdcDQYgXdzkA6PQ2fEdGTzF1RDGUeY3GKqlWN
MeYkZ9YGjfmUmjI3XsjZldrTRS93t+Y7oVsmKy/lue/iwWMBEVwt4hC+OL2IAq9v
gkclTtgvqtEyTGkT6m9aAXlEKOXQm8xtH2X4vU1e/bpaIT+Di8rabMOJR2fibjUA
b5Z4JO3UD2BhxnCRfpMJ4gx/TRMqREGo9aSUAE6aBiJpKDoxOKAtNxt1Jywow68t
hoxWAgeyXtwXGR+IeiOEcKFAACXTGwbdZxVgk7hLPda5W3xxw/pzN+CGs3Y+DgkJ
CeZbh75VN5e08ouIqQoc/UDFaR+CaBgpRQQFXTIbHOm8ARjGn6srZIY4Rx4VZhTq
EM/0L8+fcco3x9/TWPuigiiur0Rl4kNuEVmFhSsVKKWljqEkNZpWELvCR7ltToIk
e54RYSQQCMQ7fnonOac04rHqGZlydYfyAtstSPipJgI+3UfwW5LI3P2fuaI7JKHr
yLmXazC7pVrKePWw3s8UDKa/AsRkX87pnbfBo8fD9wJ8detcrnH02dCAVltPQoq8
6E3EQYD7IpISVHuiYqopG0vLox3LCt78gaRa2iGP9qtHlXkru8U2NWK1KU4uTAky
9jl8sbVUrGdubPvpBoFY6FDzzaRePSAN7o8WIJcRvq8XkI+fs22CX1Dydk/YIsSW
VUoUU0mo+98DeufIyktWe+q//T70PqChn6QHJLQbE7fZlZAZ0hcj80Vdj6XiTCTz
A37OVMNJAFOR4mwE2HKiHUbOdFNyVjmPYyWDZBre+szvV+eFi3idezPMXdUpIvuA
1qmcCsH2+fhwLjfETDb+sxJWBlDgq4y3ZtLXhkgzgetFxP6WGQ+TtfCdzf5Wrgo/
K+HRMPUcZt8xRcvnjHta2m/M1z+/hR4Q5PTre43LoovqxR4I1ftUNmQmClsmgLRU
gd8GlYC+Zu7DlLNmnSRVJVXOBAqzQyVNZD6OWa4disNk+EqRQ2hnKsySFyvnlN2j
13UIuOKzzAMlsYiuGSVd5n7oGW+Qozwki8re9zn9UzVdc8Ea1Zo/vNZ2AtKYPy2N
FNFG6j+HEUxCnjdPu77og0Kx4kvJvvXBYawEEX7hG0TlXtQNR/L3XhoxYisw7dnB
rTYif8VPEWG7GakGw5smrM281RG6MIBQDKryDeVMKuCeYzsIrPsVKZhIYkx1y83u
/sWbmyTyJPAKBlSLuIZdB0Ow9mRERb0DN7QFQNJ9xkYrG7d5d4DskmydQ08z2wo7
uL6nP3+aX8XkaKDyDEz8OVL4+nV+iUmyHDSiij2DmEtmOQldQ7P3ui7nqiTdRaUr
G9ljb4cyFaYcfr9lT5W4RpG+9oOAi3jDeWaV5ZFh9mNe9AKMP7EHE9FeC2tp2xpX
BN5qb0nXXSXlXnrlOxN4INRaJ6jJFVJdswTABUxLM2Rn6vLUhKNbzd/IajF/Fczx
rL2GSo+umMs785r4GZrdsPtvoWmeB+DIDTGzItN5qJZuoxz29qU+/KpZoMq5LjVa
sA/OtEvTMBwgkoIGAICXOQRJOx15tAYKhfprbiHyeg8+6FUAOlGSASDwFqcVVU9b
xyUl+dayigkWRaVRPc0WJg5FLf24qIknszcrDjbPrYUBd1825TiqbxGZKSRMGg98
QaTWOI3BtgkQvyCp5xG21d2BueCBAIGfJFL9gheWb2LVmYnD9c5bGeoOkK7JQ3US
pgy0ulKrd6wNqZ7HrxbGq9acqfvcj//KbaFq4510k0LhJ9QpWRK7yZDezwM6tgqC
GBRbszqYCARLBMzSLWQ0ZayYGlkx2guJCqK6Ff1GWcHKKtk6DRUexNuhQqM/bpUe
zVxC8mON6TgXpG4p3O9RK99sXzyG2swQeegjXYk2DftH2NUXuz0QlsDxBcmX/wQ/
WowMcjBK+fCnpo4Gy83MUHhPGjNlYt0qJCIJm6GRQ86EjxbEsSVv5ay3la7SlW5A
I8g1GIx0IbakbhPqXc6o8ymsmGZPjTlq3HfySXvTQ8q9kvpOlrGfmegBuF1gw60E
zXQs2cVA3eYKhT8x8ELhw49MjFT50jbPegmcHDLAFLURY5X+0tTLNC0Qi4zfjyba
dSmZoSGc8b1qQYRUE0O/bY/OGOyGYc+72MhmlJEBEdZQZDgHlBENOIFzUdcwYzj1
uLYQuGIiyutbh7YSU9OGaGnEgq1AYl3iBA7px7rnEb8yIySgDt+a9OA3s1CjYGpd
UPtqs+etk2BomNzLxZswfOi3tw/mF9DKhi1LOyu/M01TbXdUzEVjGEHqemRu+VtO
YnRoKvNd6wi/OnFVi4dG7A10QR9j826aPOLt95i3QYqnV7KQ8OMnystLXP3Q07CE
jXT2KepTKyuoZD+j7/5QuUh7O6OwNLWwLLydxrtu2rrOMP+SrieXpLmIn2ofQZ9/
wcDPX6A+5inBhBZKD1l8tgNTTFqze7A5ITxZ1Vht+u/Il5AZU7PYfIfcYFG8iN3B
6s3T9vQjTOvOvNhZCphWq/4EnX2mRJmJJCZVc14PQk6PA+Nlf+Ld/FuscmB682d2
dQmGC186kC7krvQv4c1UUONIlKk359ebsypz5UiMDM+Pda1dEkBRdLp19XkuUyg4
cbAjETfeMcPAnwIr8oq80zZO4QqXfIlZQLYDSoQI9i2km5JOMIdWjpmkaNGY9jXE
B1hzP1G3xh3ooxjzFJSzkTF8R3eyk6mJIhJAjwVFu4+bJlyNt40uvns8LT652qgz
uAlAl9RBSNtXqQUwUKY9JGHzM+jrXx7RWS/jouC7zH91FoqbGuC5ENgDTNAHqxao
YMr0xDvwz3W6vj3Qi7yZe4HRon9AG42esAXWdN3SzVXZOo/3f5V8PECJHt1/C6tf
uLEsYvznmtX01lWgbpNH3PFfy70t25oIWy57kQcszFvQvzIQYhXGMiN+uISaDlc2
VkMui+O7vXb47qqcF0dNOEfwCc0oySXqEERjWsIrIkDLgtJq3298nj9EPBJGzHfU
me1/YN5ZcfghR9qZ7hCIqK6btzvDV9qzJuVn1/HtQZkAO19lgrEcyHhh1hibUC1k
fYXerCkDcdCpu17YT0BjuL3zxdVsSm8Sr7uOywthjcv4rUYL6jSBq1Q++eHYk9+Y
sXU1J3I2lt3cjdCpubsb8I+jIgHpHV8xz6taVZHcUgHMdqejBwNGjOuj4mooLHCI
ozVloE+uUfTrj66EgROZEE/Z88Fhq5C7RdXAaMhUwHzIc0AgyX5Bf+SujDWCiA9V
kf/I2FPh2JXL10ENEAVzNVeO5PA9gAUEytQly9u05ophFH95xATOWnwCAFHP60eq
GdFj+006wMrADhOGLrh9+hVmbZFInk4gWqhbPwD+yqtpkNNzPpGmyOz4Le6JNEvd
lUGlz3LiFF3q/rI+kUWcfEyo3y3Pxgn4l6Uch2u0GXnMrecLtw49Isxz5WYUC3TH
vAKsRAZ/gZH8EGSYVa9aDq4FGUh8sYFVU3w1G1WltgCIBPBFJcTmgJ35zTPl/9G6
Q53k8Jw6dIO6mxQ3Aq5saIgG7bCkJVs+HY+NE4EVlWGJIXu6rqwMyOPsR+3vwEy6
+8GXbc8plhUZjDaHcBXBvQjljY0E/41iaD6pDbXlbsaZxEZCFx0azR3GMrWNGvk0
F2sHF20avxTZOpbMGAxK7uJvXVP/VWayLGfIo/u4MPd93Hmd7utKpGel4p+dS/OD
X2636/RzlmUGOHrDJvffOrV3cCElc3UwIg1uPApGPjc28HQxJ0l3G3yJ+xUbFas3
yK4WKSJsio32s5TTA0WeQmKiICLOHCoikt63wH4YNyoro6rxHy+ZTApElqqLJEBt
kdnsHmTS+jXSLi0fvboRYHYXMZ0oNuJMQoj79O3g2MGgnOL7jjCmgxC1qtpjvVPG
kguiyy9rdOdllr25fuxgx2jHdH5U4JFJLuVfEgKFhn1ddtMvqqRdQ2Gi3saWzBd1
ysvlAFcBKe94QEupmaTymWdUQ2q9USyIZeOt5c1bg3xyNs6sEa7inobd6iB4PntL
/NMXM7/Qy0xyaBYXkbAl+0p13V7KqOGtaqgNJ2YTxHxaQXekg+mwg09vclJxfStc
ws2K90nrPI7ZXF2XrhEQY2+XKG9A9OvNI/VK1HUcOsLdE0O0F4pU41Tu5fcBbEXZ
HqYcIktQCvt7W425b+E87agsTH8A/nwDgszpE/avhWLmJRutPp+cOgkNAyPjLYfz
uNmc9nVprbesezUxtI5spdU2NbmRu6hj3ful1XAxxsYFK8T38U4ae97crdCEzZtd
psPiocuiNjMVSEEecBPb9uBuMwCwZdLXKHq0VjOq5V5tVJQPGBspbp/CTarOjBzX
Xh4r+Lg7FpBpCpPpYt564cHPemwMNyCb5TUPwnggHSZ+6ixDAKBGUZJDImVIW4ld
rApWIFv02MA9vg8957n9mkhtf3/J7BxgIZ7neGoeX7G0PtG8TJt7ldZ8rBirzR5y
HnOkOnR6t1EuFymRS59BviJPK25XTetwn4QKli4f9bA9evtgOu4VdDW3MaU7oBJL
0e0c6i/gJQLyy9yYZU8wtQMQB5SJut9nDfBmTMH3uXzlwN7lbYsM1oRRwALjOVe4
euUWG3HvB4jXlVSpX9WIR6ebYSgq3+lEVHY9X9NQv9fuJPwbF2CNyhNtm8hQ1or5
gYnXV/zud9JA0KrpLAoBKbvCOIKUe9uurhhzEQmuovKCpjB7fxFAq91NrFxopQGb
xi/K9NOc1oQhNVcFgBm5ayKiWH3MeI55wqgsfRV1IuCeiiZrbOt7fX2ZRxK1x6wN
8ne06xHi3q72Iqu2FiQKNK0s0Xkby+cNNjD88+6evEVxwTnzrdX/M/HyLshwOLWF
fNfwuR1fFPqsAhfqz3HBdQ6Wh8I7WyoJZADBzDALncJUgALHX3P1RKNQhPgoDzfM
fSoxYxZBobnmJcwsxjJ/3oFq4UNsYNMSyQZArxrLfoCvPoaFxliYTIXQyeiwSM4D
qbNlMfhD+E3jbDr0zPorPhGRbdbZMRrhHosRaAqRjyY852/FABO8jXxemO5AtP0c
JO1pZL8GXG0xEOuwjKSi6n8axk/MMgCtxjkVLwWGTLQfn42ZXWrVprLhf6Ejo+Li
TZVt2RJS0+vPR3hIBw54C36PJeWuAunbFORnisski2Bm0fzy4dtb8DxHBOVBlEZo
80sQLGbOFvw54FiWCXmtQMfQ9wG51sG5/iLql/Dok37fjrWpIk63uJlInNWVXntS
7CqjmpSgSOSnyHuaTUf2oSlz1PW3eR8ax+AUfIsvNU5nXK7D1KnaspexOUvmDAWt
STy1Pe7RQNXdqFjjjpaPcBcS8RYAf1zZCfOwbdWC76jblLjcaZ3IVNp6G6khu/pl
XqNSXg7XwSFqyO41y2z4XeV8IHxQQaVnPzdb24wGG6rjYFr9bxVim/KX6Cjv26jz
0GZ42CT5JVKwBuLRnGYyuuDi3vz1OCe6C3y2gR4kiI9EgrJfp5nVjRYxsYacdJdJ
cVJeRz9QlSMH0cupHEX2CSxajewEl2uhqpGix+3COeJ3xKYyQUS171Tn1Snn1lHb
50+e47d50/iHfJaOC+jscabKZyJMgBajA5oPkWm5p194cOVmB/ykWsQ49SY/4Mz4
W/V1PQtoecqxNcwptFQOPzy1ClDvzCZTVvsz4bbJiL+VKqyK3ALpAeyWscHmxjeC
Kw+FX758f1TGVwy+icKPxyF0nyg9ot4kwztexspn2ucxqVvcjqDbbNvArMY8UUfb
hvu1KP3phbp2yK93Tt7Q3DY771FlPuY8NgKifxkISwfv7lPccjTacBHje5+Tj8i5
DqgQDUtSuZjOrpAD0sR+7JGiHFBugTtrBZMJHW1vkO/4Dqv27DKUNrfX/77JQgw6
zhcfabzlRGwkTfaYWTkJx7cwKi9gT0HKvUv80e5Hi/upQB8FD7ehLZrhjv86KINR
HrYOKosuxLdZxk383ODonhQQwnaIWk0IRKs40b6sbrXz0W1MSTvhBYfu/uS5UAuA
iJcwE9MIxSpSSR80o21aSu5AGUnz9En8TP/6mHvxzGWRFtmY4Me+GYboto2uho0b
oHXJhmSxhKCF/ootgRRu+jlnt4qDBOcyYCk2rEeOLxb2A7vhj//vTyNFlvNV75oZ
ChQnHLe/JdJp38y01VjbCnP5T4AlyinD483E8uYtYAPVJerkhg1sj+wTtuxu7kuX
cMDpfRqpls9rIApacCVotPpTE4R+HingJXfS/oSQcIAyYqiuB39aCCCso98XoGx1
CFcuyGaIoity8b1mRGDUs/1mkr6ndikBkAyhiIlxeWyezKhkKOTXciAeWfrQvaYI
2d3YQ7VOBfUH3pSSNFV1ESxfTsFwOoY83e+aMTH4lSMTgm07NBbHP6fGJtYyCnL+
faIfuLfE7+UcYJyJ2xAr/kGDylPfFyxMngTSgDy5qh6CyKMJUyq1ZJsKU3HZMdwb
PRvW1JMyHp3KIaPMZMFkUMHGT5I4Gbkw4IMbemmfOlFDkO1ApyDGrczW3GiXplnU
scVDINN5fSsDUm+CgI29wr9YiXtt36cQuoJsdYr+o8oQonoxzqoTXJ8gMXHBwH9m
xfg3H+6dckxSxWv73+Rl8RMTrAYv0Ahe08WeqP7pI3SnlfBqnuxyvX5/suhBpIgz
ylZzDTcXlKMIm+9Vzdgxdi+N/EaFjVniiunUJ1Rc+UADBpsx1EBcnFE0EYlE5m6A
LxnQkHIBoxfdYiQF8//hqv/sH/Maw7XWMtrBNfOeZSjeims+afRGySoIevb+ZYFq
UyUGHLwIDy9xkw2Q4EGKmnUL6Gsqi3CakqXbmTOR+hZGJDe8s+eivveTJANZMNRt
DrFrmUDU+HPaiwUsbv7xrgUEdAzU/yMRCwNbBk4i6lwLRuMhScSvKE8h4b1NTRZn
6MjC5zozn/5JTXGh4190AVHM0onnuvgTWut6nh5oBnLllBNOAxvXni5tC42JT4pA
Nj9rFJ3s7KPY2Kdbd3OH+vh9ZtkgTDkKqZOloBiXPY1ZWeKeRKyThtCgTys8WXV/
tcbPRvP+5RT7/tFwU6UzF0jySsdivX5Z7R5qs2H1QdlMmvP9tAg78u0st6eNyBLz
I6dd69zT++ACzjyUmSbVmLF1Lbbf//15zWvAMYnd+O4uwqhZQEMOzMRpucKUbtHP
XBAJnqAIGF42oEMqymxi16X/b2kM2afb1xVPSo/IaA4U3T5quvg0UN+9FsMSfACo
EC+U31dsgB78hSj6Y/SINcEiA+/cIfDrJ5NECtaQVbm1bmKX2MvBSg8hzwuViUUV
mQTr9maIrVIQGNe5QjnyKEsY07CHStHdQ/gcEuWtIaa21Mvvo6DWx6v6grOs8mSA
E4mqDGRVQnj1SJls6slmlELkMEIHB4qGxEqX21pAfTV5YJTyv+n5baaeLTpoyL3y
vm89d26KEwVAHcFi+QkxRdhUfFYCqmdUuBRj8iR2yq8qffsRq8NGrpr3x/2gV3AJ
xznJv8WUJ41VgFR5QqMoTJGJKZJwZWks92WngNKu2lLlBZG0IdYU/mnFbplJhHA7
7OlerFymiftzJ7WMWEOatfv4MmjCoYIpogSpMmyz8JGQj0CF8DdtQhCri5W8x8xM
+v+pire5R00zRPz397QD11dsd/s9Vc/8Uy3ZBzpT0ToyFRzlVhicAmhy0bcFp74d
GPstl1hC/k668vx6bpG4AXlf3OjMijkfkFmr4AF9KPB4/fYyhmJeZVoeqRAk70IJ
uf1BwB7JfLmP0X8Epv5B7KYF+c8wgoIQK58VB1JCrZ59BAPLXip/h3G2XJFeoNZg
budlRip9QujNckU4L7RJIogl6VLW30O3cDyIH9fmQ1obBSYAIp/fs4VqvRgr9g6D
sD4UYtyvmma1tI7dqGkbCi/DETsX3/vO1MLOSfy9zzq/02pr3gN5B3YFbH4uutBT
07KDp2Y8/EfbHBeKUpJmHJ2RLW26gueocaAYT6uXR2q9h+lXcwUKADEFQwMEAED0
r6HQFNMpp5xXPT0H82g7L8xCPWw1a66krFSlNhrjekUt7By5Q9R2G9Nd+X9EhAGq
amfFpMo1mS+Cro76aUB/C5Qksn6fP9qOaxLSmBTJ/FsYi/hNmorPmW46sI3QaSpA
hvEm1bFSmvo1nI7q81Rp6SwII+c0lzdsHQPRnjjkUtBxVzuPikZViuSH5vlphiP6
rhg5XX5oUJTaYFTEQVbjn6JSvBrtvGSexN+PS1IA97mVXMtNDARRe77b6n6Kstiu
ALeC9X8vcJkRg6MiqF5qG0FBSPqU20H1rMYSiN3ysHTHJVjEz9BI7hbpEg/sZKR1
HvX/7N53Qp3cFLkwzlKpzl4x9qdbAKtV5yW88eyER14lL7oeTEDZk30RGbJp3tjC
ExdeJccNBhKE9XHci6iZU6qf/ruKpmM6IsG+6HvlRc9kZdXbkhiiF5Mine9RGEcp
HA/Exom+VmePzt98R5SZWS78XyVjYPXLSLMeOZZxHLMLW/QR+QItatxts9zn3vFh
nFLSYek0dUUyihCtaQ8r/Io5IL0qrX9rHWJ0yllvqJUWVOYi+u4/zYH6mJpZAjp+
Kq7XXALCGEpg0tefkXLAAl8TQN6+CxitMCqN9xba0OB6h/tCvi6C3z62XkwkO9W9
3AYzGyqNu7oaimXYd5qT9wgDWca1nIRJwLGCIjjsg+LtUyYP7iHq/5EB3yszBYHh
N/bPJkIsEOeSCgNVrIw75eAU4PmFkGNgPmalgooZnyTjKoJNSUYwyjdO7PyOsSgs
vSSfjRHObkFocr+qxg8vpphRTYWNZ7k1DgMrBjDFI5FMHvCinUWoucX91qJDzs67
Eoi5piTxKjyknEmb+W5se8p+MzW1qBCAFhfEYNGVnZrZ84klhWr7TEq1aGRY5VIa
BJRCsg0ZJ++/gHJZG4Dwv0l7CBoXVhOG8VaO/hcacy3RVQS/4lt1tNODP1+TiI9T
ZjBvJFWzsTAa3rZD/2pogaZKzaF+qxelzgF0h9IL7sswkew/yLwecQ88F6FMZLiC
1knbohR4IsXfysU8nzVqFIDqYc90jq0aiA5fcRSh9xCn0PxcPLeXsM3ux5hmf/cG
2P2jGfI6iKunqNFuTDpuo9a5YY0qv9d/wGJzgDA2K7ntxqJZAq8H1mcj410UUT8Z
8MISRDqfn00gNhaooVCCNrAvNXCSrQa8Sf7UY8ckHENG+UPro/5bfrbEP7FGx8ho
CAfRFNMpkjyaHgahNSqKyfkSeBuChKs8AZh7zxJPdITxq5IlgpeR5Z/NUPJdwvLQ
PkryAe8ACfLaVmu9k8ZJDg7CwJBfN2Bg3atwpzY2bxZ9QMXqCIfuhRYyYf6kmkIe
rn/iYbRSAd1dTp1oVWOjXFxhy/NCADwJeyA14DICIxF/zgqd3WEROwk9ykUzVMJo
ob3WU4CN67tA7OZom7jNE44xMWtO2F4xtpRZYACwDDRTI/amXWIm/WEScuxVpx+p
0CWUMk09s32vW00Sz3830PlSbmdfE1mQTaaoH5wvJBUqjDwicXcxqTIF/CEjn/Gz
yAonlHDyPc/gVqtfYBtqjBfXY7zXwPK8vWIvGiTP5+dYq4t2VKQvcjq9MDDsUrfu
Fssz21b6q5k1SKeIsBEV4tvtY93unG8xUGsG6HgWSIU2w0DO+FbvXTpEvAV/Up8F
uzY8flXwdJB88N2NJv0kKyFnHVQ5NGI+IJx5mS5DEUzjU+52ZoHLcoG3NUBkJw06
cwRjKkszyquETP7WvJrWxT4svAEyYvAEV9ZE/Rh1XOOWWbc3vhizJuAdLL66itaE
zuse8DBOSg7DFLROaF6vxCI9pI4GRMyGrZBGrEizIeM9bp9Ms1Mk048VK3I5bwgR
uOCHekhnHtx5UOVgg9Iq9syyrflMiRwBkZtWfseKlFtKayR37ClkkldRpuaf62Es
L8bP712nrit26LXRIxzsZ5IkEAJ6S4r37O6XE6mwtRnD6ObSGpbllx8vygsakxAX
Q6nkEiHiU26qe5WlaWAyE3KEcdIU9ZKb3gIgAlBV8nOCZier7OsbdgWnbm6kc6xJ
H7cb9Ekt5igcK6q343CADyKePz202lJW52f/kisugnheAPNyBEXvLGHH478QOyJ8
AFzW3pBS4QqdghG2skG9tM27y3ZdzoJKTr7NQx9Sun2goiBSLl+K/pfP1lbSpKju
OcSzhtCDi5A7zl7rkEe7uuxIZ8/o+TTBnmPkQZNllV2Qn+wFgo+d+34epY87bQlV
vhIX/AGvjM94n3hBcuTgfNl8fJ1D4fyC8w60cwGRD2D/WzI5FOhlaYRj1ZIYiof3
/D+NxNYVWN9/pZE4yn9DZ/mod+qxRuqw2XGmc849ld6S/8exuDRrUfSm18CbTMmq
hA/cIg0uzpZ4OfFM1fY15CVYtk19D4uber9k8iBAeTtXpiKUwa6quViov+9OOx+h
N44f6/C8SWi1CrANomGpnQ8SSZX4IEGwyLt/uOnZSPVyMufareuVNhE7fxwlv71B
k/FJZ0/MLssQ1FdaO8IwmFovUQwCH2BL3Mv2EIVbyOQyH3CvFjhyAv1282dtU7fA
DJRcorurFfT0VqT2BL5xpaGVkiL5cCa4Wkc9T7B9xwCbLVRb2sMG4I1j1/sjShPS
KU/5EgE9U2tkJtBBK7uhRBeRFm68pvYcitjo2/xOUE/BnDPw5a49DwwvqQEPjQl6
s1pAdsGvHNySupNlk8EeHF6HbFGwCkBIEhT2eEDP75L3JtCgpd4f7e40B6oDVNme
FDV40qx09PTJlgCfPFfpP4fhLdrvRL9w3JJC310dihzujM8Kd0KP13kkHc8akcl/
/nTblErRAWN4GiTPfI74RW5elt9MlE/se4z1XKJuaZRNwTlaQsEIlM9Cbl8p1FnC
a2wCHY5ZPHRc1EpxrxtnBPzbb4u7YoQ4RNhMkhUT7wKiVtbo17kEoIrZwQkWxU9a
Qu9QvF+lTMpopa47I5dBCfUSIUQ5UH7TZ6rnjvDMHNLnsk4hT4c3l3w2kxmlNBmk
t1OKk+BaulljxKagHIE2Y860cAkVacKVjVvdeIQJfHe2TuxQzd8Ylk8Ta+GwvRAL
q/3LVUITGaRVtevZ9tUviu9y5pr2O3aIUedPP8NfOfXq9s+hQLP1DRjkLCy/R0pR
Wyomvj1rTTWNhV4EIIN0VntQ9kjCK7Yw0qbBcUZnVkmzkRRcWYJRdUecl0IpfIxq
Rgd9F8ufN000ZQO7tjK52ufu9hfajp54Nha8t2jY4i955DOQxu9z8nTLfDFn1jBf
dVbnAQbW1fl3V9ypAIaX/ROW3aeb+lFz314j2if5E8p3t15R00G9wKKLwsV7hf/5
CiOaRg8NXcqgKM25XLRY1f1kUEig2JrJChBT08yXMSIcU5RjAOIijG1IofjczjGU
EUCP0btusuHIzmIdvxaEvkz3jmbrgkDzblmXxmWmaIvnI/lg/vy/pJXsSVHYyvc8
GBXVGCJU3jDeqNCewUpoSqjtDHqqRuynIRWCg5C1qkH7sCjru/enHM9wrMpAbcTX
5oaLsbmB59fd0X4yeLoR38DvGBKuvTm84+z6FWoVGlQdBhx5W6K4dCAffCIArWFr
5WzAB9TM8LrMVUIBuH65p9xoHniEhZd9QLdAmKM1fSFXD5o4jP/DKRf01jaXSsqb
P/HINaVJxKDkYzySHLizuOW/O14vdl+QYSLWl9WfdUc2squrTO34iQhRjXukoVXu
Bo3ThNXCCjfQSBa2gsnAt9RHn0LA4GsX8E9lIc6M/l8T6Z1UeDkpP6C5xo3IbwcG
IcnwGVFu3t94GYjLkq0c/BiGQ2kd2+ur19IbgHMB9dTPXdRnTiYVLFHE6BRYzJJM
x542Q6bNRZu0NyPu8KXYDIIy5jqgRJrIpdpJze7n0GfGwFQsRnVu6LBRPxRWqRma
SA8WvEpGJT3vTC6iHC0xA21Z5eZI47Z5a9r/9Rjfj/vVbQQ6BXuLioGDYKuH5SqD
7528zOP8YlpL8QnFh6lSb512w6jgCIIJpl+8ZxEsb7sesC53qqhbmw8viGWdVzJp
Pm3iy7tQu64z8a+H//Fos6hDy6/BegerLgAuyBFi8k/cu9cffs1avfiEMLJmoCCk
89tWi8jSyHyP+hyHi2Qcpg/+laZba3aJbyA/slSsVQ5aSpnIvhfqBG6FVj7v5bex
57s8qR7kwEW0/OnJCqDPp3SyweukeqgBdXBR8C7KN/2lnex8wvYmQ2v3BQKe+SXa
OBk7H4JWtJRZLWBpPIdO5xJK9eUB6RjNCaMK4qSRnv6YvljNoNfoRLkHGxNTYwv1
BXoozldlnh9X4V8ddQunWmhl/1kt1pQqLe8dkEB3dZg+SNwjJ/wZ7sSQ5AvG6PPA
BAo2lSJPXTa0pG07QO6cEh4eU7XJByyUnDN9iNEGiiiMVddYSp4hCAQ9w4Nk3gJV
nj1gGIFVEDWAG38FKWwkc87DEoZBjO2z2us1YAmmkt0xPLb6arFCXUvgbUzGNwFs
KgM9ooejv7wfh9LP3h7FakYbqdUZz5+fFCuWVPaMM1ofcGDRc2k+eyTgXY/5o2Zo
+ewA4xVLPOxZYC7wncb6okflZOLqke1IG/5BD8IRWLN/1+w68upo12FrT0bZMSKs
NuI95zT5UmxmdDVf49+9paRW7Ly/yHTAU+Q2K6Bx93KHlbh1iTRJbvWSBTk7FPwE
qkptNmGIiaei8sBFuHUmyyl+ZweycQyMQCvuS0reys0jLo0jVXLH0U04CnQcJKZ2
8suo7G1eR6tPgNC9mC9lCNGYt8SsL67DV1XxU4Ek3ak+Hj1LuFIIEf5rR9AkpY7D
lcNBExVlzcw36PCH6N41uG5i05DjcTIJ6Hi02rad0Sccq2VISfxBv6U17dLwxZBt
0yKIGE4Udrxewz77G40npSY+EcWQggw+lbHIioCp894L97wCC9avGzIoD+6HUcWZ
14lTK9UVeUeGAO+AAptyf3o6iFF9JTczTVq8DytJu/1FlavtHkz6axXl+0L2FM0M
Kh3DLhcwQjkqYMJZVZjVXYPy91umv4nhb9xP/TsmoFZG5UE9azCl7lSYD2DIPKvx
IybadN8htxxXTwpvGWCU9lGWpNDK1Wwi3Vux8lZRiFPd9qAkE4OWlP84zMPL32Ha
x0GfyNcVtHdJ12X0NiMtTOUUMft9KswUR7U7PMZ2B/6pf83NbbkHfCjKGVAAMD3n
QV+wDvbgGBrOiFnW81oK5jhqa14vodv01Ys5B6c5GDwoX9fx3tqTmsGQ43I07Hms
8EmzoiLAY+5I6O9l5OLBJf6isGXTvG7NcusgubLpr7VicQn3tcm0IPRZVid9vQWZ
wdHWlxjgecNyBgp0nTQ4h90r0l3i/T+g1EICZgQ7k3vQ2uoeO90z3TLip512RrAU
S6aehLVYq/06Beok5mY4Lmc1zEf0NRdiWiBgmidWvIunPrQmqWrbPWf/bmn2kucf
zU5oX5m4jK/4xj4sVSPIz3AySbY76bNnxx61UkrQ4ARDVpjXnb3Kizdj08QiqRaQ
OQjAuNgjBb5ebGfo2e8eQZ2u3KmMq8u5hi+9jTzanca2lUYV6XxV1wzuKLQUpUUZ
WQ2d8jMh16+6cANhscI99/4t7wQukOJp/4pbKTKrc14Ymo66WxY2FZdnAHPPQZ70
3WQ72+/Nu7oTHkZZCaZx0jQPKCDT+a+aDkI9ifvJC17jhLDnVLrBpJlr7THMdfXO
9cB7Dd9Mp5o/n1Phh4pDK2Mbquu7NDiEjsa0/nxmAw8XpeUuEisBA0hH0Z9n+Mnv
NZj6hPxILkdd6F+gfjZDBNk6NEHNxZn+MQJqBdHHMPizJG5F8279d1h5c/0NcJeg
iJMi5dsCCR4WubB3+CQQK4URYL+3j3jFWth1xr9Y2GywV8pem7C3JhCahHBmA3NU
1+pjVVcolG4nAVSEGEfp/kuZDicpXxn5ir2CrNCheb7YY59T4frBxrTp6YiCIEsD
aqg8s6uhuuRq/wWyofLbuKtX/8vbGr5MK34qJbpgGovue3uPv7Ujyq6TZtIIpJYg
FgrP54iqfzzeCbhQY+1gr2cUVNK2yiuX4bEuhMela3c/NDA2NPPGTRnbQ6tDg4EN
j1j7xd5jYe0ZkqUQl6Nd7AKgyQ9yNU/P09BF1WPW2SFshQqOO/aAwwqIxE7kPE/k
jgPLHKztcELL9ulbkphcyOOldouXw7cOxO4IMEcGbWzhz2UjlhotJyYSR3yIsQs9
AbevpuByJXcWY9lb070psIinQndPAVtpOnbF9fX6Q2ZO8cUskXBYz2Fwry5WvQ9R
Fsm+D49ZenhP+iR+Zz92ft2AYiT6Jj4r5pFGzyvLb4gIKCHrs/bDZTeQnsre7Kav
BvwQ0ZoltX5VFkpW/Neo7/fk8znnv8a/rJDPNgEvIr4SF+2W1LBB/H8ZhKr0ZmYs
fPXWGGmflZ+fGlty6QazgzPljVmW6i3B8PoQOT1dOmlT09x98MDE97u+0UFtMg85
7kN7/nnPvbbTgN/MBoWTxAnLERze1gxUK/gMz0BJZTCjCMCJLIqrGukS0j2V6CW5
2TZa+4uzokE2eG2cgQVb5jBZthU7uVo06YwItq6UfmqyMTeG3iwE6l1wChEXyWSK
tBxceJh8t66FeOjRaruvokNiUAgnFTL8nwPRB6vQsSBb0B/vsYUE9KNphVNrdVWH
dzi/mbFkF4wJY7ZwSNO6K++fHudRX3caLPNgxPmFck3A3aC89DddDvisf+CgM027
xyPOulN5sIxXWSvR/LQYvgbmmQAorjupJqEuW1eYEEw0FzjR7OAp6mp/VJTdTZ+c
iHH7IcN7lh9IpiXo6MdfJ8HrRjprrKeDxTJR7ab7cczBRW36xH3xt+CQNuQvBvV4
mRl3kHmKTXVlXwjWZsSpkaz7E43qi/z2D4o4jQbRZi28qjPE0Yz4jWPIUyA08pYL
bh2uThCnobIryUEGvjGfK+TOEfEl3gvVsZ7rS6HpDSLWgSYXIB03WDp6F71/uHTw
OWlRrKBpQLKhuMz+71v9qFEtkNBkktfQrQ3WaiDL7/DLbzEpavYmkEOqTi56qFxJ
3/0XXs4FtEGb6OaXXrFK8d0vfr4VL1v9qhb4JOzQGMUR9OinKqKQ84aaCIMSIvVL
4JeZxb8BKkiMSdYQghLvsxsQ4TKAXq9xrhr+3pkBqvh3FABtaSLy61HrKNZgpyMh
kfQb61y512ZIqh9OIcqHwif8E76wzaBwS7LQcNlZyRWJevtH2+lFGiZzqiKUEWbI
s2mnjyrJdkHZeCRFemRGGM0VG9FctvzFUC/wHKeLSvc6Hm+0cGlppFxwFNLO83Ub
QzNBsd6xgVqJ8IdMuFBWgxhLARUI3PPIxTMPY4koV/3UhFRRgKerZFz0T27dCfWF
SoNavP9VrB0i0yL8hRVlR/mX6Du/t8xDqan1uUYz6DSnYeLUNQaC2vg0EhUS2fKC
fdB1SI4K+tmAZaWR5v8iMme6elWjMhqBePEflEzaPnRqFKZ45PxsXKhZLBBr3zzm
Hz1yZS2mSDowPBxA9EZbN6ZEwSjEgJVDAd19RUQ7DIFNjfBFupNkj9CjW2Vgrj2m
wJ553MXuz5QwjnMcjT7sC/k4tcuc2wEOlgA+8UTZWEJGPJktef/WK5XSOD+MaRpX
j6/1vjCW9GkirCoarmJGDTI0MkHeZTdcU9kZKna3XVbjamwCEQU0f/8TXKGLJ5Rs
b1AN/C4bG9qHjpcCRdF5osPk+y+z1K3kalezDB8Q2m3KbApqyz040zNdK1UarBjy
OOOySsVKeCqUbuEXSk57xw5kLqh0FIFEM7xsqPm2gjXc3M+T3p/n6magcabJ1hXj
crZG3agzoP69iGm9icsLt4/ZpRoCQM3i0l0eip5gd8Mbinh5+kaWu+W+nGvYvy1x
H7t30AC//oywb5ZracOe8xiockXqqf1u3e3ob5+J9ZndIr5J05TRCB3cdQW4kP4r
1n0gkWoeRqNA5aIsgMb1hw2q9r9wCkyamMDgK2OZJRyJeh0aCZlCVRSA3PRLUwa3
dQIO54/o3JJ+SxANbq6FyEbolV6yja8DBiLBBvVwW+wtcpr9BmqELJUTmzqKhZWG
IkyEvYqEH+BxNZfLplznqtLqjnemNYP21HNFSaFvuOYkCqH8RJHXgOvqLxVtG5X8
fWhxDdymGhyqeZkRMbqCj2ms9NehtdOVAfXOIVsa2tUm6sbvCPbB0mK6ueuX8Sos
inlVDv1PGAos3g61bZBtdxQndnqXAeRXWt1/Y/m1JavyCDYcYnFYDv8ghc+S/5uy
Y4pnsjLrA62Yz4ieCBPUxaH4vERYNAmsoEbDZttN/eppw3gYUjs2yrfV4mVdlsj2
97D5T5Xz3YoW8usygTqtefWNiwQulvYFiD7jyJwjMp0AIi10FyamHckQYlkeccia
MIkUskPRaxl2hB+fRQ3ci6TSP0ViXDagnD4v+jpeyU81Fk0vLAuZrughx6r5XTZ5
IttEp6TOK9bIhgH77dJyrCg5eMoF7cS76Ssd+QpoBj8KU0Ks+JurK9NXclGyzoV4
iWRa8/NPZtQ3sjOehQ44emXqKSrqiMEZGKo5pe7XQQyQIhiSBfYqeUiT3/XoI0IY
24mH86tO4n8OWKwhSvcimFL2uWKu3DWI75Hrk6aa0SV3UkzXpACdgBYlVP3YWT2Q
1h5WOE++awBx5w/LUM/o96XPRd2+ikpSpRexk5Q2p+bhbZhM6XaGgQyfrDouXuDh
ewIoN2vqHPW+azS8sDLIyfBVmOGKb+IvScBvPsA6LVBwNMEfCRuR1AbEEGadpZAS
JOLsTt8SZgdHHypM4fS/3k2nOqd0AP9PmqOqrwkROuBXDf72PFIMVh+FCk1XpoUP
ymQmcFhu3/EijS3aN1GaAjoNuCPYgA2zuWuu8REg3GbWxGKqrvOzKxJOYgAzZWjp
EpzRcXnNhWsCLHkzQUYrsrJY+gR8OWFJGex106CjDMV+pTCoAxyV2WPy1r0M+s9P
NArKy704SMPB1Kk89RX0MNtvoGFc/BJvDU9mF+c9DJcyCYYodk82I0Cu0Hf0dYV2
SqMP7wFIwyGa7VAxS0TOzdAi3iHKgnllOqiz1k/HemzHwYqfql0wDRYhiIbOg3zG
FeL+RpVUVLRTXRnByhKLLETLxFW55W3vOU6i2UkS2PfvjxsltRZdCvUf1SyKheKa
47UVAaMBX6RxN0MryDxCt/ndK/Pd1rZ1zOYARATtZhEiOCFPcmV7ivKzEzN7Dzwa
69fSJJ5qEf2TR3BfgTH46Ejc/EVzsTgDtEe18SXS3Xd2I/TjVk+w2W3xYyjS+yxE
F9IcdE3LYfgXyCgQkYGyRpWmhToPg8S8dfd9+SNIN5i92DNj+ZBAQ+KBR4HmU119
lOdrRXU79PFQIjCoM54hBmsc3IqrrIUIFzUX8r+i361ub4qzMbvJ1sggbWXAQFwm
bWyZf7CIpsuhW3n1wLzktokY1aUPDIyV2gbLwoM00Cktf0qfEbUpC5MraXhW6aiw
L5e+xB6EZG/PH0LCKrEXu19fg64t2PBJALQJtRS7SHpfjaJiGLuT97XiuLiQzZF0
GYgW7tyWaUDOrrmlD56VUhwRNdAHVBqiCWdKAh250XC3og2YVjF2F6t2D0B9xE31
AjmADswXG/jfXJCuQEyC3pCb79R1mNP9Y7G7Zb0p2r5CFLvoOS0T4j1Q53DV66ry
QmdaXq/m7Gus+QYHJd1yhxHF3ahnYdpzHu8W+R1949ZaiRp9NHQvx3kSyORTVPCd
QRDHDn52ibQV8J4K9ffvuf6qArvBjsDJICwlaQHLq6iHhSFlpuWpfzZNkWbR19Zg
2gJbL1/frcOOCWNEfCagy0DAVw2/GUGSLKgeUkXYM276Dx9im+bo/EYdGj/LNdOT
Gt/SGjya9xJXK6n8W1VVcEElj8D0+qqC8s5gQKNCmJG2XQI29zQsdC3FYDsemGIs
Ruw425IwJ+CebN+fdfrFgk89YGCxBK+f8HpVqiPrdvF/wEumCFTukjYrifOUSGdK
ynWzSADsuXG6IistBC8XGnFVgEX2lwfczv180SRmLHeB/fIdoXWpRWtrKyfavmF2
8XfJq98lZnXsEEptmRVudp48wFAT9tKx3BrqaNrpDSXpGWwYQeiNu5lXLlJhFSSO
Yp47CxDKZfWr9ti7sCbplcl2719i8zrpHMg9ykjOtLPVr6RpLMpLrWo7wpSZQfn5
YUDvo5yKy1imKoDc2Q1nhAkzXrBWSJKXMfgxgS58lPqjUhvffoDuc8ScYokYMErp
gfUcG96Npp1WPp5S+AM/bMzu9LU0DzbwsqthLXCfhbxQpm8TU+eTuwr0QVAzOmQz
8/KiQUbyPP41+R1qKUo0kwBZ+ZiAsBHpMEkkIAZQ3pvvAclRzGtQbQ2z29t8DBw4
qWhZPCjRd04BfU5wDqLPOOa6Zcaqt5S15SKFeCxqc3ATL0mUtY7Pz7nFc8TA9tYd
d9GegI7C6s7drw9QA2//QstFRHn3S9dzMLySf0JBs5ZPyQ/xBNn9g9seopvNuHVt
usaqZfh3CFThMdRcAljj7ZiakPCUqO8W2RRPLCw5pKJ1Ks5L+RUChryG6BCszGN1
0xESz+vjLgqRp67yTPR4evkrrByBEv0kpz4x9nxqZ55wjnsM0NgWy5QAlCMog+54
JVw7X9IYCxmpUQVRIUfxUdHJDzZFVopj6VhOL8ZXvnqIgNmdQzOl4W5iiIquE6Zm
h8aIxeoInaRbedylqRJkINrQIOqZSpwENCqiG8ye32RjVVo/dtK5NuYhYxjz0RC9
sm06VGwDDat8mXykSyPUs7WKUAhIHllUJdlzrPVN1o4AypZC6adEVLO+csNMBnv3
dtqLRxcpIoz/vCe3KHUebyp3ag/Kiw2StSCoZAlMdWuYX0uXWYnqCpCvINPFYie+
y+x/KXDNiJGoVpNz4UzhtV69/n51SjQFEA9HAjC4LrqoEw0YE79MMXQRGtNuQPuN
8h1eFtsMdZjGSC8aXiq+4r/hqq4HOtHhKFRtsxYa5N+xs8aXdF9cKF0bkONK236a
gfsO9R+pIlgUYBhNNJkdpsGZmf2TLdvNqLvni3QherW17f2vmNW9thWlGeIfmOQh
ll2quRVNI7xImisn9YPSS0KFHw9rvPWNzqYWKRpSFE4cvCNnEbolgRPr5eiVmEOD
kDZr76hx6AJvoBzwLd6D+4K9YgQW/b/gjf57Ios009RHfEdE4Ya6Kj94jxcW0dNp
CpitAq+HZyjyStvZ9U2xMq82Z6TqDqbqs37Zy4xP8HibGhZm5YBIWieRaze67g7u
Y4JkeRjbvOUpcC25omh8MAXo5/pfIg/Uej0V6ybcMEIoztWIKrzzAZL3niXGtwsT
sVN8MXiELsjJH7rgXEUPrhY8iCoXpTkJEpamFEAur0libfsw+Kuw3mClDQazGFaG
Jwc9IPW2qH7UWK9oguyrsP0TDyKbV0GBHnMx2JWpQ2nQslHDDLxd9dpIopdUxhLk
L/Xb6hR74I+kDL5U8+65zZQguWPFNih6Y0V6UXERdUdM73JibyFPEEMv2PZzQzjO
CAgZ7HJYXe57mBFZksnh/jFl3GXt7UsUwRxCn5rJ8VyC/KrO2PqnC0HYfUgAdEW6
ktXITw/w6VGvf3UpF5cknoR8DMBT6b0YTjxCbU+a/o+cvDuz80qvrvwigJ76IBy8
2VtPpJCfQ9KSqDuoMPj451uqugNevDtEBQ9pONeFQ+dSMm49omJ8YG9t1HE73w9v
JsdOlVL+xaLhU/0QznPXRR/O7DeSZWE/dOPzIjET5GTwQeqAKkIfFMWoS2SEplIB
WBnw2fqFg9IQXlfajsHYRshLla2i/jvo46Gifedz29Yu4yFwXWzAXnUXJ3E6fWRt
5aixlrNlbTvGr0M4cIOCyrmyI12mfytnVeZXZyiHWfbjdsuvVBGiY65AzORi5SgN
sEgv+NR6a4u97ZCilwt+5LgAvDiqVgK079U7D2gxbOBDswp1Rdub69kHOHAmUq2j
nVPJSur+6EL+PBhjoeyVrH6/a0ly04HrkFFIsLFZYLEJcYHmcqywd44KipqsL8lm
mCO58ftJKxZSmYqSuR85n67SJd4e8+EhrMJgWxC7CJf7fypXkoBAGJxRit8fgsyd
Wyqxa+IOTVLpgA9z9e/h2EGUP7qkb9UhvirYXTcYuQskVfuS73j0I8amXy5xDYW1
/0xehO0Uw2kfxCss1EtuamSsaDhvKbuJw3IDIk0YdQeSpWzttDT70IooGTP7zEsr
0trJ6j1QXEcHuME/sBafxFczIVgqyytJzlDfdHD0aTmg0O6DrPS3OcUnT1F+WRhp
ru5hlGRYG8LjWAMHeDpOMGVlQMRELTRsggS7XRAGaO0oLk7q3Xct1LOCPit1ZHsl
lLq9sEPoqu7HtrwzJ2ie4jDp1SRjebPyWexLsHkzLVPu5f80s0P4hXnZcH6y8bXm
dwwhqeDcqXc9qFiNv08kT0m6R4A/9pbpdgcg0PDlI3Fs+nDJF64Ig5jPeVTmyVIP
uBtjydEbmezxuczhYmJ1McWzWGiiIUmUWILbKKo8msaeMt78kvFSD0NZe3JeJLS8
lk3iXw2SbU6G1y8WxzBHq/dJXu1y3c4RfPNk/RMjKzx7AMp5d6YorJoL7xA5lsRO
lR/Hd2UPAvypZ5Kcwix5j30rRlGSKZmFKQTftWzTC0eCW1A3MUSrqqWifVxBsN7/
iiPzF0B2nN8MQYRnORIAj3pV26paTM+fSCybgfh/aKQOtxNq2oFqMXaBvswnF3hg
Ylm4Jn1BGAfUNQCYpoZpLTv7uw+NlbHdp9CURkcPdH6Hq+9jtR0sVAKTAP1nKrkU
U5nF0RZm1QOykYGzwOfNogXGFPWAwQXxeVhTIArp3bN4utODwSlOTALpMPpV/AUp
OMp+oW+M5CjrWYd6xW/AS+OfqV5U/MFoICaNzbVTnPJJ2J+UUD0rjUlJ/q3+HwGS
CUO/AxJDI6eJsXCnH3lgc0uCpP5X/aM4MeHMgtstDxfNiIJWHd6gp/kkK5r8lWbk
aNN02P+GNgZhmy6rlJ6zVKTOTwsbJ9IKmgVR9vFDkfUJSyA6fpMw6awmNUfvKP+9
LV5yrSL1++4WClBU+67WNSMiOuw9XErPoc3JvjNfwssk57pRSJO8wVWFinkPHXM+
PdI4lGl9sbddGuHChSzXMKb9G+x8lI5gfLMqvWY1FM1hUeR56O8DU8jChWEop5oU
f9q2YFLcpT8NdHHYu3X8rJunqxvrHa9b5vMQg5rZ1neiNtZsnjFZk1/YxqUXuUg7
Qo62OVAAONzcqOBUw8uob2dyaXVzb1Xf/p/Gk/jq7ii650FmkOzM0b8KTiavdyGi
VEZvWeX5AaMPZpgyqb4qU9gq7vhgTiszJXUEWEZYoW+xqhgCLASVUFfn1vhFsKgK
NcYLG1vSVFuvXE/cdTDMlcHKJJXqAvl6INIX23zphF92vq2O1XO7sAr/s/YR/d8H
xho49M2/eqFK+kuIrYHD5Iou3Vyo2e6MUESyVfyMzvc9XzFmgahzT5OpZGNdY66l
2f56xFU7R2o8SNmptrnR3YZ3/pdeSknntmxxUwTCezcq90Lr3/EzEdCYQgdhPSdR
MTiDdQqZvoQquExKcHwHONVJ/HlYYuIdqCK3/YZm/sq+FhqRMalUH499N4Olheg0
Tz17OXMz/eJKPoiSR+1NfDZLlJxEEBJaJCzZMrVCu/xIlMLi/vsldYQ+Wp/BsJTF
lbeHv3rN1h5WxPW+qs3xxj8UT+EZ499wDS+MnfHMSlvN1CoPv34QHIihcopLsFO3
YP/pm+kruxt+XTDnBhyE2zIw0dN62BtO28RZK40uvx3nM/wffyPg9PYJVcPyDzu4
m4ns43bWQ9E6Ilb+m+cLmEpG/6mnUTwRJyLzmJVjTLnBOK1OOGHYExThvuY31ObW
QMYGJCPqpOELlhFLpFvR+6pKYoji5Sfibsw0ykCIBtEfI5wyLQRjJiV0vTj28Fwb
aNjR8J6xHLc9+Sg2Nzg2LNxLqQV+4rD029hDGfdF9ZkGXmM/7Js2wA7jnIj406ka
UE1QOFDLiaiIOBOmu1zsxi6ZrD1hYoKnUMzEYuXS0CLm0qJ+c0nZU92YNTtkGAQg
dMmZj0Jd8brSy8YvIuE72FpWx7aNgMkKO4YqPxOWi8v2ntNz0pTujys1KNlVDztF
hf+TQ4e2aFdLz2GR0jTxMftFh3yvYzAUIeEmv2MS1Qygv4T44TxbqSmxKUk9d/W+
fs2zHecO8Dg3xPGLyt3ioMJffJuTQN0pDpv4saGmy0/kfmvev8hZj2QZ5eTLlL8K
5TxfeEkQbTQyvv7Wfke7aUUdWTIEhoG91weY7e/N2LWxNTzB2NqeIp9JwcWEln+o
yNokxFFmFSpuaZPaIQxI0SF5fc8EkOfTqXB+WuDGlr+cqQmY6psxFyelG3ZIrTD5
qrwPLOpR/P8hZACG6kjEOzHXdojHwJHU1k685pFJIvDt0fbbJtw9Oqpu+d4uE9hF
rlE12qaNXDfW+uJAvm9QmQ8TvH6BrpnGrSiWnNC6Rn121UXC2+zo3DkJi2pN5rHY
e3M5QR/c8xF3hNe+wdhgtUjcabOOSjYV8HR0PI3e7yqTRyiiCZbjP9sUm3pyvXlJ
YopcUjL3RMkuvxOAlbKDnZ5Gjfc1TKOHImF0/5Nx+o0e6x5Xb1NLqFYZW17z9Yly
2dFYPCLT2lXBkgDWfgf8O3dKt/nzYBURg94UsRxPJphPhmOT15UL12Wu9f1Tat9g
xb0sX3oowqdW0xCJuY48d8TmqtKth6WwmVQm3tYjwX9Yg/WE9rEKzvsoNuck5qhr
cE3UUG5zJRyVrZVAF/CaiilRONujawIey4hq2TxFLqIq1ioQvPdU8pVrIL3iggBb
RygDiOSbkGd+rU43/IECrRK0X66NCeHsXAbE95RXswyRov9tKuUC53hpHQUqzD2M
52snNRLaqjCgxqyeUm3kk9IkBTbsovFejmBnQjWPYRzlZxTDbile/gxa5cfs15WS
Sf08a6Zdr2U76HJdbBcpbFfsxTmWgmClj/x/Dz8WV2ygSzR9dd7TVd3JjTAlZZ+x
cQL+YSR7u04mcQXVRHPI8I4T9PCKVXf16mYlRFvvWEmRWLicerPt/c6c33EF96xy
6bbLTmezKAOsV3d/6OQfkUxqLr/K4GIN0sDEhrChUJfdMGuOR27SWy5I2MfMXz1g
RaLgnutLhJ6Xax0YYbyLzPtQwjynJuVc2nKK58Zr3UOue2Qy+bIKHsmfMD/Pgyo4
5W2gPABmf7MVKoUGMR1iOYbn8SQoip4sVL8eRUcUMLp1O06KTHw3hgi2175FMipv
Puf0maHMA2pjXqAh4UmH7N+JS54pszG79ppDTNgLxrLbB7qPNjE9MJ6xNe8J9oM/
bN3uHq+sGZsEY+3pnvo6BqRfByRVW894oDb3QlUXH/hDcX/VrvKcvk/rfp7HA6O/
P9BOHHubktaRruTFgHN6NeZsYRnbysLCm8sOlK3jULpZyrl9hVKYQUdVbAF6Te3S
mLgvo+eJYlji/k93yhjEx8oRU/Ys7LhM9nf/KUJo0afqu3pn3qhnAtH9lKLzZP6s
ESqvDKBTQKRn9zrZTWMj1ArX6H9M1NTv34dFU3VJQ94ngl/PwDlxRWgBiJRCo534
JiS50rJ7DD3YJLy/5p3QUYplZYCsN1g5O5tvuGSqaa/SBGlpmwE3aghTgul6orWM
JYS4wLGOivsYonDW0O2bMLUCp6Vqfpve8k2cT6sOqQ9HvYxBY96egkQTgUrKkeKt
Sp/MQ5EP4pVKgLwY+8yutkSuURYKTDvOYor8UOhs1uEklclAI4QbWqOzSb+tHt0Z
FmzXIBl8ZcSfr9y2um9T8ZmXraCmjRGbSVfuiAN/+jCQw8isHWAan6SucliXHSZg
o/nFXTypecu7Vdqe/9OF0UuXoHh/KVFkVEU2H8jT8vc5txrmXmFF+ZGqMxjYl9Yz
lXtKGq1sKFPKiRR34+f/mLHEXricLrJdxJ+o9/tUJjBEvWGDynT3sFDab361jRZY
S/lR5uC6qzVkyRyLfMrLf7/4I+fSMRZlASSnDARi7oU0yW9kD4OVFvVP93OswHVH
OusNix4FTGgQ++R2EkrOFEg8DU96xt5XzkA4wc92A9jcXW85K2b840yxxtOzEVGk
yIWT+wvN6S6EzInQW+XsBXoWqwRkU1qO/nto7zpf7ybHHF9VMi9fLRC/Xp89PsE7
FIGWMAgbS+2nOEs7PfOXbMwehCrjVNtV/JeCavN+B0oiRBQd9EBcEC9dapX2PmSy
6XFXIELMuFvIcvG0+urlqx6wWUdtykcklQBdfh8GCs6dD1awH2STi2ETqXJxflAZ
BwFbz+R4wLh1FwusYEKxk6u1GTSzo6qulXQ7hnD0+/Zk4x/7uBZ/lz0JA+KLt/H5
6eBXoZ2oxj4LrRbYrN2FkUAF5moqP3Rjr9DwOiXmoUNCzpex5rSD5oJ/MRimrEFk
OUIt/2jH/8TsZI/oh0v0l57A3FIX7XyfH/bRgxBZyLUAhOoyWzFM3iZPCOYcjLO1
u+chNPaMAG1N0yDbLbS9cdLufL3JZDj3/xpqANif26JLGse0vrJAhRJD7JyTIxSi
ZT+XRSByAkBI97KjUz03OhupBnmeY5cqjCnB1rrdenPSYCQrWWpURUYOJugLDrZ7
r0UizGO4fpOBgv+CIk5XhfAYMFliSs2rgRq/YN1wBmpCYARzB5jfbi+Byyq76F0q
/wkQEm5er7YeGSKHBNzYn2BjWNjVbMtbQxp64mGIXBBpkBJObhLJLxgv4HRCPrSm
PytSlcyLHUINwarbuUKtJ6IXrY0fm5KEoTJ+tjbg5Nix7QTlJ3zzOZVSsxO2xTtl
s0CeR9GJHNZgmhy2eKtmlluFM9gqNCGR3bLL14d1aripBm/DvfGHAKgGA+k+9yO9
BzZY+TmXfU5yGTpdlzQvrdyyOwvnOPUXL4FinFSXYUqA/mJd0D9Cur8yHDfy2HfU
hxVjf6JgHglXq7wnylN8l8ZuPzteQXKovWdvHLiE0SJRKh6MWgk2AkEm2qcZCMwT
YV5Ic5ypRnmAoaiazdp7F12s5kGqkfpy9zLTbjM5MsnPQYdiivO8ulLapsaBpCWD
AyjSaHnrx6GLhCEiHPm6isKSVA7Hi6qyPOb4bylu/nf6FrOYlyZLSSPbfZQxTkTC
zvyMd0CAyTOQ0s9cr1ylxBDJFajYG9B0eKH+4uZiLeQEjyGa0n4LeUV9CBLhuydR
vDAS0MIGv6Bq9okYAf6WaQ6AILhAufd71ypC7B+Eacz5w4Zw9G9dPyM9SLimngEF
40tDudKQQUvRStKd9BW5alzNw1Nx0YSYZ0NsO1pQXi0Dy7fFZbwuBcHVzLFpykGR
sOOeNcu9vwKSbA+bjJZrNzRWFXZtbOF1LS0czFOiKkr9mi0BhyCHWIfOvr1YiRU9
gYIoWKLN1E+wbDCpd6cVKkR/eJzH2G+f0m1P3ULUFXLhQzwG4np8jUdr3qGVj9Bl
CGmNzgcZ5O8R1lof9yo6gey9QLDEwg75pU8ygzzpQsjAvf6qjT0ZQZqHcex6ZA/r
1yc4cc93hgSaL60Dl33Vm42VqXKXQm7ayPEDnGG2V8w=
`protect END_PROTECTED
