`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AxwHFXUnBAP+dbFQ4ofZ4E5D4qFtpTs8UgxbDOMGYLUmrO4BflqvY6vgTfnVEpT4
orWufFZaiYAk9CpBkYQrXUGNLqrdEujkDzbUl8Zo/UVUNvnHE/oFXWEjmZGnB88/
VVS7eZ9XLjIPbJ9mOQWizUzure0siMQmWXfQOW/LBoD47s7AZSr7nuW4UZl9RKsH
ojNctZzpD+W+QctjoVIlTFg/NPcMANEr4qa30tj2G2ZZxTHge7fN4wyBGU77xsJq
TEuIvrQ5rDj6QiZXi6HeAYUppVmB/mKzVr+Wfp67eKV4qPXGEUudzJeWywksh9V8
gSsseT18FDIUjqZBklWIEa/ZASfZ39W+sPMEA3smpLpg3MDQTv62QZFoiI2DsGQl
jq9uWyZguZiMQRQeaSWIxEDlrWJbdViIzWKM4YfveWvEY2d+k8dOYb/EvYvhb0eh
gZXbsZlvkT98L2i+qsdwSbM7x/PePJ96NdBCH23ICY+XfG/xnjR+xoBfDW+hB3gm
uloc4qJPyx8KnUluwJwCIcJbb6aXTHphd5VSPaVjkkjXkqKLGOPiVdrvLqJBnsWP
HCsJ+5EuCkiJpuvmsTh1uW04U4IXqKwCWx5A6F6HfE1j7VxgQWqc/M+wdvJSJj1B
A5FsImmROncBQNJXvhjvkmc1TBHfpN2GnyqtwyeUEhyxX4WmLUjK9FW7kBwbSEZW
AREcEBdc1vykBbM+dMabv94Ovn8D3eV7dNats3kUszJkNgQ+/ulfzd53SGb0I8fq
bT9+It+siH6euQtssrSB+Wv4yZix8p+Rn4Cy/cYWlcWyDDTUew22kJDBrf39Peg6
gzKvLYffcZz+M0dztbpEPeDm0afRYYKTWJQHvny8QqJxa/fZcqBJ7tQuCPkpoTwr
aGF/t7EmLCfJsb+Rr8g6T+Z6OBaxkAnov7d1GSXG5qpgjuXE+Nd6pHWwSCirplaP
RC4JoJNiLHQlvGaB+hyRGHw4LiHoYeSxs/x5L2jSW0CZtmR6IERdxxc8DU6BXinV
By0GVHwq1efKWDOHSuYqcet+od3PXs1cvlNvMGE+btRafnBSy1D3xY5wsl1SlFba
s+N9vuyDjpoI23H+14pgfeYX3LPbADAiSqgI9NLA+V5c3jErCYhSTzUuGd9C13IC
5EENxHaOTgPUFeYlzmGTaAfYOCAF5aTi9yjjJYnSblYcPdfTSKvUAcb7jjeC9t1L
OIHVUT2gnuVpOKoOKan3y9Db7TR2suKCvn3OalAhi7j1wEqyQTV++9+9kjLTKYHI
25SuHru2BrHjT4gP1s7Vz8Hc+AIBIuS2h4zGM1M++AgRQAd1voXZ98cLTNOANKlb
4v0WzDd+jvggvG1763kb9jEsvElTG+DNq3833JRHHKLWN4qZ+pkoqKdAcLJSIfmI
z5fsM4mrWrj8F0hJeClnOv7GF7dHB9lka0TXYsZ02ymoyg+MS5OKN6nDGBOurgji
G9PyjZpOdNUUHgY8AiQk50NR50xENmDtbd4B8Iu9OJrHqibBKgyJnMeHhv+bCs23
Hd/Nw5LOewEVmw9TTVv+UDgFVW6RtDAUfKsHmvSkujPslIRSMJyUyhrq3Q8amvSR
/x4DMQqkLmVdqKKfEfgON8wmexeYcgZkZ3G8oIPajA0PcgccagWBe+rk7KKfYiTP
XZQzTlPV4NsPljMRPL93rszc9oSUfLcW7BY2Aj5OBAXE0twfHxdHwxF5BwkjNJoX
XoqP6k/ioYUcHm5umxg478gOg0NBePExh8UNdHqVfxB4gaFFmIY5obt0jq6xBQ9K
ozz/iNVXaV4ANWL3Sa3+4NLEdg2vPKjDf1dE0LpUn42d8fKO1lXTXHWLRzQTDnJP
Yfm594mh7VZStnDKaNLhWcXulOSEOSsYFthPNLmMRaK33aMREut/xhmUADjPpqGR
KW7CIMceErI5Av5enn5ZOdjABV2pL0Px+TEHviX+XxDUXpS9xeQBvHgmJYudHvjM
vJQQeibAXWtHptq1t0vMgAufY4BCsCsueGfHCIsFMrtXcTe34NpVoUNMpz4RT4ix
KHVenUDyucpKxHIrOws3jfMqP5rRJMUhbyDRigNtLZrSvvk5aX4olVxSG/g7n127
J/LMkKxyn0GguLVyFy/gIdgDFj046cIB3/XPDyXnV65IGrKmxtiAYfEhO/Tt+H1V
bB+mQOQ2YeOfKH570xCioYPriAzwwxkwx0G60VQb9gmXaETZns2Rr0z6QclbHoKB
H6G/ClHz47uC027UfRSye0XZNJz2Uf5Fl3XHgg3i8KQmDIM9ht0u2qYOn+k7inDu
aXpilc+AKhx6hMulVIbcgaBdeX8hyGzWIqcPMgOl6WQ7FBGqHwKSsGA+08FSp/ht
FqWoASD2oAYbn4HHAwlhmpYIJDrUmdu8oeJp0En15LKevzMovtkjIFrLuCeu/6XC
fEUHW8w74EdqyAcT0TInBlBZr8duPxtxJtBcSBbRHcK9q7H05570M7FTYOc6EukL
qAYhMfH6dFrDrDTAB9dZCtDmgNw1zirHKZE+p0Evy2Xt2I1DH6ZI2cMiyxxM/CJL
pHOnczV0DaC+Hbjc5OropkZfCUuasWfNDfX/wN4kvZSCsX1kx3mVw+IxjmEK1fqA
RD1iEcEa9xOmTBhX8No412oMUbt5/ywH1/MTB2TTs0ll8g8vgr3aT141EFheb1iV
FBdsG/p3hcbYYkqlXo5CpNFtmYI9DaL4rVv4BxDDfpnr75D/JiF3FdhjVbHt1tIY
N+rL5Nk3I2dIFExR37CbCqDJ0RJAsIdmk62S+bQpi3hHECxb6ywKSZ7Q1GRV6j9t
K2PzCJMJvQFXIFFHWueKDgffTMUD+x/+gQHGQ35Mr55sONkCce2bSPmaXhSHqt+M
n/oC/ln4cHcruJp+FbM9KVnbO8k2YsERm/89SHXVnLKrNedDEtrrbrEuapSmTs0S
qVyOVOulVy+3IFZfBxuWTd5SSckngpQfH2KB+mzALPMMgNxgfz56Tdxtz+hOQYY/
iMaLjvlElu/Zw2EUMWeY7byXz0yu6Uqj2A0DdbgIND37Cbu9f1ZWtOzDvp8gwtbv
VcAqRykekPe4jHymKUv23Zw/EpMyFeCIlKoG8hKQtNdHSlAboQ9Pf3L934OTNH1k
bLOxFKtylorZ84gMDSsNVYA05N++DddzfoOXr5ysI1vIg3NCEIqlq1XVnig9bo4R
KjzAvxaoSuxGl5EVxSbWiKm4Z6l39U6Vxqo2ELrvklihx+hihwXlm2I0xa6+H+LG
wv7UKUYpI5yiyTD7GDzVdSFPLVztMlt2+AcZZuWwsdlCaQHfoAvIUv9pZgATHWB1
IKB4LQPZEha5A/szSBVpu4cZAv/2/H5DyUFzXiUWqBtxXz02y/c3Acq9qirIpMco
ePRvO49n1yYe2hVN/cz72ce7mEYrWsAZ618Ok4OtW3knfAzj2iaQ5p4+BOKvXM4J
rJmSyr0JfmoTXsJnAs3y3DwTQPm7JYZC+KFwmEYafq3cl/i+Yy2HEtB/VgqkwwKh
MTeUjzLftDQjUmvyM9m52qzHrwWLRcCVpLJ7uvtoPukH0WAf4C30MfmRs29Jewtj
LobLzxY0sa4mL/MPYM1z3qItVXc9wux4A5PqOSIKjEkl00HNGnCzmGhIyF11yP5/
xIpHOYCI/4kGO53m4Vxf//OO7Op0opvbaTM/K0R3u2WapPaqyMdY+iX1UNKZUOq/
m+2Q3NTXG7O4FeJNwBviJ7V/Ef8MR0YB1S58eKpc8s/Sl6eUBexJjGcVqE1W7Dzl
DjY9E6hwlKr84uDJxOb61qIfJ5IkpMCi92Qb1/cP0XLAG3h/RrSO5UufZ/Khzb8E
KFSsDaNEjHWvFJO7Tml1zPjw482X8UlhAL0qyKZFs2j/k5ZJZASb1Hr5WgGm7OQR
WP+lkTtu8infAoEEwigskIdwwhItrMmxQEzNDg7+kgUks4l+B7ZXLb1cnvlHaFnP
Ck7BBr+dVP78wCiI+y4HtjRrsCXAaSbKORwCuBWzvdXmk9WCwle+t5JYhp6WjfN9
sdTUHOPZBGAqG3GZm2EeFv8cKV/9zFHZ76r4/DZ2iWAXerVQ4BgsgfGEO52wQkiW
H2evoh8xhGdw4LHYlfknGHRZ5xjvZiiKyISDn6Rr7DmueMDYkRnT5q5WYUeKgjmj
xmJ1dtv0Q0PVW4Bg7vMjObqbOjfdojyTZb7zev+ebv3crqdlvBOKHe4sdqWtGJos
4e8hYT4zbAQP7Y/sfdyQZwwWXfmr39pNOvUndkXEh99+AUX5bd8krEIBUr7Z9jlp
oqwgP4U3FkDWXFefu0X5MB97S3TN/WcjFwkl5E70hcdcTrAJIPr77ONJpL37K9nf
2mHobTu8WcRfAneXNDcZqJrDhLB3EAF84VjUnHLytADLHB02h+ryrNIOeZVx04K1
0Ghn+EPXGnT7WHcjGXPSUxcb+okdmgUihROl4kMoKViW7eBgE5mBebD85UWI1A69
NpgQw6VmMbtsmgPek50px8M3eUk/m5EmVx4SfT2DeP2MHz5Yr2oIjwgNkqqrQKQ/
+CUB30MlcaYHMGQ33c/eH5xD1acMVcQ9P4/AjyVAvixrJbZjKFbg88tNcsrxADiL
ohb55gYPXwAqXYepxnRdlDy+mBG8Tkakpblr+ia3aR0qeZbHbEetPzMXh+E2n206
jscwXHowfGoHDBi108kyJXX63T0aodjsOXX3+kLa0226elQ95m/Mlfz/+mEe1ijy
FI07bjeFbHcA8rw6PmXG/MJXQQHaqlNR5TqCK4eTHC/wsZunqcJWRoaqp+gf5oC8
NUeejgz9go7QGAXH7XnrWiGyw9IqWFewmQ499PNAO/JdBlsiivQln1NUkyjxf6pp
9OUFbd7LWyZS+6jt5PcYYXzYI1EMW6XcS4TQVGZbN4FODDMrS7w669tMlWvLqIFF
AI5GaEPmfgwakdblvDpEL08eAZr/K+WZ8r7Z3DeOQOv7imCWCpyLoXal9HcrfckZ
PwwK8OfLu0Ky6FfYHR9ZyLcGlpvv4nSn69jjR2uAfO3f8kr0ZTJVM6f8DMF7Sdxl
5+FsxOxgW51Q7TklUtSddGFouTdEZFNpoLJAv2aE4KxLI8GauJwZROyWB26mbR57
+msQFL+jCFGMdg6g8HRS/wpyZMTgNux4h0Zt8U7QeXLMQeKtJGAnK6ceoS4Lllme
y3y335L5KZ0YnfNCoPmn64XuxACUGhRrYCiVr9ewZcD1CTqybbo7lLCfiv+TBtb/
CxpAE1Ykc54ChotkIMFvkrXalYTxyt0gRLa3DTmd+01vjxbf/WtoBbBHRG12OvP3
h2hYqefrgjdaYIoWQu3/SbD/Xtqpk6vZpn8yg2hFg068PXSNO+62RgKl732QBjeZ
Cr6Q6fKbsoqSZi7pyP9U9mjazauKI2iGpdfdrn5tnUE3vR2fAz6WITNfMk5vi6UU
zuI26mqx4MONSJtJ0WOcS54MTk6pIDiXkfPDJJheJTPirPfd5hX+1tlMisGff8Xb
Jv8syfs4+NitneEF7m1NjkaalgC1fmtkTkuarNQBBaMRD0W5qna3L4XMSlzuW0os
DNuWuPNoNexflVz8xF2vTF9/RZuxTOqwwfQwXOmdr26tPuf+cyywwuMp3IXtyBWA
ooHQToGdF39T1z5JrunTwnsflmrjB+Wt9v9r6st8KoU=
`protect END_PROTECTED
