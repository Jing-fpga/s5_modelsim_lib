`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/sAMTr9WdemdNHfEtuMk4AikLyxmuj0NFl/XV5KaQuc0txHFkZwzrO/Quf1X0V3Z
5quH8OYDWbZUIEKcaQ2sRIQYvyMa5/+Hnhmqm4yUcOUIcG7jCkhXPw6mB8OEyIV5
xWn4MVJBmPfuSV8D1Iojy+Xj0jjj+T+6lM3nrNUuEWNusFswGeQUP+bIk4vjHdvd
JrzByIyKkGZ6JL3rpluIw65ZW81ip2tLmvhBBD3hQCzHAbqtmzEGIzv1D+S/IN19
ZY/CMeuAJvDQO4cqQGjeYYiyow+dOpIEgveZ78PzRsKxJMuaCoUC7LfH2+JcLPjv
oJNo1G+ZFtkNEJeYyHK3Sq1AnyfwePXFpCw5QACF06uz8MY2NbWbmSfWxoZz4UWS
83nINB6IKZCJTJ4DRytESOwQIkTaYiAztni4Ds1xz6RZ0t8nP9QjblwN/SFgXAeh
U0jGbaPipNRbQSljc2QOiJEIfkq78EKe8icO/+hPvQwpzydSvamF9G7j7glTb2vR
L65bgJ0qsvQufSKft+F/lJvddaBxfDR+V8dg5zKhpBeS5DQkEY+Ft25anVnBhR0/
xxYsxgL1RPBlxtX3dUd21OhmejupZsEOUJw2alMslxFlGBzcghv8G3sBi0NxjAyE
TYfrx9wx3vcQ7TGk8J43CTIIg6trenBDRoS9pX9ckfHMCmxl7xyIbmD+7wIjW2So
3Rb/a2CpIFIhA/ta44cHdU2hyWGHLDL8yuwYcrBEABbmeywreNLvnuFvKzdseo0S
MUj+cUSL7FriwmRXTya5tkANoREAnUma6Pa4XylNHU4a6mZiJH0/Qe2RyyR0uCoF
kQHWD1JuV2nQMv4x4ddWVaJTnTUF9cOoQZhn4AAiexMZLCM08diJ4CoPySjg0Nqg
SQ5uU1V7lXfeNNwu+izayRu8psibkm1JdMfxjLv+PDoRGPbf+z0MrS4O37gqzTlH
7+0DSJqV+6zd5gTcRmPPzI7nHaWb8wrDMzxgaOjWaB89ku+b6X+5QFFf/0SUd0+p
VbRZj1wk2fpC6fdWl8j/u8qD3UhCgamCZMuPC67OsBF5x/Q5bWRtYjYJC7mrwecR
jDKCk+IqifEXPAyn6wZ0KLWfQfJ+xEuJOMx51caxBCBDrDKxQTQxbpMNUn8wEVHH
nPA2sGnrXJ753yTjrlvg2gmCfQeqMn2DGOjzyIf/y3kg+cF7AGlqmn4xxIgf+0Ob
c0CzuClISC3yBH7mQucT2GNey6ELmXbOdFfCFaMNRS65RK2TUhyu6lkK7O478blj
6PjPqo7jqFsfNdvMord6eL0fNETyhz1Ie9mL2qoII7/lN1ZE5ZS8I6283yrt+Sqk
s4hcM9xxF+MsR2SDJ4mZHz8uRWpBP8A3c6QHkTiYd5lJJWaKRg82vpRutYBg/X+l
y2ZqjXVB4AKzRLgy6RdxxtgOb4EKUCk+o+WgS+15hhBc/GnfJ0LBQcfWUL5cbX5X
DcaJxiXAmDdTKSROi93fwoOZOW4TLos2rfZPfXD/FBbLdayuNFSCfEahryK80tq0
EOq7PflJF6wyuL+vYfQwVJ/A0lJdmTZ7Bh2VojyrH4BhXFoDBsNGHIoCzWa4zThF
YTacLk1EsIi3ePc5BCpBL+oVVtNhtnKJDRKpWfbYgOXwAkBZRl2aOsU2QkpPw5y6
D+pUSk4HjclOpHYy2G63oHxO7LHS5KwL7kD8HuGev5i32M8L75Tnd7nCh02qMiT2
G6PmW3qF6V8Ek5vvqUFnt0bNsGS3z5WQZ/i7q1FBUGA0nKjTl6Piaj9PPK5oThWS
zDmEuc8uz01RcIYB6UfXxlaiXWHXBCUVOzAM3WuM3NsUMg4gr+zrUii0MdivDQxZ
XLXchfXRepFX0sUaJpYKUEl37gX4tYFe9ykM0bdtqS2o82DeBJnN1EOQ0r5hMflJ
BVpfZ94jC0Dtwm30UmztUAIUaOPYvhbX/Pl5vtB2OifzrwgwlFC+R8p2zuq+Ne6Q
IkNrhWHQBkFjY3MloyrrfZUPU0FckT9J2dJc2TT9AUyC1EZ+N5BDHpKPrN5pgWY+
q2897c7HCxF2J2kMrXaQHt8CGIctg/UIV2bou2WWka/dXOhGv+3GOP8Mi2QLS2ov
tx68MxBpg73HzDAj3QXn3hArD9B9dx9+/jbQ3+5uPyTS+AbIE5d7H54Lpr3MKwqM
nqgccydys8Yi+raKhLfvZ3OnjSuxkZtPQV9Y9zmKJ+IEoo9oBo5dSTpJ+0FVamSK
KH0g7T4bGztvPo9yKkFXcrapcHbO6/ZVY44O7+Ndx7iI4ELMzMF41YrdD3AGhVps
r7z5Z6X/ibyu+LHWn4e8qQlueCfx7pww37fCf9W8f64IlaSGX6wyW+rMP9rmowuH
pz4igpnCJsQUvGVZTVRkR3UGg4KBv2XQ26wnyXGXSZ+qZ/fmqCigyro8pWdWGblf
zDHToDo846oXkVIpXG8LMn0+HF1kTUXTCK5MWg59vp/ONf3mLJhxSFP2znGuAXaY
AChA66drjcCnE77cu3dCaLCfiXqEjJ4ZK+1f/bkidnxhcP3smMWW9RWdtoyS39hR
iHOUO7ORPXZ3aqyj16GQ8VHXqo5KnJhdK3aEKnA49l4khp91PljzU3J7DN8k7+rU
oNRApaxZeDaYE7N3vy8nt9EgNRyDEfbvD4z4Zw4QLltTwEiloQvggc7VuJB/0tgR
pZy4kpUfWA7Bkcj/WwfKsPQez8oi0cNIhf/TuCwbYAh8mMb79fgikWHrotDhWgrA
FE5xFeamofQt+cD5YHUtfH49sizi+DXU/3AHaRPcxYd7crFtn+EtYNj9SMwLafNW
EoWEx40i6ESjisx5Oo/19+ueyfntG0aiU+RoRQLCUSrM3dJTpXFv/Bst3ye6cyG8
mmw8Z1b/FWe7EoJXQOiI6ISthzwqu6mRjG5LjAqVDlZIpMiB4ujWujgvdl84ZAfX
99ur/+d3P3wKqAk1CK/CpnzOW9cOOzG7aRUxwmmOcJ5nsroBTZiflP5yrjCx3GLp
IMlDWtVQZmsz6ARIifmgVM+0a4xUgJdqLzisWLIls67y3IvAfaBceKEFddMOj0Jo
fdfyB6hI0Q4tByaQHjSOqpGSw0TTr8UwNzuSwaf41pSKJBU9CPxw4rx1irxUYV3c
vrkkeu+ZkljCo25jUy9iO2kCp9Yfq7G9pXrvpbkUcCVa7OGYo/dmkMRhrigawWhU
LqGpOKx3wQIGgl18P4RkRRBukVyd5FvqPdCEDsi6bspPR3u+QBXQ1gp/dw+Qh9d0
5OcOlrC2sj/VmAYvvHvvbUUMfXtpvKu7afPgzoHV0tFtbj49dxBRa37txOBmJWYW
E3MH8VdrsrcmRP48hOGPhPxrhkrr168IGRsselqQ9jty1CSJwJj5cZj1GyRLTUT2
eG6528cflEYyR9TI7+2gU+u50I2x0MlLf4CUglmL//HfB3EzXTwPhRevfhFpjXip
IaIgXACagWlyXcvK5ZnkLZNORiQNrN9sPmePLfazT+s0S94/zDF4DHeIVBxk7OBa
wPFnrpRTbPJBVNGpCEi2vtrWJgLxzBwp+mitL8QIgiYc+5VqBtshb2pLpAu+4cTM
o2geWyjg19BlVLKM9VEVKghfWEYfIkblVMsg8/RQU3ghQdKn4sdKWXRJDtc73dYo
XAgjj9r4e6nV5Dmd158YIm6D+g3t8HJEK9w2PNIaU2LfAKRBjRj+4SKqabPiBnx4
tUAmQ+loMayPoXIoxmZ5xJj6xXuFl8xlezjB45d97CW4qcI75Qj2z+x0U8QZwjtW
676S+KvWnuPB5XqcD+ZLfFgXHQ1vtdVmPqnc89LiNdvkmf6yRwuOq4OVzubBn1Y6
IFJmihc5Ysod8mP0lj2wBUp1TahjZUBTxAT7fJH8zW7u2NgCuWn4bpYDLhRZeONm
cA4XvrhexZnf7ivI9uTP23PH5A8i7bsk1/xRnnU8RM40e6aAuPYIjorQI47l1i5Z
NHKp4muGZWJ49C9QpOv3ScvlZ6WaFZ4/yq9lra6PWNg=
`protect END_PROTECTED
