`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f9K9vaLoNgoShydUEDIOK5ZReCPzG8o2+TT4Gf0GtRFP8cuc4ISM7UUa3jy1VkzQ
e4HrpiuE56CaDhfST4dRV88cRfInqwsDgEscs6dT4NabZjleHuiDhxkwNyYWpoMA
erQ2XNqYFAd47b64NMr3fklCPjJKkhOUzO14z1OmHY08U6RvleS4ngkMZ2UlQNoA
PLPMuc/edSTpVqjdhGJBvvBnOVDl4dcsqxTOdZYSWe6tVG3QHj483CkFTnIwaTA9
pbdBjSPIq5bJGGdVeB1lmeDhcm39LhZfbM1KSeZRg1pbzoVTDzHbwh6uZqs2ToKf
V1vchNVF4vaDmXS8Yafzxgwie7hsjr8MPutwor+r6u/f7eSaPAQ9q3BxeRKqssRy
HgKoJr0aYTeYtblX/QQUn2NWnOCuPOe6IUQ+kzQ8eyrqkz5FArBl9NOPWCcFlzoX
GrX2P1FDsFD27nosnb5SJMH+jCbWQjYsxOjEhUG3PO/cFYgDavIjAtjphUUma5as
/XUaaAO7A8CMszbacOrMcSrD03MbKKMdJSgLPUBtEKpE9L8cokonPHKdvV/cOhZD
g2iNrbIWA/0AiQjKfZNCOSSNzQimRzjgcat4D4zFeAPBep2pFm89UIb7hdDpejwa
tife5MHn+2FikLqNmRJ81Wm7X2Nk+IpgHE9ef/ZjkSEQzHMITQgQ4PHbjPn3JkEH
+YxG7e08AAT6TC4Cnhe8tWLZtbW7QqAYHCe1AFicVcZuDqDMxf1AiKJSrudup985
KNAPknXoTxgiRZI+kFWNlfGyyX4qtv6PCfZLOWKY3SLRjRaRs5E1JWhBPV3Ux9rv
+oRWud5s6vjU6I6y0bIb4u/eNEGwjbRKm/py8FCYsrYkuIk6oWTcjJCZJSp86MNm
6uTE9kWgX6gxsC80X8g2b1echsf8TeH4vqNp4jzdy59M0wgOpmOQJEb+VmfuGkQI
q3/t7NzJMFPDxvA4lzkeTzjq1qCbPi11H1eTr8OK/Czs3aHzB37cxvUDMcdD+oLM
SwQbtpXYlUpvN7cN8XARA6ql+urFtSk3li2HTlka0Kews0uTKrtGziGIH38YBDyj
XvVt3a/JVBJP5AKCNrpOSGtcWzd6RAR8SPrhS2Ad5SIt00p+OgXmEzc+/RfLGsj6
MsDqh3Tfgv0L/Y4tG/+XDP7MscGNxqFIK6jPXmX8nogyl0NuZ4nf8EscpNY/HqSK
Chrb+IcsxKsbKSwbEfOo/RPBVkwq9L3lIo4P29TzaVp6p3tJjuYYfhX0fOmla3Ps
vK0sMP/AyMkdf0VyYD7rZlOSuP/4nxntm2ssboyTFl2XrLfZpgv7T1Yv9tzIfZnV
463P3r26u04wZM7KCa3ekn1Ylr1+hwt2Q658Y78gcqf0fIR2w+0Bcsmh65yuq1vb
KUsF247nGkjgbr+wurHOBGJ7XJI/T3rWVuFSr4FxlkoI8gc7mVwvz9W+kBEmOv45
l2jFblgJuut6jTDPVeheAAIeBBZZE7m0kQXU00lMs/JTwBPpSPw8Di8W6h0W+N8/
fOE1xEcMxM/yJ5YWyAjtfKbyYN/1+sTYlQw2jmQOQ3JFfENBDkUIIzpnziVrZcWb
U/ATSqFK9g8wm5P7X9W+1jTv3dmogXbQtskqSeY+db9kXWxZxS9UG0bjNm0dS+7d
iEa5YKWUvw6lJYoNy4X668YUDovFCb0QerfgXSxjf1W2JRmzKU/GAaDY1Q0FJn7g
/wvNFz9pBg9Dn0UBTAepnBjVqwRMwec5gWg3l2fuGBTiPT/f7Vc7fob5GqGN63Ft
o4GB+4NhFf9l9sUeBd01j6PNv3Bg0dk456IY7+RGEDqVr0X62JukY9sfYYsVbj3r
yq9PvggpFMvtDZZALA2pmZhlamUmmhTmmS7dJ9sOe816UbuXUCjXXr6XGAl4Phch
5mEwvY+OwW0O4c0QsXiuY5sXB0Yu2uDBkSh27M/aLzsDzDUrVtQA3CinK2gDePPC
6WtMbZNuINVbhuexi7IiJNBdR0P2OPw0evAvbJB/goPfEsN3sBBIELOTLFXmhsLh
a8KgpKm6jFHX3ggw22yhU4/VT0svbLXlwY+3cMI1cRXf69ZPjPcxS1/34QvjKSdW
CnswAnCDFKhgMafIItAvPUSIPrcs5OpmQACeqlCU2cJigvQyh9por4h2+n8OzeE9
JYBovvi67VaVyGqFhic0Ch4y7IP+FVXwWzVRzqedsw5HC6gokOZXdJLRNYO2hPyh
c+VMI9C+gIvbJ1d1VzReBfsV5V/O0gzV8pZFEaHbJjYOYoXqpNqpG/4gm0Gh7qz7
1a90ja+8mJvxY9MlswIy+CSU0WjB6uQrU04BmF8jIvJam79sWB64MsnJb16qvtes
8PhXV2PqbHb+QlL1ktZF4zjIDx2IbGUCgEWc3g5SJEitMZ/q2LwHEeg8sLGa/GkZ
k9dj42Skpg8S4UkzXYhFtlvxdIPo97xs563LyiVA2eHW5lAV6cqpGwXInW8zvmFL
k0/2BCh5y/QWiYU3YIiCLGpy45g03u4x2mdRTurtai10Y/5YyzoYao46RyjWQ9oP
ijP6yQLcGRMaN/0xFHGphwJ/ABG+AphbNfp+kY0HE3Rl6p6SjUDDGSnVjcCv6IcQ
F1Juvwnz/rmhs+iXrJEMg0kG+A3GDfGheCnqizjxsUWkdlohk60jlTosUaXDRbIH
2A78Km6f1QabpF5xDaIhKBMEvHH3wN8I8KZYqGtcZ9KRcTh4AqHwa9kA6JQJQXiN
eAw/pHma/FGijgmgsIAVrcOizyvAcPJxwWWYixkCvHHNNMOmPwPj1XtRBZZtUXNp
2Blym6N02cnvCjyR+PPSoRWJHhBxm5XBdZgupLgHkLNcoh8UG/A09+0pBwt/Ap++
nKmyP8AbCaM3AoiXdX5IB8pEc0hkiHrEvyviHM1McxVFnCEtuJMz8HjfP3GTYv4o
yt2Ka+ljSbTnO+d5HJwFjS9NOJlqMWzxBf+k5gP6EtM=
`protect END_PROTECTED
