`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K1EYWrMGVZsE/ByDyF3atlHTKpQCvnE1Xp1urPv1VJ83kSvGLbeE/AYsCDLBeOC9
igkWUK03wLQUK82V1F+UXBhPv3NbmMs9m4bqFZtrxw1g9cQM/BfBQn+2hAMhqlCC
RRHKqOJt3EJhZV1qKOiamXAAvW5RyEiXJDaP8R591W/Je6gwF3Xp5PacQThlVMCj
WjQkHjhJuOzU53PQze+Zprn0bzTOJ/w7bhaYbg1JmKKUB4Q75SYHvkoHHAyGeIHu
nOpOWoi+OCEVAWnFkDpz/XedY87kLducuiC1CcZv4I+Wumebddj/2VQDmsev1KPq
tpm6yDn5D3gcEnhkVjtC3Lk+7RRCZRiYCiAglfF3j+ETSu/thdPwRA8FZ9vsOc1l
XlVive9N0/9ZgJWN4P5BcYzCrZaFhTR5RVvLD2LTWYm8wyLeuZVwtw3Oo5hCPLSb
cETJbzLyo1bQbA5hvUZyjVgYWu2S8QE3YgAqNEKDvMjWPyofks7QEsHWpD6KeviS
57MIddqFi2064d8JJQ157FXVPC+SCxmx4TnEuszDJ0GedumSeksBZ89b3a6cQsum
j1SN++I0V7fnZzLha/qoCXr9BnMc8FlP1A8tB4Dr0IWqmvoFvNSr8Xim1TzbDzRb
iGevhA2BeNNo8MWlRDQURa7u1JHIW1a+vfoRJYeW6p1ZCMgtgPTtWu+2UAL1ZOmd
E2vkVLWM9dWOy7cv3pGGpnRQ76ibBLbvkY8qw0eq1oh41yepaPUhTKAam51HAZ3f
sdF5AyMlmvG7ljs0RqdCZ7LGggDREtKtTF0x+lV7IVKHhLpunniadj8eHA84h34i
WI7y07WKX/7gzN9BLaRO1VC1vRPP/pFBwY+3VDiKT0126Xkmsnr1N/2b7BX0wPJL
qIW55jf+9XkYQGikHZpk1uV/nUnEcHfx+bCEGv+nt8zm1BRB3TlGYfiSadF5HuDS
t+c/0eh8iplMr8HFa1M8QdiiaFcDBOYI8KY/Xqj7SZ0XRGEemyDC+K0mbph/cwVe
SLDy3nodSvkdwjmTexLduNhTfVAw9xY3xLH3I/42j8i7TfKUaQU80aS0kbY286OH
71GgKGIedg0DRHCDYOIYPVedtP8rq0enG8Gulko+3G1Ha+OPOBMGU61iHs+5xowA
XFg3mCyhnZljApPNxVUW8DpM5PtRlgJkDu714ICy/46kz+ZOSgNrPjflU5slTC1X
kHRohY4XzXUgebHF4ohkRwtPAXb4AkoMiCV8ElIoHnLCTryKttrNphDc4AXqTf83
ozCG1iqgr5UK0MRRv4g+LjQgVnTMFU1WMztJHu23pseLqVKyoCD9ETqM1wJ2m9Yw
qclmPyoUJO1SjW1Nz6knrvVNWaOb27dr0+YgjGGucOl99/JtgGKXJl/ZeOZ1GE0b
EFGPfLKPq98fqjHmVpmH7tpVsaCGigrwOs8irs7KXobn7KlrEhkeRNvkJKDkAzZY
f68fJtq6+6LQX5/YtrgnIt5VKpUUttqjzdmWmtSkFDhsa+ydtj/zsZBKSZZxU1bX
bGZJS4gzbn2L+ppReq1bm0QWSyT71bSoCknw5dHBav8aePNVkZD6MjmYqpkSZaS3
yJwBvNrY5Rva4W9D9TwCBoeYXiRg26dfw2deYnQFnDswUnu1nfilnIElq87DaOjm
mgLmIR26cKGv1KuIUbWons47qh0O44yiB1GuOTFXvlYVyC50b9+gL5+Y/yKM/SOg
BNz2JoPLSq8I/z1K+89lNLiResbwUTlT2r2/q5x+mGCfTfvVqr6Wd7PUNFI8/uji
fiKGL5dD1FotV9ls7X248FcI6rVEYVi0ztJba/GXrZWHV1I2fRoLpJ3SkZ/DwN3a
QrlEsKmg/7aL5KXIDnqMvMHO6kaT56+KupD05qH4DEhyR1k7VVZ5qijhZNIDul5H
rFUFFLgBSS+kcjynokZPMHP+eDlidC2hoHCbcnHQuUOoWgAd/IvK5rppySihFoxQ
3n0+pBJM24aK4tDHIOgQau6x0tmKRKUzLmmrt76fItYgk8kBd1aoFxFSAgSxw6sV
uDCr27Zhc2R0arC03CCIsED5rVH4BrCsGl/X3EKmHuV/WXs+ztIJQ9CToFC5cAcn
OktqHOx3Tm7Fs8jrPz9UJ6s7gEJw6z9a2bFRTC6fAJX87JSfI46hLnO4JoUBnfh9
jnzOZgMTsaNWT192Mxhc0ng5nTGNJ+Vu3f/MuMneMMOMJE00WVrN8HOhDv6pVugM
Vu4xUeCkWSGTqDcOja7EQ1+n6VquCdGIoNMxbsHqspBgV+WuYXDNyGpK5ksT+zON
Uhq0u17jnGK25/8bThCUNMYPBnyWYSvNkJX8pF8375Bycnf29F/znUaEwqF5/NzW
TDgRK5Uj4c50WoZ6FshLgD48NWG+62AF8pDIXw9PQJy8g7g47D9PKF9nZuhTNDUU
0PdJLXfb+l55NBCtY4Y4e9b8mdhalknkgokF3ei8poiyGFNfM6scSWKsrfUC0iib
XsBTGBCmqXSeDZCfELhJXDFLkc3a1+BJXIprtNX37rQeAjZR67nNxJw45v3TZB5D
SB/js9RvaX6tKw4JQfph6ldF+F3tKqZdmdpfSAdXiWssBNQj1fcSFUYTStzwozFe
eTDsnQCQmAIBYjymAHrrz7J5sAmKuyPA2nhzZBd00ukAroL92fPs/1exdUEGL04P
UFY6ZDh6G1bpZySshGJ13j27VUyp+nTpY88Q0OnjhIlggSsAYXSUBxt0PrQeOrDq
vwO63A5iP0dyR0CHjrCTJMOvn3zk7cvDi3ZHyxIIfWzKt/Bb3mwvNwRnF7ld2m9w
Vx3AJ5A+4CXipDEsUpeTDfU13NnKsUmxC+0zp+4kMIliMi1963WdXhUf2uCMETJ4
oLUZh0Z1732GoryNU+J3OfQe+m+Bivp9MgAekBtOoc1BYo/dzAcpklu7PGpe9u2W
2+HzQTEAcV8KdSczlMeae6AD5Zm6hW1Pm1ckrFOYzFUtR0ohD3Z0FBjqRR15Ejc3
t3a8ch1IpcKs9zUjjMVypzVxsCPU28y+SMst9PMPos6vG1ddhmC+YWB5349rJFba
dOJTtK/FXzTbJowGWhwtOIYG/zSom7fuYN2mzBbElB171eVfPxLeRI7LgVKY//2J
gyGQX42ktc2lVtM2AdSAlcx9UMWwmipM+x7EofOhpVagNFiENYdB65/Oalbn/0st
YFS3upT2gqPPVe0asOqixtgjept/qsTkb/OxEgbKMuNoLykMpZrvpFvlAJ4zvvZX
OaPb/9gL5bfQdCL2nSVxEzPkhX63gc0ymrTv/FLcnktFLWRqeEWWZxHgREXw+nPu
H923sEz1KlwoV9eh5pgK0noiHuZuBfqHRFsXqctrKMh83aCt2asg0auiOd27Yt7S
gcm0Q/F1/TVnhxsuDs9fCYhzKxSPiSEBs7VCnAQpCjYe1gdX/9tMD/gcfjUxF18i
Wl1kPyaaVMztrJQs4IF8g4UeGHAB/CmNfHZY0qQpqBNCyPMsk6a/VA4xWSeFGaen
txTNgFrT5cC52OYBXdoqH0GVgCFQLJf/nuA0g9+umyK/YiS2uuVcoNeEhOQlIept
dhjGs4+2GY52fTIUdsqyJsBZHkW4XP00ioi83+yk5MVfKyp1Zba7q9y49N3Z8A5b
i4Ym/j1x93sPRjDFO5ffUaemgawMUIsCaBRUQ9G7SsP31dlYXuezuD/9MId1DG1r
7gRFfFCmnCTLUeRdhU33Nm2hCY/+Ld64GHriDNde3J0yFStScYQ7YZAG+J5wpIcB
odOIMH8/sSuAAuZYSD3q1xa/lWYN0ite6qmRDfOl/f6T68cFgbuSP6AqfPJkr98n
L4KlI/Y6+57D7xDac/j2xNH53J22ebo3TNdrATyZaCQubYnoWpP1ZEkm1aGYlOHM
DQdWxpr6H7CQLvuBTtp0GuFcyrJN3kr/TUc1M8oLvcLPvTjN5o1v+n9o8wHy2QD6
W7utz3CivNiseLgnmWF0nQ2ItAbWi8QECA9O/v6tsPoteOzKNGCBNkr7HBH3ErGc
VRgYVNyUQpS2b9WSfhZVBIjkXErAKsmwBmBrb8d0qMvtWZIRkAXFMQ/CuW5FpTPd
hZVUHkB4+blvKsPHkeldui3ry/uAHozWDaeg8UZazsAiubJMgMjsBkEOyOfOtmM8
oTsTWtfSiA15eQDFDLmc0/gtSB/YD4OH9V1yeoEz6l418ZjAhVM9k9NDXP5ZRtWa
GF/Uwx+zpSop/t6z7+3/dq35e+ew/MdfbknLXUkcVzuiM5xhfy85DlmjT0pxR2VV
pPyOJnIXG8DFCIobvukiMOJLdis3EmkdA1pIKhHWwfzx6OD4kelLsRKMDc0cLxCP
3a3vFlN6xj3fK9Nho4NW0clJNdNpcH2ULF1bPDRlNXuSr7NWS9440U3uwoZr1ycB
p/1+2cl0sLy39MhlsG6WzIwhGVa8iSin9STuGQZ/6+Vgb9qAx7oTolWYkOOxP6KS
/CHeHcgwYojWyAW6wFHunmgY9vBn0eKIBxKSX8BETAC4nu+7yLFh5fmc+B/kvlBg
bYny3B0Blcy7adkTUtw3ZT2DgJ9PjJp3hbB2gfecBUVgQsQP/nDYv9/+XGIOMEf4
ptFTmYoWIA3We0F/n4eY9PMpc2Tw5ypcqFiLK1OdrVnLRpXUoFO04rN24Aek3BFR
je/RqbAEnBQS6cWEuQHkvUqwOgECuzSBRuJjp9rEHiH5UvCpFDxT3PG/Ya7VflOc
9BTYBaoMbfrbEKUs1g5NIi58m0kVyaOYZu+Q89Zy7lXJIla8x9qjayYMjDepDn6n
3XXnQNmFr6eiTAnESsSWWOeltwS7SdY7ngqDQNaO6T99+wfagzbC7+jzh+x0k3eJ
3TqDnDbkujSuc/fYrp7pRVzkDB9Dhj1JTDw3qsKnfgBxxi4lOpsbGTgsgCFbDkzh
Va9lzRz/IPPRGTPDqh6L1Hf2v6vHiYAbj/RmOJrpyiEs1m7219VdphWNHe9/cGo9
P7hrCn9pkTRqP23VtOzJOEw6y1PZh91wBhQL41XKtuOc7SJJBsukXDZucgISD26d
i3kZPL1tAWfaOwiQtdBUbphiThTnNTc3O4hyGANqzZ3US+3Yvx3kKVJ67RSnHKwF
Yby1arUKH477GxOMdcMz3ooL7D3i3qeREYriZ7X9Sj8VzoCW9jtfBOQ8sNqSGdcN
9NEHEj0CIHZMHvOSoJ6cxJzeo7hACDpeBIGccmD+4iO2jVcVWKmDaHRhYgA4P4z9
5q6hLvygrVNr/o9mhpixv4XcGH3swJY+mhTvEtl1VKO+Y/kgWvasLilKtt2AR+ds
dVNez0p4bZK1MLKIzQGHz5ogfkPit5rsvtIGokqqBPh4foLl1BQZ4yU9EXm7AkQz
lzlnfP8LJ18J+3z1CXIfHizQ+Ib8hDZ3Ghe/N3Z6A1c/9zfe9+CQ4fvu2OdImv9X
FDn/uUBL+HnS7DgshUmcTIBBXcM8xUCFsgAiZiCNXhg2FfVojNRtdi39aR/JXl9P
mj4hs9mjQHx2QZQfztD6HVtLUfb2FLxvvpqZHcw/wSiWxar1zZ8QnkZqCGHTnnW7
1NSHkiNE3ZNHtc7AmNIAEppMdT7Ub9RcfdPp9C04h+xcDeDBMdPnizk9yML/MmpO
uvGJlkApFY+M5RNy0vb70aKQ/XZ0jR1An/ZSAghMxq3MY3NimliCs3XjAIhyQGYp
NnopgAsf87e7raG1NQa0dPWSIH6AQ8y+AnybBqQ2ycSu1ht2OVBAAmLX2ZIwnde1
EcKxvGwIXqqBOVQTQ6ovGwxFr7PKSzoRA/roEtYcC5ee6zbpbSdzlD+/pyRNcsTA
BVaWMIxpHElt8e6x9oFlW2+2/1SFgE/4awPOPRqbetqCLeRNmtd+x8ebahvNNwfA
97U/5qNmCakDXzEnrhfwrd06CCkzf13YscFHLgx3id1YpSe48y47HZgGGKYBVBTC
o/rGXV5hfwu5AibvT5Y/m0CwJ3wUGBdgqlq0IRjLOi0ZHADYXXZAkL7moEq/1naF
IkIa8gypsi+x8WzIy9HJj71wdH8Ltrzr1stMs+D4Ck5jWv26IXRhmfHFD/9dkQwF
SwN4WTxp2ZlYJ1fjlQUyZJ+GYInH5W4cTnCLGOLHSWrVbMo6gFgJzUdrgq3xoL9Y
zfRCkhcvzTBkYtpKLQZiq/s9sNLLvC0gCwQrTu3RNfPUjiqFmHJmgUdgHvKCWB6s
Re82go/CT7bLp9wVw9OHH5zRjNFyqGhP8FgjEfbWleajLufHk5zw3Gdr0Ph5h0Ph
Obhq12Sv6GCqMTG3B+nGsv7HdQl6llPtIj5mq4B+rj1wVhIKYpcqMmjK6wuaL4zO
i1v2n5SggaXbPg/cX7Bn0Q12T/+Tz+Y/gSF/qg+koZ/oJ8/s76gl2Yx2Hqwke7/A
4QJ6ljbF1XRTSiMUhAWV6ts0f2JFeSQWhDtvtFicVDB6EFpKaT/FX9cf9iujwUbS
BWhOCKevDyDOysCsOH1iBzeNYr392TD8ehCzVS7YfvG7LECw50F62fWRQWbcjoUC
j+64qnJi2d3qm0AO+cftG45uQjcHywM9tyXDQh5ioKVZYwc+12hEUgVPu3D7Kaal
Lfr8TYFqvK6AZ3VhHgJaV8dWvtkbVhHs//EnubFET+UyPzXFOIk+wll5Ubv2lQgR
nnHW7nxz+fUNluHXBYrHgSVEUp9fgaIVp2YF94PTr26fww8LgcEKDJdnPft6H4nP
G+0exCbkhgmHehqduEsDBBOMc9OmcOSVZ1Wt6I8PzyVND6uMKL65KeKWsPN7g/K1
pze7VduZiT5yzaJcJNg8ouds9oRXFK8deCSEP4wS8PMWu2v90PKT18XoUw7Bb7/d
lN5AjJUzKXnF1T97rRAKHIKrIjtVTPo9MvEBP3Ha0/k6WRXxkVrVJzzkRU+AozpV
JzwaG3o1ms7FSDDdPPa3XKS2Uu43OYF11gqhCbHjSO7O09QeO43ny/h+EzbW3joe
lPZKcUbLHwz67Xa18T9rfavJ5Qaww/gwLkOdpwTkOJYxPglLmmaQF/EKbwgEj+lj
+LDKU5qkuA9BYK6Dmml41xLd+KC8Q1ghulsGHZ2mFeEbmZgW1LyzcgEOQqj6xkVd
aphaGQ9rlmqCzeFwwO6KgetBiRnD13r6alSgeN3EviYNm6PzBTVzLXi1Fijk3cKX
ZLnTGOgh6oPc+1VbIBFFJTCRVAPIuynYgxK8Dvugs1NGRazvNXIIxlrhiQ6o+zW3
PBzK0jzNfeiSNIY8TGXGVMmTi/7hob674PPLFcTFpFiAuZni+cLM1ZYtRem51HWx
HFcCHyvzo8hTQpIbMbmrhRAW8+pfCnAUCypFO2PtMtzcng4uB7cik4bkmPQed+yQ
hY09lQ2RilDNEe0AzWVEeQ+MVPnU60U7NoXZQJmamVEdedgkObhFs0OSoenCoD2B
zxtuSTLYZ3OHkwpjLPNKA5x9zpBV4YtwzPlQKziuTjRFbvEq2bYzpiZLFh7qSpCo
TOd6Ahv/7jMO50esJRz3CGNIUQbY13Wg2iaBJxlC+RBVcQch9ytkXwQs/oHD8/oE
tXrhEtEZEeFvo1XCVSO2qZLs1dEyycNiMp1YaMCFWjYsHuvRZK7POinirnDALctK
4/Pgfv5cud0nYigo3Fj6oZOU8+kMUmJ97Y+mnhrgxum/foP0OmFHWh0l/zfVH7Gy
dPAuufBu+0CRFtWcrHPvRuLDWMRpOOSsuQFA5CY5QVh6R76LlTUcYttS94Qf99DY
3VhYLg+EnXUPzyBcAyoRyo66pRGw7oHkPP4Z0NnorO7YcwsqEuyAM1+p1rEIaR9W
22W2QfDOz3GxM7IJc98gl4IOZ7F69sUadF7SXm6h2HShU8IUkz13GlXWltDt47yR
nq0/veLmFlR2rdFjLIqRieD0U65AFD9Rj5SUy2XjVzUjJQrVf2a95aeblzAa9Dwi
+g7+18nWl9MMOU/0iAszcWX17SkjrLX/SLz9Xarz3uSqw6Lx1RhF5qZib4qsUEws
fJQ0xR2ki6lkKCgFWHOZTBHWa9kl0oWXJYZ66z7WTmxRaDKZgt+antml2+94F9Pq
jlSIBvhIoPz/uvw1J3QXwdPj9NwS1EMoBBf+M25MmuF/2uLZ+O0Sqm8Nzu/gVL2N
NNyuczYtZt3xtZlEHG87d8Q24eJynpD2/Q8ZHJ9D8RHb9QA6cqmWGPLOaNZaXB6y
hU+HModV8mhRhKoMThYqAufS4LSqDDB5xURlkgUaVQO9yzgFPK5lj8vTMrlGsuXJ
7YRV7FBQqeSJ+Aj21Dg8tGeRxdx0tHAF2ZpVsk9tP3zsNw4eSsER/t+SnCoToegq
4XFcsn/yJkZMAIEDnnRkB66+AWiJfIOK1lAYkd6BwV45cMHyZ5Z3MRhNA+24qEDW
oE/Rw4lG1k8iiW/tw6HbwJ/IXBLCCGXSPo3MautF0qqzR5QzBB/WxZfF4BEICyPj
O6dfuJdxPU+jESbvNQckU7PNTVSS0XtVh+eS9aenW3O2wsjFkfODi09RdEacR5ED
krrz357Bdpc3jIb0RY4Y5R7zf0doPM/IMfUBhGqt6In7NrDybk6SafqG8/skYH8x
z9bfC/PYmN/zxsC51wOVOnpPiasu3tuha3APahV8jl+IfJf3z78Vm7H0d9NLStUB
hnlJfR5jtIyvpq4IRlIXHnSbNxRUAjQlIbemt8eegMNq73yIsTS0782+eYTBJ371
f0qk+g3mjdf6uhsZqOKFm2OH0kzVzSvFi0221sn7Ee9iuL0WYMoqOVNNNHnKUndy
DYxw4oNpba6GqYHbrW/be34BvbCy08Zc7f+y8VP9XSEpy8fg1VxZp9AqA6LasYrW
Xan7/0ByCbyte5V3y1rXXTZWUHwXpi8TWUVVu4RqXvW8decDP24OatsSFdZCXcHq
P1KYmNK9pvBcZrAmhc4C7gMxcPUH6X9gj74cOh33rX53Vi9dehOJ2Bwwi92olb8M
RH2/KRgvP0hsMKpJ9ZilJoRkymaUkf02X3RA7tsFO9kDIYwuc7sKSMvzlcdELHnR
SsVy+5RPAZTLSuDMLeF6kQnbqePD/Z3NG9fM8IA1UHfOj6vV/6r7p024bxioFqFE
3RQLi6mjw/1r8XorYtE4/ZtXsofM8Dy5IAEKLObV/y2ToTqVaUiPnTjoSo0Qeur+
tncCNNMZMlP/fgbFbO3AeF7Ew9s2p8H0jELEqWfuk8EFNvRec4RsAQVq3cCQKG9A
5KlbkhqrM4qT+KdE/kurdicSf89CELLjkMZS6fYnxNmhT7gpWvUs+7qWFb+q+Q1Z
ynnZkv0ZYJgVtQ6N28e2nT9zLWOJ0WQ0wAnG1WSnTwIjrl5urffRPOEKvIuAuiHI
zQwbla8KymISxIRhQGjdYV3TnlGE0nLkbkPRPpHWJZOsBbrWnso9YLk1FXqX/apZ
NXF20N3MOYBWw4spEIvYMNm3OCNEN3KidEIpZqdo4A+S5ZP3D8800Q3dukfNMSdN
ix+LeHlViIPChnGK9gJAL8UgjxLh1QJrOAdHrcV52M5mJjE9fqPfLpYR+yIAdras
Iy6gWfv/BQPz69OCkUOwIuS4SaVL6u8iapVol146lHqK7POIcnCWE3+PXszfFBIA
b/UreS8s7Dv+3fsOOxIsWy5nZRJIoPN9Pea+tGrIzKGvsah1u8GCjE+oabXGFkXP
VrfCiKtoJX+SDVj0aYb4W5wnwmvVGQndyaKOMs9bvdzSK0XqRvkN63XOGOCVaAXC
UlabmdTMEbhAMd9MXbXPRc1wckxTr9mEIr89sNCYQ50GsUF1heEo/6Zx4yQn+BCj
ZHHOYwUIN2/LrT7ZMhNnWtH7QF7pExqEt7ESNW0KL/lh89gM1uLb+k3mBo5hAiNz
mOF3KJwloXdB85+YR8fykMaUvqk5LMcabRJEsTDKKvlpDW7WqmGs2oeC/HZk5yj4
oycMpbjbhOVMWiR4taS9iBPo7i7H/ylVSfFmXuLpVh2ZxXTYhjBURwMPYagOyXvZ
C8MJLy2OniRjOt91xDFNDyP869CHPQhwkwzwmufooJP8eWSK0CHN71CFy/yly1+v
Dsd3tUPmLrL5ibrPZjS8PKg8dWO4oSwzYmFaJWBlnr1RC1hN8iGkh7X71ATc7HIr
ipXF1RuhbBZiXPYPDtv4nC6X+MW/rOOeZUBnQKGaylII1fszwP5nmJqz8JVl4bQ5
5r2jUv/3DA3Jm97WosX3imvfP+hIZmlLcbUi1mhMIerzZVOcI+6kkoauAYKjFNrm
fjk6b1RoHJTl7xIgU+M3jTV7qUzQ65GV3q2VLS3AcKBmj095p84aqQGABhYTrjPs
9ASI7ABSWJwvCOT4nQAz+5JPXnjSabl13whu8RWhcpUKhJ1sf3qML3nf8gL2F1DP
ErjKvByY/ns1uSyxZRBsbeRsUeyPtli9uE3onxSdtDbOTvR0Rm8HazFRiz79f2I2
tX8ysXszOY8KBElk8zWAyP5V3S4wiJa2yMK09t1Dnirl4r5hojQCvOhOjI9peeO/
AWPDUjR3yB5xKuf10dkI7xDIBWdLm4ADl3k9dpNBGBgQDFErWJVnFUjba9x7pQxr
T2AVijdf8UqjFVQiNcilBYL2jvUPtLrvVxyyZQV4U3Kp2Bx9Z62g907Djzs7Bb7b
lNFzYkmxUZuJGZG6Cv7HO/0/p0A8JwURKWTBW0AUKNS5wkZqVDCNAUt/WWV8I5Wo
fIouTeJuDr2AYwlNs3O/XFQcVRCzLZLhVtYqP2HB5buiAFm6oYlnrsugm17APj26
xxFOmMakXyxYoTkZWEStx2ttv8qktGmvMIcPhN3iCT6euXHF3YwHlLQ92S0gCvvW
4TpZnxYzzJ61bnj4pfh0+Kf2YWCSZjp7JThIP4QmA6UQxFEfX1p/fd+qtR7NlocZ
4cRCENduWRA7Ml6LN8xC61CAdIfPV/ZIiQfCiUNhJXwxRvnpVUWIdMeOh4ihoqP8
QOZk/7xXOqRMj0yG90G9jczhNiZejx3+djCxAzFXCgV0Xz6Jes7UvQ2/P20h21OO
IIYZgxYFY4uhYv7XYCW6T99zHaNijd00VVW5dfDTCLmNGNac6lUDj2n2KdArIbl9
JSDxe6DwBiOEPgb+SRD1YYvC0ghiv33GEM0yDUMn+bS3kcaZ5wbTjOBZUCNgm0sc
qAkaQ0wV8zYmF+cYfhuhq0baYHCN8gLppHe1VmF9gkzlTV+8KSLy8COHQ9RzNRmL
18s18+B93Y78F0XLgdoyPGTc688zvYJRaT3sTw+yGrRe6Sx1RCs9+Rc7xC24VX/h
QT7PT76IXFgAXFjH1AwbbD9Y2sOpSj0AUYAq82cFRt8g+M6NKGnpYoBEkrbsDDSo
98DexzytI59MN8TIQGCTw51BP4wRNhztoXsnYRhfVTVnGNtaFwyE4XysLSZ7UKW4
j2WqZj6MYuUtS4xTisUafB3+h90PDVlDg0kxwXvt1JZ/xACF5OWTrk7BPNrNwHAt
jU0dXbsgd3RqSyUCcUiyjAoUHt8A0/iFG8+G/em3PxjO/K3r9+IFEd2nRTSm4rj3
wjAw/1Wclo+dLb9qbXCyz/ygQN0EV0yiuztl0OkuTFkMstqVtxOGK1yUHyOQv211
fcdAaJzN8RkfymkeHN5L22zoPQbUPUGvD2hYdzQrBhGHcochrXqLH9mqrStV19cM
VFn5+WWFrZV3XEIZTdBlrgv5YBOW6C7GCp+I73tvD/z52PYQxyMPrQ0snBqWTvLY
jbYf3gmH2lPeffmPDJTNdWlGSyqfVhrB8nrOe1M8oTWrze+RygNzwdYnnzEsSJX5
QlK8RxquL6n7YV4iM9BZXfBcGa8gThCVVEhIfdQTpgtQvS2hIFX5VjCd2Nsj7UMt
aJ41oa4YMwRdHeetcIrdgpu7337rl8Je8UMLOm2ysyRfxSegaELyvaoZofpgx+YM
JadK3mqQX32L60YTRq0vNWr7BQfOMaK6G58x/KRlNmEpOPdeXK74mlioeaQ8cdAH
xyYdgX8hautpbq9BkW+m0JJbL5hFy9n+7FQ3xOPhUs0TxA3sG4sSfBcfaTlFI3iM
Ioop/uXU6gQpo5wzG3IhK60qlMRAZOdGoYcFH8duy8e9ssLPOmWvkquW2lHIK4CX
8rrVnARnJs2F3OgcdsbEPIMd9NCrWixOionatPMVs1zYthyqXqvPQ5RrUq5Fo+Gz
CsFGit7ouT3ywVcUj66PesKwctyi1hYzct6RYOnb1JpK8XiOROhyTdWA0S0/Vk34
Bxc8W8KkwGXuMkXzt0I0Uoi3I1IJMrmmmt1BCLq6VrTC5LvLFN4ISKzpc3qpO4nx
qBFxHrHe4Ho4/ZDxEX7nDaH4/6Gjmoa4rf3sWFhvzBXANLPE4lQ8gC9J1E+YVV/O
6JaoQd4iNojoT4yRsaGGMhFl6U7OqYTVKBYb58QiWLt+d0HR6cugq1ATN9RFcQJP
igWYKgk8/OdSRmWLlA1hObKEcjMf8RG9EQHYCr0EBvrNVC3EQXduCOM5OXQna6P8
qcP4jwoXt4sfbApmsvXDVhRHnNHBrOEt3yAGU/kQ3ItWE9JNe1A+D46OrRLZRf/o
FaALu6NDcrrdnv8S1BbmPeKOY36qNOP4Qzh6B/4dS+AmKC/wDdRHt9vekmpX4Qlu
tepa5rdWW5FHRMD6RL2Ph5eQ8K6SafU+ojNBfaU53/tkMFdNRqo3Q4ZqD0ggJuBy
5CLWq7r10rxviVuY0rhrQx9IS5B7/W9YCZFLtxL2WVYrPl/S1VbTKOVYyEN4Li3z
Dz8zgKkvUx8zG8XTd29ILJ6v0Z6aCmP5kXZLaVUWXs9amytQLHczxCjVqv6Png5r
+HSWJka6HL/1dt5r6v1xzcNVTv14H9Q5T4V7jtqStQpmt1B0LAQf06tlZ54Sx+JU
Ey3/cHCbjXAYoJijXWxmSBTRlhsyzqZmxrlgiAKggxrDQF3dDN0ZnolQ7MAcWD9D
NxzRpLXLL8IwNrE7qeiqTh9N7LrvxGtW5X//nVAbAfGmNF7vY9cvFg9jMLlDpYRh
9q70VTy9SQKcC3g61q8qwIjHp+mdvbLKbF6atnaS/brNmdtB/46Lx3Jga9FaJQkw
qVJs7HS93CTpGEPnesF7h9T7JMnAbeIzKTgr5aO8NzgkI2N9xc39ApyLiv3FXC8s
wbVdY+Clw8HzcKP3Q2OnmtE7NG43xVYJyU8R+A0nu1RRnw55PSfbPQrKHvkWqJOt
jGjl3jAA3XjOYP8cNMp6W38opqmT8I9SVtFefVFsnVSI8BQI1kI4yktGlKcm935F
TZkLB284tGyRPXhLKbIJJWwJBiMx7zDt6rRFnYHwYAbAJs9191giNuTc1QA3ZII8
y9Svr8TBeOyh3vurbWp7B6Q2//jTf450jvCTX7uk20hMZ8ezrn6DQtSzWMyEOxde
Kw+InKlby4Io+VdbgzqxdoFPrhHcvEK1/SXLZuY0HK9jIG8Joxuc9jGLP5UPPzw/
Fy2YxtdmYe8IdpE3CjQOEyPvL+7iIHXSrKkP+Ak0HNDuOqHKFDVdv6TyD9awzFa8
gHvxV52Q+0y6mfTg/8NhZjhq3Z4o4u6R78nWz1syiQKaUjK0AoauPZMbCgU/tHMD
uu9PXPxjn513dMKgZlgLGxrgJ1QRbPXUo/vg9OeHMZX2y+IIzwVbhXuKCfju/m45
BZn2W4oopwmAX65QW+FrATYyrVm1wemNWhRbAlWQ6UsAE2jOygJHXGYBLne3AlIY
p6m8r5j3psixnNz9zJOHTo23S7cFS7Ce7NW6CtDG5ShPiCWoIkslJYbTn2JzMNiX
zGOotkeKYmJ6k+vn1yKVEeT3f9FJglx4LhZwM2rhG3GrWwmqR8VS09WG5+SSMs5I
BGy0NeeM5zwPSwIDG9UWusqJavXM2eTQnGmmyVxpAAHnpVYktwxEO78sumQ+bYin
gKccg4KNd8/lf5FLLvquzt6jXr6kuwSYn77Ksg+AJTtJ061Mi2OPuwOTHN3C1MhG
/kexAgLFh4B2wp9ELHjvy1vO3djjWkavxlRExj6O0UTudj5UujpgR8fZIhTZw8HS
oflKiRdLI6nsHrWvIwBEh1wuyYvmH+UCFJEMK2gc6nGwNb83zFUHgnyeSRnZW6QO
J4F0jNvR+Ycl2PqgV+f6RhGtzecGoVn2hbK46KuWEfpXExVZ35ru2jLlKPqXynNH
ElQmmnI7SeJjMUHOU86ewoNFuxOGVkco9ojzn9Zs9ACbuMi3nUluyWYGP13B0T1Q
Ac3QHdEpaLo2FUmPPnmj2UEPEKytVIvOTDhFYH3aMA/WynKc9F9xb9eNRW0iIV2r
Xr2p6vaEqCGnS1BKFDKxMtvdmifWv3xr8IBNRdEUeOIw5QxuUj5WyQABwTNJ4pCg
IHKiEuQlNH+pUwjKpOdcGZAMmzTzD22iv4eebrHwxpBKNsA5hYwBl1UxOtWzbNa6
juWpcx1n/X93DU6OOQLszquAmkEhXCznbEwUrX/o0j3yHhn13S+gY0PPLJdCcRzZ
REwGr1i0vhv83wpLSBuFK9zeywDIVzf8KAOEmKQ9dKzjfRoHyAb7oSCyCqLxD/Ju
IdNmowAHKBchs6ScGnpiSivRkFFkl8UE8lkFg72BdtyAVLH738svGCOSaJs2S/Uv
OoST460e/lgNNdPCcbLuvY/R7pSGrU7AWSQjEJkp03vOAWFTdd3FISoW9y9kJ36t
z34wKO8WpJXoouY3N8/6Vqv99zd9FfEbeNqYV7tcUheDjE05k//TkaCJUAJtB68s
dbkTHVnuGL/UDZX5tSwsYENRUTg5NZixnCpkDHSlrop/H60evmgzdQtKReFzj0cE
YGGBF/n8oDDAyalsbLmUeB2hbCA2VwELG27+hqU71f4FC4Z0S6lI6An9hoJ86vdQ
tZV4n4FZq6iN1GuIBz8fY8GCiNDzIroUA30opNTnfSlgOMXdf2O8+Di2QfDOatcP
CEcJt6ScyJGHpkq0rZk5qG5AQ+Z3mbpAXZPGJlYL5UJhQUiRFW18T0mRezCmUQkA
V2x5kKTDmZscv+Iit+VpdW2416Xe3QAnPJhBko3oRLaSwmqVVtM+lU9FCa/SWc6i
6vX2Kd0PBdC5E6iwrj/ybdBIo8Cxs5lMNmV6i24epRQ3VfGroKw87NWbqSShJpp1
MXZUTe9eL7t+88YjL5UTKLJsEJ5FSuHML1WmN9JWnoOicQEb3eLQZVaVL58jeTUh
rHuCZX5A5ww9ks2wkWEKSK+Ss00iIlyTBJKHnXGWdMdTFR2hPW+kNcMSycLBWiWB
7QUzY2jLJj5jNbRebjtUN44wOuyqNVhFsMOOzt7E4u2b4rOfLux9SgKjbukytTVE
P3Mh5aPDOaEYMCOaguOnqo8L/oZdmazBN4epqyjCXp31lmw8VJMomaItrHD81/Dt
KeRE7Vj2R7dGzIjFdfRYO/r6+VJVFP6AMkyoKBKvOHLZFX1cTmo0wFAKDlPF2mmQ
Jz7F2QES/yqmwxyPFHwaasHV8qukneRi2nT34VpHmuMC8B2TRdWpT9laj/t5IGq7
EKjKH8T0r3j9xlMaqS/EBdxI1ZTBCnn6Y0JnS8a+x/aH51OZGogWUImpU1UeAwId
c5nZ8dlxDy4ad8OEuMzfqoFG+jXE61xxxTLUAAiHMxV1mHCk21S5gaFi+Xgoioh6
pzbPmYhULhX/6OEpOkWXiH+viI5k9h2NKbEh9lA0xg/vchqPceyEBdnDEGr2Clu3
67MPvIExoXUolgUvf0KYAE6G5xnr6frvO62vgRrXp0QOazQuE+E+Gsza96KXzD2x
fuaQp9xhkw4LZ//1pBd1jGR4qKcYO3mgBzHcZSf/SAhgLk+hZjlOtjC6Dbl0gGRa
WSqPuRlk4YMQbJO4l8yBwCxQeZ3cfMPqSh7Jg7zRmwYS4/m2WnTOlJk1rMRqFOSt
VdJLlVSOe0BQm3mddnYP7qVrps8ZXVUTejFMdM4UurNU0sIn03jkryXGYfNDOz2x
6pQfJxUMdN/zQHNqU96CafqG7OVJJIgrTqKT7jpvb4ds75wX8StAj28dU7oG+fKm
T7KVsZc5+RDZ9lCzU8vO0HhYfgFwQ02rTbQOwUtrEF3j1GJAeFmxZ/0RvIsms+VR
qADmJvtmnrKH7rlcPzpdelYE2IBkbpiEQf08xROAtQ+wCBAJAlAuhzBoNjOHfWCh
Iy698JKrTyYr17NSWWJl+nv7pacFyBbJlTlPVls4KRlIOVQhsC7S6iZbFth/kRWw
RHuNTMz0EMa1c4eQ78ngeFs1pf821BQ47OXhnM6Vlte/UynMFExc/FPXF0QIIALx
Aqi8PJysM0ZqnYvLR0nz51EDNxIP05SrmIj/NMOXgfpplku6OPEw6G1dqRroX4+i
KPx5hk1z0MN9dmkrtCLstlBW06XmuaDbKYUnHE1B/sacrHKThWgRARccV8Slp8ZA
+1AiilQbkUQDMrlc/PyIYGH5KklPPTA3OmUqGnfmKQ1XjlbWASwcTtv/JkAUN5X9
hmk7XrM1aCnc6KTDr4FAAEt4G3iXMmIxDdJAjmIGFMCax39+51A9AH6pLcSGBz4u
xzludOHJ7uzcz7eXwovSY3BOzwMbzoQhWK8FJuvjqBlAqQlyFjfOLs6dKCWyw7Vk
rRSdYQP9xeB+AlSy/8cOt/dDCOX2sLYFplPxlHpShGGdGKQD4lRkWsiSQUtl/3w/
lgrH1jaV/XDAJcJ1xwUVMJxRTdfSgipxKC71ai0UUbZitq+ryK2MZLoYypYmrOLe
zrxfzp7t/e9ldgFbYSVeOyEh+EZRE6w2ikgsyvT0qCWk9OOTbOwWOQJjYjmchtRl
HMR1A32yJ+ZQeu4kndZN0RLf7OBORVxXBB7Q4c8wmyP4/PvE37v7YBbV8+c8Q+1E
HuaP2NNs/9iDnnHpGMOfSTs/dljgtn6WnYCrYbtRe6etIqgLjLJie4Pfuq8uH9pm
rSGplIcD9nEmIJov5NxjYfd2JtiHHEtJ5pseShvqDN8jbp8XmHP65KFnz2m2DJhr
3G6b2N9orvC5iwqadOP7yAjuaQ8mpnBHPTUG1BGo55E4zUOJzT05/bWev/JU2mfp
u0uhYsv0sq/hAl8jC/Bj2wudscJ6Vlqhukd3ERGAYKgSb22ZvPWCkqIWughKL71n
lbEXd4hKQUyWQklb8M9tDaJX5uqRIsj91Hz5N7jPpIEEWdcfSHB+H/GYklVYWj26
YIsXAKT3O6cEjf3VeCIfLtjUaW1eyREgmwCIYHJlIo+cYV15z+ssIAMkYVEywd/o
IVQkYbQRGR/5lQaiw/TRZg5w2EOiWYvw1hDXUeE7UD9Nf7s/0wMPZ4SfA9hGnN2R
Z94lCOzOPPIrUp6ZVryjmJ8dkb8V+bAubSUsZYw9KOnwwcbJKxSvtdUX9/n08Ayc
9VY1ZsCD3n5/aIa/al50ZV5FqhbrMyMjuTT0S9gl5dw7RwPiVc+UeUJftoHXbUcp
U2OsD3Q1FyBcX/c2P4UZaFEDk3suC1NkO8QCUdcZxWCBehOx4O4PKUeTkfmsXgxJ
GmSqzPXnJoe+tv/TSIOHmp9p8NKUJD0Xrqb/k2a0s6O+97GpUXjzxE5UAUv+yfhB
B63TmfprAGeZK8a6Z+ijPWtDkjqpGpJKN/I/L5pEc9XNmEJFDGwZ6FbeRQuQ3oan
kWxCZ6euxxfN+eMkO6HheX4Urzx9hlfOO430T4DV37nI0MmPKjLc4Bnupi2embVU
dI/5u8JkUoy6CyvLPIgq4rUrD3u4NFP+BHy4okYVPyd0atY6lrxlX3+zhgmf+tVl
20kUywZLlxp7PKr6tZaYA56+544lSFmk/rMAg9nCDCp5onGzqb9NIItIbtb4WjiD
g7hLiMj71HFGy7X9VybuhODYyHGSdpVqQ6hEN73g8kf3COdKWemiXdq9wYh5wCXF
ATGcTs5ZM4bGfEs/9Q0EIGJDrEalgRkBWY6z2+XqtL32vgZQEL9p6FZybhM3WhqF
TzvpRlu4Iby71+UMcnG4jbavoBeNFT3GLVI4svAlA3xGyhqQUsqQBXXFm5B3M81a
y8ChICaAiSYVl3nt2s9PBAJouWhvx6EybrDa8KLhLGbzisGmml+wKHad/StXbsbq
oMVZkOAljFCipRVIcvo75NsZpyZIAPz40sLzDkbMHNMLmRG8KyGi6BzZ5+stUoWf
bB03dZps/y2Sgj3Or6qhha1jruMpezVJlks/Qqc3TGA6y9LKPVbbTkW7jKzJBezM
5dpxi2UVtS3E/KR46mpUBy5B1p8CabHdEOEqpJZd4Mrs3Ki5dYVDRqkPSXr0Xqj/
DmusbviilmcfRKhRCx25jfSXpZibW4Efz+oBZqH+PfG4SUgghWNI9trBGEC8cDoG
0oEyh9mNgjXA3loGfO6OxfMX0LeSMMa4hvMZEHZo5fiAwY/tsimwHeLsnqHs4yWu
wjoJuFveJLP+du3/YGyyn97qFw1rrePug7e02uSL11TjebYEQuXcPK3MGSf8gegd
npZd0LdZVOeBonzDpwWbMtmqkIXlA/MZGr9WCaFBqprYgh5xoydfarDKBYvTXoW7
KFeoK3tzlOhYl4V8X0zWJoSEu4vLngeR7/Rk9GIOMA/hL8Q7BZyQpEx7cMUkGNWF
OpqNtnt0vhL/gXTkRLOzIXzh5gaovNkmstPn+SqNcdyrBEaZJbnODgaH7jqNsvQg
gDExuptRsYbXbemiKDW3gryubZsM+Sv4yzKS59vV9ErEK+xo4AaNXpRUTabUZt9e
3dwboTB510AmVFFexzbk7SgmBEfs4aloFajMiQDjFY5JOZt7UaJuZ8RzGwgbMETl
uPSWzxYK/ip6PVcso9EX0zJ5zWoHF8WhVLBbqZLOOLOSvY+mBa0KA3popZxRQiPz
Uq1Pdm3M+E3U5kYZj3TaeSJ9SQqQl5VnL8LkZjNkj3w1gFUJ/4pJCcov52bNFr4z
TcfIXtpj9+6sR1DcEk3iYpu1JYsJtJoubQX8Ii2me9VUxJ9uAEDelJkQfnyZb9Q0
08hw7JJaKieIknT3SUGMuIqzCxeQXIghaoU6IY11CLio2bSzQqzUAjf3ovOD5+Ud
1lGqvsEXIGwFktAgLfJg4ZtV1ms0XpbHo+zmnGMnEa8/ewOWV2khiEvUkQenEnxl
nxd0VdK55E8zYrwIGrvy1D+b2Pbukwsv5/2EjE7g+tv8FlEmnh3kG9El1lWzVVGb
HNDinH87wwrKBlqUxaq8rkZtpyqwS+Jawfip7ZYq6+mxlmMB4g888D2tuZNvId5S
XMzL1d2ztj6N1xM/wJFaXwSAJrHq0PFMjJe047B0rnqSp+oHd1dZZhJWUjOeU6pm
ai9nzw0aB3rAqAaQuNr4e27B5EWWqCjSWvZwPLCpsewM1jFpUBN/n4TlVCq2ktmy
awLGl0bRn2jWZ/NKyGxwjfFcOxAB18kj5TcJMpphAZB9aB+jwKqqUx+DANdLrMpK
aSy4UWHUTHxkfGl9BdC0pfeyETcnhTSRPLhwMSLC9Ecbkbvpmw6Cotu4B5YQgbI+
a+mXsHY99+39rHMFAOVuk47SOFW3oNzj1XoirzUiLovuj0DL6mpf+nKjK/Q9sqCC
QYUEftWIgT/ZfTmhU/5EzwdLYeR++n9YnezM0kWxyEibuyuDTBeGlQfUzKje77ai
sGyng7/c+f3aBW3Zedf3y8MdEG7iuF0uaDZr5Y/xCuAnW/+N30dnVxC94m+tf9ID
hyoHwfVZizNupNyrIj3A8FVeGbSaAX0l+ftIkyEzo84T1sj8RiMWQlrSNLU0SL4o
77MSpnXm586PrIdIzucw6fvM7OWJ5T3ZA68+IfZsAkFDj96da1BQ2dBD/Y1JMtOI
iAIe6CpCPKqYAUdyJdGbSCzSPOcHhdNTx2MGkhX1RXXGuj3PdDMMUUcxn0a6Agfy
om9QrPWXkgI/5hNleIcsrTLsLTI/6C4Ag1q83EWNdIKNGbJGMBdNNqCq0s3E+5CP
mD0k5B+1VYP52eEIZzEWXBI2te/5zexacAgbUu8lyp4NTABgKn4fOJ1RQYdyTMwi
TfLLGHM18eONGibe4nXY2mR6fcRQic0goXH7N4CbDlUojOKbEp5nxrhUUivE7/vg
ootVKj8LJXGIXsa5qfYhT/a/GGtlGb76owEUy1e4Izr4hQoHD2+DV7O2oxJKKl+5
v7UZ0x/HoSd8JrqrDbxTvdQ5DT//Lso+LcBunY3HDKA85rIgdNYS6hHlTy2elqEx
4CSGY7tQT2jDgSnK8MP6mzl4PLoRf7D9uIFs9GRqJGpioYs+abHqUCjA9/y6Y8z+
1yQzJCcpdSp4qPcZn6DbZjVlQW1JKnGxBEqeLZj54miDz8gr7AFqKOHK75P9jwNc
kgC7PiYRSfbg/Ao8fTlpIBwXTp+nIU7CwsI5yfrflMBc2XElVD82NA0oBhcb6nsH
pjnFnjsLfUmzklHsrrobAIMnFE5uefYwS/YM/OWnlseiq4NWrL69vsQd/QutRR3S
5edJyUtfT/PW66IpYT9wZ72Vu+2RSUhk3UwFja6pf0MgnEs5XJZzAFQJgZ7V71U3
1SWiYBbvAq1XjdFitxq/scccRt2qhEnbH6W8YfrPyu6BsM9cba/pa/Pp6b/nHSH1
N+00fL0Vb4F8MBCE7VYuQBLPXZgFFKe01G1LkAHRFgiAp0NfyOaMM9R4ktbRRp5P
VPnJhV2BwEUM6c4FDKK1ItBtzxWSb8FYl/3wUkJDE5T88So5Me9PZ/g0hOBji5WM
jf5BZI1IgZ05iHBDQF7gSHfGrlamgTHX4nVwm9Z63BPgPxfXfLZbmxJyTnlpltUO
8zEFfw76BkNdLEAdhSQAYj1qNLtVY/8y3r1dbqWlR8CDh29UqyaAF6HzWFyYo/tC
JQI5FQpsLS4J+l7SLagHxj6yKh59Clxj0GkjCFB1hh5rLUkTSgoyMuXNruLX7Glu
eHG8ea+eoZz3u7MkkXRtp6EuoXIUjnQCaVQuyugP43PUW8WgzU7SoGI/ga7nf2pt
n3JgEFUFqkbUtHy4wR23Mcp5h/K3Mo9YRiyQ6r3HFYzZXw+971PycPTpUjRBLl4/
bVdysxgWzCj+Xyy34zXGTjx57REQyCZUTYvCpeYV1MLvUOLD8/JV2iq8PgI8i5Xb
GISouFl2OciRQqoCMAIvGE9FZPri2S9yXGcDhnpv23aqE0l133asWUA9S1Zw5fCY
gE51ZqUWMjf8cdfhDkmLtHCwkjghEtlGCpOJt/6mf8RD/bzdaPsNATKVP0uLeuiy
g/IUe7dI/q4D35qs5PB899fuATG4LZMq/zeyluYSp6hlvo8+nfVjK4IBOOm+Euuy
9+CJneVkNJmW2GEgbDVIGPVIxNrfLqZ+T3ZOPb+fDCE0JvlJhHVweSv6TyXl3W+g
xEQALepoLwKmwjDsPhRDELaxHIyr/3NRR0/iJhgSnhxSultu3nELt7DGmrphGxj6
JUTSuH8a7Hyq8CBxWI2UsJs0Utv/w6jRo/x9wI22oqGBX3LhFaQ7C8c4gioewENL
PqPJa9huGRPCmHoJs/68d3vn/Ll7oYHQ0puAUKmgivk5KqYEgmykRaZUI3Ob/z9y
ObH6HEBUEXBmsCDA08GX+4H63h3WDdzhZ0n46cHkRpeDuz2BHU/g0Hk8jvtE8BU5
79CjHBLRWny8bBnS0HVlo3GEvhWrmhw8/bIiD8r3PRtC9ICoGucS6dN5ju3DhUpx
3RoVxHPZBzNvfUzt06SLe3kWgYKyiy3EexjomcM0YbnqBw2yqH8u9Op6cwW3A/1l
qWLVl0/3C+PLYkRp1Pl+rf3AdaB8Fc2nmeRb3fBsvNw90ChQDmoK4MnjkagGp10Q
BTSvaegFH0nKrgJjQy1AYagaCWrNai0SHh+CttUshS6SrJRzg5yNbC3ILMtSfcHH
7rPSXToLn3MtkEZEJQFAxeoWcQSQ6EG3AHRSSS/kM5NPs75V14sB21j5weOpN3oi
GZ4z/ju/s+jZPJ6fo8XvLJ/5dzo1PKVYa+gbrPHPAzNSrOqWASkkw50JsnGPPThi
cGHzhQjz6EE1Y5YNzMGFqxNIvUzlAkgzqIN6BsjIOcLvWhBITRzDEjTqQ7f1XuCf
EnFS9eTuEV8veY+Een+139QAKhFnzBXA+yLN6CHrJhez1vVYkFAg0CAj+D4c7aB0
EyTKbMQ7v6Ef9d1z8+zFKwp6ePFHpT23X0L7nNxP9laJVQbR+2Qk4tLGxrBOhfUw
8n0JO3hPWXGaKsdQ0xHw9mmBwgmmKosW5bBRZBWnF9XNcSxCGLSxtJL/AIdM1eeh
8V05JOApDM4UW9O7Pz1mRGhmkBekR6jYCMG6bWCVr9IKqu1nytsZ/2/koNugrF9T
ucbcuVuwDpCjzHRUMDTc31R+IDNX7j6YpdR0sAHJ5b6UJNqKapUyK3QrMFawvWSw
KKJM6mY9c3xz2xVxvxQnfgz3lRGLQAfNQenUWTYKsfnWozWiixNWD3Ifqm0a3nF+
Ji2oGWNtIZLkmDK3/dlAgo09SRnpyP1k+pzUGsGqycJg+HrkkdeBHnfLDaG8zG9+
rlANbmAlgWtlD0IZG/FsXIk/AsIE5dshrP0xCyV/2tG0GgVBEu9dVRC+EnEhitO+
hG/VC+ZTc4BZxU9NucKZ9tys1VKP3imbrZUUVIY7Dykbv0ZJ2QzEbeqs8MyO0pYP
f0HAHMqlRNmn1MQrNiy8dzcEHdhpOSOU7IHK7kLMw6CPvc6GhDa4mHPnUUoD5MDB
1iR8/vXA8+iS/T7HzcTaPnhNH8QrhOH5uBd8sdkoSgLrlEpfMR1N1EcZa6yrr4dR
Q7vSadA8Eek30MUOmGCEebyz0lIEmYzonxKPtrsgx8FveiIfoZbsX/lhv/BPIw4g
KlGFUbsfdH7XEbQUnQZwj3rmncZem2erm94le5yefNM00v/O68SonNQqjsgS8Xxf
9ZbQOq0c73ZtPIETuQuMEtMDI+hgQ/ouQ9mxeo2hx5BnNe94SUiJiUAKVlaznYy1
KMMhV+jkN5PErsGg9cOzIBtFHm+AQGJgA1G9lmFKvjvh6uo6Au/Sjp5S5EDpmR7G
HapowAFlo/jeLfzbVxYAFP8fVD+TCcQpM4gIqLFDxFqeU77X/PxQFVPlj0+NYpNZ
dLq7oH0HKnRaD9+aKymfih3q/C39gu2rOMtHVrDu4OkaSuPCRGj/UfEjExKiE1nt
Je0h+HiEPDn3e6DYcNxTty6UwaBChMlS/T8t6jOeuX+3tx9A66foumXMwvaJocMi
kiCUcd4gwD3KGgBG9cud6O5tpe/TfYDhbUdAINS+dniamLbO6MmS1Ml/v58IcF3t
YTuI/XUq1mHwPjq5B6nSwoCCXpYNo6sC4TVnOojGwavR+ORTUD3tDiV+dTrX/hhV
w7FtyNaIofj1LHkLJdIJAQNXnlVZ7bOe/75HzoLrPRvrYU29MGb3YHVmMDeIRXbM
UKA6mYV+vKmomYkZ4UoMu1C4oF4rbE3vdxvziaNxAXGN+Re/RaUIDKly8MOQiOZf
d/cfSPDRVmXxqZu7uXFQtOllVl/1yWw+WcYSn+MrTr2DaHKxCEyiVrYkTkug0ksL
NHRianEJV99xwIhuMBViqZxHNFnSKUgdLVoFO+TXi/x7U7+CwyAisOjW10P5wZ/q
2wCKyejlQeS0iXNq+B20amJQKIuqlFTjbQplJWJP5xG+5I7pOTR4NmO8yEgnOBr2
BWcIqIDJKtR1HwxYuFSUq/f9pi/jIbtoGJjGX7XEBLCmDXYkRb4cWEsKhBloKskD
1DtzkuJHm6goyi8162Nm5y1Y1j07kTJSk4mvH/xo8ydvwk2n0IOvELvsgYVD6i1l
5UawNWUFeyI2wIuvIG5UzJg3b0izdypdyIlTFtPJkXAICBK35lkxYe42U0p54M5e
Cz3F+wzeLaoJ63dHKGKXGr12ng/fm7sbBTceJc1OgXqnlgE3JLxvv+8p6BjMOn+e
V8zyAz+1lFTJXZUTM+Bz2Kg4B35CIMifMlX9lekBrecH3pRn16l9tCrmqlngHMeW
WR29zo9FVzLb34Bp5KKc1GRB0gJy8lngDWg/FoZDHwePIf+wcP+2iDIbM4JjCJCb
yJNkArpg1QgD/LeZviCSZW9AyqqPHoKJ+e7FauU6EKFPaoYWweU/9RjpowrVCem2
Op3y6s2ruH2OmZpvVgbmMkfdf3Mg0k0imhrnR3rp0nEpADsh2kW1C40WSHcNBr+k
MjxHmdicSVWE3OwSmOkR3x+52THWCCtG4J9D3Egb1K8/U7BPqBZ3JW6okZWUkOjh
Zuzxa7gFZESsGFTRYksuzESq/qCh3+FUQ/0LImjmofZTyOD743ZuWLkM0aJK/eQB
S+kyaT8e3X1iEaBUxSO1XTwt3mta4oQRv/Iqy4T9luNn7GmYx8Vp9rHoxslYiXJj
rEA8z5Tej+h/t5z3vQRTfZqEgopuFyO1PQ6XExMTpJPSDjJbymdwqaQEMgTDv02l
E/knAnflykfGKsgdGj3rdLdfR6gZ4DCfX7LMEHNBIixYW76diNcLgjr0lpYXfTlX
HuJgApBgFA3tzXN0+5HlBk5qJjuuq2r86WytxVwukD5RgBMyp4JSlNsRIbdamJ7X
JGhm9ROSPxm4Uu8CEoYMrKTR385HTBmGQzdEANE8p0W8mQeIAh3znksNSLOUCoEl
4VY48TRF5Rr226eNEl5rgn3NH4e7Fi0qn7yF5ZxKq9eb2XyFBXeuLJpq9bpLqsRv
Sb8w5l+Z50upGbf4WXtntsp+i+JVRv6CjxXMZnymU0hkD2LA0L65xZiGPGUQXEBz
rdQCr6pGl2qNiXlb3l8hYzawF1ntAnNCUj7tkvFejZmyOnHd/DSlpYijfbvtaioB
LrOr1JCQLStjDbVDUyZWVRngzOsHAkPfnNsxqJ+55kweC6wpcFV0ayXYvUXGr3m2
+yvAbGTXZQKeK7OmufjcmVaZ+NirCMNf4eSVSp+khIj0xp7U3F1NxXT3DvH2K70M
vaf8BctA+XmijqX1GVzWTNCWRV5JrY1O+LPS0eUL2Gx5TGPcd9I1pCPS/xpQA93Y
9dI7FODbFxgPbNlLWYnU3LjY//LoorvDMQO+hQ/OMwwP1Dd7yjWMaW+MkayTcna7
p7CBZhDgpR84dMn6Q46O4QUEEDsykM8KMvITotP3rV8s5J7QQiajkW+GHeYSe7RL
Nikreg45CgQnyvj26ldP5xCEP+0wuKVyZ666T6eoux3SXffCaBe0G4YzpvWMhJwQ
rcNqgrsiz0EOOnQKg5vVckwWISUb4a24On3vwoRMJz4gXHTpfhWncaEuhcd58Dy+
z8MDCXTBejP1y1wWEZa3fMW6nvYsV6sPu0shJOCquikvrD32Sx/T+ZZo2lfmGN70
`protect END_PROTECTED
