`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H7gCHXrEAbuvldINYYlSJc45NKcZkaOkwD3p80L4JhtCI6GS9jGbjNFSqxyS011z
M4Ce5sI2HOM7gAupbcsAPNx5u1ueif5mvKGxRb0Mccb51zYzXxvLX/gn9y4cDOIG
rQ2bFX7RdsNBAAJuCoCCGaB8pcLFeUO/ppHTLEOvJC7Yxw2N1jAWhrNDRy9lwfdA
tJMwI0ritosmXFjTeP2crYC3hAQ63+yZI5IPV0BL/bau5AWzyz31Jvq1ULlG1RCm
NXo1lo69p4264XGlWpPpuaCD9SsKEZCQYqRqr6uFInw9c87DoTNGc5HRamKSrUFE
bLBmCjW7h6EqZzlTeXQunr2lpFIaTVwlRmq1l/HKxeCyzl6BA7NbEcMs3BldZAog
QMeFhwrwiHxpY26v6FNkEago/RWKwtmMADRH9f1bLOSa6QqyAp+R7t4m+uurpSAl
5k50eCADkS9JKmUeI/c1FR+X9JMVNrhU26XjTAeYsori0j4B9VA2z5dwPR7owSC5
Z3JKLRFM4ePukaXwxiIAY9hkfwiAXwJMMSrdfhmt9v0V2Gla02EYtshQ6dtIb3vR
cMP+Yt4kN3aGbZh0LecFRQ==
`protect END_PROTECTED
