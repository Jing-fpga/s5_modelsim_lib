`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qFvmt6TQ1SSEnU+FZHZQl4G/skZmbA7JGqQzy94ngjw0fekHWYoq7S3QzBmHqaOx
U5BfqdPbObnKohDrVX2yogt+m094Q1PrFBpc05owUT3q4x0Y5hrflQR8Y47ai7Xv
mD0R/DOv895QqsxBy1iTCJOyKcSCfPFJSzwFYVat/241gKaQ6ICAI6QUcgEsjetw
NmXt3ZS96BNpYb0tgXWy9fRD+F+BoJU+qAjvP3M5wVHYcPoyWH1PMd8tQHdBGROz
HcNRwHdu7eUkWhawzhocVL2gdzz31uvK2eu2qSnQNZr7p9I5FcBvrE8H5+n2rfYV
XyNgqVXijHjumQdYFuSomYMaZlvS5te9H/Q046/8YbV+Il6KNKn42jSfrIy1ypWk
QG570W7NtGPR5NZUGOQbKP8Vyatmz4TJZ81uCDYejxH9XCmdXyakw1rtxhhzoTd1
E/JzUZgEnf45V9cwWctBvVgGd7sqkmb/etcpso4zBrtKhIyeavSOeeURkkTVVXJO
Bsk04+uy+4QPTCgBOFq1zN7/PhGCSNflUNKW9LsDmliQsQheEY3JewIKqTq/C2cN
C7FydR7U/42JFLFi6APqy0LInXoSCCKB4cVoX4kSFbGb+bh8yaf0S6jggcwXHWgE
pu9wKh7o52H+3TqOfAa5q2Sl2AfMOBvMODMU9LZC9t4CUEp7+3/uutRL4NP5GOQX
DpJ73u9lpJQXszgqTwFhbKYYe4AIPMQRklzs0CSjkmWmXN8eYIwXvttRnqGu1MG0
3zUjjGTJpu3Oshj2iIFzBFQgpi3G+WKaFeHdgyZpZMGP1KMzSyZfyseMaRDID1ZY
b8uoOZD+t/MZVp/ADEprld2WWIhJuaxUF6wlc2+CQ94LffZiBO2CpRPsz3NxzTEr
8AZ6uo8j9vrI03aXcq9x30V7cF9edmzigLvDLarsPr7KSFFcEck5mFvaxRPu0bMl
rbBAp8wcARm7pU5SzJPfMQyUPWxe6piR60CD2roYKN6Q54S7/XpAoRErmUJQnibu
mgFiVub4jECbLFpJYWO0v74h8ViNbRq0IzT5cE7jC9kZf89vAyk6n41SEcuyP/gV
eAr3mQht1hsgEtkrId5wulsNmGKtqF0/3N1HGV6BkjkcSA8uSyu4Uudti0H+ybKA
ag5V6/Hk1QSruvC6PWQkj0plR4dhtuVjjNwhM7rFYcGZFfWSKrz9izz3Rru38pkJ
Rqb7gzImv04s8HBWSmfBrg0JWkIoRYQ2gKbriAhpKQ4hy9FuSzcTyJH9cHLkVI3h
oDQ/Kpr+xZ5arsXnvxWgtXUzlN5FN0XIAmI8Gz1m3eAFRFbCTNZN3dwbZup9jr8k
3R4hK3kRfbcCcs/2+epqXqV7nm0qF2hgcyYAwotwobgymA7VgaGIl7TaRb/2bzsy
2phMLfv9jWoy8+zw7uo2qJod+Gs4A+ot9giisbM2RG0jzx0MaWXNQW4z3nVVdC8R
TBT+oNMB9aBCxlruOTAHodd2M9Lj8SFelrZTaLIUlmu9RMSYUdNBOqpjd4OK7VU7
IVxowaQB7rVRnu/XUiqPZWrzl45mlwuEnnXDiGGxM43JOJbUiunOSmo9d3HlaWtN
VHyLK9qqdD55NYlqgMGa/0B9Yw2S1gdCnR80SlN213lR/bGz2WnofqqOf7Fai21t
VeUPSwLJuRPpE/j441Xc6NBkFS/CJiV7GVDBut3WAiWqxnE45arUvrfr3wYFllEH
kNTUscFclJP34j9El7BMWjcEGpMPItVnGvi49if8GLmxTblF3T2qmbIhw9CRE7/k
9uO6+3WrPEqymjrV6P6AOIHAZIelJ9nRgoiPTQC/MRQk9L3Y61F462+ARNRO3GsX
OTjLCnR6Gb11ABl/riBLyAWuVJhaGqQRjGL2Q0WenF6GhE30s32MSe0CryxJ6/k/
CqQKvT977ikoGLkBc4j1ualuSUqT8PHxK9evZEz58h6nWEh+0oAcMJbRoZbFMfgj
AqNFngiE5rqYSn/+23GnFcR35VSR6zaBj1NLv36elPr/ak8IW8CxAZvgape7HYKE
ltn0zFPmXb4ge+KqUzHDZ0gXf1JSOMIAaQeTDkdT1RTA8MuOekCgEeUn7GtB4tUe
jekbHkqn9zhG7Ch9PftF7aQB7FTPe1lQU0MtNrAxDz4kSuTfuIj9zaQxjEesGpCU
knV5u8DxfFTOymxLgmidpglWxRlhbU5j6gEOn1EXILnPCyiJR6E8ANBAb8l/XGfL
D794cIEA+oir9qssq5HNJWQTzi0svbObs3vtCNHwcU70hNtvJcTF+b0QhxKwofyC
7Tt0ZpafatQwhD8x0nZgwgJNOPBERLIW5uPKhJ0a/cVJzLk4B9uuo6ZGlMn56XIw
FS9F1z4FCpE2YIOC4bq7ZN3gdlSOYN/wKfTyh28H2G4DTqvfwcbaR78BVPrGrHH6
/l+bwGNEoJdmixV02ZdEswdmtVRVcgt2M6IK9En9K25aDVpGr7wEXpsw9nHzh5+m
+9AJcB4Xwuy5WYRkyaHCBH8oGYRVoY4fWgJxFXxbTnT0wbz6fLUc+EhI7bUgeViX
XzH6/4JbiXHlafGSwfUiKDwM0I1oE5EiivElSX1oClFia5F3zRDfylnngKv2q1o7
5lAtPLxK74wvGCu/EG7k+2qdu9u1TagHuxnow8HZV1z0gGuYGlsCzpK6C+NqH1C7
QKtPgp5ZCveC0m8CfZsjXJQHpWHDNwyPDuxLu+9aLd8NbqvMtbfFmB1OM+6YcQwU
ZwpqOiKPwYox4rZrLz3yGjmnz3BvdggD55ne/IYGoWdvUkems+5oe9n0jOowRtQO
Rrg9HnyyZpOjSVLmh4upsvW45QVwfIR4eSr/lcpg//78imG8PtOaDQbPpQniAfwX
zlRkS76xMdgP4O9nA4gnNlBfO641GUavGqfgxV7Hz4IRo1B4zUeMcpu4FzHJ9Q+8
jSzNA6Bg130zH6rFefPCrfbQteBI5BpTSls7a3lj+N8=
`protect END_PROTECTED
