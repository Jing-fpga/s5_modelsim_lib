`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HjZpqRPyqAOG6TFVdCJygo1dPDGSIklm/jKhOClDjLIV0zXU/jGAycQIcumgEkjU
NnvoBnBAey0KsnL0epzjxhOV9xRttxGkDJg/3Wo3UsG1fAKn4U8CdJFq1g82QFyF
o30PfJJIVKN2vQLQmujN+ErPzn8es2qT89tf7L0MkRd3BmXi6N72cDukPHF+d/RD
QUc/yeenmsWLgERF4BLOarqiaSAWHbpVXLd/qk0CEWch8JjS5/azdjNi1NlQBBmg
KnLkeB1nY1l42+HQoRB44PJEne1AUcZbT07/WQhoFd4DLdB8ioOGR5n4CJjmzYXQ
7CQl+E4vbI/bh0SbVYi0nabwRjkGMuSYacAfX+JijcR9W57bJdBHYT9BRQZp3B4H
1E+571SHoX2inQ9Zmwv2ijaeC9hnlvccYAAgj4QvRnIz7650Yoof2k1Dep9kDxVB
d5Ru/upuNqEVDwZh6foeqY13cBzjVz0x6H2y6XLyKiWagMZmRXQwofTJwf19BozY
qI4GPzgBI159locgwTM4hWGigC90X0hU7kMRSnkVqehAl5DGt55gZWsTGwXIF+Mx
M8g/DZUq3+E3quT7cOuPI9369k+7sDL3V+dRTWGhyMFpE9tu/OXnVI5cKgBp7K2K
MUj1XyOxC7HGUOLeyLxM+UB3UC8kNxnGg0SkXScjcVqorR+E3mjxqUQPO4vELzUF
ZIS71wIEBHcJe2iYVL4TrO8iY7hzwjFDmnet1soi6vQ7VyH4odKOSdNNicKolTSL
z56CklscScZNnW1kKC3IMzpqJxLNfal4RSmmaINNnMuUQqZJJlT3j50WP8XMFyLB
tajJCLtrzFfnQhd4Ofd+B94mpQFRZiuliYIAwicAdLhJZgMDWsh9RSAntolT2xui
oTAekxqKf0E5QZLk+VeHfd8lRcGJyCcLGl2XnTQXhX0wbcFt9VxZU+2Npa/OtKvN
aUUV9ubM04CjkA/iS7pjs4XOG2JfbX2xpCiMVQ945OsUdQa/Brj25BgdSnuRY+Zt
xxHFFPuMHOtsxyYUSgqFpCRqlYuyQ/l+sx1+8LUv+M/fbtEXlICrS2y+vmIBKcCZ
luhfMz0NnmblUbE2cdk2yBxlUXLrR37jJlt113iZbr9wS1ZfOV287CfnwvuDhrlX
XaIMlTInI1ocqn/nTknBw3O4G0k870EFK1B5lAzcbhXLhsP+DSwnnS13N4euF9Fc
dmHekblyy2Svl/fdXB3C9S5MK90QnrICtE9NHzMGMSpq0dZxgjVjKarH7nJnpVmH
cTScWJAn44zVaQkL3pv169PuC0zCxikx5fhKaYRuC3p+jk39uNG+MuneubMOYy8V
mkiiPXW22BhFEy2mxY2LeL5fieS4YJEBWEk5R1MHWYPdz5SyYYKfoykiyK+FZb6c
DHXxnAnV2hQtzk+3vLOxTgx+nt92tcWQdryC4y60WbL9E4iQhSqKc/B4Clthg3Po
qyWeWnEo4MJRqI7ej84fEPP1EMGJ3z31o8QCIxkyRjWPQkKrA6Mjbx0lFBSx50/Q
rr1j8cvf3YQykyKQijKy+K1iAZepaGAoO/mqPjibcyzh8ay+WzpXl3NNPl5A+3lZ
KGUb7PqKej5/fjb+CH7bZ8m98TdDtBIVMVVL/jQdkBmx+ov+UcY7NF3NJCK6m3eY
5IgKQpabfHXVP0M/Zh218//pUq4CGXjKzwfwdwRM2wQwrKXIqxDfpNvS2WB0TNsX
gzvVbGonbz1GQF/Xj1o4UY2twZf+whUaKQP66BHmXDBJ5VwiXqqTK0djj4rYhxuD
iISyuHes600j2n3R4X3TSA6M4XwfTk2AKZ8JzjJaECEWO7yRNMRWok10VZ93lBEK
hw+FLoaba9L/H0knm01ils7teARVqSfH7yNQqt+i0of1MeRnSr1amK/+qQzYeTK+
BD2IAlgvhKHwwOOWmI+3exWPUy8ZuPqZG98WVK4bWpTDCjiTx+8KQOu9XM2bz5lE
`protect END_PROTECTED
