`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v+uYOX83AKIwXOqrv6fB4heyQiGkBMqzwu1xFTVAN83RunYJtQnoaj1cezsTg9ZM
PW2t8FO9ih2vWibm8C2ycDl+ZEmnkiUZvSQfSwB0CEWrLTcSr5UbsL8E0DiyT3HH
tTnpoKqY/mQ1Kfi9ij7KxNHqyPP8oJOQfkueWe3oPQFZGO6xL+B0idh1jgaN0JAL
S7grFVRQxqjE48UaJ6Jdz1OZGoNUYIwjHiLrPro1iCI3+7T2UvFO2qJSHH/tuAeE
8q0VVoQmB6A/R/DcnyKPYulrcpJ/PLCBflyu7S6DxBHrbTNyGhk8Tl8x1OsbEn1C
L2MVqBe8LUzdWO+9rafEgZW3VxnKUKyUHoAtX1iyaBc3irI3Vrj8b5E+2qBublfT
VdALO3mXr5BcG/ktD0TuI7lIz/14UsKsjI0spSQS8EvblmspOXEmneN/HEnM71+8
DCNc3CfwvpKxW603kRKH2HBJtUmVpjlvSKfrY+SuPAA4jw+KGjQ2MJfxeHhwHZwj
AixUWlPMd3mMV+AoDgZCQYDqHdgCQbyBlOZDW9kk3WQy7IAgAkyDRfIgIrP2lH/r
5DaT1kgT5vVnti+klvg3qQYWt9ZOpYpGPoClCafhswzasMzwwQpoMwSY5mULDWWC
R6yN+ggz43S4sGgU7wjMwmxjT2ffWLVT1G59pbeECW70IRHCg2G/76vHXMo/8OIG
4LzAMYTIxZMtiJgNRH5lbN6ItWQxiz6XSQ0CNQECEh4eK3/f8tciFf2kHKQz4N6p
ESry0W8X8uXL1UiOwEBMj7Sk862ELaCgJdfesZ9ru0rtG6TwkSM+lZzn5Ntb8hFB
mXpTdm38yqTyNj1F5DCcAZbl+VcEBuuiVZMvTeuQMM8=
`protect END_PROTECTED
