`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+qaJ+CPdCa3rpPVXvrzSgsja8M78LrXlBzzPCWowbtgB8l77fS72MQmf4Tt9r4qd
3igEWbmDFChNARbYp7kQrZN1GNfijRlLhqwjTtn1OVYqfo2w+5CemLZ/GGgnw26C
OHeGRljljZHLnYQJlf5wKQJkHKhmLn02IQw2gXbd5UTzIdyB9W4/X2yugkPwX1Hl
EzZ+Iai1HiN/3dZhDS7/VtARtO5H3fC+/sTeRAnWYVfIhyBLjJsGIr63W8gM74eI
+m3jY0az9vB4KaDkvhF8e+XJWOhTHWNrgf90GEU4DOr2ffP/upD16sXH2TKU8Jzk
9EOVKtNFzARlUGK6KnlZfH8e+am+aCpOjaEoBQmSmONWhGzDhAfa9UJuL4Nyp8Nw
ocy+5wp4usTTpJtesHXNAeuLl9rnwPoU33BQC2A5U1WoC83qXlTHE+wEqhfc2pMV
Y9E2HfQl/ZyHHPZd52fMLryOXhkhTi0on8Z4Ixup/+OpMRGw9+z05kFE9JpPgxNa
zlvrjgCIJJNFUEV8JGcVlU0eD04Eey/tpx354foOXfxhGuJfI9DkdX9UOWweZ8lB
6QLt+VKx6MuAbCLJFan5K9aw/NiY0DNREr3b0AQqdDXW3U9IvMsxUMyZYWa4jUkt
QgZ8Hch196WjGOmYQ2ILNglP/sgRRJdYuQquTrjk5aYX4BhaZ0UxJRc3KZpW/f/s
vgOqClthPw5WQqvc3VUr+Kuml1QEekJdq/Uv+j6cvvAL7AUU48vCkqFVTwYbb+pb
u74LUJhjJdYBZ7wX3PKwoG62bezECSht96g3XIMM7n1+GHgOIbVToKx9FTmhMNyh
NgEdyKhjOzO4RfM7Zq2oLSkcHd4B6uZslz+F4sARK/o+60/46OUo32Pq8gVIgJyD
M5bOaPeL3HMqZXGlL/+27BJQoDBml//KQ7bZl5wizsLmg04hTVE5zaucvgLzb61A
hANcpcXBek2riH4Z+1Miovm5ylqStFTr6pVebVYSPSgCwrMuvgJ4V8v+2O050xTx
oIXb2Afh0rz9eGNAKh2wHKtw0MxHceOUMxSzlR4/CbDZITR6+VFiB4/5r0yI7cje
AoTYiaY/jYPpJxVMprpWJHi62XJY00ZK0iBeXtFMk/KIrQTaWZ0fBi7d/aWA1CDz
AZYptVGxS46bMOWJ2mF+TZEBI8pw5ESETpLFnsx9rpA2ZmRo21wFW2VW8tCcNEAH
RY4+PhhtvpAZd0ZfBbkDNtURgkwUNkpk/SKZ0dj2qFYQa9QrCl3aDgfe4l0ryfaQ
1fzjZJr9eTLHC7KdTE7np2rOj64x+SFOEGQggaoo5rI+8VsCmfprm/xAX4aGuszo
qYF8zIzGD9KDq/MR2kuFM3P/FP2zV62yhr43B4twA6dZbp0owi4vXOq/D4+B99CF
p8LfguiznNaX/GUBRRfht6B+dfrJVdSIuzPuhesb5lGvZHEzZh9++vdyN8E8ZC8Q
jkBfL9N6JqO0+1SXG/G3XnjMCTudfgb8zPXDBhQIauTYFo5AtXtZiITsjAPOu9ZU
tMrNEChO9346MnpE1fAb7Fay3Q6r4WbhVf09Uuej2FtE56/qt3lW1anQVGhAz71G
mJf/9uvZyVt8cQOcE7JoujRpLMzpshWATjEzbfi6LYSGOLin4lsgBHCKML//ezEX
VgnV8JWI867JeHnHVQTTW35qYpLPA+92MQ8Vn4PEGFgNL1AH7m+eXPKraMkDxT7w
loilaF2HABJ7z3U3feXGRbpxuEIMqM4LECaHCqU3IJodGqOXgNbEdnBv52v2bYlo
Yc5imKp7n+NYjm8wP69jEElyhXCFTw5eJ6RU09Tq+ND5xvyPDqZ4AcfPAcyvlPuB
OaMk/rnOOcZxGYBO4JZRz9g09/rFtfUDtGjIqy/AaCfzNUlK6wU3vCCL6iM7DE7g
ZCzMH4aN73/Ii0h9ObERFvHk/0whTZjGQP8MuYZmD5lpuVmgwoCm1z2PUhEzO4UR
S+SEt72w0ad5eqqo3teJVquJGQy1AALuviApEIyOfkEIhT17yyahsLOZUSE/aV+W
wGgq1Sn5pd3by85h7BodvIuHr+impyRlOaJ1NrblJnc+pHKIObmCVef3Ee0/fsyN
MSV76b8RdJTJcBfhvngojsj9Sc2U6jLJrnO7/eOezpPjfjg+c9+rQL1AUHX2Wtgp
VU3R6pN5QPdAwKkZ0XxzcDh4musTMEKfV4cy4otIwwOGUZaGhxJbU43jNuNkHuHC
jhOO5/Pf8FV2QWPD9pd5FXCCPqghym5VptEXKrF9DRrfO+YyEnl/At3NodCzPRvH
x/ha1E1lb03MHusbsWtTTsdjpO205sRnxb7HcGqGPiH/Rrx9DJdofhf1v5zPrZZW
YABW8BDg8n3NksmlXpZIvm5OvOY43S3R7RyYqsy1KyZXOZQJfQDV+kCdrTHZPWIA
gLY/doTp7GfqBSRbAMoH1oqR/kV7ybjzCGPKGCLh5T9SYfMEZJnFam++Nd3eitE8
lsVzuIvJisobZ5zNXBlSe8pMA75w/NtZr7QP4wr15RPwV5Yoke1gS6dWYqAiyC6Q
dzObd/MaQJ2x/i28GeFSRZ7W5KV0VO57I8pvdACvmW7KtyyMtIc+lzs7f7Hs2IG8
ojJXeabL9Zb/j7RcVgZfqwKlOhDWjiEoKMpFoye4k0C+YJ72+uPoNzRhlRKocrYr
c8FkMbBlD8QfEOFQcdtxahcl2Eur5FrZo4kgC9C1B+JxddYKYZGPUSjU6z8BqYcj
m0qTedwpXyFD8ctgQty8S0NBdXJ9eAuKju2SEigFmLCc5pxn2LTPjbvsbDpLHzmq
khebIZSxzaaSrnetI7mgcII2kTQlRVqlI+gV2Bqoxp8d+TSq/RS3O2nyCQ/7hA8H
K2LBrFq7bgULHr1HYfzGO8o+1lB9KjIHVbKosCyVF6e6zwTvB7aQNtJGnzLAMyEa
Zl2QQnOoG2LJyQ4G2mkV7TVJeMvjqPndxjKy2LjJMhPTC6010FRW4A2Eema6JhBY
pm28ZgikagNQrLH4LitprmdhMx6BAiBW3Ea7vrMg01LeRLLTwYwBo3a2iWxkg6Sd
zobXIGThI2LRUjRuwiQPVErZTKocKKKFUDGYZP+KIa0nIJgUVWZ9+SwM7PIx8O43
LHXvoJlmI6ClrqYmZhO4mXsj2cifrNzz77CiMoExM9cmVVYIpSPrKaQZElN9gvFt
5qbjJeW4FbCCav64TfwHb2pjE0ahLS4pCBwmkx8szNyQEhaoYmKVl/RcAFfdruli
g0Wgsr6tsaGi/ZNWxg5U4IyrElhJsPIoetK9UhFbN6IpquDqtuu57S40ii6Zma3v
NQt1aA8Q+YuRsZ0awaDesy/JEcoVJcq0ZlGDB7bE6NLU4sl6VXYQZNdWHiP+xAmf
8dV1IX2OptOQZgb0oc9NjIlsDRBjuLbGOEaEg6tap6+NnJM//3Sq4wAo5EpaoD5N
RbsxHw64KYXEp6JZ1RHpBXl/0dQlbbv9JPIi96hHnRJJS+SGU+PJbhRV8ZZOw8Ew
d0yrI2Tzx7kLft1uTfv1gHQHOJl+qMVwGBZSdmRlgeAGzPiRKvf46JiFhz6Jf2ms
ay/fgajk+PwcN4oxFKqH04RJ6wPwYZndBArHAuPfY3lfD5nPgDUfcQhaD/pLbNQL
v2DYCIKgMr8jodwByZmox3XSAWMg0lp9cFB35kk8NjSMBmQoV3A049Wa48kEUkhG
s4ER2yKllgc/6iAzrrPgdoqjuJiOqrc4jyXiAm9X5aoU4XJeISHP6OgOYTj/0jwP
x6RcPXx5oFs4u8a/pNOnGGHV1pVeuXijfD7WagE9yL4CeZxj891dPyaWFw5CDl8j
0ombCNj7xTq9QhEBBjr/eH1J4f280ASvsz9zXkqhcrVKvjmcrKr2ykjuhApVHWBS
DhPhRxrTSyTqU8D9MtYMC+OaeKnAogbivfg9tZtrKeKwaIzXU6MsFlbResHqTLYY
UWveG0HjDLy2U5nKSGasU30nw2loKgYmnKY9NMlwD5u/X+anCAhwFhREb/VTOoqd
lAW6UwYYCrlFI+CVicMxu7O6v5ORhH04ICCfl4yEL+gHjNUT9fgLaMR1MWOv7hoJ
P3/RxtO+zuQ3kkHuSEv/hdy3Asygp5sBJ9S6Arj6KQl9N3AP6Z0Nf1fheg2wa8Jm
WrwYu02GJ/oVpTVajuUbLZD212Mpo+IDQ8SlQcq47Y7+J+FLqMi8qZ3kd57bTegY
qQsohZcp6J/mX2oOrhf4bUWCw53HtimkpCQHcEnqM59mEj2Lj51tSpLXnD8quC8l
Yxn5AE10RgNSFFxKyco1mh3MIQ3AJuC8oOpzaFjSa1utT722GndfEL9Dx+TnLc0X
YCyX/zzwD8yUlqGxXcRnfHE+8NoDC8iaqfJuVcfiDdeU2pE/8zWYGtBA5jbO/Ztu
TSlk1MXWZzZTz4sXfTPh/DCr3JxdHHqAXWmD9mPNVHYGvZ86Zvv6+ZGkXLgQyLZx
mTth4yZSFJbEiXt+UpRphHlc/rhr/QGm2/OsXngYwvjYen2vZb9OP90rR+KagzBD
M/x9X7/dhcPTWCfLZhdpQk8/UpXk6atMpOtXCn97HPOOlRWl5Afv8N07fvAwUZDR
Ap8Ee0lkT78DUwjcXBL9qTUQaQAE6Kp7499xnHshM1rTlRebBSXBP5rIAMOBF5sJ
vUzIwoS+ZduIH8MWaPVF7vcnT2f5pfakU/QvXQeCB9YJ24OfXfTyF+tNQqQwyvPt
+Nbuae0deCEiQ1YvIQqLRm81Bi2j5tUBcI0QrJKNLj+7rlaX/Ko2h5vRHN6FiO1p
HGsBT2yjlGBZf7gERHiJlti+6egyz6rZWxH7VHxwTlSuIZoPV8YZbB/0ZuygfPFl
xSHK9Ogh4/lJ6BqaFmvqYS/Wv3i+czBWgjHQul3t0Mpx+loTdraii1C52LtdyKjC
J1lDIq6x6IO6igxGuZ9nBQd6Z1zMp4Rv0R++nrcm+DqRjDe3Jvc8IlUx+gajoHmc
yWjNGfcQZuBhynVra548GvturQ1gmXpy4Hse9dNBqWzAK16/aXNgrJ2Sh93xYoHJ
rINY5ZIAwzfIC0q6ElXnFWw+RUacW0NFCw5qwA2GIO2qDehNNEhR72QFHDoaVgvI
D+BoAft5Ppecf8xt1CxjXdtYTRf4Pm6u9cRz97d/fGHKhQVHH2uA6zGbDI2/10wU
cEzIsf4Uusm+D/h74NW+6+LbP23vyhfB/serA66oBmB+SyLr7QpwBSdnyXXVA/If
C2FA+FsCHPyQ6+uUjDQ0sf8lA4R8Ud/8e3ELCnjbxYc512X3bxH47T+MSCQTu96Z
+0ZZkl5P1Nb4zSGF0IGZHgf9SFDcKJzTkBUIe1YnX0lvgHjF+jDT0sa4BGutBF0B
oQEES/ffzC9O0wGZUE8J3spREsqztytK25I68RGc/oScFYLsgvlu5IToC4YWjyfw
0KP6WAlCYki5aWgrsCPEStauiN6cbWOg4BUiviIUKTwDRDcti85KARYnm6LlyQdw
2ybVKI7k4msYppcmwuncP9wdZDAq+Zzd7LhpLtY23ADqNSzSVF4LHI31Tgosvl1B
g4p1B0iD6NPhw4f3surWWZj4BxIT0a/oSppqez1DPJxTReYrsa7vVpoRSF18pgN2
uD3/3E+TPsGgu9cLcw7s2rafxC9LYZz+13q1RnEPL6e11HuuLOPwts4DhL9I34qX
Vc+8EYZd8g6Fc1r5yiWMwAd+Vbzin4iaQzkcKzvJuPu548I4U6EM2gxcX7p8K+LC
7RL/s4xFIkBqTX3EzFDqYml4f71HfJQ8k1vPvIPPrJC/NSXrmM/gMV+jS8M3m/Q4
oPTU7m+3iysZ8ItwQR8RL4H89N2U6TvsXB3Z0z1Ubp+Mi+UKnPwj3iIyGoHEFDiN
clUFqiliA7tDDGeOsV6Qe56/3NrkvPnUDThm7NaWOPAMKDzblrw3V7pgJjWnwE2i
jt8OmZfTO7oCF6N735cho4TEmZqttCbMQb3t8WycTz92xZJRu8vX4aNqKD9U8IzI
hNMUcTOf3z8hEzS7ENWmvuxDFOqmHl6XkZF9REUDTiGJtgeSjq+zQ5RUbnp5kUy2
Qt53EjIkXoTuZTBNnOalFpQ+J3a2K+5s2ADbPR265Eg5yg+Bk0W7SQEUXe2rTHxl
DVRYM4Zy1vXjqVYIU1/97SNL+jXFOpuoGNfqbh8O85GN8qCdNL5mc/v8mrVpSoW1
/tUd+B8w2AEHE6kuDqc2aSQH4xAVDJMXbiVFn1YUMqlb/WwoU2FP4zGmcdMOyTyJ
KyseBd1NCyLhL2R6i6cghYnDTbx6h6dT/kuee66c0jhXgrogCcxmvzEGuV31t/+V
dSOpXWg5xJMFXJxijnfSq5AV1IN+oYTkKeRw8A3WmzpPspZ/JPzy/sTZN2trlh5P
E/T27+v+jUjOBsiZQrOV7RsjcZYW22ZAdl1UR/vYoodsFDPA9orp0AgEc7PKFEBQ
puUhJFTx1X3pnZxxNklvhioizr/5CrIs7551dvRYz75gJ/soK15ywJDrQKLulIh5
jMOWb7N+9C4rwsM2F6hql+S8ZedN+tJ/bIf/C4qudKeErzTua3qlVnHFmbcph4xn
qo5HaVpchLa7xuWZywjEjJFF8fu10GxtkvX7TVJZpzaTAaFv6FQVJtRcfrUEJeIG
JlPiVuzWfKSja4znJix1P12yDVf4GG0UGpnsJMfFzp2v5AiZmod6ZOpqR/r40XA6
ds0CzCrzBTrCZx6E5aeJmF2rIxqzzWuFEwJSVdPT5U5yHTAOxeHMBB/WS8W/Exs0
+N5MfsvaM3Sx2Oxx6pFDJueIYzEwtIEDodoSwiqUtyMNIlow4RKGm+BfSF3qWCfV
ZkYhhOH9W6FbodHZUkVB+aJPTEyj5fJ+wOS6otndY2rHKmNQgKXcCniav4l93vuv
kOEeGVGLbCNnkUCJY60vWAkKYFG71Br/0PP0KBqOz0DUGFt869QB7TgBwqYMPR5h
HtadRWoREwGCFo9OYIP3XDlpAu3pfKZykLZSHSod386NJ28UpGw0bvCKyGBV2Ap0
xhn5vEW4zF2xjqxIjQ/4BwzqwVjH6+d7ERsnMDbY2HqldmeAks2JQmuH7jdmI8Gz
nT8XOmg3UxBHbLo6ZWRh5ztboDTbA9OVpyTTgFXY9mVvCt2LYSlv7upMTHM7e462
ahzJ2jlNx6iWDT3nj+c7c5Blv41A0xeUOfhNnzbJKc+QFcOGKhPKUrEpHuu0PmgK
lnhpKTxgQgCd9D+Kh8RPIqttfwemZYLKc8SuIeoWFgwWtw7Ulkxdh4GXZms9DzhY
kWTzMTwhY82NSkJ/xwck8bkQ0SSv2uBLQAAvp7+kUe9nN6VaJK7NE3armcI8z0En
LKVnGyDD+HGvRNuSU+HWn2339uv5CiUlDzLPhny65HT5pHKLcqm3HLPUcBtu1ysL
cwlAMZEk2hcgEteyYicuCFezYYi0dckl/15A0Yr43vLZa8aTMIwDTq6hgveAecPq
mKP3YsIdr6Mhy4I47/ctdvRHWCdaVgaJ8PRbMpFnyzvfI34FrrpRiVR+EBGMowmE
H6ON3Xj5wLI4DqqM4nYfNONyHt9H7SEMXzZKv7vY4tRMXhWEHv6DrcyHQqGr9AcE
NoHJzqCJVsXbCjzrvUALw7pxKzawJShSxqAdO/sUXO41nhH0wFhCCPeUHUjov+mj
O89y5ZDiZuEbezXydxE8qA629S5TaQHki6lYJVbtPts+FbL6st1pe688eRuAuB9L
NFfrSwFjQm06RvnyA4IyySf6tBAh9g2bl7DbbD8t9zlvGTsiWezcHa0A7rhS4/f/
r3iOah9aMblRU1AWF7GW5LekjDd2FapeE1gFsd+fWhqXfZfZ5CsuxbJwydrtPIQg
56W2XTFAEucHfVQI2FUbuq0oau0IvfEQhd7cPnlqVQZ16cMEoMgBVl/A8v4A5DYW
H9VftqLjne3fQXVcqZT5AfeFWCUnjSTH96GUkg4w/t8fU57S4BM4EjLFkZXkAksG
qeZnS5TzoLJEhGj6tcnOOO1fvjKHAi4ysCn10zUjm/T9QFzCQQJz9l4We+OyHNNY
BUjTgNqB94tYH0yHi8Hw7WXyei/ba+6YmDtAV4LpX6KQyKyUqkdsv1h/S8Q3YXfF
K5iAAax1LIGGYu1IH/6KLVkq/TQUUEun+o8RxbiYfJw1baofScJoKPvUOpGke9bq
tHuXuBW+PLyXUTcu8de7daFUugATsllTReU8ohGpOdb3n7pgb4DMpZptVGqCp/Hz
FDZqm9UTw34Z2e0F6520A+sdVU/fd0lh2Dz+fXleiwUULKWEFI1bRe3DyLNhcVlq
D2J+pYKbiwX8heRPMeRQ5GYP9KImJYCyD/nLQ5GJH2rhjR3mRFoMU78rZN2empQF
5fiRcJSiFpgylY2JuIYTxn9CAEWHyXw5QP3IMIU46MKYCC/G8r/RtDTHZrh5n7DE
LTkVXWMkumWavXT4L+ZJX461jD/PeS1Dpz3nGNPu0JavOjmHX7YXxfGYcjEyN1F2
JdDi372/d1thPcU8CTAEG3xknZrPDM+vJ9tqmqx5Cq4oqL8gwQRz3kYuljUuobbF
yAFGPTj2XuEvLFDYZ+bitOmT1rd5PL+tTYa8HYCjO609imMLDC2Bu+OprvJqdQ4k
wKuNCfD3Bgx4eSKN77wH7n889/R0t4SuvtfmZ8Bpqz1Qjl8n9ZVjNDDxPdVgcppi
aSOgPFj4/agvwNAponTxBoOp7EnDxZgg3AEI4xUL1ysTFLG8Wv6pwcH8HJkggwal
+yRgB6gb1IEUg/nZNfTv+ai+iGKKYgRMgq8KVYFtnhhOpG6KnmQVjRpZZzApwk3Y
XQC4gmfxdgAgiH4I2J+X0+LlAcpzk9oaRiSYCm84qoRCrN/aA5CulNj4fnDITIsJ
Me9JJdgS/Iec5ZGQvpED7TVICMYhqAfXNs7aK3HP4Y9vs3m4k5ilLln0CeopUISC
HH1QQaUUeCdBl7ZUdc4YiBblxiDrplrBX16ASm3w6D6jLRvkSJk9fcThNAty9tqQ
goTnDKrE+2wlGyQuwEx3vbtdOPDBEDATRxYoTFxABIdnH6F2mvWdCOU2r4KMFl04
agcqTPrpm9WXlKPtlKSeYFfqAhDMmX76TOvqg8Jl6zgI6zvjKHHDj01oS0HAZA7e
RhP5bkVGxtoAFDNfB7P0t4MY6bad1cNJaqH75Gh5SfpOx4lNkbRfu6blMmwIcFlV
HtjV/VF5VofXz1DnnDP/OjGRLKmHcrt/Q2oqQL8uDXuOxVUL+aFWHKLZ7eGRDI3Q
Ca/Cq8Fu7hW0aiRCIqstFFhT2RNcs0VGTUz1e1Y8wGxsL2IgTW+y8iOWWwA/YzwL
TilBciW/l8qgUdEO2A4C3V8KejU2h15d3zdwJ8b7A3gzAUhKFU75ofv2d8F2ee6E
zcpIfeP+zkREtpBQ9bejNZTB5jo5sJKUYyQvfl8xTjOZnzb3MrVyq0G6EzFcAjlM
oVSYRwAwhlyRtfsEmxkVyjoF4FqKOj5rm2K5L5OPTJlHR96KLNbzQVRHO4Jy08PT
Io4/qnZEL0JtGUXxc9LbKYGGonPmgw3sLRo2L44JVXwgKllRdE0vI3So7vWIWgj8
qxoHtVr9IM36b7FWHuw9XhCUGYm+2/Vyt5FRlSBlo/43KeYgDhEta+/OMb7W+NQc
r4LzopWNjHUQMXpkzmZBpbKPNnYfr+Pb5GfjtnC6vKHgN6+95EjWNqrFEg2wwW+p
UMkvQLQFODswQbzIWUyw/fGTrCXyeGNg7iBXq8DmhYZ1Z1h/UX99BP+6empGRGt2
uKPPGDC6zFUG3T01+87nayCSEvOuQQHsQEcL8J3nuque2SBqcQdCfdHHH8YjsKEn
39Nrb/nWZz3ZjfdtofS87+NJaBNmYYvi+fLd26i1uhPF7EO5GmPSyThlw+bYSLQp
QFq8N3nTIMiFv6HmSHE3ZabkLL6a2lQnX2v2mEHnS/w96pKSXvq1/IfqflbALrgH
eeqG17LtO2yNkwhD8tf50rLY9yL/y0gUmcKlXcysITXqM81xYrsajyQxuGlcwTiM
Lj0f6cVBDa94nGBzUaZBikyXl0SLt21egjVtZpREEDsvlpRF7ASfgR+KpHcb06nu
xtnSvg50edE16SyXWIfZn4VHavM5+b8lUthzZsJB1k8VeiU7OsdYyl0IZs4e8ymk
t/as8/PWdhcbA46Va+U2k4uJ8yX82x6Nbey/sZ3+/vaDPeLd1e+39eLm2k+iq1NK
J1S+EYw1mreeU9fjVE+1MGb0liOsaleTEx6s77JcXiJv0jaTuUsnKM3Du2Hlypm5
rv51NN0UqT9Utwo+RpvAcRLcs5GxI+NMoavvobiKb/4acBBdUIQ6h7LmRCzo1pBh
3jmJR2ScXMD7T2uCDJYcgAOQMpL2oYe/inElRuzvJBQLAIrpFnNgkn9Pt1xQthuJ
zzzsAKXlDu9kUAZ/XnHtbqNMJOYLXAcqLEVPHRc9PbPailZnv001Y+WicqMABkF7
i3YSZ4QMYEi0FNe9bzFgVUV+IIkcMTI7JWX3l30yDcDG3H1Iw/usjL2ziNv/wTfo
9ELOrjqdTRMaIxDFVqYga6pf8LhcPJSu2b/TXoqP90DjezqCvXpyWtcJrcLYDWiQ
/x4ledEOJmun1YtxAeybN+qQ/AMC98zzE1y48EfDZBIVnojvgYS4DZNuZfb8RwuY
zO69lyC2pcyUEn6X7nL87d06h9cXT0W9VV/K8tJG/+UL+2PQbymzBFCHD0OlZQ5L
6Kvp2fT6FjdrB3nswUxLPkwJA/4ZPgjewl83Xyqb+u/EsP3rCOLRm6UXkqqjWI22
akQnNHUKm+JD+aQIhvLXAxLp6RtKcethtQ/aQL34tt2UXJmcfQILil8uhR2D84ln
JgmZpknbFBXLXYmTuyYO3dc5Amvn7dkOBn6wuz6LHyS9CSb+f1E50LQGzUMCOUTe
uyowy48AizUQy8BcfOaBmHpxN+yIHUGxj0Ih2W0xgHTUjsv3gDmCnd87/sYjWBcq
/fzsK2FHB3yBv8slqV3WMhcdYCmBZ2zkHcpmcEKF4j+MgZvtA76GG9fqTTFAE/vc
pZNR3s0UNWFHL4AwINfoH7saLY9WwK5X0Pd+XoQJN3jvCjPtd24SAyQB9ycu08k+
sTk3GYWM0aEw+0ZkElBu+/OSekrEXkWVFAgPORBXhpyP/oaKQye4WNMcrhQ5tqo3
jh8sxTi7UJ6wHATyVAybCmrm0/5YBRv79yy13hWzcaiDNKLtcBq6FQ48h7D92+vm
gHBAXqrWN7PNpG1EAy3ObMJGZWBCDO2QZkoJnUVn3XllKpTKHvynKitfytTA+SbL
CmQNuXxaEH/v2/HsLVZK0olAHwZSkyWpOb8wq1nUyI7iP8mnzAUoJnT285XeadHB
ACqG6Gqwbrm2k2+KevRXuwpICn3COXYxGycN4Sg2OofobiNWychuC8AB3r8h9ZRT
1+rzwgw9QVoPEp9Y2mbY2r9pyQzFYNYQxBBggLoxDb/9W7+8EZjXbpgt5vfojvym
22rmYrSCSTo1D3D/amKzU+zH9TM2Xxub5X7c9YiSt3v6ppiyEod7ZIRJxr2S9dnJ
yP2dPjI3G/DX/y33pbaJLBczecYnqdvBStx66J9CRuT/J8mzyspBQbBG1lfo03Zm
qtrV1MWUSloxZE2Ffhxy6smb5hMN2jKRZr5ABZf51yJB0jagSuWfXyUUNvFTsyF2
EC3D41gQHZ1dwSgKjlFZ+ZP7iiUiK++FRIyW32EIqe/lvkaIeygbQ0Gho23T+5yD
Fxh3P7tGozCBYfvOHnpGFiRi45bdFma1h461gSVwxPkzlQzPLgtL/5PXCuyweNtQ
mtlqe8pdeNV7G2+bSlolTRpqoyqrr3+YQXkaC7V9qbkpDfJUxkKAdnVTZwlmpmgQ
z8n2X+B9zt22I2aAVtiN1uS6ILCp9Vt2kC520BxkXqk0blwNFACEtql8IeDGvH/d
bgyrtr28H6qgXGlzYPxQRBfe92RWofDXNcEcDtFzurOYyfvB9Ry791f+yUx8NLt6
E9ZFAWzspfUJUjVeYrlcyxjfuZiF90deGxxSOIwVsQyP04EC0H1J0bRD3NhMrnmW
Eg1/vEgQVkuzqZ3ACPRyfjGvf1gp2p0rXjiLGu+/yyZTL9eKm8MKD3eMSHZRmfCZ
9iKxFyMhxj93lJk0ixFwVHZi1qkvQi6kpJhCR8+jpB9/M31zC3he9xJkC82QcLAH
HbWr7lfWZWVJGdn2kFkAA8QBfeSOBXSFVVUKX46a8crg3lMW2MxWNWAUCmnjkp3H
Z3FN4GMA0z8GUzN1u8c9OxETO96efE4QLnm2J8CWncd2yYK33F+33EFqqbpQf+zi
CnZvyEfHvI49CFnrrhGTLa4shxSNPPLeubBGrTZLoBPJ9wJyyMQ7Y557jm3CxeAg
GDqp/Fk1GXzrubyMkLpyP9W0SkXmjB+Jsotw4i7NnwefJvaOY/rD9GM0kHJZWYKD
PXx9e0vAtOP8vinRLPF4vyJHLThR9OTUty4n1/QLr9HVRvrK0+jiwQVBtSDtjye+
++wkjOIEyuvaibE7gVNExRdMQYObtlIUqatoZgk16+w9a1JdVPpWpguzkVPj8/Ya
wu6CRu2Mmkgd0r/i6x/3ZQiVZ1acF30O1FMEJzQnh1z6ccpOETz5uNyfa2C6rN1Q
BKYLLPHNBE21aK9rR674wIZn3ByKT5wIkSQTecvIbE/9XmwSekCuVN11Xf1+sdu1
E7pP6tyHgQOLv5sIkb47Hx+HtARjQIL3NogpOcwhLAo8w26/wrlTwRxN7IwNLS2x
SOv5SeW/zsoklBhq/xaE4PcwX4ivKnR1NlM+6WZ+3/h2jLnqx4DzlFIszGcHDi4p
V33iVppAwhNrXM5z8gY2PT5Yslgql86IAIFu1jd449b+vaZU8s3AZmO72lLgmpGr
476Tv3QcQJQ37mgwCcv8xBNNyEl5Vy2v3HoK87Kcw54ePweyXlRP/cCxkMWqh58T
u23DNs84rOZd695jgwhsReR5F0tE6r1iUcUFw/o93Ev3HYHpg0YOVrPUM+n8Sl/X
uq5X/Fu/waURq1f5gWRn+x6kGtZ79rH/q/XvmDnLzs/B8S1Xp0UH8Qp/2gNfnj/P
0wkMVrZ/NzjinaJ9Jq54Si3kOA0Nd7fMENpv75AgpAZeJPuo4+eK+4FXc7Wn5eWE
SU06aZ9njq4dgffe5BTcVeefNdNbXak9ZD6KBx2oDiXjV8KAbPddDlxd4i0e9xGb
JlYyZGidCVdSYY5nY/vFliFyh/+xiOsz+0IwW+RkHldedUXm06oAVnFc9TrhxtoH
41tQMZ1kcXSMzeBr9L4GV6riKnPU/HVKnmIFjkU4J8E3Ejhr51psezhB/Z8P8jo7
OCkZSLEWALVdC/6Rrp6Oz3pRqcqwleb42nimpcdzNgnd5Qyo4n6XMcEWf3dg7oj0
Z38iR3/iBdRMcSrEwJpUWen/ZfC9bQwq1HCHusvxaaxoy3uq8TjogHp0hjb7NWFQ
cmMFlp49XVjdHGtkTSzOdKAruz/TSCol2OZda9loPlx/I+X/w64oYL8nQ/QQqzFt
3OnoBMSkrlXcqIhd7Lq43Yi05Z55iKSzgM5u/sHGRmcMWrO2LGI1OG5Ob7tu8/Q6
v0rhNumnGghFNxvCdzecXA==
`protect END_PROTECTED
