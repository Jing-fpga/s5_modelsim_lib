`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dIrkdVcMYKizoY6TY9644RdZoW5OE7AroAvvDkpAUBadck6uKIQNiXj/d4PrX4VH
GvQm6rfGbKKvEy8MP5uFj37Mr/aUWTwIPmJ9Zd3IYnJP6zDceXr4JOAvlX51r/oG
am50hu7r0d1NVoHtc2T8BY3UsmRbWinnGRTMpv+YR4KUETgI39jgq4m0De1XTVFx
I7dMV10CEbE85PFFTJvJCBCOlWZ4A6pMMrw2ZYfF+YypYqhPL28p9rlhNvPB+IHO
kt8OfHECdfICq8t5lTxcYKyYllD5dlMmo2J/s1k/5vY+v/d0f99b3jtS3yQBxDfa
+xLEbZdDvdnZ3/s++kh/bvctcuDDiAB2LWDaBm4sAYvzCFQXx+fXny8qW+/kwcTd
uQimxyY5+1aKUD527jg4DwXV5aAVjRn5NkaXgAUcp8mngObrYr2AbAQI/gdhKo46
JZSYZZLg48rD4cAFyAG89unN3Er7eKm3VOaSv62+WJwEEiQvIebUicLLuQ726mvd
pswx4Cf9FuRurmSnivcCShZVsOp6gRyIAeSu8uMBCNegDNGJiUJi1rwmfue7psFt
L8QiydYrOb3a07gjupUo/qtvHGXwMkaXBSrWLm7DnpSKqPa5Sx0jsh9+D1FbyMzR
74Z5qqfBJzCX/7Rd2+2eWxSdAzAgm7GnD/8RW7ftvmG/596jq58c2oSNKWaGw/PC
NgCic3gE26YbTrLHdK9Bz/9a1dYuKk1hA5ntv8EQSN7PWqZdNuPnaT4YAoezcPzs
v/2mQDjU7loBZiIbqbTZYJvv64gl4929t9Wc3DLkrFGIeke1cG5Q1R0mOPYw2XLO
W5CtTupcm13ZpWE42t4y923OdcikG6ru0TlGZv6Nocf2Sb62K0yurhzZEeL5Vw+V
`protect END_PROTECTED
