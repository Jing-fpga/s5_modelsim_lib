`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
reOQ47AByBZWVO7rn6Hd3qLl2LwP8pYjUqz1XzUQ+4AkkVvxF0HZkXk6sJAi8HQ4
tNDL2snaxqxfOMYb3EojVgZ79gZ63oVdQwSeumpaVpIy/tVnrD83ai/Y/9wpsoW6
TJ/ccNcI1R7PiMBSNSBqAoyxhnhX+JMbm4GLaK+P822RX+VOilNC0x0gh9IXntoc
mcLAUXI4BGFN3rooH9g2CkTJqfZYwp+Gjk1/1bxoWSmHPHPWm1FsekYbDAJajkQD
b1p6s4Jl93b50Lx0f+yWDoPaLTImtmMZs4zxHE3BW2MkTlfEgHLbfsJfAD91Gg2N
JUmj1x7WEfq8i9yM58wSEwMwCzmnpe6KDPEnBxjOQ8tZ4//sZZ0AFr3wgSpZZC7z
JTES2f3x/83DMf62CudcHIwAYmpd3TpfwkRnTwBDxY478ugZHnjtcPkpterwkm/1
1CDuWJTQVt69+xmlbLE2CUiBNo76eWuMvQU3gy6qonKU98ypK47tM4cQo9ssmGzJ
SBWEYfax5kyQiw+jXspgZQukewwiPkG4R6Aj9AB2svBYHzVqsCnNWo/0KyfoweH8
pOGaEhPLvpw5/Ji8N2mcpQgrNgnly91QTHgxe6362Q0NfxyyQa9paPa0DU/b5FoW
43IZ3W4i/2nt0PZBAJGvlrhdpXQNorKii5VrnIjb7mGVUI7lgOgYaHzRSCpDa0W9
pAcEufWhcpOzaZFuhuMQsNz1p3MGaPjm7WdL18nCDkKipn8FmRiZBcPjmncGswVm
Ekje2VZS0Jb0jivt8HuNVnzC1FTXK9WSejND0Nyz22X98pkYimz0rgA9AcLp//Pk
AzO4+AGTxZeldWnWum02azv5KPzSot7JTVjLsKyHvutceUPdkOSSfAoorz+mgMAI
QoNvFl8p+uGsVKtG+9IpiAt43VvDVNy15a0rr5e6OjQw6u/BHzxM72n2scZLYZCH
8Knp2ea+R+6bbHWvThugOs2AbHv/4xwsE4JYCb8piwzFrl4soJT9pdmzOscFaKHy
YmExXAykaXPJlS4YORTxahNASjjjGacxCUazTm49T+L2fC4Jv3XG5ZJpO1w1i413
GOKxETbwW9WZAIA6Lj9kihCBBIjfaXgM6amnqb5MdcECjOOS/U5QdXvWm6gSngYL
DlQv4OzSwpTofINC5qfg7yDhHMqPkBVy/3NaqTkRca2hsS9jm6AugR4tTaI/fzaS
IHqIJRo5BPQql51YUuKuHtv113SIqWZ+zUBZf6nkVPNrmV3xJF5OAWQnec6pmCOw
kA7pI57UmCQ1rxEp1sxWm8S9zJyvZSt9B06G8/6OxzlTG6szc0MEQzecoaLdJ8JC
z4FCBgr/eXqSYSZXnElXBVl5mXiZl+ZnoweQDT8zyqWVzOgkRa8JJ1+idA9W84uP
mj1oNoldwZ6edRMFJsJpme8K+UTGcpc+2kztepGUhtLXEp/RwTFaLlLa+AMvVhMB
PGTxRP55u7n1CW9bEq/R0789Jc1PN8EzzPgTN8HKNPksbKmn2k56kAAiWITSLD3W
/qsBJQpZW6TNVGcr39/5bquwKklYxZ4hrWnj0yo2zSuzsqNYRYeTTUM9hOAYBDW5
JbepaIJ6kZdw0kClQ30qzzpwFmPrMg93pv+bpg8O9yv+IUM94AyYGH5G+l/Fq34s
1ZR4DJh+Q2zARmy/x0829B3vyT8BWoA3Zh7kcop/g8OenQCXowjqzWXfa9feaXQJ
azuLbacvDgLl0g4sLUNZL14pyubCvptNkn3sbQpSZP+0azO+pRAy+CeIz9HNrckl
0T5GYjo77pCzJYzhT6N5t9aw84zzwajIE3WXS+TeW37v3rKIdRiAPLNOXgISh7sH
pzjCa1IntV+dw3CltLuQ4sLgV+m5i1izYLHcDDP1pfuQjK1gprKcbnNz9F/i82N+
1Aen4Tc0F/nkT/ZHHdy6/Q9RDrk+E+R4fZjN5VClUgODvwYBLMpf6slU0rBY2Gx9
9E9qssXmJiPMHdktk8HQBhDYlxDZGHp2P4WQpndhRbKqNIJS5nyts/SVq1l9WLO7
D5kYFICiNnqCDYtuPClHkTjPp2XcnUmwdogJ0z49zptXgNagc50U+U5pv5opisNM
Syfdy55zaDiBeau8wcwUFQ==
`protect END_PROTECTED
