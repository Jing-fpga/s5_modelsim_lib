`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1IgTEmM7T7T8VCUV3WJ49LGUUNQsb9uJcyb639+Ie1zBRjY8AU8m8+226Ko3xohK
84d7ENZ8C/fES1XYYpzd/b27uqGaKG8sKMQhdfTdsMjTZjexdIvnPRng92pKDKCx
JswRCCESOdU4e9lf6s6Ji1BvO4D+RXn6ifk1Q+zDNj1huReJ8t4ZzOOxUBHHmiGt
cGR4tnjzYEuasgJUGdLZVwFtT7lAdtY7CRxEz2ivUUnki3/YCgxsUl6Cg+QgspUv
iMRpXBLrY3aBqLgQgb8x+1eITrI8lHv7F4P4NAEYgKi/NbfT95wT/zcLW4G75Wyo
kd8ArPdTYAu8vmGAzOUhW3FsB+e3FCRZJYiDqcP3jK++KeCPQbJTOHjto99qfYpj
+cPKGbKQx1AfQefMhh0WMeAbCuMnLDMIK5v1sRIapBpCtr66K+KO4AJR5Mk6JmBs
uuEJjv2p0Cgz3xotT6c9NY94Aaz2rsV8stM+WAZORZ6FcRv/zykOjVdOZ9NUdCr3
Z2WwPh25Uzw9WXeM+D3CpBec/AscFmDA6yWfux/9+C5LKjDs5CXavlZMk4fgt287
kn0kJ8dcxfxzD3RSTlovI63U4tHHnLD1A21VxaOsvaPb9tX9CZvpBNuTOSf+hyse
HgqT+G0hilptrKVPNC+lMMrqjPtMDfKl4tr4V75YzA3WFrSz6c8YOl0kEA0vtzwl
414gMxVqJVRAh2SvLNoTyvu9Oq7ZIQoBNojN22FwIT7YLNIiRi3o5+Fn6u/ygZ9y
Je5XRMmo1bRanR5AfYrc8RcvBwyIK1eUag2c/L2QxAjETW1BcxmMPAKXX5lNe94l
1F7H80AoEk7D4w687ItcI5021axrrPx60OPpzEwjzo8uOx1ZXeIAbUGHB4t3ptn3
bgMuKwDE2mx94FY2dBrwRL70HErV28yQDj2s5fqV0DN9fqfJnlfjcID9tjDgCYwh
DfYuBPTeZ2eLLa53oDvOVViTa1qqFXzWM0rpA3les9t6riWdLn0Hgzks39Aeb742
Fex3SQ7NCciPvISMzaSTorMwuWsw5fBc4pW05lTYCNpntXCe6cfAbyzfMlRX5QxP
NZ/uclcBoNRP4+WeHho31ynpIL8RrRouIBVwDKYsFnsH9n9uHklidE6N3xmtolAt
qTK3ogV3tJtHZAi99lcxLTZZm+VgME7nkP7TOeiPa4oW5icD0KLGDUE7kyCGS3Uf
p1Wd7mCLd+GVpXoXOamoJ3fxxPzOAkn+NoB2Xj3m62eA28WeoAzybs0lEXPLn/c+
SsMD37ViwfnLbS5cd6J4vDE1+alXvK+WWlWvwXWnQ8G5I0BceCtcNPGIEJIcA3VE
ghmdaUW1vaH5VzTkXQy5jdMnFAwjkPGlmX30NJIhKDx5MSvlkYOjCdcBWXjf39/v
HKyp/gBfjFOu+VyucdYC/MBaasMkV00j0N+WsqfO4il9gO2cNQ4ZuCfEKN7nekqn
Ockgbbr1pgi2QHh8hVWr84cNnDRaIyKgSLrNrC3dHjKWT6sD37sVdS9x2A+Q/w+S
JWlsvQ4mW6JAODcGTiz/WRm9G/Cp+0IfhsNxf7h8XA6oyOsfnb3sHWbzLIOIS9uA
iWvPuvwQ3c1ydBfwbdFbWnGAXZ5vMpdk9nrNHOW90WUGbqjs1YRnScD4X3ArfCQ9
Bzadqee/JfqWOOiP0+z5yHkIPsc4ztCzjJJp9c5xKBUIl63igCv6qLx6+XjErBtb
akXDDv3/sbbE+st7GZ4aWIScGf49hhEBJug6yMZ6MWaF6H310IxiqCOpBsDDbBzg
JGMud9bm7ofjj6TOApL2NSbqjLoRKtQOEWupsaLKyZFsV+kB0TvyJEKo3lgXUUzL
30PLLzE3MvWDLRS8cRa+b3qBs0SPErzFhLWPfLB85m0Wjkvdbf+IksT/JXNMyTWx
X+hwCtjaEkUi5ccCKxixMYwdhMobQ07BYNDdPcC4POhNtwpydCLzEqfaXN08Ke2l
PaA23kAmtRYOwUpfmTpV8GW3m/WDopSLW2l2FCCInfQjqilVuMiwAFbynWcDqG1G
sMv8S+E9mDHb/BrJSm+xSWAeO/W1XwsxRIzOOp1k2/6ojbG2usNZCtSjSD+CahSg
n9g/DRlU6Kg5zAxP6oyirFnQ3RxjNozVqNezl/g6p6lR1Fl/BvMXIe1OyR/rVl0K
BI9s7JZNwZqlHvOyJ+1K9YcfvdMmOyv0WDX6OksVteOQ1ccTo2yql3u46fM9aak4
iNAzo6X16WlxlOybArQJBpmOk2/i78qC6S3gOn8jedQ57VnJIG4IxXAA18J5qvSl
my8UtTzuJgj30suGwXZ4ysuA6YzOii4e74XlN62yTZQ=
`protect END_PROTECTED
