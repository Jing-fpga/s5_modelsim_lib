`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S/MRGPyu3SDqh6pR0drjvS2CByTty32jK5q7ya/rjgrxeG9fZBu6o0g7bLww9MKI
UBwbVhcUpHeSAYJSNqiiloSoTkhm0yKqyrmMtjb7Bfj8fixYkQA++oE/FvPDM/6b
gbzZ0fp92RrxDIHJMmh7ec2XVAbRLU/fMQR8wbXnTeu/onJg5XxsKaIpnhlU6fpb
rFsp7KllNYGgjHzf9GYoWMODdALjtXSEk4VFdt01xTq/NPjJxGbko8q/feB31lpT
gm9UI38dOg5biBQxsjr7JpphdsKm63zW/KKmHX40Q4WlCsUEd+vVgXBYUS1aEDm1
+Las0igtNdz5Wv1EieUzXA==
`protect END_PROTECTED
