`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6I1cSkFiTXwhblRkU+vKcCktqL7pSN9IhATObh8tVhsq6uvjnk7cfwXZRVv9WWGT
ZTGScHQuQjqLjT3AXB7Ytk5IUw8pmQ0FwXMp9WED1fvK6nLuxiqgYELqfVuZLYmu
kxZJapvr7fLwVAusLBqTctOkq1kuUWWRbJCEPVJmUWD80A7ixlKVflrJl8H8UDLb
xkS/XIrdk5WPOsOt7F8EXgbMV7tXH0Xo10N0/NX21/GSlUrIKi7ZvgAGwtCjPm5H
M2o7AVrG8/HDX1WlUKHJA0o0nIdZ5SnbH0+geBZuWMBLcE60A7ZXbmD5j/w4Y8a8
WqH30oqqf4JYFi6vFqeIySqf1+W7IxzSTX9hamdUoJHINHQiMy+29HQgPYkKTta4
mJ6oTduQsAz1ulO5D56BLmMlatZ3wG/B9F4XJBH37iJ1MxqJoQZyU7oP3SiQUOU/
LPtHiAV9xklbnd63tnDxG9FYDzvrhU3VT3EAYT2HHm02PQ5RQNdYit1gPXKH0crJ
b+wwJoFXv+Wnoa/2MSSDO3sjYpu/GgLdG2lq3Z4OBfpD7RUEoW6Hr8RBgh2H1NL3
4AROV2sWVHmeaMaYYdY6gGH3BxdEZTjVVZ/Kj6QxdmICBMXTi2K/k/7N44qeXUQu
HsFVhWJSuxYdj9wyfx6eqs8da9g2rKO/NM0eAYy9ffm1/AtKjWi33+cabNVjdE1S
NEGtHptJk0lPJ70FfJTOKguUjkZwbKbPFmE7+AQ5mWAoqL8d3vIjiSw1TfaTc5iJ
t8NVh+1EF/9IAiV2jDE8oTUtFWLbmE31eP2ULy/FSm74sZthlrZE8n45XAeXIdzX
JvUzWYX3ByUiXbckfwIH89f3h2w/8unbtqCEnk2OZit6HdvLPvHY5+wy+M3A6kzQ
SPE7Bpb8R6nDfbrGx2OcKJCOs/jzEzTsjAB2jxsVg3mDqzK6MwjTIgtWMr4Kmh2e
/byoxofmnBBo47fVF1xLMZVE35V8Bj/ykLF3bkjMvz505rKDcGvyIhXIEqV1lDBk
XiIkiA/+tRj0aREU7fQXHBXeULk2JAzKz8r9i3aSs2HJWsxB8ChEaGQpTwsArg1L
kvfpvi5w53S/Rcgz/3iQEwNdGfU+T0AcGgJDmbiDYNTPokfXKJ4ui6yDLT60gLuf
QMUx8JGc9ybriKq32OZnGaFTbVPbZtqfGfa2scctc+Uog2Axy6YS4ScWrN1ANOEL
VTmgxNyG4Dp6il9sXVV8tvelGclUm8Scd22ZwJHi2WMVQFrJVgKIsw0sGcSQXB3m
WnVKuMB2UDX1C8JboibIn4pdjgebHdCgsCSc3VOHA5qIZ3VwDUXjfSJ53sOJwiBZ
Cb1wRoJ4gbpyhhS+L0BNU2b6ja1BG7UDLnN3u29jq1sCwd9BgL2JsB80+woFb790
8mjmivAPMUs8uyYbIHClvbT/KAQuqbAKwjbT/U67jh2Qs8J7Fua9LxZbhlEvupui
AWcLVDk/iUiV+FGPfakFl1rNQU1ordS6ug2OYiJ3TQvJoqOU4V+TVS4yIEku+j3O
As7lb/MfaKg8dQ7HVcikZFhQcwOVxGJgmjnceSZVK41UH1WdNAZnLcQ3prk7jSmI
g6HjsWjKxzyq8fK9J7+L0J2NsFu5iGo5IfSpcMQYcNyz2D6mBeBYp+oD8yoOZ0la
rmFofETnUiZgbqdmS3G2M6oBDtfOZHXnG4juxhRKeMCwS21/bTpdM958IeIPj50J
yzPJ5PVvzt63x6AtZq+O58hORvWyTX9V54/doK3gyGDm0KrdBp/Vp1AfU75fLI02
+Ll4KEIxE6zZ/feX7iIaHdAA6dWzO5Bl9xC2e718J51Wqk2Gr5Tqu9wLpapuO13E
WTBGCzNKuiBw9jxGDJv1BFYM3+KiQk7/wqa0x60TvbKglfpNdMSd692KoFBOoWDa
IeyHN8zq+/ZmVoreL/eG77aZ1cIv82qVj4tX2Z4eGupjKRepSrb2CLDsYdpLdm1t
FAsGTol9sfvkV4jcE0icD06b19AkcXO7qfQlj0mFDelmSAX42iuydScmr2pI8Gt5
yUxUFIx+RhtZC5e+jUlOBSna3GpCfiZYhwQ6c/HVuPlBwzzDLx9JA1V8H1/VAEu1
k19zYIVX5mS4ZLeLNnYc67w63ve3D4UCwLvhofuauSc79wZnz+l+9mKxJe8gcmZo
4E7zBuhZzm2hSIegyl91NT5ylR7azRMnWQm/yBhl6LaJ4fMTBCfwodRLeSC4OYwL
IbXwfljOI7QQj4p9C50XRkYEZIzXO9kn3qHtOmpd1g5zEKkaST93ONHVh+M+wu+c
/Vo9vfrC9G5uJNdFgi7+I2992tQhNU7xCO1PYq/pv1KC0Ssu+pGqKeS40DOVGRf2
7iZqMWo5AHZ84Q2h/XJFLo0ETlQUuxuYQYglfxmes1YYnlNGlndeO5OLrAFtftsK
qqN5/wT+ZCwcSTWB5MWQYYWaUt3CEVGFpORFb0/i4gxRk2k22eP620cw1FF3jt0T
0KTshESDy18nUcnX/Mm/+MVREoXvAz5bIa1qKUl8/AG6eKZk3DBaorxK7i49BuMH
/qnTmUFFE8BiiAKr6dxZkrRZMDgJvhqMba2w8g22hQ0Hp26HLlxjgXOmsHbB7ijY
qtLyV4kvZIRYX+tKCNW+VQfcHWU2EUFJfIjcNKH2n1wCCnSgbp8qyBN2rH2eIx0w
s+wI26ZdEnstyXvtKr1mZSzLpPf2FBSqM5VuIw2xll6aWoypDd+zUAHbthHxW3lN
wpdy2qhsjAveAK0lFDy9WlcZwVDvCWAvMFCsttfM4XoOfybitjSqkaxmuAf73WsE
wynRPbt4wAdUw95g8Z/gASjLA4IcGaHiQAtWKpwVGDnEK5qZDxQMapQh+pKqAeYO
5hmTdEydg0jOt4xqlfy4z6N/ExesBq0P1lQV8m7Sfc/XlKFbzKU4F7JePUSpIo5i
vUnREQV6iC4u3WKHRenC6fHOpCttEFcolqTmqCavrvlgDlWkK2mYgRYXtaPqtFUj
S3dIjXrTD3lXmLwpDfszMTtp84pLLtyMnK/noiZbRcJHqdId+nutn6rEWMqzYu76
xUDa7QO/RpGdKedrulAm3DRpnxvuQ0a+VhVon7dSkNynYrTtpoTwPTghuZhY06bs
P+rvVrVip46wVwqc+5GiUO+qBJ7EBW7ntoDXESBSgMFq6Y/yjcycP52yFB2qKrVu
SoVpoEVm7U26eo5e5QSBHcckj2bwA3BnaibOMJVERlzbNOgPMN4zhErxaPsPgYSO
w/bPVggdEkZv+W7bDMm6T+2OVtFFgvT8lgf/RpFFuDOh6CB7hO/OZW7wnGpL/QEP
fxbyC57owb92EShomsR+gAuwIEmSI3g3kY+s91MfSLVltKuggQgjLXoXPiy21glw
UXDUIE0LHARFoNa4GA+HLmkNYRzA806CgsbW1KfRdGuDMdjxpyUU84zxfcDVvsWy
cxSFQKbU5l5IIwqLJxDQt+TdB/+xtH6knNxsyI4jYo2y+fT7EfxTqwEYsz/M97KV
3IOryCHaTNMepk+y4SndxbHZqRtMwF8Mqt2Xj+3sZPjYrnmPVFysx8WTvnIYZ95u
jxNAjOHDE9F7CHJADeQsHeefB1URAodJYJOAgltVnADt47nlAMEzBTEuj/a6jDmY
xKA5HoHMRoIOkssuPrtIXU551DBCrQTrRd5f13ocFO6EKQeS+AMqPpYAfid0Sv77
tVHEeIbI3ayy4G17rbE6w9MttnXtxPoasdt1CzQ0J2sHeXbkrm/Fo1YeRZP4sXXQ
mD9D/4t+4XGMK4QDjV5992NBUcPXCRr9fJlFp0ziU0RJUbpURPSL9i7eOpQ4iFOn
Fv4lo/3Nbr8c4PbwGrmA9c0iD6RFcN63jfxeJ15EMx2AVM/7RQbe/VySHPLKB1c2
hTUKmTjSaiX39BWr/TpYJ5GP5OyNmTxnoSsygGuEPt/AvNG2q0WxFw6itYB2/Kr5
Ud2+fXSgRFlom0WCrMf9rRHHO4zAQsnyAFIHIANXPsZlJP3fBCJU+EGnCR1uSIzs
s3ccM0WbGR3x16VHOae22Lq2vgU7CtIJ1jPV7gJtndWCAFxH7V5UhFIT9b2O4AKD
WYz9LjLG5goo0NUS36dBI9q3CNHC8b5sXXvKRyeeNofiojkWkwEFZ0rbe40dPBOC
s1GM8bYZ8Mcqlf3qQMHSAoGgI6JlOaqU/Y4ENPQhBOCazbsowpaBcUJ7ovIu6px8
pen63wLN1vh/L9HGC2czN+jEra7a8MRVInZ37p88rN26Ib3EI6LO4qtREa2DSm7k
gNzbFHUH+HcdpVxCVQMPa/xSC+Agxt5+26Z6dpyEt/2WZvH1mzyk0Mwnzu0sX5gY
3aeJSf8rh3GJx+0qipzBx+dXXeeMRFlylFDMnIGV+aBBTOjzLRHX2R6Nff6lxXEK
dmQb7Sy9CidNqjvM+MVz9gviUsctKT700642NpYk2XGsZBsqZBXMtJ6cPUGgfV+n
GeVpSoqqfkwxbP/IwiHM4dXI/Ma9SDtl1BslAQM2erdhzJGlF0H7d+EMFeqBTj0a
3njZtJtw2TvZdg5qpOMrpdmUSeiiO9i/pc28VJO+WQi5N2QdsbVX8rHqQebH3oPS
Wakx7qOtpCsLDcGMzMwMsn/wP2lhAijIxZqgsa7+sGyCWTeTd3HbwM1/mnkQ3CkM
pU7k6vWmBl1VZ7hbwWX7Om0O+3XwI83giVHHLqRQTXioPb091t6iimjvbUfXI7+I
pXyyI5a+C5bPVios15DXKsVKjnPMa2wpzFxXFMEzPAPFSpOrJMf1NZHc94fw1l2Y
i/dLvfGj+t6phr3v5H2RHen5w8z1oPk5ZLzupiDqyIuZW9MLwjvEW5IOtVfaKTis
ID3zDExU4/tlCXsAWnXvuGNhLLWcyRYLHsgZymx44vjPAJ+drRcuDnU5G17b31jz
QnI7PRmCRjOERbRe402mIpYIr5EUzPdCRfFLE6kbHS+7Tmjf0sagB7bfAcC34NHr
/lL0tKdn775kfutZ7YfOA07EjtZAKbtCeSN0rfOYUaQMfeFPpFLjpvKlb5FnSdh3
K3OmWoLY49jzq1hdBMl0vLfv6UUaDxT59qiKqz8KT3en97hTdPwKSzH3CZi9+LO6
CAbSGv6XgtmLHC1sVcYLPGEHIbz0mpMVw+KkNlKanTXj3nNVANXQZERJFqIM80aR
DuLfqMhy1mSC/77GPhb72/EOXB1VgoTUD78etBfnOksChIZsCcRq0Xq+bUg3EqnC
N3a81Xr9QSrTkEBvKoxImoHiRW2MXqlc7TIf884Cw9aliZ12lFnf5li7lac2FKcZ
LY8y83fxGO7lfJ5ZJoFoSrheMQH2h/SoK+54inrAmRKXmM4SEEcZZq719qJ8CwBL
hPv5SRgv0egORkGfIbdga7F+7L5LkLXYwEOF2PS1cRjSj9ehey4ucYF6evgglNuk
9AmTa2VKmXjtah3yrP32csr8H87ner/ovYhVXkVZNl7ofZ9XuqR8p+QqOwgIeVeX
NfhMX+3U8EW7wG9Z3ke9ohzXeuEMHWum37TK3sw7Fd/3/pPL5r1Cv6RAno8ygNU5
T+A7Zc672+gQLOMeCLpwHUgNlO+aG27R/sHz7LtyGjKddkpSmOQuLeb/jzo/pFF8
xE0LP+akEfZRVKaZae+GQrvMlVu9tggHf3Ls6oqoyF51WrSoP4qjiXt9srRQ+wTt
h/j2ABaTFSEWwZw8O/yLm6GOzYnkJtCUCz23FQmI0NT7e7WM9+10qREpWCwLxaq4
CmqQZVwoXyP54c/9x8EmtTu2kjao+XaMI/cDfqJZ3wEWyazlUeAN9RWUGhpSutfD
J05SoAbj+p3vcN0cttzel3zeZDFA5jc8lR5WhOvufSrgVD41ulnl6giuHQZHr9mZ
GGYiP3t71hoQ6cnI1qjMYAPk13eWDD+jpHmsEmG0l/JUm2/U5bs++7vIZzN1Eec/
jiRVw9iZNU52nVdoOk3c268yP4hCRr/sEJnPhD5q1B4ekVzankeoFFPCS3OLlIwc
9UEe1kTlzJJ4kOFy61Y6xVGWBvzPjqlwfKY1wyOP5ZDUBuyhpf29tRQxckXnPbq8
4OEhJbFHc+Yd2ZV5NmJESS68ZYoSu2BN6M1SbTqH8axg+djmgEJcuY6KHpyEDSjY
6NFnosP6vukenanXofo0a5Gs5KKjKDJA162+tv/aU4haGLCyiKo375m4qpypyvju
AfAEhSZCZIBwCTJCf1O5a1NHGqQ8eflJOKK2snamj8ehGXmbuGYRENRIRq900NMW
44eUjz3IX93yzYywJ+jVyzCDV4RMnVtfjcduxTJXUd/9V0hKehTitnWq/0BKImrd
PtdlLkttPZn8IGWwmYYxirdJrR7v5WnM2yDjjxB5/j/u5G7KEYaM1nIEoMb3cRgR
MWtupC7iUXM2BoO7rSzfis2oayVZ5niK9aiXy3liw+epCLDxG3GoFA8gx+sNhmlU
ZQeCCEE/7PdXWApzaWwb2hSptdKpKrp+HDPLDQhRE2luc8MGtqVzXGyeNRWw2o7Q
Ha/9s9iJV35f14n8Ylw+fW/swAgTeOJcjPHyjudRv4lGGVLoltRxCPDioQGxtmG1
2pP72ohcYKMGKzlONclN72Cs9YmwiJt0JYdaVEOg4ZA1fkT2bHBpRROOvYLg2V27
3kWSSQMxdF7HeCvjinFW9OBnuFWGkGJbMk5m+g1r+AeasngYf/hcq7yeiEmexsSS
nHXsGkUulTVFsVclMpjIgTRXhFWQozlXhPv8/ukewSXzR1W1pT8kM8j3KI5rnUIt
d+6iQ8eCgxmlLtIy01VP8sEwiuvDnaeqICtPRTv9ZlS9t4baGynQjs/xvn4uQmQt
IHJI+gIUDVV3/iYX1eAXfHx4CQCLR4Lc7BlU0zFd2jifaoZSNWkp3jHBMvvGc0L1
MGdGaonJo0hGOSRTJyyAtA/oVi5x4OpHNjXZR2Rtau9rNp82GMNHlOMGiblWAkI0
Ju8+sGZdE0CksyWO4cLiy8jeE8KuDxG86nepGmCwyDZvKSUOY5NjOC1uovWKT9IB
BPjt7dx9EVtM/LEo6zz/vLsyJuiwip+PCeTm+ZUTS77/tWh1efs9nT0rQoGj9rXe
aR3JdINVqu1BnoH+xaM2NrXZAPJhXUDXHDn357eagf7cCOcjh2UcTT7uxjk4+dm5
6NGbGnKSFGmS9o206yXgDiaoAU7/ugyZCW5vVRmPIHLHZwUGMRuVcn3Sr15jjOaH
tNs+L+WaWtu7YbnsvLuthMG0uinG0AjwsUtzp1fJ4+dRn33NFXGDVAeOXAOZPqfR
F2KmBCNeBVI/WevRGodu8wWfXamBg3W1CCqanwGp+ne3sWQk+c9N59S1mGzOAxcA
NDWmdvTty2trdK+UmBhKwSGn7olwE0L2Dq3w9rvzO7nVin3GhqNwIiUZq/cdRXYj
hPLX/nn9+ivbYjQkJFZHVqxGNSDJO/ohBMj2rCLxx23BdleDJlc6h5LmTWGxvhLG
ghHl7JuXcOxw0HPGj8dcIg==
`protect END_PROTECTED
