`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CIgtzc/6guqTXduVFYQ3Q6vWjO4zSfS2lAK8a6TC0Y+9TGTRSwULPBRRE5MH+9kv
DQ2+o6PSXySLxutRpJWgKcBa3dNzvMoA0bFBJAOTufrY6cIPEWkfUmV2NDDohr19
6USg6Z7118S+Tsvt9SWnv/iRmk0S+MaWHIOKa3EL0ZyA8ZO6kiELg2Pq1JxRIBCj
W3pn0hIXjuyh99/u4haR75s3Ce/RSdT3kU2a0wqTTp6dVbRgXQnT/cm52MiGdwbl
Y6lTNrAn8qyh1botWObdnmFg6d4EucK0RTxSN0ackLb4qXyHuvkKkyhvoww5hfiL
zcC+lPAIrT1QWqGBHG7v4fLRqihk1StIHXB20xV6AecLiQkDbU85YkC2ObS5EE+k
`protect END_PROTECTED
