`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
evzxfb7a/nz+Bm53AfKbRbnEPb8IP5KjeI0B2m3XZWOBYCKTNxBCSBp7x1bP/2pT
MPLoydwhTbZBUN/hgCHyQ6lGGq24G/1ZiIL3o+ifnROIoss8As8/ABa2BJmqiHNc
Fa62cy0CmQ9rkHOK/uhBYH195pfXXflKero5y6AgCB94QzXG6wul3fYE9JS3Ibe5
fGwUlELdp/wV2fjLhzV/KT3+tZPcgQu981pRFW8AiB/uiAnDaAgRUdzbZR+ABnMs
AWfKhRj/ikuv0ioAZvr3fQbhYZcWBb9K6pPYiMCCQCkdgN1nZZTytEwe4qQVfycL
HKzoEL0OCQuXLKP7kH407kn5TBrnrpt4VfyADvZm4haoV6N6yfctx/MWkx+JbTWa
vG84FgEdpKtybrriIi1PtA78gPPGUUOOBqL5/Yj4oxf+WIH8GN4m1kJzJQD/iHiU
QsMG2N+DzdU5OB1IVETZ7uC6/JtPxZic/GqdT5XOZMQ0PebqiaJ/RLl3uGKsJ7b+
g2JC/qoGcMqNb2Tmzq4ISBKaaorpMlc3SvZUeck/5U07I1+x+uuFMwPkKVQC8f1C
TvYS9SiP1sdIq0PWyN5vE++i5u5lqhOzYLmmspn42Gn9c331tZYHS7tz/DBIz9dS
EYJDf9IFTQo8FFyFDTI2gcT1Kmii+nJ5eOQR5Yf3Y08+iwZGty73uIF/ghlJ4ur5
x7mTd3eKfFomXnl4fvkcl5pwdxueWlf5bR6K2xNiDKoLMAJIU2zm5JrcgU8Kcgbm
6s0GwCDbnG5Cp1nE/ZoS6k2Ph+YFBsO18FDCjwDaVoZcLEwd/ge/TdGYlIT/i4vX
WOWP1KzPuPRjdB1pPSZqkOfxtcyCXdG0oTop8d3jisb8uET6eQVIHBjGcdfHgLV4
hXILZ97NfplBZXIxXuUlIz0CufxIqjtVsdZ4UJLJZZzfYwUwtquFgyo9J0xpxkL3
TEDECu7KN3DdzfCMy9g9IBILvu2rUkPCKIKOwzPm5jWoUMLfs/vsrB+JOf/8kSyl
kW4jPThl6IqV7Qd4YXJE2lLFjcgbJDTIUSbx+380Ued124Fvm4YbP8Fnf9d/+YXr
UqpFtdANZRtUH+9d6Yb633ju+bQ+fq0I/irf8DgqSg7BYRgKdYVGgRcsr0YG75ol
rOH25Rp3lKvuE9G1RF4RIpgZkpSzpwcvWbSYNYAgQQ6EQxwVmefBK3DblHYkO2Fe
dQh6w04mrotkLe1pYxEHvpNsv7LGgqN807ezIh65WGSh/kQnuyGZQOdG3qZwJZT5
rYMS4frI7R2oZ19bqaW8qcY6vxLIBZbWFVsaGFmgomlhTC9R6fahjQztLYjxXTz3
ea/CZ5TpPvwyd2/mBIuHvqniJwmqA5c/1/44n+Qs4e0iZkIV5RA4+A4S7lAPLbQa
SDDnAF4OmP+xiEXAhrFnOU9xwZhJwxOj6K7bIaJ7XkQZMSrL6ZAqzHT4rXq4swZ+
lU6fLEHnJyNKcQBrCoMM/AFOjAOQJyjIZpnvp3zGmiPBsEfyX39r7O8JIiQN+tX5
FBLINhv/JXfFL6q5MDe0gAOk194yABK9dHCNqvTNHlG+GCOyf/S4cEVe1D30VyfN
PmpIY/sB9RiR6OUwwRiG4MwTjz5EwRqeHD/xlvGHizgHnzu8iD/OCmbEUX0gCY4K
DEoEcaHqUreEKzCdw0WWoo/Fjgv2L4haxZwhRDwk3QaBBP6chcoevIDRx/bg6aiH
A+dCUU49L+KjZYHSu+2KCp0H/a4sQC9QUjxvf+45ZfE+Y7CPWt2klbAdim2K6Wrd
KC9wRZ0+vTx1UcWeVv+c4S4astpEDNuqoO/jeRPNweRroU3cV42w7XsARukFKIDL
zMzlBk8zvQG5DZ3OHyS7CL81jNk+3nGUyB8Ek3+7cAAaWF32YDfPVuQ2YMoK+m15
EC9dhupPaS+EcQTAZ5suxhGAePMqVLr9N1UbRyi3e9JXBNj9T4vg/ymbJIrwrzyP
ux6SCACUtzhr4iniFr0vtta0rZdqo4loah7MZNSYgiFzszqxvAAwyhtveRMJtVEG
HBVHoN1s1BxXfgtNj5BALDqiloxbMjyrD0Q4E4DahyUWdmzBKDZOtL1Vqh3/+2Sa
uPDZVy5Ew9NmtMRO4SIj8yd+sIb9sYeGMuBmYnPtk7JBN5BMHjtSLgRqLqBkAPx5
qKKakstOCCwmHjjT6eH3GjwFhtTd7VuYfSMisof6pDx/0/c4ylcJwaJd4t2OEnSx
4QlRXvmoBHeaFXmB9j65VqAl7oPo85UTNEM2HC5LrNjznMoG10AjZ9aBoGFI9UNi
jzSl5CHY13ArFBy53pLmqgkKVEcGTvlnMGmRtIoe4892zIzdOsnF2apgwHdGwP/6
h/h4DZPmwC/1kYqIjEQhOXRcS94fTJ/bNhHA9RdLosTDwflz5MRzyi2srhiHM8rl
H6UCAU5PlNr3VqF5ZimhTg8nuEsHEIsezGhmhPRvcSuUZmNu94FZis1ibrUfQzPX
rdYvr+8WS3v3XSWEZL18jrDs0Sn9ZC2yvqqkbSxgWS/iYV0gl1YcY5X5G3umWvu8
AelsKBh8hG6Llvmbhr9reDJWvlICZVnVaIVgslK6MNoEB9YWhA91iHbjDH3V2ciI
R5/mgQ90S/Osu6zvCnVMQcHsVIYSpt/aUs1Ep7uUBVlnfyAYpt85JOsuMhcrJXJ6
jtW5Xa5jUeMO6FIMj9i48gjBS8L9tYloCKgI2r+v5r/9tFfA4F9uBhFRTCpgOydI
dU0p0EP3eFhdt/E83irg7/9uHGE/xdhZ0AODx4Ibkst1lK2hxrtA1sIaA3lNKi4N
jSpzIp8fSLUjm5glC5v95BPl8XkTAps3CbOMIk2XXjzbaC+iwb+TBzZ+k9e9J30k
EL72TQYmL2kcZIw9nMjKm4/yvtNOFmlVtCVwAd61qabREY9ao+MDYQo2w7gMxizG
1IGyh42kifFM6qVk4C/eksx451bH9SH7rqb+aqbAYtbjs97zhIcYeMG5+mGGmRCA
0eQe2CZi1ww7py0ezFGVb0riVwB/azVTRPEGUO/9xqEDRe2VypNudhvfb7warMlP
/tx0bfK0JRs48383dsYTZouCbeQ8OmDZucre1pWGDBL6cFikuQdRF3uUUoNj7MGT
UIdUw9jGcpAk2EeJVtoiA6MfaVUN0hghxHVjoHjSXNQketqpYbtdH2s00nGisA9w
8uYvS+AMuk6w+wi+b/yjjM+jPoh6dDKOCtTnjsnfrinlVLsrpDs72K5W2RxkkyVr
GuCA8JaxFOSm1c1zS3W4Dc1QhS3a2v7Q/LohP1hk8fUliRKHqkrjjjqY6yMyXUW9
kh3DuTrsgLd+DDv/lmHYyxJ2BUWPorKzbXTPvfUbKro2bO0f6+HVkuydsM1OR1CG
/fHPPeKIYBMvPWhTdHPEaC70lGy0sV52KvO5g5NSYmPv/SB9Uqn0CmzBzddzXnmI
iXes/qqhvXE3Hfp83WEvyHWmTcuVXL56WX5TyK6pFwQklRubrV/uTjJAYfvOdQKK
jniyutbXeBztFA3BXHTDxystnTbg3wtzQvB3A6ZcsjfihlpRynckh0CTH25Tw38W
BT176tBD/mEpFJEZFcZ1Pciheda7CDfQ8Rl4SPdNcvcxYuv89k1oXGUoOUKVKM/n
jmnkyARiYtKMwmuDk247Aek9cW2KYSFsavSQGJy4lIiE/6HUUxV1aQzR5eztvMbX
hWrjcqiLirqaLBIJlz9xUbgTnmvc8EfBALVNXVqF10XjO9EOjD7WNgOOtLF5WFqA
DaR2asuBKsG+e+6WpVPNfVlTT5RroJ+We/liFmSbrYEz5/nkMB6melj2BV8cl3Zr
BXkIRYY98JQfmOCa1G2hbaQipNWn6TiKqXQnwJln1/RA2CNzirlPsNz683OR9Z0i
NB0eYITxmHQrBMnoknbYpveP3tYeMzZb9/ovsQA3Q6wahKaDdGSyLTY3hszLyoM/
VwCCjP+ncbkdeVCPZ1xCEs1bHPv2Rd43lYhS4X0oUqMm/q6y3tzyhOfVNGjcIigK
18wX1F2zTzDZX8vIj+6iJdi1gLwfwrhkT4IRQR7z8I0Y9gf7Y1oi/RsXCU5zW3zG
pWOpcaW480EgcjTmVGB/DYDpasODSdGYCLYR/bLriuGGRIfX+hauOKFCU4bNTtD4
RQtE8xUaj0fMMsfMgkniI9XBNzbdCer5yV3mkyuptIrxa44u8D5d7orP1zM1dyDB
YO+yc4YuDWvE1VeCdfb1p1a6YRzwvf43yZl2ykG1+7ECCql+SvyGX85afeJjjZDf
Immm3WSMmSqsk2QfwzatkQgFNwmQ9APXlNXDJuX8U0ebBwCDLjbg5+C8YC4S2Xsc
QDAnerQ+oWFNXPfNg8kHl/PSxGIPfGF6u/y+kM6SWvwE3Fvtrw0A07mmVBb9rH6q
5y2VuMoWlSvbX0ZWkuLlqcWJGZ/butoqLFfHI0hFfNmFcZNZiD05gGjW4JPdU1bH
cAfllVFg5Kn1LDC7hqD5FrkaMprJ5tDuGyQcevPZYRW5m3dhxbd0pUlOhjHz/lfq
3c/MOWhPIHtO/VpT5To9OFGZ/1tjqnV9LNRmW3VbK5VPXXo5Bra/SvQllWWFlMah
lrk7i5ANvntUdOjMYaoGHu3pQyWB3BDJFs0PGIFPJDPRrW1UGnSdU7f70j0sEIeY
8IOGEcfV5OI/KQ1+FhABjmOwbrseUXGb79oHT0bWi9W5v9LHQ2fNOYr+r/ZplKke
BKQMPnLbAyS4UHgulxlmKr9aCf0/PJ6+8tRu267TpxTLz5s4PaD98Tkvu80PDgCJ
goyDPtuMJRInkappCSnPxee/3crH0FCcoddlhoyGKwfdO7vKtq55ELHjgtv3UVD/
UOkN6B1c5ePZz1zfe3LW/w+0UYPGM5Kyw1ZHrlNk6Dy3SlJN66T3NnTG5I5HNWro
x9z4cHeQ3U/MMbzcyqq/2VW1lBI/gbRgaGfxO3pCNadTNwIgkBjUv59i/lzGRvyX
A61APPPk/PcFKTyzyqjR1KGzQoLFhKUDZxb4YoTkXnTy+IcRdUg2l7nY7ZDSJGlC
+sQI8RuREO95N3fQbxddLR1CL5fYe6ACtUMFtQ+0Qur+F/7ylUWnvpq/eamTfGo6
dyR+Qx/1zAL8SnzMWvgHxahcj7DKJgerhCs/yFHISjr9OmDIbkscWrG4c71aH5CL
rF4ysIhkE0GfC3VLpWTuRcrM3LfgXd2GvmNoCyHmDwSVw1eQvgAZzhi/NdEBf1Ql
N1umFbBcrKly4704xoOLR8QegEEjmVjh1xtgJ7calkKokxcrs7zSzoIipt+VkK2W
DxoJ87KlmmvqvKYL3m3EDZYKp7PYLHbFg6ak/rJkKTtlna7BkC72wPpW0IhI0+4R
vUW5PI2mXu3RDTmACjPgdeWfGHqJMF1M3oikDoWMxKi/lhNaitNts+NZjDqjm0No
XdjtvYFUjKvhVCWvHibf3vLp8FImJC/2tBBTsXhbaW4BNHTolNqHay5zAEE4bi3L
458ojioIfsktcKK0Di2XYUx0lX1gqiuyhuNLTvFIEjyNsi5w3nvS/LPV0ZKv+Evj
1ahIVXTO9/Y8pxCYpZ9OHQuGKA9z0foaTNLkLJedjV+HOpRVSnEPXfT1SZ4pRab9
IJchmS2DAG+0ftFIn1lHvi8PQR4VRPqm2beIozuyxmLjKUppsvz4MeLb+nGw9eIL
KKbX2DqoIgvzoVC8m11zPaGOa9h0Y9QjHLEAaSAS6EsL2IJNbtBDM0i7gjHxzcL6
7y29tjuwBhc7wSkuhb3Qp4QU74VCuRKrFPT1fUKgxiBeXRaU52fbppkXRZkE0Eee
HBQYR7hWV4j+XtMkyyI3ErF8sc72VUQIbYewlKejuETkPf6tpqUNcbn70MVUgmxR
MuIz7+2WTUOV0pkC+DxtStJai5GM6s9YnqDO3CvV49uKd1ZA60Q1dAaaM3+fsNjt
JzK58x3hBeENTufSIp8+o4F5D4dQYSZjJPRC4nDJkJsdedinAf84gq1IkzttBkTZ
A93wQ6EVy4iwx3W6tlVok0NUcHOSPKxzqeuPu65ccbRi1zRLm+jSoctHEtcDN8is
vUdKrR+BV4GXwZvDpe59CYFgCrxZrb+fpMm4o316Hms8Am39TqEOgzNWPXdcoVF+
qb5SnigQKgQ/BvLq3EslDdzTGfh6PtgwNiansJAScvw1Qwwfw+2lVv7y6UCqLuhH
CdRavHrZb5s24YnPskX7rzy5k9TRdfrMHvWEzB6j6AGW04C0UDQCvgFYJqQ/y+Yr
F2hwCWxL/itwvaTazWZHYdCmz9hBKZP0KHGKYpa+Vyh2mEo5zQooa/jEllZEygHZ
IcxCvLZI8gqwLHK3kVRUnzPVAs/2ViYkQVed8NH5/kQsnB/6qSSOFVCz/VktUDwC
L7R2Rv9tZpmSofHqcPgdp5LcYLxs83WwAReDBrC72K+vUsmrin9xbabuV5JffWby
t1f0eCxjwR7//OhzfYHyTcL5IF33Uo1lxZYjaMGwsELkLaWnXki4xAbCohzofECG
KQEMK+fysNMsxYJ+lQiXIhQfwpwbsi9EpwhKPlJ/zyv6sdz8FOz57TVyLnpVS7+0
WxkDuYCC+N8HweB4OZVRS7h+Y0AlLACZDPGp/RdFWNZ3fLtgNrGlJnD5S5tTaDy6
ml+fpQsx1s1uSPQpbJTrtjhUpX9gEvdM0ZIktospZlk03BIXTJx5dV+n86CQTdhR
qwgW0LrhQkpzqmLVAoAO/IY6USTTa/4UUbsAxUkvJA+YSqRbRpNIawu3l1L79bT9
Pn6wcat0PRlgEC72fsD2HYQNxjZ+5Kg6ZLi6iBujQz9h4XOR6OOGpNqcFmr9TiUz
KhUfnc/iu8LQ4jOwVI+sNhU/g6yktyMFEVfOaDcB+QB4Ql/ZhY7y70lxWVZdcjs1
9M6i11Izvafi9omnMKyEPj/TNRilnIKn/Fr5rKWNogY7zqhD5a/B7HZyITRLiu6t
LD3jsQWkh+cXhnocMCDKc1a4S6zjm0J3/vFNPhPx/6sa/fXUhk5Tk9H0/1kM7Uy9
RrUKnSBJLFBjLsxBVj5P/kZm8V9O9M9NDQpX8XsDCz5maynsQoKzjel4zot5qpG2
FicYlINXfh85CP4YLg71QqjImi/CT4iEOHnb7W0g+BFhTT0T/3pI8cy0BRzWDTZh
Ov2dWd1eFSC4CCNlDXDpU5BoVdUcd/yH+EMxnd0Jbw271w1565wfbkG6xJ//6bEh
iJIxaC/oCohQ/LEIAtzemWveJgWKbUn5bfRo9NTkXzRnK4d2GzMoj4bAW6jjrOmK
LHb0Et0Bpv7aTyN6DKkwHHxDbKj5pCj/RjV6wpszzUXK5qztRKEceYIdGQLA/VwZ
uBndQCf7f8dPhocT1zJD/Ys4HLNVCFJdZqHR4awkCY/s56JM7kEqeQwdudUGMCvU
iuCO77hPLeoLu2sCyRwxvFPSiAOuf8FPNFttjNzOte8FYRYhju88QvRtzcEyrbZI
ecL4I4uftyHbpHD1unDSIsQ2OTstU+XBUEoBkT6SQNdN+Px8KHU8KI4gH+ZQ6cH/
6PymUewIpVAU6a+th4QVyQWukgdtdMGAezmsKc11sI1Yz62buATWf0hznRXKAbXW
W98RGRIFaIVBwCWkCblZaMq8KHo5qxckeGhecGtwaNxRLIHDXm55OoYyxs2cA8ma
5PE1mVyDf9SQwSBaWgxZRWCsFQgCUBgbYPAUAZM2Hgaw/5lb/fqVn29HgDHrmh7F
BLOcKKeBm3z4G3BSRBVBbVOdingpFJWNf0AmOdwaW/7BYouc9vqndD4kCKXUYyrb
iu+8inPvoKzbYdEkv+zyE24Hdj5cqe07Hgrc7CKCHcbcAG4ReN7S95AFHdY6cVXT
GTbcx3PtjnWEad+TaUBJeWND8GgvpPkYMCX7ewhbiocWiGHlKuSV2YxoZkgeX+bo
jAkHtQ3KA7wtXaH55r3CqlW6pkVHVpgIeDVCB/7yO8bM01DPQF17t/Gu/NmxT8np
UYMX8mhgHgc0qbh8uvZRvCgGlm3KY5HZ4BH4QDVMbvc/MmlQOfucWV4tO7gFmBqa
xcmxJd9M4BmHmbdtvUuzFmdwkP7YtwjqYHyIrp1q2h4zzWQ60QuggPaMhGdZtB4m
zpE4e2MsGscVnHdFd9+qXbZvDj76T1G1TlmS/8HuyCtTPstmoGMRbDw3Hu+AwYRm
y0EsvJi9gPp8AXuoc6tBRdP1/PviDglCuXtNyd7tAX1c1kWzb4ic4/4Ay+7OZoLi
D3ulQP3MiEwnw3jLjTr7L5wB+/deGEzG9yRfZEj5tc0BfpzEYha3RcIgja70pcT8
MZnKw6T/VonZYA5P64A6jjHD4kAqEXVar2AXTrDl7p1Y5xxcZBeNqHiw/gzn5n1s
1COOJP8AM8OUbH15midUm4sE7Xp/es0LYl+ubkvFJa+w5eEvzwZ4JfO3HXKGPfqX
+37oXhYGgKzyET4h7jXmRXHlMzLEXC2/+lXRM3Gje3T84UneJOdxetiOZWMbX3+6
i1+G1liqDnIi0iEWeKemzaTlrYvg+R0KaTPTNskWY/M4HpKWc+3xzajcnL793zQ3
r1VdFYQKuMo0bvHYUEWR/EObQraHp6TqnOwdLdFa9ctXO+5m1+8KcgEYpTIqtxgQ
J1ohe7POung61MRgaMVPrEp2k4etfbOn+Bn9Q2johZlwZv+U47mbu8qsSKiCLXXm
mYMG9G8tj1kyKKB0UEZFgLvm3xVqyDciOubFIoe83oyi8AQJBCllhqsmuN9V9r71
FYjv+Z/eHs4N9PEYe6BcRMiUxj/Qg+noXHJtnpLsfG+rZTTVf5WQ4i6O5uX354Za
rNr0uhvBAGwmwfCiAo5jIVDVaA0kzxN0j9P+CyHbK3PGHXs3sgDXt2QrdUdC3plR
BYn0A1/8YX7UmI2AzH8NsSRnBvISYDYGXXoVZNTBxE23iZW+UVYx7iCTVQwAXiRK
5RjVUGOdom4VysRsOuaILdJ1HhrachWU3k4K8oWMKLY/c1o6dA0zwzPjyNG7Oc63
9flWRRKh0ti7VJFkUdjK8vG0iHOphKx+Kd++gdgdshuftft/wmZ4rF/tTnsR4aob
yiF6uaqfGzssLNwXp34Rwcj/k+JQ1JmlsD9vccx3h2bm4Ttsw6p0BrPySuy26SpU
EzFN2toPKIAAhKLDxx56YMRHfhrxlObv7zk0BbOq3Y9v3vnceKuSoKVQ9C4VXHya
tTIhdB3H7FZfY45DpNyIdufM80Mt1evMb1k738U49KV45WZLQMMfhd/zdQKx2v7/
eSLj0F7iwPX5Fmf1PeWhPLlNweFN6aRlgW42z6ORNikxPlU2QiNn09vkg/heHtMr
IoL1VegKmDiU0P3oNPAkzX4OD9bA6fHWNw1jVCNnVWnl4fzP8LGw0vaSdZS/2A+7
1jEMabBTP/cgXAKeHqzQs8GKhEJ1RYHtiE6p+8aqf299eh57+GqvuzaQSJfSIQTS
05IYBlnph7vSwfVPit6Fiy0vsBGiXL/vB1shq/ORM8UZO8xJ7c8e+rdRiJnsEE0L
KUzjq1vMYQBGf9VSeddrY/cjc0Jd7rFAbR/aNfvwi3YLGARFuuTZQXoD7eWn6ITg
mEDhHUMQJGqobHlVa4U/yDRQix83UIeya1AdRK/hAUFvqwfr5oQmzNZzqtHxVpc3
BXiCL3D1jlq0hM98PwJGl8rQVJARo0WKfdpQYLAvZevD326IEak25DdrtdLN+UKS
YkIjW9LEoQ3IStr+YFRRHdU/pwW38WZ9fO/fQhDncnZLvB3N+/KKLeSfE264JMye
wEYT5B9fyw90xAbGGt/pUydsDT/b6R6161lnCsIlSnUKdL63wu46DL5V4r/azcSV
KDnA/DhDcutosjkKs+n45QM3NJegS24jWAdKjbsf1O0+6Z3e8jic/xyZ64sf1sKc
8mJBj/RTwvZVDusfwFRj+H4QbYgwtgKdMXQ5IHJeDCSuEPbSxQ90eXxbywPb8tFX
ISSpYej6XsHTkQbsvaj95OwZu2cBLUiGwuRn+2JXcLSWL5SYGkTDaw3O1SQr8biu
4mmET6cuFBaAL9pROgWnEBUS+/E9m1rc+VBFVEKCgiHmzD/+CR3IQHHa6tO7dzW7
3kyd+Sf6uM/Jid+2M0dhLXdMMr9kMmIv4FRgvXEmL9/ntzEEpKAQT38SxpCGQQrP
RNzdLbIdEN0xVc6XfzmjvdRQd7HgUA7nrR9ePlAM2N32+5GE7+xe0k3TLVOB1t2P
yWWhOLRdkg9IxYxlUipNL50RP/M/pE5JbqPllO35XUwovA3sYxerDwnggc1rzLwh
yWlUmBTdgGVGngZJ8apS2vdS711z7N9CZ/9VGSPJVRiiC0jaRtqVhgSTJ5uvOwvw
poJIVZ5Ka9oScGl53BT7vSqu0i8jOmcBsxBeUcWlc/gW3B4eLnFnQ21cK2kdkMAV
hbXwD0bOFTWtLmlAb5Pd1ttU9Iq6Syf46U+WgpkbDWS/wvG8V3+CXWw9wauu4geM
Jt0C45Ne9QC+txwNMBeAf2rHI38gfkSVlUHgZuvypnbDkTd2u7b96WdJvq67btaU
3Q1EU8wV4ezX+xqMm35ST5qlq47/fhJaoRpV71d3ZgkmcnY+Ig3Rdg/wJvqxA7oE
5UiFSX6MredVKVw3YCIncnVba3/IDQ3a51xk0cxh/9tWtbduwZj3+3z9oG/KbGRh
Y9BymD/4Qdd50jJ3+lvualJK4fYI38AV+zQ1R0SZ/gS13dJSz4oJyCpevkHNzoHw
Cr8Y/xsmWRxo9HKFDbvfbRVFxWj/SnfWAOqLkSthUbFKwpaM5B4fYwpR+dF1oToy
ewz4urWcGN1gMvMdSxIfb6WNlf2BzVhXpfkKoubOT3C74sZ7Les8FycBdZ5FEtJp
bhvyMenWIqF+j7kdRmW2KbXMGRMlZY+fCT5RFUAcOO8nnlBZX56bJk/lnfAy5ACx
V84vo9Li1q2pz/Vq/qTrEIefkenZhsbWU1KXyGOunx6Ryz5fNWkkKPvkIzdXCePW
D3hjS1JpLhIvbmp7sesCBaQz0iQpcvyLXuQ2RuuLIxA+gBtlUvi8njMKXftRjDr9
ts6s0oBcTFFVORQyH/NJFS0qF+hP2kcmjGkCM/8whVl8c4sMXv+lSWJo4IrU5Weg
YHmvdyQnOlNRhf4o6xSlPPqNnYmbe6woZDfWgUpO9Cr11baPULMLKUiD+Owgzp3B
mPqx4Dr/xy07zt8g0gl16fzi5tDIS1SjTf3yEqVgzW4ZW8l97E2tM6qm1PLGU4/V
BN+FWugCjZxZmWnbOOZFwMWPozEWNBrd4nA3gKGovwLbvNC8BSCSMk1CQWT2RIVa
nPSKggT05bU9ZH1pn/uMFE5UCoK+rj9KWaI30TEB7fp/Wg1HYQ+OHcMNyyRZa40V
HLnRmSHHQ8IvBX9X8n5Vzw8vlFfEaZ0kMKoLFtrm18SFxhjJ8jmzqNFXm4AOVcyO
Nn9s8JqYC6LwU9zzk8Y9C8hU9QDpUIobDCJd0WbqjFur1YuKAXEBNSTEfAWkIz7c
Om9fhDDvChk2ViihGPDDPOX0HYvZcOTkonMPOiAr3lEti9o1JUWXQ3ia13Hr+wA8
bi57lbIEvS6pjLZ82rU2HqT5/VsOIE7pHeNtjsNDm1Q63lJPsQAzkQYeL+Iecg0k
kSYMvzG1dtWHJHssTfIfLZ3Xqp+CFxkyiBMoHE0eEf1QYWjracc33FRFH5Fxn0do
T5se0J1AGDIFdDw4y5wGpvFVNGiFU2N+hyWTQAcaixrYLnlZCxc/9YL+YtLgLxJN
7eVv4JCqnYrm4JB4+daY6bcijPA4+exLtPcUsLe7CB9JCGO/P9HSECDkT2myFpjW
AGaGqdWF1lmKWn/qNiH0y7zh9V3lOzaoepjW2HIEFHYbpDEcvGG8GgKStEKIs5yi
KOPsO5TKKy64CFZ6/A8yb7l7qR3nkUpII+1k0mYrIYyhcC8ODBDCuB8RmQLNbQIL
y1VUvU8C1hlupCXGKmbrbSLtRdI5+CW1doW+9AdF6+MNSX++x8KeDzxgkQHutTkr
Lzj3GW3wZ6KAbYf+4vXMQAPBtGY6ZgJ66UFaoa8OgUMTkU7eLppT5nS5/o7e73P0
MfEZE38RvuuEksPXLKE2UDjQR/Tft3G4zig3zxmZaTpuo7rzdo2gR0v+18bXEO7F
gHUYjSpMocvLvSUOUVAcAuzVAeanMm2fD+z+BsBABi6HHRN388qk7ijTf2uzhnne
8B8zR1vBU4UEoYNU6ufLottVA9NLWO4EOUUQF3gfsen7VisY/fgjNUOpBx5VsHbU
2n4nTnfIU1Bk5xWxlYnQ4eI2QTlVDVUW+/ldx3kQ7bx8wdKiGnN2haq07Liieczn
ixXyUjnog7LdiwaHK/yJ+tZoXNk8FUWH+WBS71rUhaw81+wEh+N4aKPOWgrWRZW/
ykd1EOOIbAGl3payqUPTuNi8Arqxr8Hg5tWMczAvd+dH8eCGAI8Mmwbv2l5cJsfx
RbyOlBsG4khX4gsbr1ga6EeF+KnUEguf+TG/ox6+U7lkiMWpXBbzleG/kGZQ4mGo
6N+epXFzwHhjU8uXx2/9+G3CoVPYMtbkmMhde5EICrx3neB4VJIdPu1GxnLe0+j7
CLvqx6O0NlXfgACA1KgIEkw5D7C8nzcAL0VC8n91yHN/eynpFrVkovBX73QhVutt
+xuOHb4YThltPhIpmklnfoK+lghc67x9pwdWEhabKpwl/tKg9kjMuWFS18GJi5Bv
uXwOm9jOVSPCMB9lbPpqqqxmvDhzAtkVJkC1iYQM1Nojhu2s9E6k1zC18GeieDUG
CigaFaOGvJq70ajUQunDwkaKWME2OxiRt4x0pSYPi+wFL8kbJ0JZTnXwNXbtR509
wIp8mq3E/87QrJJonuqSgI2d7E80KW+bpF+xeEiAfz5noxqiKVZ15fSKSI7mAQFF
mJAT7r75p7TWIuHS/ehPsIvLNAe3lEs2cgoDW24edHxVM6vj1bXA2+Z2/4vZsPT/
79dsvU/Z63wJmULtkN4h2qlXb0jIWWRuuKUe9hiK5x0+Sj+shjAhdhjsAZqnKD8Y
CePxrv7EX4dhSQb4VOG0kiFDnS26ULW5nNtiCHtHvT3MRNTM9ilOthiBWDsnNDwr
1Jfmsspob4kN58i7/zEz+X1aNBFm7IvmJ7E8/g2ff3S3l1gy21NarKnjzPdYb26L
pu07No5J4oghmUclbC6bxoGNabvYZ6d/TAbHqv+ksVErF0odrearSnr3vzLjxCNk
fdpXKPZk7UBcvOU9nWYaeqLvnW0rXcFhh21JDb4omTPZjY31gJJW2rp2tXhiou3n
/SxlUBhgd320wyYGcFYrA4nqiBr68ZU8YGd9P3l8UCJsXsSNRaIRCxwG3q04T5GS
GwMQYHzvGzVta5/VQ72H7BrKPkUi67sYvACnd2Gc4Zk0Jj0iEVIO/jk5+0CkOUJ0
pP8pWTKrdaEQOBiFWbMqwZl0Yh9miqubv1hRDXy8VjeUMdMo5RBUs/6O7qGMJC+o
tio6YqXGcXJj/FEOkptALML3FCm19lBLpszFWvrrvDqxPJCoSV4CjSqtNexUaCQh
3RJfvc5jp/ziTKVPr72YHVJgRq99aCTe3ApZiYXm8h+I9A9Xt5fj2HSNU5n1Ejh7
6QY6dkOLp2M535iPq1IVeWuBhQzRRlwXtIqMJknIrZLcSJ9UAsHa2Df2iiV0CKD4
hiwNU14gZH7wkMKGZ7Pl9fbCeFyCO9KRR3IIGT/7rPPlG0TVcEdwKTcWFqjQoc6t
OpVl8d1cSIBgNSB3SPEcMQaWsL3kjttIP7dh9YGL0UK7ovyND8KGfW2slNSZ+50G
13A8A3CW5SqH7vbOvExG4S5HPsAO1VoCugJzdJQLH6gu8c8kZTpGcpfhlOYwom3h
zS/TKGSol5tvm3JU1ghBy9iFXlczs0211d3zF+QTH39W1Il+nJ0pXVeuFlJoycqC
kG7RVt8bmMkKEKXTYEb2Zbyx/QPuC+SvA9oGiJ/l0pwnhcaW4AV4mvk2O9DnEkj6
Y2wAwFniam5dPw3d9VJhSvApffS+kZnzwmbp0uLkwDP/btE5bXW9r9cbgiUiBYW4
JzGEFZ0d4eayqgjZOHvov6vjteXvzcLNpUVeLCtbTMqpjscqjpn7U6khzmL5XSAo
Rts41raeB7vzPXNaZxDGYSJmiQPWlgAxIduaiEqlZW860QKSgIfhVrSOXXt9L06i
LiAqH2u/WmogucD8ccBsIFOe1QBA1+73H2OUZ7I7SqTDX6ZVobO1ctjcn85g/p7/
3KPfSRriK2HY9VOeCVDLw/rf807uM0L+bZQqFJo3na4oMPKtUeSHfTfdxb7VTDmI
qqJ3F4NHhLtHSIUsvfasqHTT/16KHpyKa7rdzJWns8d6IgGGOIJrioUuDtWPZoNM
xzWx03MP7SjPpBIw6czeNxMdvHdqupji/sQxFSVVO9N5rf0hzFvsFTgmeO1qk+Zf
WBjzGkyrkS5Y1myATLSvqmu69UPuKyJ9ZLV4vBkrffWGAwLLgxhYcrCUrSoI4cei
4LtEMlc+VNqiRDodyqdQi3BB9DtfLvdKA0bISR/E4HhUyKjr6Aa3q2tR1rl5iPI1
hm4YKoYCF6K1QXUq0Zh+M4/1zGepGV3EU/bBTIi50YBTgW+bI5FbaT24HFBDppUZ
PnGQMaz7Ti/zJFkb0Rc1zj6gAj4KYsEVv69YDw+XmlFAQbAK/Id+tMjF9ELFZLqe
hK53aEgoc19qvxeMIyuys0opK2lC9weOIezKNE9PM2gkY+X3lkwBCuIco6LwXvwi
fHOYDds/2LUInUe9IQcf7on+DtOR2eq0JnwtMk3cimvcoqNej9axibOQ6Gxcp99P
QN7JIgI1yclDg5wgCnRDVrr+aAEAcHcmdGlS3FOCfaZ37qhWvEcD3qWMxOjA8kGb
88jyY6ovdE3OgLFuiJfqdwjtbPIbEJyEeIpf6oqwtnfzTj1TwNZKaTjIgindkl4E
MQ3gxTHBEgatdo3aJCKIB2fwCWyKptCH44pMKnf+aB8EOC3Cpg3g2CnnZmMp+5fm
J0liiQ433ztk84FVle2ScBM/nWhOUoPTciEnVhIqhlEDy2SgRF7wfvzFNiY6j/y3
bhL2DpycC/M84hKTGMTolgbBrQUwyuZZgl/OiXsGpOxLLhbvcQqldUZxInJBc6T0
y0yS4tTNu+9XeNVcIvYuHr6F4hY0E/Liz/9P9bbAXHiLSonEJzyxV5r+k6ct2jqM
mh29/IBzZJ7/Tf6lupjkOE1Hi73nX5BR9NdO8oOJtBVMcXXayq6gRP+BA1iO39OG
v0YuE7ZR6SllwZsapF66rZB83wInsFMRkyxz+IFSzcLnEsSONQKDnNDIvEhOhVUG
9ZIUrTQyAjWcPogIc8plJgGN38GPBzNhHdZE7TGgQSRd8e4xdCH8Iv5FhRrTisE5
6JsniAxJyni2ElLoP1VRbR+GJiML5XYmsIs2QZoCDahyFgZeG/o8Sncc1LzUJ2Ah
sbfD8oim1sr+yeGgAgv+Pf/MrzZBajfMVmyS/i1n+QoHyMBQy7gXapMgj5g4Wx8f
GYR+kJO6B9TItsZniOJBoVGtoCnAHWYlxoKw0hV4dpuGZyrWSs1tusQ/0okygB/h
S1MBqVyKaENoQ8o3J2dBRuSBegpwaiQalddreLM+nhJSj5FIRsUldK4tbGDM7IhA
wYhPoWX5KmbWxbGjhTRsZqqPzPYNsEfIU036jXdalJVP9dg/O+PxXvQ2V2qxtKof
mSI9kIM9iYyUUUnxrC0UPaPfalxSlgmTLhHVZj7Y6IB5ohksX+anDpBjOJuA1BTP
vRPRdlcIIdCxuElbQTiDnV0Ox3PxHofRzFQt3vWffQM/oppj1WBhdHSZH83cH+Pj
pBB9ne9JyWmnyJjVw9+qX7wChs8OAUt8D2nZqlFuKAKcTKHvHvov4jlmjxom69OJ
aLXar8dXSkaj1SAAQJJ/ja78IhgwyeWjSU5JCWRp0LHe9KtG6mWjLnsBCn3q+geI
iSRuDVqs1WEIMS5+SwZkSTZpRTtLKaZJ1ySypA22U76vwx+R72oqFQ0rYlmdm+pq
4b9w7mwanws0QmMcqC50nPIVjOmPvJYIQHOzLfs/AlGRDMIpkRtyJ3HteTDhs6gO
+8zPZrYYCPqDr+ldgD9N58ZtVuSisMXMbPEw+4xjNkSHGshIagk8DAvB3luFeTbx
gZTmoTwC1eNmbbl52Ilng50BW8mxOzNqlM1Y/rniKsxu/Hb6XdRHsqwfKeHwjGET
7c1e/NP1hRvVbFYYCwv3+VwFN3g6JtONROPafQ1Gah8qtQ7epSPWUOLdSe+ceL+j
rWmPsmFJBHgRF85yqnJMLYMVs8S5FcEf9RYUPXQOccfgH6HXoD9cuMTSwYeCYPN2
BdXYj3VK6aWPeZOappqDXInQbw3+Ckhh/u6HU6l4ER1PSl7zaHNr1h7A0GYgJJjf
sByb6arMEz8MLbv+8zM3EjfwZYIq9uuULdkj1bJA4JXeDmg2CZmy06gIguFirisV
qdNrGCM/q8gvZUi6kI90OJ96+nLxexW+nty/mnC42xeAe9bHGZ4IXeB48U5apsmj
3i+P40X1ngnY4avBOY7T9vCxbiQQHXvk+ENK3k/mps45M89bIp7u90l/kWz8TMwY
o74sIhHxnKeIDqsn1n3qB3JmzosqmDKZUl2nyJ6vm0CXngHm0bZjWC7mB3lJWS05
v2RI7uA0oeo2MMulD12AyUEM0JQU3xR1SjtlnKysps5CFkVeUYIfl8xZ2KD0FD9+
sLhfwZzCS/cyD8rN0j7+bYDFnsECuimTNquOfmzGg3rCIC5RW5LsZ/XqR3P55YPL
jRPpIdBvHGlcyGtGnvZIaMgO5nV9kuPRdXfreJdi1rSoOg0AT4T/TGczXNoOltNR
KJ1QCRrfasOdhrLMDd5Ooh198QttftIqtSi08AuwZRS96C/tswP/Z6eb7jcK/vnu
dGGPQir5Ad7zSpGg0SKE5/hj0zc6K/B3VOQ9ZtVaSlhwHvU49U3DKZhnzGGv9jDL
7BGZwv9anFsz9V0DI+M0h0OIzBXJWjCJat7lg+pvhqfzezXEtr3a9sIbxgFGo0rC
CuSvEsYMEdVjfvO0GkRmjtVrFlYU2SXTm8FHfcxQvpGvSFOcgLl+xvVDwFFy+k/N
gZO+2OCit1A2wuTy7R9MJh1YIq33de6L8Uf8FnGwrouvCXJHJTZsRRg4cd7JqlfE
sUNiCoaVACkjGbu8dFWrJbFG+nV+6v6YQgwAiarabXIEc4ok0Mazu5ESXJTe0dNE
DIySV9r/tB4DyO5A4oh13/vRecxL3p0pG5b7iL2LI7KqaJmZ0VU6CKlHdVhlUR+2
K34zRoBOsvMZb8V1qd5RP8Ur6rP88C02ef4IRfJsYnKOsIasYNfuVCY5teG2+Kxg
G+aUuGV3HXTzfr2k4jycmfGFpiqGmX8EnYgS9XoOMUiYez6o/601wFcf7PvlVuiy
rdZeHPccYecST05psQBqUypeyNdsu55WocsaMircqLCz6036WS0eFv0PPE1gjefv
7MAtPYYmAJk4tQyXnE1KLrEpoy3wn+ghZu5FVzGDb2wET0cfZn0RZES0jdAyPHrX
pkcVzeXJWjrXPcvEn45Sxf6KLXHJxaM83UXj1BeMaLKXMyxDmAnkIWRSvDRXQA4r
6efa5JGNzHD2sqdbGTwZoBB3m4T0eGqChLnQwjt187BzvChian9GhrHBlBChJKYq
3U/JKgxwbtkuJ5umhl9wOHo9mB6y0k2WRUfnMe8kQtm2BkPQh8Xaz3+EdA8qHzzN
RTchNVwk4RtxE5Nf0VYUq/jG07x0uEberX5dfQfxNBgAkMA7bAluA6oLkvmw7xa6
1sI0224P1VbbnlwLzoIyIhX/Lbq12Sr8br1tMv52s2Ur1XSPNh+c4KG4HGYcfEmQ
eAEfTqd/gIYietuuJZDEbXrbnoHFN6a1LPM/6e4CBXEgUHVPcu/SQXF+4spzlNTz
DO7/gySaCJqr4qGEiNk+8PVMMudUEzk56EmAw2krOWIfK2P7Kgv15+e5H4uXDRwA
P+o5YwAZiLoH8J5VvWrzdJ4nTjedoYfGo0yz9/mHXXLJppzNeTQWxcN0AJujhuiG
pcxM/r3I0Vg+cVmSJ1Mzmf6aNfYXxod8yHk14oficX4+LRhyxMRQVAOYpm0bmZi1
Bgu/WkM1U4IhAwq8EgqiAiDJOpeUqvJIwOGDMftOUWrAyrn2tejB+TSBoMYQu8eT
6EhDcIvZeN5/KaDLkaev5WxqnmctKOjBhB8x+zSnwtJpobqP2oE096J1xvMygahF
f/KRwf+jh59gavYShpdmGXp3wQFbm8dCZSnOckVhDKr/yQP6n+JGiYUqfHDda0h8
LJBjdBe7K4oV5hqVTq1+Wu0By8u4wPFx101SuknlAhOzhmVMX1eMnxQ10+1HZPmD
tT8j3mvjxBlyvNOnMSHMLPutWQBYM89XSh9VI9D5TBuVhJSIkS9l6HuSSVVg+O5Q
LYoUS8icU/fvFr8rdYbt7Zxe0V9DLZMLJUK0it1niiMHqf0bAyXNhFREMqcEIoPT
OUSrUBD0hDKp2bCScHBNvIV/pJUIYYJkOrANdVq5Uk2hz1ntB/Qocg75rINrAWyd
1WbWqX3fCOVzeAlMgDiKovWNLrGaZel9MpVMZjPv5Ga4FRUnwv7uXfjoRBgwIt7M
sGxoVd1Ij6gxQSS8jDA3j2Hwuv4dW98xhk86KjIrVynfmHSEEFtK3qrBFYAEa3yT
o5rhTfllfN1o68JE9OesqsiXT0lIs2e7Wt+b4E+oo4M1yWom8+h3x+5tzgnTqzF0
nAYB+pS0p5jPvGfA/xDTnmnUIO3Ue7M9ePAXhQtghaqV/+RhsnY2bExTFxgm49kY
+oYNBLDXOa68VUaXO9HUhtr7ODISqltUSCG3faQqWY+y1KNG7LdEVYzZbziZd1dt
kvRryC8IIUrToXVKmDvkSnxyEbdca1PeO1A4WL5fvXZO3VA6GvMnG2nOwty4z7AE
SCAVU7mnqyvVuBRn8Hgj8a17+6vluigxqAMOaKS9cs65klq3TT8MKUFdgPVGtBhO
L+WtNwLK8OJQJkv8BwNnNDEm4JsvETQAzJn1H0RirsyO4N5spEtAMS/KmTFqMFoM
XZrPS4SV175nmpvz1ZriYuE1aU+Z3svbed5azBCAeGb5HaekFdT4r7o9L5LadOR8
BeWgwM6Y8IU69ouJdwdMeH5zJR93Yu9vsijcuqWiek4JuNW4CO2W4W3asBFEI5U+
v6X6vZUQZb/5wJEvs2t0dSyCS736hSQEWnv1KbDhQWTR0d5b5e90eNB+tn0//iKy
iIOsPgik2byDMKoOLZEeU+03/jOtYGeELhkCOo+QZkt96IZqFC2g5JD1ri1/NQlQ
ygyrkN3y8dOVfzctBzRNLuEWbfX8Y9v155EaZidybB46x+dbbZYj1lTSPjt1NU4F
16g8G4fGwxLocF0OXcRfAd88pxQVcF9b268ah1dIjbwj6/gWJVfRYlk+yMEqZVcL
AArBM7R9xfVFSUuMbayqvRxrkGHJP/bS1g86tbFBBf4hEaIeud2q0YgPZK/sS7Lt
DoXwxNqiZ/oTkXSvjSe4BEheqNavKvZX/rlqX9AMHfV5OixxbDxHHYAN2P853b11
KsYOOm3FZLZDYScg7+6g2LpcKA2XWqiMzguunk3NSx5UOsG6eOO1pQSgv2Qke0r0
7uTnK4d0/EGp/23PCL3Y7Gco8IrY/qRwCHAfeqsISPABeg1U47/Y2hgdeOw0c2Do
S6uZsRDG3bEsvhs8UjWdTSIKfX+M3L35PDSqPJ4WUza5w7frxEaJf7TtxKePQbIr
lqXamPKpIyhd6JGBSB19XqKrpVnyVU9F/yFro1HoYD9PqQhphSOuH3UGASX6zZY6
DHVel8xddH5MvMXZkgstc/XTHjhqcsTEsc/OoQBJmw/tIO1NNEc7G13vweImivnQ
ciGRR/7sQJYpBWIhNJweR0/BDS2EmEIZYTjsCE7Cn0vpSUhOc3n4seTlceFmw4u6
oAX9AB6hKQylnEreXGnypbd/cHBFrA3yy3jwhmi0Z+mUk6z1n6ZLksZEgYuVbx5N
+Q6BiNvm8A4+YhqoEFi4gdTlTjkfw/uGCdugNInTD+7Z0J9KmO/Qp/2yZXwec9uH
3+WJq57ujIDDlLlWaVDI0UE8YfDqObHLAy2eMoNPdtYpqtPzQIJ7fguatVWyIE5u
eBwUllgPLXo3be7nMa7ax0gmWfoWPJZGMyK37bqGdsAaAsIH/TLYFo6bqic+WgGD
xcEfrpjjnkGpkL6SfH8J6Aodh1OVDfsPPKpUlkibXfFauMa3DsPMj6j+xvAsHQxW
Mmy+t+J4vBrU+cST743J9tgJnJikJKK+DYZuq96KnJzgA2N/qwfCToiaDV62R5OK
rnmJAImcSEkXVOsOkJ2QPOvyUZ6pIrwJtqABufhnDMyR1iTZHy6pBjbnRFs4cege
np+MoBVgIikDbbuGJ3vjSZ2egPrGTlcOCgNScm9/n0KOEvubdJBcSQPtL761AnP/
lawXeTifx4OfNa6S/xDJJzE7WJ3ZJvXvY3XmxcaHR/DneJ/dJ0f5u0VFGid508rR
Quth6p8FT+Ssi/ovVNlZ12f7SOMei0DYlGwJqZnBjr8rxl4nd0drAflwMO6JnPhq
ZSzN4fMbkhJLcC9/M9sqwVKRAFZMTbg6INMIfulBqBi7bU8dd5L/6TURZGmtiHdJ
qTCmYQd7MbbsWqf/TqIP2ld7U3EvG108lY6gwHYu8P7yKpmvUPLyITnSYdn9DbOm
pjBlxuWMtJ9AO25XEWf+N/+QZGDNVSt0jlPBTYcUGinGLxcRppOqeeLg95yS+JfR
t6Xmlj9GpkF5jzFSM/GmLAARQpEHTr36CYJoyTMg1oo9IFHAPWlZQgnXa8R90a/L
FLRVwdgBKCIkfFcKwRk1tkKkLP99ipyp+zb86cQnmYEYVRwe2J2SCvMzZorX/fIH
lNqWidartMfqtwCzPleuXtS8dR7sEY5ArYaRkqcbPaahruYWNA9QUqbre5puHyuB
GaoiGyw0gm7MyQ0fy28Lc9QyF6m9yTmrqj5h6GCU9ObhceXh1ECldH0O43JbN6+t
+LqJO/pk9t7Lu0Hi1sLBaSKoGCWt6bFS1/klqVV82RC9dRiBdZJGTDIjmL9OOjzl
uLyNVgehS7rHM20ArAglDVoaq2Cwixe9QeVBy3sp5HyTYT2SQiLRxC9NPJBiJvPW
4HCRFeiWAqrYfOs8UJ7V/w5BfkuzuMT3mzJ/8FrTGULhJeQMrQUoOCVXVxMTg6VO
H/HFygtpqPxN1vZdEVp5XulMDpd1Dpt2oorDhOmtgLpEcoXc78DzUcmdspZz/AC6
LOL0qjg/4Hr/svCAYwFs04UVWykkPZ9I7EjNWdg4LhhmiqyPou5YAQGYXFP9EMEJ
kJx6W6NHn25kW26jQyWUeKZuPN8DklJ1hSaKknNKYZDBBlaycD7ygdll0CUYPSPB
95EHdXU15QOYJ9ZOR/jxd5EL+1cY3BeO+kUaLfHnXmKcF5CGDzxhIwgV0fQPsc2G
D1HSvTySBlio31rz0msRyeu4fwCdTv4si7S1Yj0DzDzVTpPMGthv3V+LI/zolfOQ
8AJNMG03pHsanFEGq3lqHGKpDI8sIJKjuQvT7AETMWRWd8Cy+1dADJc/Yo71DCTO
M3ZuXM+jbCk9cM9be0gNU9Mn0a8T3Kk6bUPsuPqipNlZuNzw057FksiS8EuVfGVa
mDopVH7y5lnpNETd8DzkEpiHG3iwY2SGQBzUaCT9maWle0LL4AFhLU/IY7RInHy1
+Uzi9DWIEG8REhMt43THuwSZjVjU265XLDzxh9cBv2ydkizh4huy2e5DCGJmQIBR
NhJsw7MWd3g0QqJoDaywmAg2YiU/4vb2x2cTH+xC/T7teN3IpdEMr+wgoHJrrkXU
OeGP7myHaqdYYlQCoEXW2cJpRg3YwdeNPSTVYbm5LTbRMteM/XozQ5NE+++OySDj
nVTT4VZ8geP6MCd4vAQrSF0C9NEqsFG3fsl3yGbrTzhshYcAe/zONUJrt7ScblF9
RhNC07hF7uYc5PSB8I5icp6DzdYlzd6KyKvlwHrZhAx6gqqvMPeKjhE0vQ7dFAO3
dgqEcoohZq7Azzgma8Xx8xQuB7Zra3gdyzrDIdlMK/7Umk6y1twCDgCcsDWQAOcQ
3Gg11z4r2V470qAVutYbrtveIluQNfJuVyjj92Kq7mej/4Ispm5JC5cn1Y/FQ2WZ
YnBfX/ybjTGeWFFkYz56yQ==
`protect END_PROTECTED
