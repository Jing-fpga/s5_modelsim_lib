`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WGaTu5YFdwsrnxSsnw8S5UqNqtcj3QB3T13j2eeAAkUzGPGjlwTCYOneRXNfYbmR
ck5j5g4vkoTHN9pP07gaVbf2EyN2g1YQQ4zZsl3XOKpQl7BuepY7Tv90O8BVnenv
/sPCt7H3U6ctTHYKIqEuz2HGQ+4CIb1G3TPtNqpw2Q5teec+Uew3zXCAuR5E4Egh
WqEBzMzks1i2PPsFPxt3z/UuTb8Gx99wwAyW2kieJhd6MCTOQMy+iz5CEzXAIySB
oUd4Uql6kjU8UTVmgFErIhHTHJAgo0UEh90PAksa6wXNG/EjB1gDKnRDZfZiwbD/
9H1hfZkijXBI5A8BPNwLSrdGJdppz8Q5aGYsQFeW0AtekK2773iba6qNOGqHMsAx
Yde5P8sJ8hhFH5KFDK6SoZiO5v4f8+M3xOFq1hctwAymM13OC5bUG67LOoUQd1Rz
304iezj6lvCmgGfC2+C8q5UWCrorqCInkm6DkquRJe4lnTdW4FeBf73TitKtpHhG
UgH30yfuDYzgxszsxxkX4nZJgHX6Cp+X6PDr25OinzrDRa5t552YcZS5PTYa5WCN
Fq5p2Xicbkf1OPJ5HjoxcsnR1gONid9aTyDIIfjxINYbTPpRoJu8JvLz8BqBTxpk
1MUEYbu4u2LhHtGIIMQDIQhWaXt4CejYnBPBHkzwsKd7jQB3qVjyze5KY6zs/+P+
IPHnEUPXjAPiHGFcum4jTI/ign7bbd9YTx+WOHT8O+k/5nq1zDjK0xMLiN0j7yN6
u26tLx/TQRxobu2RgTasnasBk0J5gcLTLj1U70DXs1GHuUE1sbU38yNmk6waToDm
buBG38BzBnZDyQjeLCBLoXnJXkT0CnCZUMrsWd9jlkBHzFMq60UY5KXae9mP01O0
7O+pSwcTx8LZq7qap6cJWHnJj03MyXv0YrSSXajL/YRitkktNG0/eDf7ssZWuu6x
ppaAVyhGmS09I5Gzxr+UNRdp4RQJ/b5MfqoJPRFBG8v4TAqDBOWnF4d9cH4QnWzo
CvoZhYZSBkK5PIwfvlnOYaVTA4d25aM0G4KkrbAAELQjwbJmmjoPyNYOYy0HDajG
HWGadC60hSzOJtC7Hi5uRpkNxWTw12Adrt0cJMEDbXho4yXykUUbW7ddlD3XAoI2
u/NwbpOjOi6xW9fgsVmyYqzpWIDJKd9WIsSy0Y/wQ5J5UT4hADSEexgG50ZOHz8S
HF6Tw14xW0CRzh6fTqkWy5ixJ+rduVSOQJOtIs0bi2kLK45DwWmmeJPyvllh5W9P
XU5dEJstmFdEGgZiOUaPJIII2zrcNEtUW9+HXkdi9Q6kT527IVlH2L4yv2dr0vye
UTPGDO3qPZH1XYTIegfXZt0MANQmNVNAWVfuKqeEOpoOEZoqh9v9BsKFI0sacppF
zEN4tlJptPebC926AW0pWfSuyMPP7GppkPSAzbvAN/h0hgBeMr/jY+cMhfg69af4
Mcc+yIV0JekFxOEfo46CuLDqDGZWQwRc4f5SGXR7wIt+tFDEL3WEArdxjc7VC3sA
amr3N4055o9xCZamd9qkxCDJm7VfxtRj+oMpEars8d275CBaHkT7B+lJRwaeI+ZK
MBHQ+REePB7g2QDYKnd0RpaygcVFPN+05hATEWtIuwjZAMtw4ZrVy0E/PZcgD102
Dqxo+4SVjggPDNilFnkhmw==
`protect END_PROTECTED
