`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XzYH5maM3/LCdRPbenIr7x/zCrqkBlGnISRG8OOWXt1n64QgdTv5bAIJbEqA6Y2g
sBG/wNlYzfV4ziv/jYsetpbmmJb/5Gq+tyO145JiqWHUJMYj3XC+sxqzkvp05/Jh
fjbgx7whzsd9w7464/wwJKU3wvXnadICdLYBBSuC20/YvL/ulmmrTYfzP7i1C+Yq
i86H7gMS3xyCPSNKi+2n7cZj/QIXiO3KpN6/YKiQk5oeVm1ct3L54kmYql/3D8z6
AEAYwpbVMMcJqie3pQltqnK5/91gRK2lqwNpL/6vG42Z9BXZsLfVxN3+gxYCEErK
2EY2bDs+5za3IhnetKnxInWAfHXgbqFT9TG8e1e5ptmS8GA7qTbznRlaQQ0ge6mt
9M8LTxJwOgRL024y4VsGJW5uqTYoQkZhg+X6+7Ph9eYIsPKx+3tRgp6699xrAT5G
0PS+YfLEokx/aOj8cKquUNS6CEqA1GfG1UoJ9C/ivFeeCkaczYrH4g/S2eC7VU3G
LXM+TfYgV03htbTDMQPrSJSrpLXaoSxGBCvBjjq4fivz5tFhhMArh0hLGr1fjT6r
sXB/4cZ6kMlWB7xAAVLPPxn4kiKnvaCSozMsgPi3xh5eqJmnc8DYhzNMmdzsEig6
G14lM7lIAEJ33IcCApUPpY7dj/LtE6eQX620qAICwPlWyjwoSkFJi9CGMOoCS4xj
VN34It+Sf6s8GcubwXaCO5gb7cUyGB8Oqkt1JJcLQHxLw47Ord6MnfNbLqRsXum5
Cv12n/G6HCNtpPMAk3o+e8YUygd0S9u4UJhrsGMjP4Kek3BpuXXNI1x+ZE3Vhqw7
3BdhEJCViAPSNZuAWG/nKZZNCDQBc4AbNMtVI8v942OeDD1IaW2RJSQlCG4pZGR0
eYwpt0UvSRrl19Mh5i9rIS12cwXKN0Jvsgqp3BQk7E/cMFzzUldBSK0CsqoKZXZI
XtqVxV5mol2wh0ii5BFF9uLPkClBZruzDhyopXV7z951SIYGdiGruTQvtMMYkI6p
AOXbgKuagyD71jqm8K4VU9ktQUP/pw5QCXFWI1mNTDem6gecuj1fiq7EyBMp/pG6
ObVpcrlge3fs1leZ/TTB6SBw5DqCj8BIHFgGQQXqOyTvYBMs0obrZ8w7EFih+ItU
FWRWVqI7xZcWC/5JWgDenh8bdY+QHtAkphTn494cSO845fh77p/IAgSy2/zHK6Ic
tbPHz4Fa/tynE1Ak/hbqL2KuiWFvwmUOqviAholwQx/nWW+lPrwlIaAZ3DSH6frr
E182tPva4v50t0Deoy6IxRZRBdWQa5apW4tnIlOXqZ+zgToX8DkMso0VwPHxzJIR
HQJrsPXQ6tst+VRbeALrTRWJ0qV+282UPdQp0pNAt77GTGixINTSBD9KYVCt95q4
pgC45qydNB02I+Bva8DXr9Zss0dbG2YfpSTCulwW19/gHTEmztpgQdAsEnyjho4A
PRMIkE0SPbT66QySFdYOkj4mUZrfek9eStWt5V1k74A=
`protect END_PROTECTED
