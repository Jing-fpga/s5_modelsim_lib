`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FgYvPkFWcDxzBEIi3u9sBC/dV2xP/jLCKOJ2kB/cuZQFHukgrlcta+25eb0htr5Y
oEr487hu62Vs8U7q/cFIC17mnXhuKNE2mj6GHWoW+CmCWNniurS15MhZN/GrFvmZ
dvTKRXO8REMvTj4cQXszBTUqOEQH77NDGfj8Tdtzw0nN3/HGHC/EfWcpSuCO7qz2
jkMdyg8JLOcvwG4ql+gjb5Ub3PKx5rQ/5Wb3weRxGwl5Z2IVpM0pkAvpl9CBi7Ll
Kqoti6KJovtrBJHEqropkiOySZod7KATgsw2n+7haj4XsDWK5MFfARGSnhojMVM6
jXn8hQKEsFwfVTb0z10n9xPFqorzQpf1vs+MZT9n0haFhBQugCKzg5dz7jAuHeDv
V2Oa2xNo88g5ZXTzLf+cgF16gFBJWxdA8QzC8+CGQ0FboiCkuxzSboGgFhmpDisZ
WE4TsOZCosDVOr7sqwJBorq85QiZ5A094AZY2/SJhFp6Z7y2+xeXElBKOl233+MW
3UVvtfMAZdpc31ohaOSHw5pw0H6LylO6ZTK7dgTRE7OMWytHyJ9lzO2+fgKOSR/u
g8b3n0yOG/RHpEQpRi/lllGCw2LwgShyMhbq6KEs13OUJXSsUKdevbHOGv4HoZii
lc3tovQc6CRkVEtZ6tSMsDq3ZmTQKIk+TzPJpLd0NQhxhWkvJfiKerVnFRt6tqKq
3KDGC0Akp86lyr2nCp1LR/yyvq6Ibxq0DKwdPmcxqQxAY/Pm6XF/uPzktGrijHCn
YCxoVmzU+lKbXy+oFTwOhq1ZwyWECxFxbXdPEvg3qXThS/BYmN560jtE1pct0Wil
sl9b+HbOAvykGQi2JRAj3bvdlftiuY8QuizssBk1mWa66wSSiFQws79nHqpCTGVD
jwurxT+bN/NuCJ/9i1dYfUsu4oJfXjikadVpGtTiyTjUvk8pDzzOuaNmWG+Vb6Mv
hxpTIEs5l9vNhkOhE/geV6MGk9pA+ggkXdbeSquOjl0XqDnutt5TMY6fE3L1DuCQ
BUFRJBRRpRrc2jmdWPwNjsT/DnuWk7b728MotTTbGPnho6/n3MlRqRxmgap3KmBd
VpUlvPoA+4Qlh9yAGr3w93FyGJZrY/+wNEvsnJgi+7czdlGY70CXKRt0zV3DaDvN
cchfiJ+GyVSU1If3Gm9saJSIe/6n8BoPnEdKpyws8Z8JB0H5Frtowq/a0VsMVWPl
GcM9oWEK9LJcyyK690Gms8WAozIvLUuuRfFLB41TbbogQUWPmVJ3gi32hUJwg5Gq
fQYnSmaIRM26dOuD02pJd+88o9yxtDV/+7c52BxcdeA=
`protect END_PROTECTED
