`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fnRsGkXSoECnRpqHw+A2dT7Rd7Oh06pd5f0+Va/MuoAHLyIVJ37VC1G87+BGNlRV
KkmzvDE4pQMKLAT2Gwky+DiVOvjruG9vvNNRSDP61GytIPS7StvZeZgpcWmDvInW
z+msErDNrGZ+JIJw8pt5sOaP1JUguQVXnUIYfwUV01VMoMRrAnmRPXKz8RNW5vQH
3kzl4U1CxZw5UhiL3tcyTbYr3XQBsztxJVlus2CyuwNReOPS2evsIl4iKdK0aTHC
spy5imVAuJhDb46w2NBruIaqvxOGOhx0MenZufSGpUu/A6bVb84yWqdVankv+C6h
y6TA9GCvE31Ja2GdJDC3c4F70E6rpdlldAU6o8Xzvuc675U37RsOFucY8uquo2mC
hsWGaLLkeg/RVDy1z5XN0YW2rs0+SW8USQGN/ysAgmbDOPaftDXHCqcJZVXYcStW
qosQpiCTFl+SfZFXGrXrbA0nlcybPncWp/ysSDSRtnkeDjNN+YwW/PfDJPIbqYgf
0l6ZF0JZCcUZla+zi0dNVuhoorjkbLuxYqi7+fqDcPq80hE6aKEqwq8aOb14XUtv
95yS8/thCcIyjdvpQuH0iBiqUnlUHlN75o9JWMKUGTkK/qLb6RQ0kXlkkm/vZUEE
+UOUOIsQqmmEj6PfhsyTN0NV1b/EW/Hi4kznd+si+d16ycKyPYG7x/VMpqUvqqqR
LPcnR5PclSbg/DxqfmcNEBVi6HUjyFOyIBOR5smcDZspYi9p6RrPL9FYSW52wBA0
bvNbgMkSsgZIzR898Ngd2UDxDS4nXSC7ptdVwh6qYe1MnPWfcqwQljkwIl1xCw7M
juHmyepfHmPzyylMvwdT8aYrPRSQEB0BfjCxC+Y9CwnwCWTFKy2Me96RQ02fbGm1
6dUzVTDjdRgzSFV2u0cuX9q8+iDNlR+5z9PcGcXy1U4SPW9iYYU0WCMmzLeIgLAQ
iIe5IFr8/QqnOD8FzVaE5IRQEvRm75qxnH0qFLk/M91uVvMXPc2V0qsMoWHI9K3e
aWz4FYqZOGBv9jcYWKRxAcl/f4U8Q0Wnkt/Zsh8ZVUbj8hcItLIzaa731UxX/kcA
tYVOd8KaR0wbVjymWKOtmjZsI10yZ4Rdf1duA0aoihqIDIPcA5bWyzYT5QwunXlI
OR5GfykiWPsUnlpJFyrr6mbxwefhycsyCJDXDhox84BLLnO2Biyd68mjkRB1tPyE
vXIxlGrbJRpjdfUPoj3njjhC/7rcazmER6qXYDIU3JKN3kQ5zV1lHjjvmMZwW/L1
ABZK/bkIa7ny1X0rCl2rROtRGN9tccIxzu8/9yQZwxVOlgfzPpvYrAsDWf+OumiQ
8en8VAkTidB6OmjJZLRSNVZG80oOpvJUb1nnTPhG58+Rn+ftNWdXD7O+mdSMdCml
YpR0bgN1GVIsjmBw/y0osQuV0GtmH/x9NJRNR4wptkKVfvESWJ80zN53Tl99/Ppw
sSZCsZpkT0fGziEsYCuPgUsfdxwAn0I/ZBkZ31JvM6Qf8ZMyjOaKJdTezkaDnIDD
k/7vg8MuQ8QVby0agY5mgnNs8hzqFwTJzmsVGejaXt90K9ipL7kyiWlwRhzisX6r
6Y4qAk53sZFQwQfq8rkJJLwUksBANmh3c5V4Z/eiLhdRWZcYg2brym5IfIGHnvOx
S0jwhcK3O8ZsmpC2zO0PX7Ki+ZF8enxDfnuEy+HY946Ss1b07ZKgE8YdfK7BmA5e
WqrWN7a3sYU94juA6NOkgm2c6hjQU4h+eV5CMY1/3LJQHh77MfqZvTG9vQamShGB
2N8N8X1yR96AnnYw+LQTXYh/2ocSgL46awDpesYHLwk23wWGV2jat4z3SaMQLccA
/1r/Zgh2DEmVE9OW1QqqA+06nnc5QjJ+YcfPMfS3/LFCczO4EuO4xENkstqHB9JI
mYzmPTI5om8BlwJSJbfWGnulpcHT5EF2Pfk+C6lgAJVyFwbCCymNTRuQ/U7iFOgv
6pnuYTYIg/o1N2jSV+ldUXGux8hkJYZQZOH8qFt8tMY4bd2nu8tgcRIFQs8SxPXo
yl1/xRxPGkNRZ9P7PoyiqqhWRepJ8TZDOyNy58SN/ukbx5Z3baLCYduRivtZXIX0
ATUIlgxAssMAJSke8gS7cZcnJ0LfML6K0DTiAkJvw3+v74/q1myWoZ00o+3zEYy6
T5ioUXVDWYUQgOhYPD7lVpB3qivQ3Kt8Sag9Sc6Zr9LVfDDrrfhHLK6V7xJZeydW
vV/nqJaNnfiagosMy2CfLspMQkPIrdv4bz/Ll+raq+VVmckshlhiNY2NZ9jlsBwF
0zGQ7KUXbXa07ZTMxj0CkIqanZKqxn68np9VcdpnnUEGPXsbZgj86+1RrK/aFulY
0CAmSW8OtrUYLuS6NOksl4//lYsojAAas2uget+PLfLsQ0cNYKHPhHJVRJ4H+wp9
E/oLJ5UpMekCx5RsA1bnj6t3jZrhXcWvKDfeA67PApARCY9k8ze+EB69aLYyKoP2
vRqRL1vL8Oeh/X90U1BNEfMlkVfl1h3fmqufsdXRR7yx3/Ez2sHRbRhsLqYI4yOu
OW7eku0Nvk8X6iCum4X10lGNWSt5pE0fLrxee/lupg7MmaCK+XjCmZDrNBaI1Q7e
rObxSnSZEUG6J7GEEsTfRvOVODoJ2BPEVzUdUkyo/OiYUFcurcGMKB7tVT8GMeMc
vVhW7B1xmSfrduwOcaEblb5XehAQa2xwFv++nMkfSPmU47vcaQKMzWhoJYGuy6pb
fLp3IvcS5zAhyVOgIVrK/6/KO8mczyuw8LDd1fOfuCTh54yMvvYRW8Bpzcrpb7OT
lKOaNiBBrqGi4MSlGEBk7hwJjMaE/4nWZ9IrhxqIfXMLpXf4dl62HfcniXLH8E5B
xhbdHelz3kXRbYKmQW/2Ahr/2BrY6UnrcEMDWDYB/wXw21qbga1wC4OROK7XtkXK
awh6V0hnYYBDvmrtt0PyKneKF9cqv6z6E8nj3YFdVaS5UIcpgHE7HCDEhG+MvCEl
ktMy0yWBBsR89AZuq1iiStpYjtM2Eey+2XQ8+hb/M5Ek2gX1KmjICmqpHt0yM+za
Fq3DktC6dOSkveFsyTTvP2iahC8/sAi97oALRaoTkPrFhzVENwRZq2zZqNANEGBw
g+11hObkam4bYfeTW2n2ULHdBFgf+NVEafh67Gf9NbIHXEhcC7FXBV7C3S9cZvJn
N6MQd4EyEO+UIh4wOk7Tn+hw8VmRjR0hlqZyX2QsPTe7RHYFgp69dxSHlOymTMVM
wJtdg3NMTpK0bReBa4nNOmf5LID4QdDkGYJnPbTNqvxbOxrphOD5YuWmsxPSwp/D
7l7ee5D8ysvBa4GI8ZXxXKtHZTgDuW3Ph22hCfkMC3xNrmLoGVIa4QBHeD2/XhM4
1TJJXbuqbP+ehrqGNkAmzrTp4fzCrv0xKj8msCLL13WLKxJ5txx0I7t/JEvlcsUS
Wkwg/cL7Olcsx72iDtRfxYtyfzaBu799xipSD6PlkZ9+tQ2oXYqSXTvnB85Rnyva
3sfX+7S1VOMHFTOeFYqPmWgs7WczzfrSn6pPLRc8KFUIoGDL7RPEjq8jfsO28Kna
btzMdYTV+jj1yX/PjbWTQGfcfZZnR0B8tFqdSt/WN7YiHwjMlSDpHvzySC7J6mEd
32O5x+t0mNBLxjF1zVMXVHinCxG/IEiMdsbj39TmdKWYLaAgVTz1fQnvM+0+UpEi
wfEWdxu1DKg7Z91X4czj/687ASTkYI5l5dw1qfv+wV05YbFmNjMZVULOpEjKJRSY
Z2QpjgRVFUtfk/buxK+pIV5q/g7Qco0fsxtmjN1XJl+gKinegFYGad5VxE3vTwzi
vy8V0tKImbvYtH9soJnaByUMzj7Dv8k4UrjApL5W1ad/hutj50LxsRuDHHLQ+GmG
72JXT13uTh9nqVi5ZgETK0cb/3KUfJO0VOs7zS8BrLT/NQAQVzMiWJB8L8tV+ysh
`protect END_PROTECTED
