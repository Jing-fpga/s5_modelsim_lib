`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
11hKqUt/h/xGGATg7ZMPIf/DZxuGEUlK6iV0FeXADmfgyL1YYyjfp2sh2cwDlnbK
T1PeiAlEV394rI9bkKFZGKyBrey5zEsyggkBFcj2n71biFP5rK8bgXIJJzRC70BU
Y+oZSs1OAqYIQrZM6h8CLWogWD8C7scLUXRpZlxENZmEJ0kZnj7Ye8X8mQi2IU82
bgLEhqhC2T6e7n+9LpGN8pgU5A656XDMHSLTprJ6yt7XNx9RSG0ZjQuC14WlCsIh
r8RGPGM6jbnh9kFSQLx3Da7gJQnfuGNx8JvkyO+isfIRKO+HxE4ZO3in+OceXGQp
BV568xqyqYGUo+8HkVSekPO26UApRou2St2KvXIPpL55ym7PhDscoVbMgot7wP2A
GzK8lIpFXvnfWEJ/OQ1XyOBPEiDqcfE4YyWfSOEvxl6A7a6x06KCyNbO7PuQEduO
ULguPWUPeoXh6tzgvw7oyFyIbFDa3fKEI4MI3qal+Sg9WRH/GVKzbDOYaupcHHNK
JSqg2eK53XcS9f7oOE+xjxar0nlrCnkwAFmjb0d3VMSzzWoxCdVr37IQB1kTT4U5
lw4UlaooE9LdflNGp70CaoA5Mk69s6wp2zfRLXOOkk0eeJQOaOHxik72x6nCN7t+
js4sXZSgQJoAqRh8h7yi8V05Vb1j2KJhrwJdf7FBBOUdg89J58fcUUAAkR1hLWKD
rqGiFIVuncPebJihygM/SI0gLcbhdZZ7caQnYfOlg5wh2/bIBuI9Kp4R6ifV5sAK
28XRzo8Vy3iBxYSgzovl0aBvCtlIQpzGTD5meEokFprzED4HL7/TWDydj4szKbYe
iosy9AL5601NsYjgwzkiYlX/2MAss+TpZdtd9fejh1qQL7QOt1u0764XwH/eXlgG
Or/IpMXstti41EZrCGN5qyxaYlP9IpoRXrQ8fIDbkbiu/jo64W0hDia1F1fh6THt
elri8mU0kxgNJF5xVTvABkcdqBlGgbGaSjIw3WjddxQBTRnSsFvhGLymLy0kYITi
ciE/37i98OvXwtsw5k+Sui9kjvLyyFloS+Bh5Jlo5buK87pP7vrxbOEUaG6SSMn1
TgYnAx8vhSspF56whxa1G259Q4SKvzIntsM7/N//UpkhBWvwkppleD3txeLjduiD
kX3cTYFwd/OVV0++py9IFhd4H0QcWlZH+ndx0KYvGqpZI8xjbaH1pSIZWvhAaLYI
o+8ZEJKn3Ar3/oKkzGJ9WD4yEN4tuYjG0g2yovtCmTonLlMF6YMmzV0kNp4T8kKC
PiHwYLXrlC64kK/T89zm1py0nf3+rBzd3JvGacULpf9XC6OqsQAz6t8ityzoPMES
K43xmD2i+TDSBGoCAQSxVSikvPv+e0eg0QJhucBN0Qq9ELXQYn7Z7nKM9jY40+4n
YxVHcTpKBtEAk46Yr2VxkcDvx4HSGuMRpFQ8E/wbCm4/WDnNiXmdT3O9MtwEcB+d
y/5KRJphbbwup5WhCYqXNYk97mWCe+bw9JJWdsnPBxTRCLnWcPHnM8hfLOgp1OKu
SxMDaWKbDJf7mL5WNfkv0btYnKQD6Iuc9OYpIJGuPEyxWhNKhF7jVirnl7nZLsvn
bOYDnOdYGGRVpsqujrEzP9UmGeW4iFJGItYBzIzNYUpYk3KMnbGSrUK9fG1/pl03
3LpvJDkSHaBZusLCNbj4qRKhxwY1dYp6CPzpsuzgKupz/bktMxAyvmmu2rowyutJ
XNen8RDyZacgy4ITdHS8TRjn3ZAfFnWhB8AKIIOdkMBgHw2gaodU+fez/08NGf+J
fpTOUM+VQRoCxZecGTzoclnKnQjut26ymcEa5t6eHAay64/sHc7Nyfi0m/+O/RIv
hnxRYEXqVBGMco1afzX2m/b9uWCKUwkB/5QhV4qmQPPzc6Hu3OPUiz8tbkUC4i+C
IrOiwHmrJfyhXT9paJAcSZaNdvNG58zFzJCsuwOHNhA7wunVC9MCUDjrtLNzIk9l
58olo8lNVvWRXvshM2dnV5g0M/7uYQc25ZucBajOM6KSOmRtvSRCMDeT0OWWQEXv
MYjH9KGnzDM/CdGC3s+PM1djdhX0RZfmvybQ01NSkx8Ie4pZDCD9gbdN1LPJAIrf
yBuD3A5mDvG29Ovl6ZNBMTIuyNq11ue7BfXZhdN1Kd8voC6l1S+MuAfmXxqcY1rX
8rENJsXCGoKB+A5hbKEwOngFw+xEPUnzvp3tekwQFtAcUKQtLc4UjoGKyaimGtMv
YrTnAOaKO7TKaB2aVSw4VCrVhTq6mrNCgTBq/UfNGeFQPvnt9WejjpTLvgj8PbMU
qbuWUC5tT556wAzY0YKMyEESVWXpn78fVNhCLuk+8820pZjOq2HmFqUnrSHAqmdm
oF2mYA7iQK9nagvQMpbdDQFubYxDNfev6+GU2+Z63svMGIggPrdWBUi8PwoGX5Mm
+Qxa9BEIQTlZ+g4OZXMXDM++gX1+MEfbOBBm3jRDsAv5YLltdZoak+f9dEghZjU9
r3Y4g1hWzA3vlsr0Ss9gIIiRTIAAFYe81TRWULi32AsDn1G2+0Y2+y2FrUxdcJN+
v63p/cgqX05SKN3QvSGGDwixo8VQEZ8rkqQbClscebx1lrV+VvK6dudjFa/RfYkE
WYM3XHC4b+WUodz4m5ccCfsr7+bYyCvSzyAfS7ayhiwub/mUZQ4xcdHzVlYLnMW4
8qXUoC5NITvSx7ZQQcSouiiOql+P6pAG9hH9TOlQmHHVVdmfyBJ/Bie7ug37Pj6d
KsIjFUAxofQXJkmJx3pAhzV74C+eOxf5B0EBZCu0TYe+YKoyjY/9mZcvYiHfhhIg
FNE6BOSLDPTX5TQ4gYrbCgFC7Y3TGzd8+FSNmt+0sX2y0Vs/+pwTibyMUFmtBjjI
y0033U6Mtk1Ph+mQWqgOvLMDYRzIcvYqDmEAmVy1B9Cx7pme3inwoKSBFraglRyf
hz8jv6vVv7duiipAEFeMC/9bARDmhha/ncYSBRiYcHiN9rlR3vN059X3i6vhLM0d
K5CZZTcR1qO9aM53Qv9nLoaoltZLpp3Mm0EXct9ozzFpiWhEha/FiSF12vGfnJpD
T3Zex4s4aG0pSYp+a1Vx1cdz798QrVSDR9Epkbub4uAjORUd7ja5dzxKbPrf/wuk
YG+FiN/Xl7jHAIthZGKfCg/jRfMYkOK0zZrOKeiM1DbjzQmusNpmdxa9jmFceP65
dKCeP+8qRp/IRVJ/iOcMKPH6DAw6b88iw+asIB+DHRSRgCNnZg8IPXqABhF+MBEL
xGIKDZZnPCAEzbmEal1gIhGxH6z0nV3Dv6NgGAClUL/M1QjkdFpSGrxiC7Dcnd9a
g7lLfgUrACjsoecpVGMKS/vL1R0V2EXrg+4CKZiGzai3iooJF6S1vTUsRDTudSgj
7T/l5Covk0P9EMHIbnTtu0WOnixX7aCX0DlKlf6IskdbwEPSndWgTKZSLqxf/d/h
JxYr9fdnjfgtI3NWLRiMN5y5Avgr4LKv8UOJkcrUw1UImEVg16h30nM4mHwEHDX6
VmmRlKdtFCianUthoq2TAJZ85T6aUYvJz3Jx2R/C3VPMTtsJrFTBjg34bUIo7NPZ
Fr10KxiBsbC0EuWHAsKDqH61RsGqPmC7r+ePDVY4ub3gyGUHlC4VmN5fVqRyqlBT
HyCU8BPX9MdfNFEr5/qHjo4qVRbrq/8/eS/mc/Eylg0JMw29bgMOQFfbvRk1ecQs
E0rfGdlNQoulLe1PKwcUPCWIDbTGVyUggRqaOJaoYkk2Ha7YLXh6l0cOTwiZSwbW
caHyZU4/PSdztFU39eBF454cl63rht+bnxU8HG5nLmnHIbS5H7ELFmuwYd3R3aG/
Ia4yLc/nWmkfgnMvxJOYRa1shjlEM6EAraAPEcoDVDwaFLlyjMUFJmUVGGt2gP0Z
i4oE7s68nfvUrPNWupWO58mgd58USzo1r0GaueP+f7zcD4Nsnb1umgBo4Aupqbmr
M16Ge9c7YQHqncGZp0V7pywt0IHUFSmpxF4lWHLaYGpz9oU0jnFIgl68TxPrSIhO
iisHd1/scyeW8RZqUxhMenQVMFbgNk5B5Gnqjl7UVqVTlAoJZQLDnmz8wAuXje23
Hm/nhFGO6U+h/azIJWWgtiFpOyCP86mrQMzFz/QhzRBYTKCB4bhTSQs6biE1xovU
6Pgvdf9GOCa/3VQhuhQTQfW1ak9DeI3Lt5z/KjrQh+CQ2Z+Rg3lO3ATqQXSIOhar
kQYgqI6u/UrCsKz/J1R3W2ikMJgiiO73PJlGdLjjTjOwFT60OehispMoGtcdZAP5
lN+BuV05ebq87FFeCBWDygT3Cm2ucNhWoiiEcvGbG5lPvGg1+l1EH5nIgXcsKBrd
ritqNXK1hLG1Y8BwH9mgTLBc2H0JQdHVZFWqUQwrE+rn1vitsnRNZKyzK5BDZZSj
5oJIBOhpZ2OWw2MDse6pDOf0dPsS3XEQdhatBytirvWx0QcH5BqAQ8MpiidEkZ+2
DKulNrRtUsiTKaQ/q1syMbE2bvm1mT1b20r8wP+dHIIqxCv4l7nyWxzkbzsZ7yRE
LwfmMXjWWBeRChaGiSuKpirhT3cKdKHzzu/5qOI3Rf6B2xdYxKl6zcEdias5Pddz
UUDKfvfGKFqzxFJu4SU6B7pJSpJJoGyDFABSfGQmWcK7WN6gEBPFF7hx974JJHKH
rmJK715hbDtLP75PFMSQPraFShNL04jli3SZoerOAAkXnr4brpDlNpzoI6jDVCFN
lImhcLHyEKVIJlWGjjwzkIpyc5JytvS4l5ZARWPhbny1lLrM+FAIntI47PbLhKFk
PmfPhn7qxxTBDD6HKIqTB/T0LnmKnAPdI59so9eZNBUVMpO/ywbGhzCqjVy1nzs9
JFjcB/vHpENI+tS6SCVuncAQm+Rz1vstBNYguEaQpj23ZVVcoXEg69vyvIDAL9qT
KdxoUe8iMAct9SgV6mj8EvKjrq+0vzZx9mPU+1WH+ZUmx2Pcs5np69jOaLSAZDDO
EWfcn16buXVYvlH2TT/8pDX8/Fm+K9rW695yrEPpZaLgfJ7E9ySQXFPoewu4OIsP
5zscJ73PNJmtnecgSp3Xyr1EoAdN2ykd1BKplWtKBFd4iLiUk/R0+GKcvspAii7h
pZ6iRlDivpa5HQ6/vKU2adO4QUl1dIFmZn20LQ4TdeKbtuoH/kP0NzkgPuerYc0U
7ucJqe8p/q0oUXXnkcaRTOz1vYlq/anijYt7Uqa2jkxGmz+YpMkROowqOVZmglxU
PFVrVxoB2zkIir9z5PLU/h/nDuw6gpBzzniRKoX5u7VeMyf685d95Hj6B7YTz6kX
GauY1Q1BR9s2Fc6ii8m/W/2lTSqq9ZPmd+bZUl/u8dqeJjcsUU7mnDx7nGa9bgob
UK7JdeRxOOybsgYpLY750N6UTQCrJFwOUiOpSWq9B541go1rr3z/yWslQBDbZ85+
giGPg39h5korz3eB6ep2IYpMmVm2Hchua5aDS2MR4KYDV9Luh9SpapVWu6QIG0hg
nXCg6mDOhndjzKo7M6lBfXRfvWx7ftE075lShsGexzN53wWHs2ZzQUptESnbjhl/
b2SihnZKGVHpN737EupXR3pYovsJa4rsUJJrGO2VYB7Z80AP7Fd+GicaHLZUu2K5
Iz1trtg4DLeai2yhknhdpXW73tqWZ/W7vQ0YUuGCyUebaIF1KvHIsdfGlaiiDSGs
zsYlWZkMALL7CBoDujIqO/UblZRpRqg2c0KrDy8bH/Y7ARWH57FYRRCDfJdOCIpY
9sP7O5afQ70OJwxkMKHzscyx8Zs6ULn/gbfXYHKsOXbVJhyyZmPyAmoV//19jykz
AjVmUmdg5ibmVuhNjwUxr/+/d/WvnwXrlOZQRi9QNq2lFTWkTYrogpqb4lpQ3NZg
suYS3+flXiLV7vusCzX7VquNuA38FH0KVM7O14YgL2tkkq9nCrXiTjefsugkKSZy
RnYM4Urod6gd/L51Lg9yThKVUf/MbTWazkHuRJ9xdbWFuxVZXgk1chE+MujRWtkR
XgiXeke8yfDZ1whSYXhluyHs1wCFYAPsoiG2rr3VCB5IhUWYCksS3lUhJsY/5FXW
hszL+MXx1S/3UBHu5vT7Vmu8D39xG9iVhgNRhW3RC6SBCVNRGy9bmq36/8fYOBaz
tmFTS6GhBETDGSqpZYHEV8bvATI0ZeCTx8txNGJWkLQOwMJEMUb1cE0xpY/jjWpT
7SnVNN+PjxUZRe5D7w6j+sbHBiKz7W9CMKdquonXuCVbWiygfZks77mdEEIYtLOt
2BPYBB72Yo0zYuhg3fpQXclxvVoSf7+O8SdcJ/CgrSkTZd0kqmtIkwxTjmAdYdlP
BjDdPHyYNS3f8zKOyPkQtaDO1iJwD+01wlqG38TE2NI3pzpV/d2z/VbNbpF5IBO6
R6KTuEM7EHLlryODJzlOkHC0krrloIEI7bkEEQfsyZB23FUaRO8fN8+ymEzah7rK
pcB2gi5ZwgF6PBnHod2lLVFKbK7NoxiLI+3YOTMk8+/+czRYZFNjtraNia0a0iyY
cQLsONqtdm/KRJY9YMa0RB4c9Uab92W/PNrYWQJCCScq/oXeett/ILlZLR5Y3G7u
K9guhGmXKtVnIZsFtw3xoPo4wCEXDXgnFx5OOad3ge+tOU7druFgASJORXCRjypG
ufrYq9N87faPk6hjyvKQQ9bdSQ2K5rVh+XRaq28lzw5epPH2aKboXmv7odOoeEkH
SaDXrbmpkBuP7pstGJBDhLb2wlqn0T6cJ+5ml8IKK2x1/E0dnn8az+bBFy9CQRyk
CA6SQM/a8w4XlDUp3pIAZxUVaq36aTeZsxPv/AKZb98Xw+lu3Q3js1CRph6krygq
0jEM+WSokTTstvokcdegN53TNvCrJE8EbGwK0PzpoCMHKoEJK/QRO0cmMvb33Yft
7qfEReNhtRiCRyjzrV1DT5GkeYJ2KkGHjTyyoea8WNBxTKjMsZBUF6QDoywVt18N
ZNqAeChFDQ8hKKqE+hDTc1xbjpU3FE0dk/Qmc5Si0iw1BbSQ6fvxo/vzSGDBZMq2
EFqKOYi5UMkm/mkD6JYpOhYyPXGliR//V/OaLE1wbheU5qhnvFN803J7Pc1su+oO
HMMWcQtvLallUxrfJJnyRcvdaxDTa0VZSrMvLuFASnHmbGvqsf682OKQdCFIslT3
hGjB3xw3x804C2ZP5eIYClKH2ge1D299AuJW4+GhCihaq7tlwvz36L/pxioayBOb
SxEGojp4NMZvKf2+zHzBfrK+AZRtiWC3jSYYvbnBCh6Deu0owH8MYemE9kGFmirk
4kGxMqkEC8MqnL7bq3SoiCH3uCH6D+hmCThcSCMsnSn0I7exASVII3ft43SsFdoN
2COtfBSrlLUCC4zGkjASM0uuCu1DF7crgecmuUg7fZ8v408IYuS4RR3KWqQikLrI
rvxfTjPJiUpGB4J9283HN7ebUIG2nPB7P/dWbd8Gwh1ZS0LI4F9CQLhVMfmavrP1
nI7X9F249/Sc0gLLQGriMIHWfE7xkLKMmKb2DFBNKfAqxFxWyx9G8TQym+ERli8W
BJryixqNvE+T/2aNCn56sYgByLaUKwJJr84YU0g06TQcso0ZS00usWiOKnv+gixu
b+wZ3ivcQcntkxvQ3q8jm3iCUnoDDUz2VHmchbmP5CfF5H2eN+Lm3Npr8cpJju4T
8x2favf/DQ8p25nWad/iCEhALBg6SVMBXbWoeknrrvQusMAxAErAnYzN9KrQjS6A
myyAZKhnwXDUTS6O4w7D5JHB9YDGKsSAD+hxtHTX/Bin7uq4HB5kGMUjPOh0xym9
ogxr+tEn3+CGx/cz3TK+/foGLUUo1Y4x8rbJfLYQC5rCZPQKwr5K81Qx9LqI5OI2
7I8ettH+TVlOjTDoybrVQgZsC3h6QGdzqIx5AwMDaBJyza+fCwNE0H/IwdJa2j64
Vt2ypX0rDkvc+byjxg+JbfNKPIPZ1c9KPqwxScaYYn7xJjGxqjAL1ffi5TKK4OYj
33q/0VaIH+7A0vQVn70A6JGwXUfGQRZMypb5P1WYAUStiUX6IpUjnxXDaSs+u6Xg
W4eidZNrhqNLAlGjIYN3tLeJKPaxOOAPCQcDX6JFg3ukKbhnxQGa/5SVsED2Pk+B
lGxeCILHBNmh6xT8cfQYlGVb086/bnulH+9kA62iNmVvQfB5lz0lY2gfyec5SyPK
VPVv5CVrPpHjmNhEWD3Hu1YvrEuAiNo8Q7886YBNEpjMmeLGjP0NH5OqpI0R4+wv
c+v66jo0ej2uaybthQSqrPtAjmaKmtdhKnoSct3yBTZTvHhZeMJUDoLh/jCdCqjS
o0ejpsByXgDgXlJCOxBurUnAKtaUxkTH7Xaw0SRywGzDAcJHCyxVWfizbNuOMiI8
6bK2n1HKtWj03+5NQp2Pg5tHXV4/vKk5jIFWCOIK3snOnvjIpZxASg4EoO+TsX+/
YJ6Tzr+SHaiVQTpAX0/r9gfghqsmH6M4fkJiqGsrq7u7wb873/A+fW05394ty7Fr
01EzyBjDHwyJwH4B0Xbhux/f8TJWg9dSqBFDOaoD2pBXcgL5PilDzqdzA01qGaq5
PZ9GarMY27StaQipEqvdzvZnQKg59qj/Unn+HEMDc5H4MFDROXyaAMM71ViQqN3k
`protect END_PROTECTED
