`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tFk5Rmzf2s4kfEUfbhA4HvNOEO4l/FSqWs5+OZZgHmyBOnK4umXB0sOeBoxSabhN
BA58QvkYFwZeW1gr5K0cNhBH/TxT/z9cY9j8Q9OXhAbxlh2jUdRP+0v4APIEt3o+
/l1DOw7iAhyYp4bgdvECb6t46qmOUM1ufQV9DMaJMuGujrKAzyXcHUn/lIZCcfDL
9cvnXtEqqzZRCgGKoCduqlZvrteJvwE86RPDOqjaTq8l7vU4x383gW/DVibkK/HW
cntiqcptqGD1U5GxUBVPuICbTjnax0heDT/PaP1tXCLDyoYQ1GLKplawEZX8Co1C
PkDcXqnslwbfTIreiDNn6vHQcnF6opYOwStIRYvM9btQg1kfeSQ49LAT9MiuVMoT
bMJrKu1ydNanecGEMxtCyaMd1MYlGsBRd5ExasI4/o+ddlASvi6M2E1266nmz1P7
PZglpe5J0pFqdkvuo2Khrpqx/UZ0pxpcXCMiYNC528fzayO/ySdym1CQylZfA3M5
dhz9kn+2B12Zd0kj22fA66CoH/WmYql926OOkUtUvaNhDAhlGmd76UeyXdEGC/a4
TJohVZuMQvN7Pi9oFBG8LZ4bxA0JNpxUVg8PF/tizdr8YHEzvynItB+NQazNIugN
F/iRD3Tl/SbK+zxgV0vywuROnenV/hLTE6L87O2+swxNWUM0FlmrOepx3iBCu+h8
iejbboAT/yZlZ55CYwboEJnVNOPsENJ32yoV3y0Xgrjvl0CuFKos6QzQvAMzUfiL
NKKcomqiDkr2CR2hUymmTJA+ev+05g5XWcpJKdizvyZMXTMWu+C5XpzwqJmxKsom
qvGF+gg+ckNJIrqyMpcyRDxvkTqClm7J26FltPZ+DmQAPpslCshFyMC+16/V80cT
fubrG612g2/8sT0QkhPD1EHne+pfUU8rKSNQjDbTFLJoCnx1MK0omfnMxPcmzgA1
BKGfba0jx3daGEkOEIwwcO8S3rqKG4/B5uQ9KFz1aLI3zI/F2DHDs9XOZlyaNiDD
W4hr1UYWTujJzHjGI6NYen5i3KLOFxRk1iWOFGk3HAT19gl554nKxItlKGm1CRVF
REfm83XBLloeSq4X4U8bKjINwartv5Zae55s3gg8n/f5AaXK2Lxi7OHNny3zh0Wl
urJ+qlAnFQrqNWvwbNPiZwMShX5SYG3sN/ll/jm5doSwthm70mQQm1ey5ywlcDd0
7GEpoEXnphOsZ9wsfGK6mBaf9C8fpxxb8uY8+J5j/DTC/IS3Sb23x4ZuwM0FGj9I
YfqjmODpcSKTDIUJNRd6TkZhIDZzPeTDxGCYYo3UOhFWyxYxDg1Q18Il1IqPmjOV
MnN0r2KYELkFrgBA1kVPDkKIIHknzgMViEk3m+B7GtsdWx2lAAjC5h9KzQW3Md1X
jecwlNuxyg5VxebLLC+wz42tMhdTBi5oGGtFTCssfNW7AekrIDw/CpEAif9yKpXi
+tmutjZh+6mF0wjDOPHIZXC4gfgWBNS4QKn1tnRhT32F4Up8ukFYx7mVzWX7HutO
f61VE5WvUbNCiQUYrfqwbFMeL+qz/Jyui1GNt0W0lWopQL5fKtu7v183XqMyHXQu
yLyL8wYiUelfBhgarA+lCA+/iX/aLb1rNlbXNW6VNvFaOOm4n+Vfdjn6TfJMq10y
1zUrbqnnUOMs5mz5m7F8flcqzw7BGpLMze6dnr564TOa2ck+dxGL7TpmsSDje+yg
1OatX+wHcoa64naPXPqYcsJIqK9Ei2VoQPkbocAjS0TgPDfCI7jVXCEd8FRlNewR
lxbAf5H9gK0Vj8952J7OEn+XlMAis/gIfSZudSLozmMsSVGQZmrQenuWsrpxD5+0
8myzqf1w1+TDNHFlOskP90nEg7608/17U7I8QIo+TjFiU+zNqRpcrQEISN8sFKuC
Z+m+cydtebKEVeSDy513VaT2Rbknc6GqIZos9rB3AF0JIZ0put1xrpjFdBeNUn5b
WhnCDlErt1pyfbKOhUgZMLywCNR3Ef8+NG7kdA6g8of25Kn9u8RA0wP7QblEA+IZ
EE6a03EwBFVvTsYrg1hD3f1KqCKkfHJ6BR5wMB6OoAP3V4jQ5P92V8QnymKNu25e
mDIdvJd6tpT2wLsZV/o10Q==
`protect END_PROTECTED
