`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wUgGA/em3maxhc2VqDcFAfAoiI2dGNm2iNLt0aEJfa5t3rguOwkzJphoOhsAPHv9
HjfwYAWeNnmGSwd0cH+dXpWN/6M1wVJ7itJkSMfLL2hzDOMYErmNND8oOK3s1ds2
6uIg1RLm1Mx7hWVW+rWsRvjZ4U5OAdwxRaZbM1N26s7Rvfb6N42MiNcSlhGWve7w
tbH/2RW1tsEineejxTXNc6ep44+/35FzCHLoiDlg5iYIFPgfAu+i4CKBKhcS4EuF
kT41fCipMPDohfSyH2S0MSTEby5zeks41GfArBr3hredIY+WggZXEci2zrTzoNCw
Ya/i86uD5yMqFrapiW6lX+3lBMQp3pTZFUxNYkrq86LIwWtyRtAuc7qgXdZMXpCD
EtP71USFSYhP+U/sxGwJxPgs2pLOa/obpcickUMOhKJEjymYYzegppoDsMfxSIQW
1WnfA7nFJN0zkSE4sQX4JK4R+O7J1eDffWuDqLO01WakSeNk6d1UXhkR6p6qOthV
z53Xy8AyTbS8g2KXpxN6qgCYLdtCEa/rq+tozrGuSkJsaZVHNWzQB+Kvg/exF+2E
`protect END_PROTECTED
