`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rQLzcP5Ttq4c5THHDe9p///QJZLDM7tZowYDgeNYnRGQjGaT2TUl88q1w94ANcU3
2n+uPyQJTkbJrqaIwy3c7ac2tZp0A40iHSYFVGvJWdfRQKKC2VfoYWYDIpJME6kq
49Imswuhcde/FoRMBegu9OZ74T5dca4GzcS0lyaMPpvE2nJbzJY5qlm20MdqX3G2
B7sMdNKNoUqzorRz7x9V+z4Ew6DtXzi8Nt09DeZf1XjP7ooVe32vBTZ/3fbgXRcq
a5C5KZQ5RSFO/LE9/bGDX0PFjMcHGMGl15269qq+gMiao+esVXGqzKlUSrC3JiQh
/jGSPQmBhhRtH+v15yA4coKsdqYwrtcMXOjRkNoZ37evHLD13+8hgp3iEJQRIEqv
VOIiSGvpJjYObfqAECdrw5BIE5zA7WagGM49uIdI0UIcBWawb2/P+GiX/oompCuY
Z2pdEwNWXKXPsxq9z9suOT37+SpGYz2kctN5fzLX1UkJdf2d5Nuft3vmsm13fgAA
L/MvL46R0EJHLsewWOc0+z6E6a3xPmcGfYZPbpJjttmTiubrdjaCHXMynUKLeopD
3eCHw5aDmLywjibsqgmUDdVjwvYbD9godf83HT9HBv9mbdGXY1muTUI2zrZJXGbY
YoLIKhMj6/C6/0qobztuzjU6FuKGRRPEtBOEgy+HkWhuSHWl0K8Xsmx+qjzHWYCr
E4DfWyud9bBto76ByP+l9PnHCBgh1pI97Xx4Qno2fho3MgNtCCrXgurDA5yE66PS
SZIGtdGGCAz320fZRLg4h5ZPSCb8uy8vpgez2wy/+nGgu2SQ/E0577NpZQ950PrS
Xhk6BEi6rXlGjfXFz+DYeCatRnfYEjSNeUKBbbkyUg4xXcdUYjOTSdq753at8LN8
QTWNNCRKXjI364KaEcf4Ofy96gpkDFTKqxqy1vJaWrhRi2cpbUipAxBMEaKRZmz5
ZmWs0STJ5G4vqZElNSc+Rm5+bTndgY9HTWT56bYyv5oSY+HtHpzUJbNqqti0HktI
4auijjBEuG6xR09fcBc2mpOaWp2DCLc6koan/07N6CrjpX1z+hcPwmRuVI/Y3SsP
PzddPSuX2PldzVq+s0W6FqG+PLYvpoAK/M+7LQkkQB2SBNci6CLwWF8oTcsYKXhi
CiN5S5EcHl9LfgXqiBw41L0ck7rxSFTOBtsCyo4euEMp7IHB2i4fEM7guCsdWL3c
2gfCHgu76JzUc8treuiOS32YFembxoqZeyMmhjSRd6vTs2bJsyZN++ZEcTebOvbK
KY/cR8jwGIU7BcYFXXO6HuCdkCGz4Q22F5hPDXuB48BkxIpncmNRj+INezSJkI5f
rkmnvvwM9muakf0Johvaspiui8y3UwM/I8bEAvIuGrHN2bav+18NzBw8/bcgXyS3
dDcjHhobLSZfrxzQVRqj44jWXgW3NzaZw/5t7qk2IfM9tZd2wbgFdI+sGI8W4pVT
S1GkLGUu4u6bHjn6viIpz9vywVYa0DYPvEVlO45g1CcquoA6UsIF/dfuhxEi8z+N
0pfGcrzt5r1cPyzvkIZZuxfC5No0Ee9bwHYGNWhtafLDemAIffECEuNDHLceXAJc
8kslsEqCq3StoEv7qk/KL35JzQgxb3o++dTeJNUScHQLnusNzJF5+qtuvkC3fmi2
3AeJucY2EvS0fgzysZWlSpN2nzHOWYusWZQ1KRtwN+lj4Zbc3C4lp0TcZ0cUWqYV
tlg1MUGh5hT/iiUDxGMG/gawWz8ALYixAO0NjjTE2tRjUuZXomasfnJcUK9ftCC5
xHjaEoI2FPZrX6XZN+kBRu+1zk3/IBDwlLtldvCRCBZp9daDgTHKowMiLjT5spfw
KqAl1RmCxaT+UA7f+7pVtygpJHiEwzNy3TEcl9uZohhhnq1UFEJl5r2PeWYEDTTd
UNcYEFCA3pm7hCMbrqnc+MNND39GI+9qiafbBdfNkTmOsg/VNZnAEiarU4MstiUX
/7ciP380kI1PDXTBvOeTKmVMzvVSiHHsngycXx0GRmf+J5hSj0nOEsAvwzgwcCOq
3Ek2rTkO9wkwI4475fk0crmxDHa0FAemZQoPT0Ub9TeRuQW9+Gi/q1H4BjMr7qiV
jhBIGrkvTJVaZ/M2Y/HKXW8N+N50qv+/BuihhW/zDfYwrTnwOTA4afuvbqMmUKsE
J951NYKfYkVkfofeS0Wq0VNB8NyXPC0+eCRHhrB5USdpXTW0SviySipU5mdcNpFm
ISDhbM/snew6kz3BDy+ZLl7GPKp1vrcGNaojQBXfZrYhDzAKq7nZRBczxvVOYd0H
qKZlHqfxUeXEnvKiUa7xNQYy8Lw0DrFtBqt3r8RNrb/AaG4LkYPuEXdGgE7acfk1
XSguOPCELVWsUeWT3cmG1SfinNIKH43bchBzLjs88kFMGiXq9dI8yTz+FX+V1sl0
5U3uX06TJdvz8sOi8HlO50WIKYcl8Q9kAoJlU62/n2tJcYrR5C++dmUHgmt+2wyv
EAzepXrGLp+kRMvPEjRoWEFN8xZaAIlcK1FJJUJluKqxQnNLX8RKItcpbFavuH3U
y+3WC4mXP2ngZT4bbvkQ88tVOjcvg2Jhnj4ocZ+m7b1st04enYv+9XOv6nlcHWcw
77HKisy5yxxzmMdAaYbpDOWKTpfO214BpUAr3rMDMJUbtX03bxLyB6RGJ9cf4D5q
hLdgxISDPFeocRfpqyk3nVPMCZjLyoHEJYmiIztUJP1wyhYdUFIPsgHOoofshJsT
yoCWIvkKfnVwI/5zCXoVaAMmPapW0cQx7xe0GO0w1ynKv4NnUKpxumY74JB1ro+4
RcDf4PHZ0UbOz1V8/1Ssx0bWCAdd75T1ZuqCrhAaX9nG69/tT3aqSDHIsob/U1OK
2kkSrmiXv/sj4YACABkd/4i9Wlk74sN0pAP++YedCnHifhB7PdT4IA4Hk1YnhPC3
dy+kal0mZ7CKu2FMc8VjTVhvVlkNZUTYrIRrR+5V/8avVDBT7btZgaUWLnHkL//p
YM1LG9ggDZ92bDzfugn/2cYc5ZlZQUXBrMu+zZeUafQS/DQ8gevgbxJ8dFzXBpJq
NvF/2l9Ob8KV7QVeLGRj+afw45kWkVa8lpITsnaKbPccr+wk5cItQJ3Vft+hvbWh
6IGcyXraoS0sNqMgL6HTR6O3LiFgOPcuAJEF2VWmS+fjLImDgz1bbUmzTWdBx+YG
6nAC/tENn6yg2T3Jqoj17kQxXgVae6q16Po5htHAXZlj/8zTmDkwZfsx/WCttOGk
hvsAsispNmJGrvSJL1tT3PR3xxoN74t82xjhDs0YIgm01prlC/3ybnI5E77gdPRx
rLDOdv3rK6f9ucCgYhnVB72qZOWQ1tKUqf0VQA9+pIkHym/qqBtP3kHvksOfQGl4
InlrToW2FXxkO9A3IjWrvihd3fq92F0bvsKeMYUNGXcjWx9j2IITNaPsIGTXx85H
s/4ccSI2Tqi7TRJdc+WqhCTM4VU0NK7rN/LWmt+9eKAY5cbOeA3FDQkWlhqx2WLt
HmV5gOgrLclFpPYPE9CSed+DaZxyZGOIX35+UFcup9wmr6ZwkOrHKTkwwf7SADYC
+lGFMhSarIJxI8vdgU6rjoW9aP4Dr6S34TiaggfVGTk94tFCSNB3xJxXA04J5cT4
ECHxoluq01PoZK2Bgz58CutbMmO9Y3VNzLfp5KmXJb5+cWmu0VVWZTc6OGfl570j
NAWuq2+YJsIH1kdQssGzlwtVR60+kFLbbYnBd/j2AAYfpMuHW7VuLfoZEyMW0DMj
DZVoAylNU0/KLhQqd8FxsbYfSwFVJ9tUnAKKhtsAdRLBWBVQWFLdUyRZacB1BiYU
CGwfwtay/UmnC5n09PuqWcRrd+MincPzZS6uxSlXM35xrodnSbVamiDh2QAP0E4k
gGRfP2y2kWPnwche6eh4AFbMazzTuYNsT2zya14AzZaLht9h6vzmyzuvHW/426up
6tVjWqhbJLUWCaEhCMJeRimzaZRuDT9DdvP24KRziX3FRLKLVDAb01vklWJU+xov
ZVdtebn6B7+RzKqUKhMhSmb+LekckgTq/QOS0DaZwsU3bN5okccg1TfEZUBXhYV6
4W/KryHj9v3BgqHtWfJ818FnDDqUwiK6vMjl+l0nzypViKnxngpGMQe8vUS6pvI7
Bkt75PCMk9p4+QnJQISf0xwGQra5coQOY1r2F+zjzmw/D2YLwrkUn6WDAp9CBw++
9HUaGQ9nD6zuIjeMlN8kTC6JfwSoMq9jFni26/rYtIGJXUaygLyUtDd6I1PmWTAS
JV12ajtNatrdgkaFoXsUlREuK915HfWK8ev5mHPtYiuHxCB+C6F66zaC0GloWBEe
QNtoOvZWBqFjDnoiqe6kMgsJZcOYpu5J8dLNLlfuvUYPw6/meXigFDGwMKr06UE1
+zAx2itLNOiNOty1lzxcjT/NC4Opvsve5vKxZWkQjqH24KdUsJRA+JPsCli/pw4x
jUT3DP5zc9EvD1voHkttLTHSkGBaoE99u2wFuJiLRAF6mltUbpK5rp4wf8UJlbYz
GPc8Guzl7sPbJjl1QixSRIqH9Zi7duXCNb6Z7Ig+9eA9TzPS5E/4OKHtOMo/PGHr
skK5Xtudhj19KMN9NHFX5sALB0yMvSkL3DMV4XAfea+zsub+33seesHJM0tm9xEG
ghDKJBFhuilJMJPmYsv3K42HL7TgczMmGXSmoR96W3Scr6os5SAC4lnRcGdXVd4o
Tthne3PVsFOW4foankgq1P3d5r5fgN1KUSw4VYS9Zo0API4UTBgAVmX3A/oVmfCy
LBY2ch75oyCco1G7ewRl1pq/dkP/7gQxwn1aCHL0Mven5CMOmDv8+p7sUo5oF3lj
koa7S2R8J676gV9nU365YYlKNStRM6zqIVabSA7rRCsnism75w2EmkLAI1XsPCY9
Viue4Wp5Ju8+OLCMw4ANPQBBCeyveoHj3yfuPnWgcTlQtvwHd/Ns0/REd5r9dgfo
4lLp23hcxehRN0OYyOUPr4o953/HnwiX9idjRaBS6qfL0E9TpC/3QGDjRZFI5dza
x1aduOuJnlZ6/ZcD01KnoxKiUoI+GqmN6Ujp9KjzCi/7FzwNbxvJ/LsPwOZmj32f
moiPt3iPjW9skX7+3t9CrwC/9OmuzDz5CUs0NyEzL8dbIWeOjk3j+V9ENw1zECGW
lMlV9jezM8bjcDKbgIQa6W5yqMoDVTjvroDsw+pxtLhotfmy52s7v7heAaPG5geu
ujkTOlTcWNzOPbZ85RTpCiEu/L2LeYTNPrkWsp30XDZaU07RssDXDFu/gSGgVkct
T09nXjChl+oIPqJjVcXPUVe8Ij+gVv86DKH7l88KZBY9yPZRMnyEeOgsFWswOKV8
9jkRkJPe5slwdAY645Uuc8+/jZ9FqdYtjkJ4hs+2seR0qPLMWk5DY/IGqoSGNu4V
TqoaIEGUOGqyNOQ8NrjlwCfqiily7Lim8QqWEQM4gi9ySzT/F+PTyRKzt10wOgCX
U5j3Z1vTtZxOXrgCYM3Kq3pyjJgb7TGIoqfTpBitq30zm7fImCOeH2799NTYoRu6
QL7q4AlhmvnylXTKASrkx5Em2626eZNkFEFhIDOlDQM9OpKZ5yWI0/T2hCpBOPhy
TTBe3DgQiYGVVW14VlaqXba5hZIPSDj6p4awL02T7jN1SFyZXIwvslG97PRRkVus
Nh0hyeK/JG1i0XZqKeMzkCBczdJVi7/XxOl3xFmijeMqyIlRL+5hG8ouEoP616w7
ixg1RuSmvlXJ+OiLYsMvg1NAJ3RjOHOghWRyAn+YToEJBBtTTCfrSDFwWf+ayHDr
ku1fbMwhtWi+Il8t6ed4UV45Uf7OukhKmUH7wfzGuHhD4iInSIpzsJ0W5ebqFAG6
uLbKF9wKhxfpxVxJ5+4G1ie+tvZcwdbIyLczEtIeQpC9IvJgbGEsWYJwoccA/bkk
zg6JOFfR1/Smuz9zkHzl1t78RR2oT6hmjysR/kxY3iRy79FudZbBYgTJNM/m2ZBJ
wfiDEcxZX86Y/DRydhJ3zL7rFBFvXB4mBuwvARhovppRZEsekVV/Zq1WPD+maCy5
cJn7PjF9NfE9LQUB6ULDggx9S5p2FprvUFkwjDjsfwx+FiARM+M2nIjp03/LU2ft
8ovcOjyxwEhlkCGqxsXkHjEoOxuFtWs6TFqOW5DG7JBEq0huSIIUOZ4mhsu2UfKS
fu85eTemPsR7/X92RzdBh+eMu74J2J7KqmwljHcn8LHhkGu4GpBM4f63o57jLBFI
DBMEGLX9efi4MDpL4dQ+NT3VtpF/bmwk+MHp+uOfwU7wgnnmdQ3I2iNBv1F8N9wm
74uij+G/WnaG5onZzGRPuoXoei3PzCUTxMt3Q48pplwh53eP5WSb2MZ9wTX2cKI6
hR5ZG7WGwA83EhLuvNGF2XbIeUaJNnZ7c9f1cUtklxvT91DL0iyuEQLPwhbBHu/T
l5BMP15zewhtb5VOFvHGy//b+29fkqKtVxM9jhyNbBIS+9bBI1FGu2mvPucE9kkk
TKBAwDlbU4OJtxcMb0WFwanxoFi7fqi+nk79uxz5R6fZXkSXhRjrEAtpotm+HhqJ
wsw6QVLx0ASMkrpmsHb+yn+W3caURmRThG7LNl/soviRljtR+gITtmGHyJr4fLT7
ciomT0LFyuPUfgMSqEx63ayYMbQeC8gZXJpSg52E9OOm/RFkjM7uyCkMlD/ceh9Y
EIXEKXlmh3QO2ZhTTKP8+pJS6AiECvzWCZFlzJaE3EEsX+O2SNkfSZ0CiIUrzS+A
aFqepgUMewbueX2WVB1bhY2SlSm+8mcDmfzCA++bIHG4F1Npqv1ZKJAyRq/0XDIe
dUuqGr4OIxIv5U3qqbOkIV1+YJav0XiioeSOT8tZyrkw5DPBVYpb5CBlta71ykDG
qS5F7PGHW4/Jacq5h8ZwE8k7ioxmtQqSgLRoUFDVDJC12xJDIGNMyJlJ2CXqHoxK
KVWUchtLoKK0t49bqWA7SFuDgEj9stEI9gkHYvc1Ol4zvWFXETQYEhA0t+mslo0V
Wt7iJPc+mZFNe89u9EUqd1aQGblg2MelV+Smz42oV3f0vXU8B9LgxmMBTUXmcytb
xXCYp/v5nXrp66wH5KzWXn38jl2uUC6dQ6GD9R6PyIv1tkf4qNUbDDLxi+FXIe/w
F9hU3UAb44k+0BSCePbSM41mA629beeiYG2DGN7h9E8k+eClD8WeLmM5qcCUcj+0
g1HV+Mj9QKtrbyRDDmOYbNODBNzESlGojLi/6NqC6kpp56l3G8Kj9k63PS8/cwEf
tmWWsfQ0VxCXx22uDz8o1Pwz3DwEhzDQUHG0J/pvLqv4byklZsZCbXMQH/b9Qalh
gJhjR8QefSVVWrj9tFgKMvEW52dVF7WaNFslgTzoejRbZTw2ZkQpdHieNod9PsBn
kXhxAGjn45AOCFXx+CtKgYEX30SSUDZyaxS3eJVP1FFDWhR/CVEb3Rgf2NZ20f/q
FFjqXVX29yfSQvc1KReFva83q4gcy24Y4Ur29UC5b39PSVQXB89jGYY61nxYeJSZ
DgWSr9A1zX6DHPbKEbNZ1OjoLbRPhqcWCCSngHL1POyKLP0ErGo+7GsiM5FpeXbJ
6tsoDR7rHFQ1QpJc86sVb5QTF4gT4xKbBEtAewPIBOnvbewzpaehkK+OhRse+s7A
4VheNuCJIOA0VnVaJfrpWt+JxlQEVgRnkzg0MlP0JNPh8nA3CJu7mEKDjGYW+EDj
HMIMoRwjpsyDCgyQqYypnikFmAzun8K0CEwW275jN41scVU5OP3mLkHPdmqZWTbp
1dG8z7LkpPI14vzHL2orOgufVWPxAFCfkJYt9tqiOhOlibhBU078CzN11qS9n3cy
uZVUrIQhET7nTICIRUeSjLVxqyy3pvJZgBUIkrhioaSOrp6taDYkiqD5SQVUCQB3
AYcMo6/RJ9/eURJXh2fFZCmMxQoKUL2u/IfOtzNvCObVXJnpKBdjl1QCx56kcDrm
qlilpUZeyQbNamxZTNnmdz480yPHZD4X3Mo1/oXCNviqsnt2ttLOeGJs5b15mRt9
AuesvqhoDD7JoLaMpXk8wZdenwBhkQnL0n0k8SUSi1AngZcY8Qw6c5TsxEvboa9a
PDJ0xl/gjWEe279fMlT7Tk9O++6s6CXBZr1GPwW8wTmAUr6PGnaAjaV1Opc6bNTz
N395Q2EedpZdVzi3FYMwoggR+L8mj/g0Fbb3F3hsVBwvT0R8whednRUCKwgO0wHY
klbBUhHbFVMCrjF1YXJABPaqiiTaKUqzrGWhFIB5Y0xBcxPPe8hITvPM+A9E7+eu
dIAauXwipi20caNMOICqfAT39EUPRX2+UWFEGYdZuhpiQSiB5be+e4GeiV9QJTHE
XPJAl6ZOdZmAncMj+qESW1vpOgIncrxGBKmiYtFC1CYQsdTf3n0y/VntN773+J4P
6/XB2Mb1NG2tJRzIEGxLGWFh+a+xhTcilA+WqmpVruNGPAad7ZZIqRdqtcMte0/E
mAHvwLSCmihQYCmiZWT9mgrpy4rbudQLknbadbNLy3/gXY/BQ27pUDTBeY66tvJC
ky/VlHMyUqSJU9a504WUBv3JCI00MTvDT3f5VE5Q4cBzJdIIrmCAJxnGWdeDhgoE
eKwo6r14muPLq2HAdrb47wOAdq14nyClYj5Tu+EakkAgBqgww/2WypqfmPVx4Uhr
8P850KsODlxOdgctunDPJ2IU5QQnOKE5+w4akM9APU+5OzE49063PEss8diA5Z/D
upS7ftFRlZdq67LraxXk1tJ4kk+Fl2WBbCxD0g2Aie6m5dcr+di/YS3lMrfakZkd
e7XGiAoP8kgoP0KEaNAte0XzyJKLzJ4ZLDIKqkm8w/gXq2IeZ2aA18dYhDyVx4nD
cjtLEbiMeKjcLUNioee8LG7HCBQzSczspIbPz4kUkW1YVuP0nrspcFjY6IYpDcWT
4O/5OMmFORNQNmNSUJy0yIzPmYrHhKSYXskSsN3ede0vCRFlgl2+A14Oq34kmtfQ
u/9RSxgbJp/VQ8DKRmG92J1EW+kKvml+XiHHZdA7HHj4eSw8Pa5gTIsqIf1ZJWFv
udRQYXzWNi5SsBnh+o7gCrrPC/dI+eeWZ0Hq2phJEyuu1Y8JZSRAaCSfMdJR936r
mP1TAVaeQJTKrWzxJQ+g8gYlKQVbJytyodxLU3l+mrUaYu304juWpLR6Lw8ChK3f
pqG1MyQ5HF2LgnkrKMIy6+ReGNsPmxcl46DWG67Dcbiw9GYz3wF20dc+qfcoUyaj
jiL+TH78FSWXhKDQsoQC+cjQbXOsB/H10ekITUvaCBIX8aOcMO7lKZXFK0dh3dgr
RRRV5OmuV20RefwIj/C+OkcEE8qEu8jEp8RPLJpCsaTF83fjHlAuAqahuvwt9iol
GO1FOA9H8ZKk6ZKqq0R0umQKRgcJY+DpJOzrtl9uYS4AUxsmRzxQaJ+GiZx/AcVX
+8qNPU4VCdYRdHlwQBAZ5nuVaEl7ZSX1L3PboJHg+2+eHdkTXG9FReUnHOZxl+NH
Vy2/XQ7cxpTZTZ9o96jpB6d918ABdD4WHkbavxhArnflINjXPYvApOEqAbgGSYgI
131oJ7yw7yYNbOibtJuD4ybFcr+V/vrCvlup7PVlX66jmlGcqMDAZAqzr6EW7CSR
WPm6GAJiUZ+6uancyd7FX8ZVoLuuX0e8Zr5tCMu79gDync5yG3dkZcIKll7JXFdA
SyGl09Bj1CT1VeiJbi2t5X/dNWTcyOFrfuOnsH7jHjgvzVIzjHh0T15tfCPtLPHK
rVyoWq4uqhMFC06hMOiqkVw6K4608Cyu6ueJFD+R59qMaRU6O/W9fZl6b6sGu4z9
OQ7RixeB/Go+/xFIaikXGwpTx6rtQAf9hunT9btAUZ5qZP75Z6xLyF1Bfyzt7a+0
Sius/N1KNpoN8i50xBbiEoJDeZ3esPVK8ZsaPYDIuUgKqp4fmWJT+8+A66XUJduY
Scc+P4/Q/U8lcFJ3IsxzH+/TZhdN+Fg+IIooYdfrScRp+rNAmkmYk3FZBt04BMR3
lfXo/Y4EXWTqfamfvg+dgl+GGJxqgZQwHTlZa8N9Ez4RRRRHyyKTZNeLBMpynRp5
+jaOs9ZBe0vn1rIoVhBl2ioVlNmxOaQLQKdQHFm0yn9xvztx+tyHwhCKDWHJ4dUu
Eqjamtf5IEW3+kAPTCWgXyDLdT/owUxxOY4YTymT7aAvVacSc3/ZX2klO0wZpDll
xAP7+rMZZ7uWwyJS3ndybd8lL0gKBCCgVKu9XwRLGtgfyi+u4BAsAsVDiCIx2afQ
LnfKDbEIKhEB5kIYE3QT7UAdgXLqmn7p3lEpz1fFPFfUFuBO8jThyvcUkWUZStqE
vWRdVewmOOchgiIwe5h8Fr58bCbw3oXj5PqiobnTjeOd+qd7h5DKIitVKFMjuYlP
3PLnT5noiQyZYPeW9MQj28tLeXbUjGb9gYfjiC+vH59KEt/vA1GRycmeTgGr41ka
pfSqBhAqh6wepXxtzAkUMTHS8+azN2h/a0ZwwBx+VClAjDYZRrej4oorJe3nrPU7
4VVDILfNR+5j7uq2xafYn/9ab8rRc7hXa/r+kSnNiuVB347Wy0MjBvKtHWqcDFW7
DMROSoPI47+mIyqjRfBr00X5N7Nqjggl1y6I2WXjhldtI6EIJJd4WmhiV4+9xsAi
s2Rxjq8zICW9iUPaq7k6gi1PjABeM9NnbwrymngPS7B65MBh0eiCxssOVo5zQcQ9
qijUjfoNMuhR6r0XnwkUaUorXHxMSYQ/6ZEElPOVC5MEuCzcs1kbyHeKEo1MCEmv
YfGtpsMF8+9FHULv0WzM8UtS6KhgTRji8y0NFesr6UHz1mfpy3CtVYRFCbkaHBgj
HGKegLgWs7OXjW9W4/POlZjxS8dw7xP0vL0S+ElxGyvlltL+5oGEa06GXVyauBP2
nTCRqZ6sovYbDfaKu0ZpMmD8Oqf+zdOCziDF98pt8ot5OdP3oAGGD77raY8rOEMW
7XWP4xyZiM6pxjTwdiBOOu2s+sQmlIydouCqmLOltMi/o63UgJyMnST3z3DG0D58
p4pfJw4G479yCcRnAJz2Y8GrZrDqnxe0McFqdKUUPI/SqmlMpYJhZq5iDBCWOFcH
sYTqLkj5hEPYOz3Cg+n+4JrvejaMHPw8Q9C5ImrgL+ECwi3PVc/IeLBo8ClyxfCy
kTWeLzrydjdtN3wdBKTr1gf+yt8cIoogMeBFbUfO9TuPeTLwdDY56e5Vf5xLvm/w
mYaJKZWIejDBFAePV4KFY2FeMYcGxa6QIO2OfgWrMyZAjlRn4xrsTKhdHqyr4HG2
oj5DERPqUID0XNm+Y8aqoC6Gb6QtRKElFcwrL8VxbMxEMoLWfpP6PU8YXsH4/s+U
IzwVUxUDkjPNb6nrGKw4vn+KkDsTJ6k9ibG1iNjwSh1Ot/PlGhJ23ot40b24+eBM
NDnME25NZQv2UDjX0iveYTJV7EZLWZydrxXDgfNt4yEkAo4yUW8qPN2FFaogcaeo
+Y+lUWKaKc5HusBnhd2NEkMVL/GoS4w9cIJi3kmTo+TjTaxr3g9gNuhAhJG5Rk+8
xh4zCFWWTIm1zbbv2kDpvkuffef2cjvHB4N5Z0YaRQjBrZhvIaYFibC1cV3roAEC
+9t5pP3rGCHJY8IvFqbAPLOB1MbjciPaVypbJi5n+N6L4R0KuZ0E315TdjiWmADC
aMBEUHsJPtTyMvdZetZjchQ+Dq/EOGS7d7LZEHvVLew4pdJrKtufS0NzfB4YEZY8
PzL62/oTFl5W5+DmvvaEOHKqjLxGAQ2pHM5Hwfpb7UdW9M1CSLovxmFy6h4WoLNT
ogSdTVVBKuE0QhEnFgWlpAtx6Lt72tPDkT3nYB5nIQkRsqzaelULp46p8h4116rm
ako8fib+Mg44vSop7rf8G8ziI7LqrmxBJKIrzZ/ksmFSRgFOLIaEjkzTrPj9hMHj
HR8EG2QysoHhhoeEeM5b4CT9sXFCxqpGiSepPJ3zOODmlcNBHn8ARp4MBbxtdmxO
a2sySij/HB1MknXsd81KHUaclMC3MqTbgy5OJhuQF0IVjK6sAsw5Er1/PmXmDMA/
qIhjkl/7yriH+DSL9ykwp02YGrwY565un4gXp+ezM/LZc8/vcKxD2qmaK50D47tr
Wk0fQIQJepFgdPdwRsOCEFla9opgkG6HoZfNfS0FhObUVrIATTwgH2lI90PpPWUY
57vGaMc4ecCkC5nrdA8DzvX/8ul6prvcMD18Nsp67IzTFk/iotSNzVV3FafrdCCv
TGNX4XNYKtqOAJ6KxA4xC6CVo3SCVuDkAf/G4spSRhWhiKl/oV32aMHCagWiPpG0
uxh32EXJchLaa+VDtaHY0fQzvSZ/vBzJIhwE9Zh86b9Oq9CkD6cnTN9QWtqRwkel
G6dWAidOQUWnzum5DhGaWa4EgKIovu65Wh6I/ZTPOLW3KnC437WT4Mb7zAhJjKA9
qFjjFLnAM1hn6Mj9+u2aebDOMkr76ogNaR8LObKB8/r3DZk278vG/pCUQMD3r2BY
TwnQvDRbz9DecemEYdD4FtvRaoG14Uqtf4aeqoVEHYGKHXzc3nEOnV3YhUokC3PJ
N52j2CeHm0VWP3InzHj5gftsfO4F9B/Xl+eiN65e1f9oYL39RHCyMORqCjYsm1m+
NGMrqZl1oTLdoafw1JsrXUkkHIdItm+nuPrrsPpBqFsJbo/TrUinQP8AK+UvAvqU
xiDBMdL9Ly3jxOf3pWTnQ0DnPf+0GMu0dKmFyMSgw0rY/LiokhvjdFcPWHhK1C71
EClcrNUaVXvfJ0nEycXg/rrAnocyngiakbWWpYrw8T24keVwv6l8c7n+P+Xdl7/u
72vaAUh9DaPN2rbFFLhqxkcgj7bEeZzRmbBLvwHeUimxJKp9fkDVHXuwlaTD4CvL
jcigdPVY0t3CzuhcTmU4/g8uIuMFZoXaxCYWLoP2z9omZzyVuUoUYjIsQD3B+qp3
Jr4DYUDkzmU7UGDDIqBpsYqkrZSHn6tH+TrKDgcZDsjYf6FYmpDTBeJZkwnS8dzR
rhSMiOQZwm4YZxpftLPBzgocuJdwTr1rn73/mi9LI+bXJLVQdGyOxvzLhq8/FesF
LqN2JanpTTfUiHOiXspKTvzAkk78IAaLA4NBjlE9BC7pJvltO9gLls2VzILLsViG
/qfRhFIIJaJEcEVhwkmyrMxOevrTcnMnednQo24II0FUnMM9oYXdWVXcSfAEHSyX
3HrPPEkFZBzvHy64rQIaakqE8BA29hnNR2kLjZmXHMuKjYnibJLFyg/iiEf59ehj
vZ1Xlfa7hHd9CqF32i12s+hSwBWRECVOUbcpt7565TBwG0ZQnprEU/wpl678zWgp
58ruNywKlW6MLXTte00/tpdenT27i/P9CrZ6/LjYtZ+e/gd1c+kOFFjl3O/IhGLA
sis6WaJhmQ7sr57mNB+21elvem/vJ4SDK7vhEeDnwqivAUyPhXjFTFrmnzwF3Zkm
rFQZlZXT6npFntUQN66hTePaCJwoqLAWBZuNBO/gDU4pau8mw/i6viU9xmnK4MRv
dpwaxcc6+f0fcjvbtYaN9YW+rmeAgpiP6FOxSXAxp2mAMYIm6tnZEXsKWfQkl4lC
tFFoZDZk/UJBrh8LXBUhboxri7H4hRhB/Lt/TR8ew1kcaKEaE7Fwzcctxnla5nhN
o2JB0RzCFoOxhR9PifnsDq8adOUApcwq2Urx8Dzp2kK4cAXrHjlbme0uGx1JLjG8
mnGIhKYL8Kz8oLVCnlhryw1VMk2t9TNfmnnVH1ISIqB91TyZntWbITQOR2GiMN7+
4S90GCaBTDngV46EYdGKyJEfbX/LqAwBoRDFmSfBeWq4RPtIrUPV/DpjV5kGMb1O
AhEPwOXwbs/yeuSElPdh3y3g8zTksPlUY+BczWQeeHP9q7sG8+E0B1Gr5Bn6Xz4c
v6M92mLXCqRz++tLujQw2Tx5CDVnjNGUj9GGOVb09mPhVuLyII9yMVIRhFv1WTz4
LgqM3vNgZnwIaMKWGO49+liAkZUmT4lhDWU3eHkzrJ8aMbTq+zDUd8bnkjh2cXsV
492/uuvpFpnmqwn3mymHUrnRuY+UTsRhi4vKkVA/Rf8xjp0nm7d+U+aZIf8acf5J
K0+Q4z1FDUSdoHp86lIbBc/xHp65mDh+c438OsApEjK5CQzxLulcABPgiFaT2NWQ
9xS6cOAIfUZpePtuBGyiQAu5jtkRq0apDQ8EOhURtw/u8WGr/X2o0PWK5NTitZf9
KR7GfJpkSh5IwvYdmMdoukUeEuw8wn7qn/dZ8WeumLFSgst/r5Hv6x3JZYVdCN4b
IWRKf29SwtSWzsQYBWYAibG/TqrBHHa072ydUjg6tExOmH1Ywyixl4ezgw3sdfNC
nfS5S0ZenizMAmDPR2IhSV7SwMkKx52ON/99E0uXxPTmSMLpXjtUNLZKwxeRLEKp
FkjtMeKucEmxCtxCJY3208iNxLxogpAHOqjirLgvIg973WYEWNMfl+vmnrGAd0i2
RcsBIDTQy7FHMTeqStYWgpOv8qoT4z9ZhzLeOceSikexnUjhVKzqS9CLENyJukgO
VaOfaXhsKS/tRGLgAerEoKwNgkaysTiRiGVM41EWNULR3R0JdPIvmrvBm2xUCyGv
hfA2+HGuUVzSeMV03Q/G8pbOqBdbuOCygFGsdTU6Lk4Wwm2uDipQfaJLrn3Qi4UH
`protect END_PROTECTED
