`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qNJW5OHZdCo8ELjDGtERsZiQhkoaCArYbWzCpF3MI7nNNqycEmrsC7e4ewVYRT5x
OHjQnHfyK2A+wsI3RClD2m1Xttgw3kuvcQccObc4v+WEHXYr2P1K1LtWmLExyQmQ
LeNTnLZuA3WpdlhXy7N+VDA8ZlUYp0elssJA4dV/jv8lJ2ADAVtNescSayxUmY0A
dAZSjZH2Im2Qvd6F+sYAZj0mFbCOCFKKx2IUtu4apM2po8/D4poaEKbw79Skz6dd
CI/yQ9Rtevf0b3asvAriGlxVPuBFVk6A2V7nvxtDo4x1Q2LIAVg+pdBdIvYg6OaT
39YSWwqt7lmjfOSyjTgNIwISyO8tiL9qJ5h8xM/IWW6uwtj2wJm7PdK/kyHVh+ht
2pcrmmJEwnLx/jiJMGseQq2kaf63NDUZ1dgTDLaWEIah/NoIr0Onba+Z48tlqZED
pJKx8HRYlBKs26TowEMA+cixFeUV6+WLIV8Ko8CHoKI7DaXVJpgLVg+TPQAx9HhS
r69nyv/BCJ+9nfVI5ODFtBajUBxOQczfHF+owiPgEytwA7FcRChtRFVvAiPKfonR
uauRpZTjx/bs1CxSTcTLNDa95sT9XKWPzfA+fqTgfwVCBgpwhVsO3iWtFLoCKH0H
bOpYITDXQbhFZNHr2UL9955RvO9D+yHpKIvrljw2CBlXycf9mcL3QvHqMEogkPHV
QGhtOnatG8oC6Q5kV2NXJM0oaQjK8cVZ8V6AJWC3szj0hHKnrTouUYb5TYW93Kyq
3HPZSfyWFhZ1wN5XtA/4CKL0c6jaam/+zY8w2KKGOTOfYmpRTw/8vWZi6yloOd51
k7bWnKzFXsvbYArfQBB2NcDr6Dgn6k5uXAFiuME1bX88c+w+z4tauVYu70Y92RvD
Gz4duCUno1nlscavbt2yfS9ggrURvrUCA2vV1LnWwBtdXP5R+DzqTX5IC+bsk3VN
en6FR7D6nSmhn+mr4jk+ysDYn+SduDGwplIzKaLbI8CvRfPGD5ZtSX094nzrbjm+
1mmiFgj8d9cihSQz0JNwZIum4Yec6f1dIgpwowHM1Gi1GZwYpYIPcJWHuDGABT5I
sTwnoha0qZTZ26YYPANMw+g26AyfSNy3/en6RzNUitv+/qWz60LyDlM37v8JaWq/
22Um14wDU+nQG59sHQD6AUXxoMGvNYkl//OocR7xWNXKpX6a1Rvz9VwO5xtQx3gl
ah70TQVXI6uPydCTS3NjLw==
`protect END_PROTECTED
