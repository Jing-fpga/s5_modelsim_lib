`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kHRtYlwci3R3esbk/BH660EfVrTbf404haaugC4yQbbKHJ2SAjeoIgrypB5cX+v/
KzUPm2IIFlPaMLvlHDL2c1Wxr8OFOP9DLjug5IwjNxtcABq7VSd33eamRN1ezwPX
yVeeoP4bD0ct4+qAnqoNY5CVTt4kJ65L3iWE+14uoDYpCv9CCi+Hvr+4wbHuA+Sp
EByV+8c9uZeRtyxOG4vXAmER2w+Su98Hq0DcQBiBDMIYY7vXmhXofXMBZ10m25L4
DlXYOaKi0HmETadCVgSGHyV7QT9Qeq8qqryhhujI/ExI/nTKv9d09kq2uASKZtDt
bOf0rzLbiL+IBC1wxyGqFLJEZgtThn1poWnWtNlZrj3eGYnoD0WujyI9a/sC9t1Z
nc3DvLBMyPAp7zFBgl78g9PRRTrb4W/HpKkb/38DAFsoHanU/a1+1MsnSScDCnA9
ssWWkjveZTtiwSDlSjU5lJIwrvB15lSU/x7U5JpO086/9UeRl3N5aCnxvUbz+SZc
ere6ajRqrKsL554sSIUhnmIEHmVoDWwlHw0yWLLSCMRhaVwbCnePUgY3BL2kmiI0
isnU9rf2gs3Tz8Hm+vQT+5tojbBQguaVRI/M6ioqxGzZVuqswR3TvA4rivafNF9a
lPBHzUgXNpjepXZUoERJd6+hmcKcR9jhUdkGC76uBxVz/AulZ2Q48Mlx27SPkNM+
N1MeUanzpKQaM+dJSgaw9JyoxluNreKj6k2jsxq4VN5oeOPCcWJt4ZSo0Xrh2yR+
MFI5sJEXu0FidRkz2YPOcrh62+vLSH4UkxFNsZVxKw1bmXYy6hQuJetlS6B3SlEA
N3kgq64LS76jpJBMiG0iH5hkcR0ajbZ3HGGrzVn/tO7hrSxthhpJ8p712uL5D0PC
d3JEdCANgTSA6DHmhYDspY7CIFObgLi29ssKc38/eNvy7DjvvhYQrE/egfCfHxN7
22Qm5JUO1i9eGH62HjxSD7gx5iDsYQl0akD6VTyDju/MX0cSfXi9ZRiXJJh24HrB
iHNxye6vb0O2kdpy4NTv6nM659X/mS8RKO1kBI/0sZzqxkXlq6ZnJ/mkCi9MFWY/
tzPRl6DRow055Wft4yxVQtKyNItuAioUSgKi3p2Dw6hghRGtF7yNIglu/mwsX76T
ROtxSYWcySocYQJ4c6fMT89GFfwZTYqTnBw294mQWKTY7Pi7CZks+NdwjA6DemMW
6ZPlbkjeaB+MmuYnm1ar5g==
`protect END_PROTECTED
