`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6vgAUNMUnxwbKRxpIDmMMlxmd+5U4RAFC3zPy3e1AIsNYH2aojb0Cbx9pSoVKPb2
ea5Vdy0fdxV+nvULe3C6ZoU64jsfLLHD8usr+KT5QkXX489iQfbcjGzvuh5dweDf
FDxwaDbDJQmRaW7lPHZFVhUCFq/L1y5L/U3toj9ncRqqSdKx+GojRGgrSNKrBzE1
j6BSNjGYp7iMt6GA7R7qDud9px2gfwhTxL2J3SEazCTTttOLPq7kIe9IddwJOxu1
wEogbgvWD9lI861bYx6jLDbmYCYXX4cGR+8gazxxTHLzn5iVHrTwJirhZg1gqB+u
OtUPNlbC+mmFxRm/vehdY6K/+3vMkI1SEbbwznUg+dkhfjKd0Ib2aR6mWWu3OR8Y
kaDDU3diNwZdWLvhZVERcyOSDx1wYodENb69KgWstEHgR1tNF7LW7brpU/vKk79O
t049tBqH6MP1wDDrT2ERgE61EzJUxa7m1gY1uzcrmjlNKEaUR1KoN5mRM9ZEe44U
OsebrBqaotF+vqi51t9yz2A13YfrI/1345nIoLdbz0MAtZZkNRsyuTbCYa99S9Ad
kzQqGbIcTSrFw40AZQHB1M77IK4EAyUi9UoYakw+NIVsc/WjIRegFxhYz88Q9WCk
aeCoq5JNXab3ZgqymY96oOBXX2Cy7CXStj5Bu+HyyY6thnR/TZCuLBrftDUKQBJL
EXurlRzKR4xXigA1xL3j9UJKljCQYJWIpLOm8dxuoyWT9L6wZn0fQe7eToLn6vnL
oxvqY70iCEUI/nRxMircCPm8+L+XensCJPL3F9EypXdWhsz2LnMlXZqDjiUKOEV1
KrO0dGsHisCf1V9PkPXh8Y/BEHY844oRE2rLDivii6LthMEeiyys8skkT1xiZ+j0
Giq2LhLEt464v+E6yB1glYbR5YP55gYOlqXnp2hBSI1CP0t7yXwdj1Wxjh9X0VQF
raJkmdX18pzDt8E268v/jhcsd5ZZb9hkhe8/hSOWNMx4Gj8U0+G6LE5hDYvWuu2t
X2QK0HBIVkAVpI/zTO1yytN9OhIfp7xn+QBAzvxSKf+spARpdtjxXTjkDX1hcugx
TDOETnQsK/JS+yeUprNZPgPM/Y4pPk2sqpyb/TNRM1oeSr+raF2F/rqh4FDUdWtv
40hByCt5zjLeJMLxhwBrkIF9PvFGwkB2YxyyBR6s/VjBGGbiHRRbsBXxORmW31UP
uTbryNxut6Maklyghe6ATCsp0B1hSbZAzbFSs+q9BUxsNcvXv+xInt/64G0ybJpz
KS4WrlR6zHvyO+ZqbIi/GK0K79FrCo3z4ej0XymrW2LRNQpO6C873Sg9WfWhkOd+
RP9EYhha1haqKTDNBuR1eXZ4FVq0XldNWUQlroT9BRGh5kVrmEzfiTLPaqze58Zg
9gwj+3yVTh2hu/yBPfgnSSNey195UNhSJo28NpSsxaD5XSLUbtJhHm2dO6cUdPcU
UOQn9lsg6PyL/yojLDDzMk0i6ce+mjbpsbbCqedjJj+0VC31wPj5jbBWoqzMUuuZ
D+/cwZkhi+NotYTpU69I8U54pI2/IRG2fuBA8k3eSPBJAiUfGrK16omjCU59lwZL
CILPHfwkpLs3RGwRGjPRYbcROIyki3MDcPXSDFP80j8CxR47+Gbb+f3Eff6G+1Fa
MylLawN/qrQtaITPWjIGnKn6fRGluK++XQ8kPKdZSJFW1x5l51xsNohgJQdeN3UZ
VPV2U0wjuOiuiukTtXwAii2AqmnXzsR38I7ebi7TqjN04B5sq+IVeJ8zXQj05Qs/
nk9n02lFeeg89ms5gcmypZt/L27nIWQhkHEiaBd/uw8NISPiAgXs6XhBGI9xVh5a
t/MsjzCj8IwGiH5/1MPkGwMbgChfaD5uROEOQfJFc98Ao4ZxOgf9Iztjd1ypawjt
4wQBnTL+1ka0YlosADLuh8nL9VPc5xOWAfgtR7dhItPmmdBXEytPmLp2q6Q5NUit
fKurky8tIGEe2znsDrW08mSj2lEXXL0xICeJE+7qjQwjlbSiRDUE8Vi9y6HKk55s
BG7KsBdNI3rsTjbSryC1jPcXddDoCpAeKbdZx4CBofjjTxJXho0KqJMLEJEr95Su
zEwEbUYhhSyugk5X+BhmMqkBprX8E03gSOIBoi6XdiS3KSpStbmjw3oBBnZuQILP
sRhAwbKxLCXg/q9rtvO1yRPbfHW3odq0cE46yJMrz9PY06oRGgGmmGzZHgtXGm8H
6tignMhlu5sWAnr7JcrXZX0LolwWKKHiqrqRerhEN8As4jVV3LTcRJnN6wEp4m8n
FnpAW34B213i6kq1+Z+4zuHrm5Z+YCZyvfucd6dlKwvZr4ngMTq6qJtda2iOnARy
yxnn0/Jv8s8QfKMb6XsrtEU1YIIyAzVlQGpzArcH4RcmoSHNdmBTH4z9fkiwWgNV
grHwVUU++6pU0hWWXVuhcY5I1Z7jO9SBfLX2XBDhCYWHgLbrkRWLylljk3GY6iYL
IyovMfFWh60L8ubBmLDvfGlGsn1M8shXYqs+3JuzUY/RzZHyfJtI68JGrZgxuBPV
TRCI0Rzw1gnIpv/U0WkMOIfTDlnRxJa2IFS28IzPQTC6Uzs2jfT0+AgwwBXhMxJL
TALh5KvlVKElFTeVY6UXjDf8TKDExQpKmxJ3vwMgBagBNKkNVLOQZd37Y2AkerZo
jwIq6HLSXVdqkBVKwokzJb+au+kvWL0J/40XDAspupNy9/+X9s6hv3nuzdh2YvlN
MSSyNXQSCBbWjClraCGK1xluhDvD4doR/RYjCPrNeGqgjww6oQfW+XWr4RYX5DqL
As8xX/EjkF44VJY7mzLk8sycvBHJ6zPfHMrIjCMdr544/Wsy3fTRemxU0n2u7ANo
0704TKuUmgMeHtHGQ/9amtQ+xAm8zaNAI1ADR56p327BcJ4yPuyEAc3uRvWH2qU6
oTgH0+OKArExTc+zTq+ptkZQi7QuggdowTj+FdkmAsRzdk52/qXYBHucT6nTWZCp
+P8BuPP6XyR6oUsHLOlsgEZhE/q3aM1/tx8XXaBqDUWgzAJUDctpeRO33hhken36
4Yeu/Rrwg5tqIlEuTqM2vQKu4tFOiadAOv63+GQdzgFDVi4ES4XbvyBJFKQcBL6K
HNFbzzNB+AKEF4X/ZLOZJsfNNFSHJVYiPbVeHd557rvVd9xk0SHAuKLJG2OhXyN1
DwlFokoBYO4wAMgbWYqTYos2+sxCxGNWncPbojYvcVj4xT+4Q9PJsSIqo4e71Q0N
K/m6qfOvOBYcwr/3t8OXQsOo91299oeri4hr4WihaZ8pQ7Udq6uBsKZxfmtMjves
9TiLvFNav/20KIWNVxB48WLHQePihtNfYvMeW5KUKNDSnujZf/tEsriMXcNIVLKR
g88vtcMV+XYZebUcX3JMUS/hjzE4uLg9GMPfaQz71EQB2HPo1qneBojXN1y/RT+G
M3sq6m+hT8rL2jZqn5dR9OlOOOeHCOUcaOIygetvAVbo8dq5tcHNpWfwMuv8/YQ5
3MJCLkfcI6k6hdF7RFLxhHPUS67SXn2vD42TUGHxtR4cbJ27DgkGX1qyucklh9o0
VuT/3oXcHu0rmy/hCCcAOQd6iAwV71d5ujZueRVGbTEqlOZoSAZ5c/fGyNxVwa4W
desyBqi2LbMSyo9iUR/+pA/zvNf/vN2x6qgDYCA1w2VJoYYeo/ObJbHJNeH/7BeA
37Yh7DHnd1O5tjssNeTPVpNhxnv2OGFzQj1paCZXKxcoD07GNNtLfO7sROQyc+Be
opzcWFxKMXcEIsb62Gwlrv+VX0W2wR4Jxe1Vce6EfDwc1OEtGc89po/46gU6TvlG
CfoLwU9W4Y3VuXBpE8u0xc1TUZsHLsEQ2NVcgBdkWS7X18Ies7AKeiSRtO47x0gG
LKXbrPwer08iYT7zoNWItDNzM2MAE0/UM12Jx4uk9enZvL1BzCSejY6GIYflHrO/
5shG8ISZtUgzVRZskj3xVXGVxvf7NK7fw7h7ceQpyB8NIKs89ZRA47R7qUXfrVId
KkUJANqbTYpSw9S9TlTLD7Sgy3jjb0Xht8DoF0z0qA1B+j4ab04W2zMsWwGKMV3O
RhHCll+eTFsyhop6tNnnlEUhGLcQsmu3tNDNTtCdDGaVpDoFjTv0yb5pxRHuGwGf
5NwVLTdG4GsQQuDrA3UWjvIp7RMfEOy6PXt77tY266sTAqe59nO+rRi+THOpjvXG
ihvyAspddopbGb6gslqKxq+n67tkz4aqUopfhOB5iVVFynsBXbroTAoeEzL+3YnL
9g2jOoQHpM6jYWxD7G9967kHaOTcmiHLGPDzxFsWLFSdEeTxIXNAjLiXeXMvumLS
LhW4T7EDbybM+CDRWkPxFtTlxn/HYpAgCA1DWO4wa0J/1KAVHaa2EN1u6KCqlz55
XlqmehYT0wMxNC0lsUxZARJvSH7E0UtXYNEiyIJAx84/BtfVy+4go9KgDJo8WiBG
LRuEN+VKSEgIV7jmsxrbRI1SEGDSDLXd33XDkzgYAABNBJqk17IKfzcQ/n5lR/4W
bdoBBcsg0l6H3s90XpttWrf4QeQjl3B0EmLM/G/cv6l4fO0vQbg7CwDPK66N9yr3
nmYDqgvmVRMI342u+I55Jf1jluvovcG20uuW7FNSo/rI8BewqCNfDjjyHjfYXaqw
mSTzNYZfeWS+TCReYboTQIaAC9v3NGW+PNEOQLyukBt65bquDtoH8HuNPwTc7Rax
lFCM+w5iu5lNq+S9FrhD/xIyAx0xlmucZMG6T9Lu/rw9su15+gdtpXd8tuLCRq20
eTtJZ8+LE20rvwOsaK6o3PRQMUtxGgTp9SApdXrsrglcGL5LXIcTNW0r90ckrVf+
p6wAQfcvJ160Bc7T+SuZvJdFYc6nNHqlDrAwqWruiqvMkMhntrQG5pCGy4HWhmeo
+NFp7CykqBaf9gT1gv8OAE9hMdB1lGvpda+ZXT7AnV6Xnpz+Ccd+ns1x1Jf2LSR3
xBpyfQkejbLcwIPyL8jICvZenvAlXlcvndltdxXfYmPHssAheNFwOm3prdh/tctc
JoQI1rzKpSiOBiX2xhA40K7L+vX3gKycp2rTMtw4IwYJgQCb7lpO2Yky9A9I/Q84
8hWO8xUeeFxppwwWkQH35n9mtNc/APE6n9/mQDrVn/5L0KCM7YgbKEq8ZrwNwZnE
55hwsBKn3jEINaAK5uVzMzb7UBqOeCUCggqhA8spwN3HMLva/Pn3uNeZWTaOyMwv
s9ZQuRZWHZo1i58RAArMsPtJ7HKm/tfkbNYifRU5NQLKAzifxL76dyRG9ojCQOYU
Fyxoo8b+AbjvXOAPYax3tXarJAHne+/yVkP/QMICVxFn8vfukwpdDCkdIusqwe2O
L4LJlhZwego72Zr+QcbePEdEXRtk/1Or+/cEm3Voip5w/FC7eCG47iS3MaPT7hQ3
k7WLF0OfFn/fZ7ZQuNlyXLcns4n8M55xPdrgEhNyo2sG+WYywyhgxPD4+rw/78q2
Iq0ra7RPXazOEPeWdoKZloiTNrigGeMkpiwv5jqOXfAzWsZteamvyEW8T53z3K7z
CCTS00aLLgmzeUq7Z90EHEQpdjkk4bChSTQRIcJUArNV5V0w9mjlGvpXwOXgveNG
1ONi+Fxm7BOTX4iC0hcV7wSMoQFqahNRY6rHv6iMHmSMJda8QO3ZGO7h7urRA91R
xy8+jzEt8LEJHcSiCw9Zt23mLfoKH45M198e7Bnr5gEZ5wnnfkvIICQH7UZlJojp
2pgtqZAY/YkTtrWd1aOt/sRDGIMNvafsLiBGwGFxKYjnK8LgDs1KrSBx88UsMBl6
2wrVRMZLuHtXXBuEqBOtLVQyUSe4/1p3F8myQILj9zCTCOabLYOs7ygJ86pn4ugU
TyekqhbTOyDWcdB+cgRvCE0DyQriTBR8YMZpz6K9zfouW0lD2yw6xkT5LP5MiHNx
3dE9eWwJXg55eFLG+rcNufbNzhdwWHunNxyftvMte8b0CK1DieVse8DgVj6DN8pH
wV2Bpt26xPyvA51Ai3+H8wVq4Hy2TI/xHjsDBSV0IJlIrfWF9KOAkQRdVIQLhq5b
v/MasZsKI9b9HcGttE7bw7lwFp387F4D0e5tdfv6g1JTqmEbgB4sx+5BeKveNC8s
k+VoBJKXhdzreEP6/i0s5OmI0bC8v0YN8sYQtNhWDt6CMo6DyD4cO99tUdHRUEad
ysu5NT4/yGfVKf6v1IHtrE2rVKpjzWfWLoVR3XWBDwF3wVgBIny47PllwC5Me+y3
g+CvSWnf4KmDYUm7BCt0t5dBzuoAGnRrmU4/MNdEDhHz2bK5WNiJXRotKhNi0PVu
pbmEYvidr+k+vtzEBOsvYLyN1Lfy+/UHLx5L5JnUb+dHDELRsO/LoTT5Dg2/y+gh
fgbBK7A1rgDLqoVhTc3nuOTCKCNos+rbW1+9o4NhOpYk0q6nD7gn5HmgUlmBc3uc
wy3Lal3XjewzTptVyKYWGekjmZBjOzDx7nfLUo0Wf5zrV4M59TBWfNYdUixSPs0z
PN0vAnBlHDVK5aWg8rYEUY3Q664EHDLh2d3f5db4PLg4WLrS4iQB6lYo9RXCZFGn
jPdXKRrvaB7eDwd9wl98IABGZWOVkme8KQ7jz8LqGgQ39+wd9Jwx4D5EIczlj2hz
UfewvdLfbQrC4v5Sj7jD50Z0TYxLxed1uOhSpN8DHCVfBzNQLVa/aMZDCy2mVQ/q
B+epEns9ziutRJ5W9Wdyk/c8AzQIrLa2fq2dQUBf1Y6ONfzBEPDZ3UfyUMDWBQ7s
MGlhCpy4vcc3F+3mqFlB8eUEVsXBcTWb+O/FUxL/QU3FNINaD42hceIpNraT4pAR
8v3RPhQwWxial7NH9KR9XoE0ntVHd8jE0F+QS42qfAeb1Dn/7umwoCYE3Snp9AY7
QLvvH8ZrmChdLreBNvPuR0g1FH/o7Bep6fX/wPgE6lUj0OPkz1dRj3WfW+0hKtBo
6XPbcOd24hIVIQ3q+IsPEtqMT5r706vwybVpxOo6Im5mROGQ92WXCMPa3eKINpuA
l0ESlqXRTvhFk2yBUwTiOh+ghLOHyceLUnVlLikhFw/zpH9Nz9YoNo92lO4FktjH
wm4pverwC9YEIKhgOSeyo+15YXjAaV6hiDs/DtKFskO9rJ7QeN10bBxLMC0FAeMh
he0GUMHQgjY7UcxofajS73X+A0JjflJo6pwrKwvkKSzGrF218Y455yahpuk05wVI
+B0Ygb3bLdRUdTWI8O0cReFiGkc7lIlPpJ57rzdbGgvPg6ukqVFp2pCwbaBJdIcK
xhPbV0UybUcFk4layDa2+GOWlMY8pH1JQStelwAJA9urMNUe9nVgRQE76YGtFaxl
r3xo4Lwxkx4hjkWT+yN4zeAtMnLuDhwshbc2jd0QphHO/MGOteP9vtqtdIeIXqj3
gPAspUhkMxg7x/wV8F7Trvm/YXcJ54uqNxLJdXTYWGxPBDfLYj1wJg9uqPaZ+4aQ
hF4o+Teqefjc2vDxcSrJYjhMW/fPg9C/RSKPYaVy8fymJTGtbdEkjth+6O+hfJcT
zS7rn68uK9qQPlXov4o1X2XTZil1rlSkwdmEmfaDwVrW2ze2mAB5YA3I2umyCVJu
dqIxh6geGrY3NRO3X+R5IdChl8nn/QhdZa/xbKEI44zlQA3HghzV2VogoSREJ5FU
uMMkxkIFdxIEBY50V+ThEmYJI1Ei4dsv6Zny1NCK4agbNa1yHdGEtiRFOLXN4Sv/
XXZF9j8OusidtzKmzEgywjtUprgW+xNU0A0cH4S6tmY736vEtSyII1595qg38+tm
cZMLh7Z5cC7+6QkaX2/PAqtz8uZj4kFoeZYlXVCn5LXwLpfG1lOP7hvmHHLOaZ9z
PGYejRgXfa2lcagk30UnlQyOr2tGpibz4jCMl3J6mMpU2kqHeNhuyCfLOSEHDVDH
2G0rI/fA+87KfLK3+PT5f2PuuQCr6d/GPwsaaOoQsGXp55//bhmY2IUzLimAYEpr
h1cqiOnl2fIepTOHR1OdS0g6mrOWXS0K3HBIkFtfgXVwrwGscyzl9uJb+CDQbSB4
clfIILX6xgVzw5JB8FySwxuaDcWHL8v/VAZJ3TmGkTS/28xrAFQ068zgaXq59D6s
ldohaveE1hOnfafTWTUUOak11IvKnb3JULnenJqR1qHOVrb6E6Kvq/6FCNUe1Btp
SIAkjaWZsGcAb/T2u4yv96oWvxrgET6fjR6dDGFf/p8ORW4K4GyfavR1KEeUsnFp
m0J0J3cjTHZltwIuv4CH2ce2SC9ejycGp2sIlxzDlqyZItCvv466mwZzsnLKwKpX
bDnSDTsoMO+JZeOnZGfBmT8AS+Fp0IIxu/4cs1NC3/kfQWbApHdpwI6xEU+yzSM6
k+A5MqC8e4WVANo8z2cXdchHGQGU/uoOeqxdg1hfZKovqVEo6m6rkC+cxJZLJ2wo
Ku367ouhwUbth5bQ//ylRgSltHmWxZ/Oe3Br3goimNAget4jDEBJXqzm/ygI7sU9
sOcWGKHYpnrgyZtjphUVLxe3MuZONYLvMOnpDnqfJ3mbOmRQEARKUcfY4ZozNxEJ
Z6aKyhsUk8/oTcH+UULoF2XfW7N0cXrTR+wfJZmnMli7j6A1a9OtIt152O7LzFTZ
CFwaAnI5IVvculA0Gamd4FdxA9o2ct5rXucqEPswvima5jfUUXy+CO2mTBjyt2KP
rAPQWLaHQb65BeqeEseLDc5B7HVRMtdFhwZNNuqmcUciS1Jzin/9FL0uAiBAngEj
Rlncxj2rvKZ/U0OJS1dBpPo3Nyu0v7uGxLL/0Qz8prh5xjNopZvB8aO94LwHh8vt
iQNkYCsjXt1cpNQ1zaXhG+dkUk4u+3ieGirGnGNSCG8JcRpDx755iYjX0HzoJoDq
6OYi+WNCpJ7g2AKmyj+Bc6cnaPmYIxPsoy8LrEOiExT8UZNAm1llKnLibC3GGJvB
zyxZlxgPpsPmL1rC7St63Ktak+UVWceklhgtTsQYH/u0D7uPtJVWLkKGT1O+C9Mc
Ld0m1WUDUo9x+ZWc52oXipo5OEcfv9MPgzH99jg02quphJsHxBjPhYiYSWaIsE0w
bsXbeJixbqOgSPVoFFsxRVRF89g1sBLSe4tTFKjU+u9FQQoCAt8pTvhIDVgqpQzb
u8uKPia+lOrRM3iCqyYviJ2P6ck00G/Jz6OXcCShc+tQGryURhYQO+kP3sRnsuaS
w8HE+hxAMZAO09KX+hIoo9na8q5G1SkYhCo7XjLdCUJwwdiSoulAOnZ/vdqQ1UeA
s4lTQJVgctuYpH8iBNAAmXc+z1AA1cTxrJspkHWhGQYrx4hWDXd1SrpDPCzn08cv
9iCQlt3Ms8AbuS6+gew3hVP2LTGs9umoZ3XuLPxG3e4hdxJA6nht2YThzTK5bF/k
/KgIjk1+XWxv9WrCurmGeJZPZuI2fkQu24QDnZt4bxfYMz5BpTL9DQOCybzlsZuA
0yK0pRomCDfB9UmFTlvjBQR+n6OlJVhnsEWR1aDX6k1mMusoaGWVQxWO3zKgZQEF
/N1EGsb2J3CB1eCmnNoWtMULFmvB4WsnSEn6GCqR/l79VL8yiYCoNab2XW8Jk/sl
3+LSUq536lt/jetTzKPVGb1+3zUva2ZZQR8TRCnwl1T6PYP7uxRGSRC2DvTAQeQr
nUsnOEzB31Hx+9Dx3iRQl9KRHYWhmVi4Tqc79gt9X9D01kI6oyV5cIdDdW3dAo3v
qHN8lsMC1kUmf8i5scmvI95D0a/sg6SdNS9vhIipyx4AJ0LEerT4tDk/6GkIQf4E
YGLHD69wpaBWHqfzsAxEDAITIA5NU/vBahx/RWUusX8xI9iQS/JPFTUO4qhhkGVH
7aQcRWSGa9KG7OpA6VmQnaSGm1Ma1H5SYYp0ddB6/vuJ/uYnSc3FIDD/8ieEMa02
EnYYtctTgROzrk2IOQvplzSB5Ba/K1PdxfmBOu8nlgbr0M0atPJ7JLxjEASEaln/
hhYi9EN3MPX+lr9ajT2fxU9M6q5ARSNXgvXJsr3qhwGZj1rvAdzNJF56zuhKxWt2
laAUj4T6sIM5pYk0GODI4CaQqprbPokry5WIAqdlwqO//RW62eeaU2xVyvhYo0rw
Rx23+iwCmRtSQ092sIiAgdM/F3JbKxEwzt87FYgyNomfvqhyibUr/G3NJoIKCNxp
CVBn7amrTEntm4K0i23MHlBZWj9/3WxxPllthh4DXsG4ej7dKUUDUWZzKpSAZbR6
jtBM+9NusMGsvuuZakZ5MzdA2BcSzjST7HGK7kKzzmzbU4Rw5MHDdANXFwjn7Sj/
XCtduStjBNrwtYrhw7Fx1HTE9MIfzH6ANanOHT06qK4e/QlL43TErG2iR5kMzdtI
o3Jj53K2Yup++SDrgFIoSNocaYYZ8DOOsuVRFgYsKzNdga9Ddew09z+nMhBO03At
aYZyy2aJQZUaKvTZKmndlGWfbei0EwC3zjOtSp8n0dpFMUGVDiwFvMEHiPJWHHSi
C18ypB+fJ7KgjIhxUW6/QCqlz9TbekLQNdhLYvBrK108zA52fDuQHvuFzZjx+KxV
XLnewMKuzkRz/Tv770DCPYutdwnp+8uAfPg+1YjvpOugZ3CXLr6Rgc6RL6K/bYJ7
YTjmzLR023OLO3JrtPXOZTBYegDVuqzxdEHS/Z9chAnUh35EHQU6Cho9HMWyphn1
CdKoslllqe7YYdcI+/gcTud9PGANYwUz0O4VwxNMzTtxekBT3yf0CGp5fHS28JsZ
on2SX3rIpK93vKmP0XIcKXSUcRzWQDe+3ivUqUcxYARQoEWBLXLHLbIl1VmL4u7+
+YtSbYXLO/zHIQsifHnR5EcrAanjhZKzV9fffLFNgidMVk46g/Hwxt/hBdfuPJlr
y9z22yipYoCQYTEcaL2djJkp8gUs8qW5noab9RnPdyvdagHxXNk5yAMDxkizt2EJ
bquuyBM2KG89qy31skVMODfGTeLMCgDN4AfpL3a4d7kLQKi0aL85j2YUWAtmnhDj
1Bgyr/5XKjc4TDf8pbj6DEZXhD9w3CgzJZteN4CMldvsEuHYChXDpjqgPtAgrQDT
+tfD0Qp+omfmgK3dXwADLB7y2jKq0ku0BnphQfjlgSZAgT7oKk3JGBtpkClvcgTU
Un5DvdBv+PqfK9XFv8WGIJ0zQQuX18aDOElx5FYsuqMo2sjkvHsIHziFGSDHkpNx
lHyA9RlzSeJJCDrH2B0rVdweeKwE9Z9NuFT7OVmDr11YFFJIt3qRiq4kg0+/TnAJ
vsz9RF8Y5RysaZ52oN7hz4Y3aW8+LC8VMT4F/bnTo37L/6THmPg5JZNZQep6WHSy
muw0JZliW717fpEeuHL9AfUGFAM3/7wps3/e7DD6jee0fggWuXFKLLQGxw4keAFJ
Tbx8kpob1vX8DkKcBicF6fuExum5d6UZSh/0ODcqBN8HnkRrE2BJs0OlLYfJfkB2
4EdZGzKWuw9pJhckU2kBcPVHsJUeGQNfnwmFNNgxRufcgaxNTBJYtdBe4iZ+w78I
gqP/saOuCzYS2ANU85qfEu2pqHl04jrg4QjwTKpUBxtWhus1s3cO+MNbp9Uw29EF
yIUoFzn4Vxbvqzps97wZW8HeqgWKsloPYP21Zo9cr+m/illgJnJPT2CubnIBey1s
L/nowe9v0jPXG3DeUFS3HxVpfrZ3f/Kf4Oztt5e/e+K4JOgh1m9JGPTyLBNyWnjf
yrGsMGu9wI+n4JOml/tG7J2lY9sB2hz3ec7d5Yg2UdgBW4gaXW+yxs7sdVMWwON8
DMGzo6hR/bEwmTyhblCxDAJkcWBmCNdf784jfB+sZuqP5rICz0+MMBqS2/X+MoYm
4cH/Mazf6ouYeOTDKnLAWD2pWehNtFyz3+ftjeD2tcJxYsp6zox4ULW+Prs2Jec0
QfvDHmA+cD60tr5euVL9r2e50hftYRu+csUg4RHiMkytwcQWNZgUWp/Xo+aphlOD
2EaasTp4hUFSDxbGdTn+BSTmhMVhBLHHIbQUKPoU0uLZHwwI9n+igGpmL1rmTlXi
03+UyrFEsJxX9s1RI+T2Fk3KmLH4K2OPAYIhPkDzHps/HY6xYQgVcykoXpbSkf94
3XDaxWZQyfBD9liCxqW7Yf9dbPvUUE4CtmRMPKp2Kh9t9iC6nm577lm645k/y055
DOj05lq6537+hQ0XRUsw7ia67ilHQLAzuI0FhQqxs8jhsKLsTdDRTGDKo1k3J/TX
XJLIEjH4+OHhTpESi27LYI4u1oK3yKPdqvrqQw9ZKhMh+O5zBVvsqtZDxdJ9cU6c
aXG2YYbbqwl6qu9Bczl590vpB1m1UBw48iAUJ7BrtUapdU0ys1aE3Rt/MZHqfy+l
33AzJ0HO1qj5dOXL+PIS8ZwW2nVSExD1kBo3wgEOs+p8loeiRWIOAcp++cm26d8E
aMXShBwoIR89MI8i1KC0bkM1hJYdjJwAj5+rlBd+7j9qAXlIpExHMzS80txtaFAy
0TBxsbIoQLK6lClbmLx138nVWvT5Wjf7uBEzTY5mhqfO+y3XI+ATz+JDIo3qB14j
D+OWZ+X+AiHaDumkPWjeGy6nyn7MfuZZWgnXQPALJn4vWR9IkxPPLnVexJr9zyCQ
+l2hDEJt/NHSio+F8fuaqCkxlJ0as35+FxnKQpN+gOpQ9SSx39nwrVefBVoast7a
kcXKw5YhyuO76Pb/bwpCNpOT8O3jP1HQ8aEF/jWpwOuah+JLeySeRFg+0vwslDUg
cmmK90IqQBxWgDLI4nAfltyk57F/Id0Uhc2Ry/Wgj8Yfp9IWTv10mpzoxm4Im0CO
BuuH1vcupG2Jr4DqvRvBaU+YxcIgt1YeejN86UkaVTKhg0Oo3QtpBWDDHjDJrGJG
aer1Gxp29rYVIegdLjs1ladrWnA3LWuWSzpj9/dh0FGu80M+2aEdS7EbNmOWDHHu
g0ZEsurblfd0oQoLsJ9aGeZ9JrJob0FEFf/sMF0BY5DY/3qFzujzu5se47y10bSG
3UAqYZz/Rt+DInlyN9SXws2LIAcHZlLCseDXkAXCr3ydeyULBIBnlE4ByGc+ajvG
/7iWeQAQLABXbLv7KXr3d5PTzNqTHFcUcAR+Mcuj6YM7DX32X3+wp7wfRRlAirGQ
l6t0AQBl46ujdYhjsHAizG7yJVSSNICsa4RbnX2G9sC4n0Fz2QConeoAv0v7er51
uGb7DXuyjANYFNDSevYB3S2R3aLNK3TKoMbC0cNWjJBs7P6jwSk9f181Nxj7cYKm
71WKTlayoRnJkTB6ZKTxCrCRfoGw7FJhASZMjYL9BLROew5IEfgSy2qztmtkXfsr
yPGL+5D6071RpHKf1XAyOvvCNYxYfg+W9A7Md4DLc8JRasUPSrWCdPX28b8Pd+Dq
rbTBqs9OTA+hzMOXJYmS9Qd91piIWPbfNhGC66f18ON9nxpLt62675cYw7Rj5GX6
zyxMy59xLZMO/jctW+vx9JdAlkx5TLZym7ktNP6QE+rimrsOzeOC1cCD4yCmua4+
1RtC0ugtQk8vhbTLe7wTEfWqqFtSwKZjGtcQ7fcn6BeJ0TDBehwyMKS4g5c5R2pD
sXrNGD7beiZnB/vAZdXgPaNh2oNoAMW7nWdZ1l9lVVc1P5yjfBE7ZjiIpZ+YWWye
zNgmf9cKAoHCuTRusGmYydScjs7xzRDMAAbo+denGd4kO+nHRaooByv+vfKi1D4d
q4uw6KWtSI/1zEIJ0EbLrqMu/S9NXRAsMwk9rqGbRDtCGrsbS07PUM1lTgoZsIzs
PYMQQMxsdIN51qKO0iCULbIBqBpHu50j0MEU1KclAGaZR5w2fL8jualFe9HyCpnd
ozGM37NHXG15TEExy9fkIPKIi8u/5QX6PvDgX9l+cnzaUbbJBkFs7kr79gToCRBz
nm14/jdgnGARBmPtpzrYSDIj7XA3RascnsgBstPxouhlbF44wRfaBefjBa+nF+wr
DlbFoRRnxxdYQNjTaSBo0oLn+/3L70m8PkF9jij9gYGljsjID60Q1zMv7BjQrimM
lfbPIFM79RPD+55DY7leMqjOuuz4kVQRp1txe8SNygL7xAdYDxpM8otMfxczTkkO
LKcRc+0xOC/X1E7b/8EqQskWVZmsqsoGk2Os+Iba9qjxInR4mjEYgyDO+SSkVBfj
IDgv/mytbFTBRCKQK+tQBtEhTRo2lkIOY3pcUY6C04TzKultwV8p/7yMhvnSrUJi
WSH4q3P8/SyX1Z2LpJmXoKUbFm9BAWavWsIqrZO1PsXgoPBHg4iMmC5wnI+vtvNl
l/9RDw7bd9ACWQPuO/NSM0syzE5Fgs17ovUWPFA+xvE6d/lyzuWlgtLDpBo74lN3
qZuxAgJOdMydav96tB2wOkx0+j+vkwfzvqcXhD9x2CCRsAoK+9jnbLXjeRyFXctu
0HQRIAs9G4K2rjcXveM0xgB90hl0tcUJL+f6GmTzxaGuMRwPBAWg826AlbrMJVWr
ou6gaqmsGcZWgT3z+bnRtgGyeQf14c/gtlQ0X9hg5Da7m+CWqYo027aQcjSX1hzf
YcjDiowZLRzQkVNrEr0SlS2K/zl6SxsBIHeOJdahqdJ+aRGC7TX2m+gOIaM1Qw+l
3VhpcwdIdn4yi6+xk9eSeDZMN0CBP2HOI1BnSwAOS/16GcOyo+pSJn6L4vn7cc3m
hNLIBud7pBqKxzMjmWHDPOvxm9FXQgnU6LtNB5YYy3EQh/1ARiHmbnLNzmgl1X4L
RPVmQbZwBV5jOCXNt0jn6NrV0UM54fe1F90WaDWzluuGPwwH8tDmuBpatqpg/+p5
OeV8kKiAZTNFuMyblXzyMtmxgM1XTZfUT5uEu44UKpqCUBYIuBmeBUhELhE+n1nF
6vWH/qRuWsLZR57BEnvMxlTT757kw6eBvRt4fgvtxCeSRvMfDdq+ww0sgTSvodzf
44p9qzPx17t2EdclXZr8Ye4WjLxCKMBLrPZGxJCK92YefosJeujmF4y8uG4t0IrO
xR3dJEyhaiNS53VSDIG5MbbqQ3ozbLmQcoP8e+r7tCN0xitgIpjYJ4uTKkvDTm8c
z94Tk4AVBZDUTzY7JefF3842ff19hlrMBwWuUwnh0FGdBk8M+BWrIpHBO799HVvl
oio7s5Ma/wCgFppG3wOntqI5X9Z1aJcu8DLoPHY3hiSI9vgeT+g9/Z3g6cYDeEzV
SN46Q0FSAPsXSLocsb8qYaS/SlADCMTVDHfCQt/jeyduxFAaIXNt9gTn0QMqcQLj
07cT32JUURyLCWJELQJ6QYZKlICJr3GK9KdV1+qNzifkinGm+iW/bbhEO2+vI7ky
OPC1vrNS26h+tPigE4QesfNbF5TRFovjoH/2ad8zGi0fPGOtrMqEUn/XTTtn6akS
BZsHR8b+yLpCwjNYBiCsnShBcR22rXlDYUBQjyperFp3zPrEomWUUeGGQWCpWnzY
NIGCSXO9ry/+lo6CvwSW9KGAerFpL69mgzSTL1ga5+84mGOfmZjOgp7yYu+yGI2Y
f73MpiyD3OHxRz8C6T8wp2Nzq9kKl9ZHxAN7HpqoOWYAzHCaa4pMRuctxOG+EBi7
ouAIhRuoWFTZ/o2fNJVosaAZiqGd0QKAPFExlzAPQjTOnXtaFixqSmNtmh7NAwOU
Sd8aJ6XCzcs1JyFWw+wI1oH4TH94pwDdGbffSNftQM+YPN96ZuEO9SYBEUlzwepc
fFqQyrRgbuxTITLedetrcnbdzklUv4kYLoJWY8cdwpJjr9Qn4LO/zARXVZlDnw46
1jJS6UL8DgZ6mEdk5swcI6CyqIr5+7j24r0F9zBoeS+BR6cspzOaLS1BJQ8dWojT
fvPuZpR8+rr9kTejD4Lbre3cb4pIPQsaZf3sxzYR3U8VZg/EnYC2UQzz6b0zjR/f
XZ6QuZ1xdXTDYdfEh0olIj7Cry9dupA+/yzBez6dZEK0kLwhGswZbPTM317WSl04
rvXO6gTwEBo/Ec+gE09IRSqqTpP/j4PuHH91/Q2f0QaRFBCvem30MyjIpikf2qgz
0S09NqzW2X7ok66f4oqF3BOoCfquCEP09Rf34Jd0KL5Yx8O6P0Z9rDI/ec98wysk
frAuLbMRN8HIafDxUm50Z54hAs3oZs54rvYeZBSvzCeAI8qzwGQyzyjgaeZ6F9dB
KCms2LkPikiKCgNSYoYBqQheRpJ7R3D/WcgFGrUnK8U6P28PCB/RrwKOECTaCmKO
+8aDOXs8yWePmV30e8cOAOq5CfP0x/t/S8ZmhfFnB0F1EVEwDvgVQXBurybYn0w6
aAqkdGZRTIxwMfN7ZK3tZPJoR9T1VoR8ShcVjhdN3aBIqHgnT5eQK+xnwicjfaQU
8uPyD8G0P46VxMsvoCDBHf1o72vfqwYUbOBpEi/osNCf5bYSbqzWxqLEZXUfGP79
d2Qk17cgUzR7POIAlkg0YMvZK2TB39rmkfhKPQYtgJ89Xz9iNNYy7ZxUDNOk0nSA
z7+RHGG1WI5Iho/vU8Zc9dgSun9r2cQyuwdjENoPmVvh73w33n67AS1yC8BksAu2
iPFOqLDia7/UDAYX3aa6LGonwyYX4oCGwPJfGUB/igrW/adHwM+mQuNc9v9BNl2G
8vdq3D1By/iNRT0l/2SlOhS/iaAp5tQY/X7DZlACUrF7Edtl7CaxbC4nXFLhf8pt
TkVklHYt1+lxZZm8HiBjFe1Wj9U3lh8GaeYI3FP08mKJxxmEIw0a/bfwtSWJsWEo
LunTtCbdu/qbl7gqCowS7vNq8LAARFtz/VxSclWn0YZceGTI3yCvJ0bZ3eatAMx5
kGEqzJhdPNzIYuuE3EQ5v6kRAar1YyseHaCEsA8wFjJEekt3oKM0Nc+S8KJ2Xdg1
Pdxbrn/vd7LQSLDILnr0+KclthohZlNvdZqYSEtbNZXqVww6eiQwzApeCMERWzAF
UUsGUd2PnGrfdo+71GPbrioPZcBjiBWJK831pPin+56GN0xygwsJhwFOZBm0J7fs
b1xm8Zi/YqH4yOaAFJADdXNpHjNDcfAyJNbCD9BqlYqIriQLghqzomgmB5yuxNNP
8ubkOZwTCNXPPkdX2p/u+r2UGDYnoXbjE/bP5k1GBqOZR7q5UPHuiUxmc5bkCpuN
jv+0O0ulKGnEMFq3ZMgFoAxRmAhntYSF5UB2rU95QOmgQ8kYo2Uac1ODr66pb4jA
O6YL/EZi6I0HrNWlMAhoZM9JLN3soKRaaEwXXuFXza+jsv+sPqsoNvhRDD67568Q
LtJ0EM3MY5ip464PAH6WQ89slndEY73liOMmxBKGc+lOCm/w7RUe5KEur5kbrxpV
BdqvFjEKxK9fzRfes6eYppoNlr6QzRk6QBCOGPWOc/hct6e4EHv0Il6dgy4h8ohG
wkBCr8YViEJcRXoQ5qJzMQRDskn0mz1G78LgClVxaPRUmTgM/V8n65YCBf7oTW34
bchskzsomJK1eosmwLXmExW/S4MiUR6umgz/DcAEGTdYPD5T050zVqx2OF3KrF+r
6X0/Wt/+Cku1ix9dsDVED7eRySqVslgPb3qAyYYtlq80LEmw326yyMUMxUQfkFAV
sECWUtAl2uzMqRbYQlnrt8B25sinYiB62eNr1//EbCaSLAVwm1LKb68mj21tObyI
527l1qpwtZwHS/8Mfd8lBkZHCZA9ONj0T4+PL/g9m9AWyzfRjcvh33D6vZPq8DEt
5xTAFV2pMLQsmvpziSi2PBaSISKN4jQLJqvVyDb7/3tPxqrHVV9wOKL0C4RJsJQn
MuUv1IJ8V7UdzBdYAqe2EXPiFYhN/A24MpG5FFvbrmVkaV5B6h5tX6HOby7Ww1cC
/lkDa/IbxiFKgn0A3XrcQfrg9xjcnyyjnKvOgm5XwSgRDIX5Nvwis2L1BG/TVXxR
9hhW4/8IC5QxSwrzNaPLQ2UlFXcPUNoeUO3YZ2uJWcuS9r8ioc5KHVEElYWlk3fY
CKSDnDzb5tzAC2TSaIXwMQoWQM3poW94WWp1gTOZntgoGH1//bvHe9OA04kZVmjP
8nPa5tCoAwM7N2kFYKUecEIroyrMwh7HDd5RGWQBA4fc8czx+VZWD1uFTkdyTStB
vrFP9DvDYZOPIxBoX2MZGPTyDzEkGLnBQKSZ0DE+v2Zy9Z6/JpRY31wPQkzHz8RP
SOQvumWGbXSfiQTWrgSrAvhumVtrKr3RaUaPRF7x8MsQAjJMIXFPm64MMc9iygc5
rkvzvpGBWZeGqf60i5/AqjCT/MiUCR9pQB2Oy1IzpeRAXvgzfH5hu6qRvtVbXIlP
zibUY1NAT+yZvhXxaL20N9USgzEvSJOfWn9KDNBtn24E8Vzw618fVtsRYnwzxoPj
rDTMXx+4zIiiC/HqafZrAXmKvpCHQcnkMdh37TqbySA837gzq9WPicbI4ASdtYBa
0yJBHNrrqS3vPmvAkzfPYPTLWR5EgkUmg05XAWJgmOd8LhQBDbCTYmlUnMI9wbNI
Xx+H6NJZ1kFU2lOuoQnQYJ191LhNzzRoApn7BqL8dH5q+FhbeLmfH6huJxmT7peA
tU6IaHTuFVlqnTQjoCYU00g7LCh8JQxVu9j2OuLRDbSqId3FdvbT7vRZTrgg76hg
rWjGOjEsNGlgxVvqpQywi+hgPdMutn8zfZWy4ISFVPSl90uLiVER5LWLnC94HSix
d0ZGxZWVVy8nwFCodDoIc+sl9deFKysy/xWsUfIBgVx8vAqeh7I+OOvYqXJleZKh
LmmKddM+LUZAYwPnCMq6Nm8B71R1H1eiFhzhA/mP0JwpcQn1vqluIaAioRsCWYWA
gRXXzGyKXt9NXMUGj+pdTkYHoGIiznXppcJldvECBtD/8LOWNyeDb5r7tVj3w81L
YWVd1ouH2CkFamHi+euKBlYLXE+MLaV22bc2pMpEZpODP+8VOTuLmrTcDS3GgGhT
hCU7jL7jbBk688K0mJFJSmDDuHXHmlHs20ULAGOX2ULjTdjKAHXvOAswZ8BLDzva
GZtukt97F7mEjZ4jeouxp7dfeg4YRM9ugG45cPHrJsr4g+z8ScFr2Ad8m56bv3hr
+f05GNiag7Q3kiCM1uSAxyR1+yJbWsy7D9uJDVuMkrdU0sU46qcq2AN18MtOWn0n
ljz7zzx4FxhDrHz67ZGiE4/1uatUJnzshj20YpoWvRsc5pl0Qf2HCqP6wtD6iarr
awxHLCzifjEoY5z7Oprx6OOqriDCB2Zko3cYyY5WkVunkDiE1hGBM0XAVOFXbKit
BMWaef3LcH8omGepTAGGQAw/1EO/0THEsUTPfCYRTbKA54y0hntz5vNWJg9J4qK3
8m0n7ip5WVHai2lPZkgkTNCNLrlRwRRVUCKqLFlKRcAoYloA3bePdMbWoU9IAgPe
rF9gNlLN7Uc+psPTUYElCBu/+HLSqaVA+IdB+soRvKmdKSHvSlr2ofs4XVmbTfHA
SffL/g9YJoujnrw/eIwDgKzdz+eaKP2ZW9HX3/EIYDqgOIuKTHjrn/np5U1bZFLi
nQRQBlcwMKq94Ew9YoUWSfRv1YrspiLAeTbmCXPa4O7BU46tnzBU+msNsyM5ksDJ
X8uVnC+oHTPCvklIg+40manFcwJGTKEe5TriyUQpT52avjhrXmQOFFnuS/p597X5
k/7OBsc99hLEgjJSz1pjVjoNmIduTDja3ehRnFg+02NMpfl1jW5QPWfbweUWJ09S
BrZX8LbTREYfT7U54++lSH8vZBmmFEndTNFiBSsTlRrcp2lGhKtWRdVDuZ5BARNU
2xCLERQCC2b2aPeYW5Z5E7kKzkNMFsVF2DAL6tQWLuRGtPsk8UT7fMtL21pswRCX
zq6zYL52V3R2rcuUqs7cTM/yyP+opj204si73C2BZ7pvcsqCkfM//+Tw159hqdr9
bqR35FoUfpitPW8xrIc2ww==
`protect END_PROTECTED
