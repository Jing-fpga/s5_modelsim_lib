`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lYKFlXZlU7CJQV2hNdBlic3kWS1D4VBSrrkbU56zlVlsa47rwzY+LF5Y54zxrlBI
/l02B8GscB3cMAwgCuSQ/hl8RF6HoiXg+PQdfh+3Ju7t8BC5neS2Q1FiIs9HIQoT
kD+6GvFFDJ5CKsXGjTbhrcPvOOsqnlQ2D2fGigENWeBxnEG+INhYwyOvTipy1Ez0
TKxmUTvuSyMoL268kQnPh/AN04+pvU3K1BFQ+fu+auirTOrgvAkbDqoPCgAw31Vs
n7VQ14K4OlDooPZNmx2apbftZ/K+uyv6A/tX7Yq/OdhmjFaupVMDRBnVEP+J+A6U
KAxowbcW2N7yLldG7XiEOqsTjxphJ9Bf0HgbUyUaa7ZWxpuH2tx+kXLVuwF+NwiN
QUGkdB8DbiekAoHho7CqxbAorHye3JuHGsaKAmXm/C1xlUnjiOcz7UMMLCm9KCTk
cMYAaODPlrv2/YUcGgdMOqKHhKHcdbZ3CXRY4bq1tDLZd44e7li4WkrbIIp5J0eL
/pwX0od0wkU+HXhL/gYbYsOd93LoKSmHfZOWmNNE52PLykmB2tvPNx83V1sCw9SG
b4EWvgdvc/LXmQ7CEUi+GvEnL1OwgQ0VSpmj0lIy/Zc1sJkQtIe5gAgnFOgeRZ0c
g9QzAdob5+7KdFi4lXT4fAAbPJ1CA1Y0QuZPs3uOKWTKw9bEsyEWoTRANJD4aVab
cfD0e2sGl0zcS1z+5OkHu1N5CpsPQsw11f5mI93/belfylRDRm1KCCwXowPcSyug
wqppvdsa/KbO5ULmHQdNXLsaqRINQbR6xEnEVQrQmTgd3i2ken8e+L0jAxdsK2yu
CNQbeI8CpNeW50JLKQEKSUY+U58UFFhIu0K+ZT1cd9c+QNCwiYdq0YQCNKIm1qFm
w6Z+RZ75dqd7Ogy4pZq9l768YdsbdsD37pouT+eJCtIKmKGjHozVnaZn3AIF49uS
B/YvjiXnYuNUK3LoA+36UbIU31OGFGPoe6VfPrq9CTQ6ISZrsFEn+Y7J0JXrvz7G
QQzwm82Z+JLF+nGcDHaEJ+xGR84SYubkZXyuZhIhH72T5L/H9eTbhHdgq8zFOa7N
Mg+FEiYSNnG3GdD+etE8S+swn392s/Xoj3nd6tzE1Dof9ZhCL4y3GEnvEGPRYDjb
sJjbP7JC/zg0wxHhPE/f8bSJZh/Y3VQBCpkM2YFg1MU0AFTTZZqg3Kh0WfYq/wbj
uXL6YgFJm+CZyNc6yb8XfIOfBx4NqJ7SG4A0HGPK5uYtS78TUAV7b2o6KDVqceAF
DxhRvmf08L60z7OMx7t4ha9WdW+a49EUwO/ePG4I9EFWUrLij6UgwdmGqiOvYRj4
OW2Opd/2myS99xGXBlz3D79W/eSJG+MEBee2827u22jAf97SPL+yexT+sZvqkosZ
SS3vNlFax3zjPe3h9ukBFr5dWTpPSP7W60O8mi+cVhrZ9bSM4aJJGKkYwtEP860W
6+RHPy4DlCryMDMSmd8/2wEuTh4OpQ/E1Hgoz2HJYKWv9ppvKB2FNFrRRla0AGSq
CC89nitjTs5FNC7mW2GajKHKVKLB3g7NBEKY1b2t7tNeT6y9uExhcBfr0uffc5dm
kY+Ee90LbOIXR6AvIWEv5tYWHi6aB5XmcWBO+DFl6CM4pt4CFS0XN/0Temb9ptFA
y9aKUBFxip8MHGLCQ0KR8DgzgaTaOt+Z1MYcmo53DID8qL3zOouichhzJlNOjotM
D12RCQXsvNJgFJJKnuJu/h8HiQcpqUlOER979TDJq1WQ5PXAO6AxXq7feo8y58xZ
oITk9mT1AvNtdgNiYkVvn1GeZbwaJTorj2Ld5BG0ASw4QqzFnCqtT/y54cdAqgKA
5JNXIGBAC0fIWVeodK/pNZ12CaAvy+SP0uTusaT9jk8torqN2LcsTiLBLZG/bQJE
Z6T8vmCQyenlz9JHQ0FdA3/8MYIEyO0yDfanY5FYWc7UsZggxYQ4hquySIiHO9YI
4syP8sdj8JZFMdB0vjIl1Hbu71aawaYoVqfKB6cq5mRtXZDqik5a3NH/5LjWgTN6
RDBPqIhly8W3wXKmjkFvNmC7+cpe0cLpE5QFOrwOKf4zVgrdTywyZsT51wh5aoE2
CxW5OQcViK1FTaofQJ52qrkUn8ci75WJVZlIzdSqEkVJamG5fSFutpODCsnHbRJi
fIey1lK+tJCajbMQUHDJpw2I/WDyiD4hF2kgybsFZADGW8WHbdNcNUneMJMmIv+d
MWFvzJL3ouRnOozqDE+Qcwiye9HlcIJkDixokkVHfgjdTpm4vkB2bKfBYlSONGSD
RCJvimut48H5Um9GWICel0f4BmBFIQXWxacm0w80G3G+75JjMveqogV43Wo+hzNw
gOWZgLhddjWN3RXYgJ30mQyqWbOL8FyDQ3Od6mx2N2UgeJVmG4m3gYmcM2f0JAxE
l6EVtnJQ08LSNVuho06T9dwD75kf55bV8GJ7wfCnfU37pyth71uXJ0fqh2Z/Sg3V
nFEN2ftPpF40JFrXZXKsnq3xawEU8Eq6+FORNAtmTBLf9bNBJN81XD8ADH+vPHWe
UCyIR5vY65IxVCSvxgBxbSheRll7gYI+Do295NepTjVuCBXkCsZlZ4rHwfWe6iU9
aCj26DDK9il1YOeD5g6PgRV9WCgHXiJ6weKzgp9qS8d+Lbw9IhBTFGAAr0PqhdvN
Mz4j/sE+cAbzsEJowjOpzjrj9Aw5gGtv2FM8o5S6Fxa05k7V2dos6pnw3V2luUeB
uE2ess5QpaoLEXC0qDRWLcB6LkfADehMSUqkyzwxHP1yNYF5m4MaRzfy6Hbd7jvq
M8XloyGKFyf5HBkIhHVbQptLo3yQ+8k9P+594QExWrSXNeCe+cBShKwe60thIdEz
s9gvS7voMLntRL59JfbeJIy78UFNQZBpPYVqUEHzvzAh3m9t6NHBLE/5cpEjaike
mEoGuon6ZByWM73fNLeEVr1Nm6swHkJNA6/AJiDM0MZgoSVaNzgQk/cOGmiqqAHW
L7zXhkdKnblDl/QHQXKAZId+mQvp2tj6pbaSTlUzVZaKZZ+4WqHfEv0WX7meSNJb
PVJFcmB8jpPSiZ6yEoheISDUWCqolxwY084zJK4nsNZltRN9p9Mt9yC1Lx36OUl4
0VG1OrQ3SgWonbHLlUnlNpwbTPXYRa6wDCWcbKdTUHN9ZCKuo/C3F91bovitVzOM
PQejD56NR54kZ8OnT1MN51SNtdSvKHcj+/56co0v1PNiJtYN97L9hPt/y61nMy1p
+J2mbfwk7ykm+96YN5xuWGow+z/3z4ujLx+iG6kcPrZKkkbGGkWYLO5fDsX9Ryja
WcEDZQw5glaeXpuZxu+E1MRoG0nYOH7ipV9YAcrVoRL+X4Q0CzBRBWyct8qXmKiS
CLT06UQfZ6HV2GbMJrTV7SHp5aavOKsbT6X5O7UTtfiURkAA03PigAeai5ZJ3BtB
3C5xu3kujz9A/ObloyZsbbOUTL74UKXf+yD2lOcdKnIW1hh1TiqJpPrGq1GpvuWq
W/r2aHFi2IV+QLTSI2CcYDRRA/ygpWpjQ6x136HUb4LKBxbFBib0zJPsUrQ0aH6p
4MBXV38XKG2qL05J5GSykEzJG0znL0wdeBclLZBNPgW1MsKBtud14t7GrPxSmXzE
1U1StMMhm2cfRHvk7dkLTacn4dQX0xlsh4MMRZGZpSFg0jS+QvBh+jhSxojurczl
qBUgM4qAH53XcaX4WG1tkOmg6FrlKZl3T7jxu+FUe8KO2Yc+Gw72mmEfRlezZKAe
eZVDdeaU44tZRRZ593d2Um5Vzr/sfNqCN36QHwHbANYkG8I/GyE+8IUqPzgpaWhs
/z4akm09o1N62UocML16NsRvbfgma46a2awVgpqXQ8OD3SPtpqCJFfJw1m7JGvsO
3j9LxDQfIQzBR4uE709o1ZhbIhW40xhTQ5HrgJP3JUEFvCnX7n5G8hX65HdTKRTb
HGLsZ7eGPwmGNDfzNTMNRq7+R5ryrsBoGrgeUy60wxrHokRH4XfYkGK6gT4/znHP
ZJT2R92kXw9mXbva1I3rebFTNNQ6iTUInvOZqYieFu4qQLexlpiL8d8Uo2n1wkRD
9MD22EzBOr12XhhyQWykBh/fUnxnIdAndZS/nT11FvtZgJv24kPwytAJTG0Ar9Mu
Im1HndLArDG8D/0HjOwmSAR+PV5+Wl3tenCK1UAoBBvMz+naxDpiJvvTaYkicMD3
rqWfYSzp4EvlZyh1Vc6uivPt+GzudlzkVcfjLxb/XvpE5wGd7Hs6PgE/KmEOCcX2
/oL3qJl7ZHWUY7Resqs8VHoOZ9GcC3sKnrAdeJSSNolQ0b1BmATObuu8I54AUNj8
i06wLqSFCCepLyE2xTSshm/93u3bo5Pe/Nc+V6kiNC1ps5SMUJJqwwNGsBtg3NC4
`protect END_PROTECTED
