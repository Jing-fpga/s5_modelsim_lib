`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gcOvST2l+DoxVBGwOf0HiHm8Y+L+qNpwX/feQZEhpsoeqQEaeD8CGarkma5K2Mor
4JYpY0MWqymQxw7GSDbukuTFnrXKw6fh6wsMbrI20Aba58c7/zHd2Vxj0rvVZOQr
kCessNZ3xEqGfjKH2/mh7yT/kyZ3rNILx2ozdtmCmRZ5Bog2sFpI4BcLe/7HwFZA
DYWheJYYDFo/5ZKN6G3VvEb2QUAW69byKHzn4mGjK9eHdysIusv3DxqWdhNTZP+6
Eacyl8+Lh4wlfgQ1Sp+snY3WRZ+iQuTAb02E08Rr36ESG78ybNKkCUmgL0ACSwVe
UhxkPoqJuOpWD6RBz2qExV0EXXmPkN+XKObwjmVO7JssrRzg0U8Uazn2dCD4Tvmr
NBh/xeZVk/63JAOm7YKr6dm6RyF20VSPQLipno42knE8e+447k3lz8d6K3I4JLoe
veib5I1nqq5Z3lf/zZpL8ek684piMwb89IzOqNC4vf3oQkush1fsExns3Wvlx0RM
w1B2iqyNLC6Eu4oolBs0RJJ5v3jrtSzWKu/QRCAnUQXwy/FENwuj12koVO4uZ61K
0YhJnjVIEVhmTVCbJdXRnzNV/TQBNBBSGH26L5eVyjT2O3ki99L37dY3nPixH9BC
`protect END_PROTECTED
