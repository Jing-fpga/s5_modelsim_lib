library verilog;
use verilog.vl_types.all;
entity fast_analysis is
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        rx_rdy          : out    vl_logic;
        rx_sop          : in     vl_logic;
        rx_eop          : in     vl_logic;
        rx_valid        : in     vl_logic;
        rx_data         : in     vl_logic_vector(63 downto 0);
        rx_valid_byte   : in     vl_logic_vector(2 downto 0);
        rx_msg_type     : in     vl_logic_vector(2 downto 0);
        dst_rdy         : in     vl_logic;
        fast_mkt_sop    : out    vl_logic;
        fast_mkt_eop    : out    vl_logic;
        fast_mkt_valid  : out    vl_logic;
        fast_mkt_data   : out    vl_logic_vector(63 downto 0);
        fast_mkt_valid_bytes: out    vl_logic_vector(2 downto 0);
        fast_mkt_port_map: out    vl_logic_vector(15 downto 0);
        fast_mkt_decml_place: out    vl_logic_vector(3 downto 0);
        fast_mkt_op_type: out    vl_logic_vector(3 downto 0);
        fast_mkt_data_type: out    vl_logic_vector(3 downto 0);
        cpu_xml_waddr   : in     vl_logic_vector(8 downto 0);
        cpu_xml_wren    : in     vl_logic;
        cpu_xml_wdata   : in     vl_logic_vector(31 downto 0);
        cpu_xml_wr_done : in     vl_logic;
        cpu_rd_ram_req  : in     vl_logic;
        cpu_xml_raddr   : in     vl_logic_vector(8 downto 0);
        cpu_xml_rden    : in     vl_logic;
        cpu_xml_rdata   : out    vl_logic_vector(31 downto 0);
        csr_fsm_restart : in     vl_logic;
        mkt_none_bit    : in     vl_logic_vector(63 downto 0);
        vir_none_bit    : in     vl_logic_vector(63 downto 0);
        index_none_bit  : in     vl_logic_vector(63 downto 0);
        totl_none_bit   : in     vl_logic_vector(63 downto 0);
        one_none_bit    : in     vl_logic_vector(63 downto 0);
        idx_base_addr   : in     vl_logic_vector(8 downto 0);
        vir_base_addr   : in     vl_logic_vector(8 downto 0);
        totl_base_addr  : in     vl_logic_vector(8 downto 0);
        one_base_addr   : in     vl_logic_vector(8 downto 0);
        mkt_base_addr   : in     vl_logic_vector(8 downto 0);
        no_bid_level_base_addr: in     vl_logic_vector(8 downto 0);
        bid_no_orders_base_addr: in     vl_logic_vector(8 downto 0);
        no_offer_level_base_addr: in     vl_logic_vector(8 downto 0);
        offer_no_orders_base_addr: in     vl_logic_vector(8 downto 0);
        fast_fsm_state  : out    vl_logic_vector(31 downto 0);
        stop_decode_err_cnt: out    vl_logic_vector(7 downto 0);
        totl_fast_sop_cnt: out    vl_logic_vector(63 downto 0);
        totl_fast_eop_cnt: out    vl_logic_vector(63 downto 0);
        mkt_sop_cnt     : out    vl_logic_vector(31 downto 0);
        mkt_eop_cnt     : out    vl_logic_vector(31 downto 0);
        idx_sop_cnt     : out    vl_logic_vector(31 downto 0);
        idx_eop_cnt     : out    vl_logic_vector(31 downto 0);
        vir_sop_cnt     : out    vl_logic_vector(31 downto 0);
        vir_eop_cnt     : out    vl_logic_vector(31 downto 0);
        one_sop_cnt     : out    vl_logic_vector(31 downto 0);
        one_eop_cnt     : out    vl_logic_vector(31 downto 0);
        totl_sop_cnt    : out    vl_logic_vector(31 downto 0);
        totl_eop_cnt    : out    vl_logic_vector(31 downto 0);
        msg_type        : out    vl_logic_vector(2 downto 0)
    );
end fast_analysis;
