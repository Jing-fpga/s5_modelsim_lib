`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NH3aFKbccwRnyN1BX36Z1KhAWontvSELalrLaJPJfMgVQ6rAUfrFD5gIWISauq8N
B70YLvqVRmcrJs5d75JHj33E4aNPhl8IQ/GAFzGiUeJSF1iFCbOhUsi9EfHNeL6+
/nnABoGiot4X0jK/SaXcoE8+mNKmgIv8OgaISEmBCu7y9cOpddowLwixaUAxtRHA
QTcZ0q2IfwxrUsU0dd64BcLOHrxFe22LcrG1/ilBa12LjpPJuqfpvAEFpalunSyH
uRtOV3w2j6yE+WC4k7wdVts0A7sfqO/B/lmqj/B44XER+u6YeWq+CMYbOvNRzyOt
INovY6kRdcHLOME5yFMS+9R9PqX22Yn22Ymuey5Sf8gVb3Ke9rF7bOqkw1zsK6my
OWtf1y3xfdfLHbI7WnwlY1/PlNaQjqKaRCZl7CBpMJNyEtLuZCnczR9c64sI5w0P
3sezcu34X5ucNqb9ErkKk010p6Bg4fNA/SDAQ7Jg8nStivp7/VgAKmluqa01ELKT
dhNlfytizdSM7ZneNYuIt7wx1czKdf6vEEtAXOipI0rQeOFEhA14QovR1ABh9VHY
HhwjuBNQdOjVXCYnm5NA+cWeCQqhJB6M0e0HZETi4Tbp0physYZoVNHt2glIFQ2Q
vSFWfqVaLqfQ3JysWTdYUoB1vDQney5mUpQ/Em9Qk+XkB6OGPW4ki2Uk0ZGsO+4Y
flLZqEauWErBwuHeJpWBoKWTwOC+4+TT8KKaqFczp5R3nBer4+WxXQ7BdVUmVHPX
cBtZTAstLPRMe9miA8rICMGYub4Ij8a0TRQ+jqASzKZmVjzv9t++f4dau8Arve3o
t+bz/IKeaRJB2DiRufnVcn0YksG3COkmDwJ0GO054raH2J5I9QiLEqSvabIZ7FbA
XJoOzO4sxCcfrZMjrW5IqA==
`protect END_PROTECTED
