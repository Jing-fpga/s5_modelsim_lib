`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6DK9J5qPP44LA9e7Hct2E+aX2E69/o1/N+4qYN8PMFwj9VlnIMoGU9+TmtYdcENV
ZpgfFCumvgj93+4ZrEMzdWyOJEo65u8yAXQF7+IBVSloRt6ao6BFS3VB11spX+1Y
EfmRu27+AyXZ7fYbjEfVRbUxVVmmQBfDzptYEGXKTS4rbVHNNI1N67NkB4jelVaQ
OGK+azzXD27hqMLlP26fXl0y63dVn0vLH7B09WgC3azyodlL8Y7HFqKOCOoKHk+7
o0zcNurgFl8e9OSY37XLwiXUu1jOFJxHeAtdW1oqQ/2jfZcXZGO6/oJXTsw6TGdX
OV1oXormdaaOaknb3RJCUNiiCqYnZ0d9xWioBRWurc4ZmlHcKHLigCkfvnwvoTQb
iyeGDGE+hsmj0yUTDzFRJSweTgHARdLvGxguuTGdqL22qz0wLnpKk0ciaetem5SM
2A0/0vP3nuNBrreH1ANODe+nl3gZN+tU/nqayWJDF/DGdlzO3VoxKR0HmEQMbKW4
duzoi19siSg3YNvhw5iRQkUJ0asbobibSMpJaAeUhOXy9V8SFMMroYnvnXQ6KJgw
IjpyhEyWuXOxRXNupjQ525IqPwOvPO8o5XDV082IzFeg8eII/1qo6Zs9t9LQkZ33
LIB8eU3jiUi4+RTGXI8sgu4BIFqnCw2nIQrIdVcG6VuQPUf2lzIKXeH4t0NDiq90
VH1qrg2AmkXxlrRKTqBI0IOh49qyOfmEaBCOgSEcZ0j0WkkJKYwhSuvkE0qmV1Pd
5Rt+6e61tXCxT13xv9KH+KAxVah2aRE0PMfVlFf1sGFtfWqCteJOdzADoShnRkD+
QApBa3HZ8SMPumEkShEuwkSnFuDlIO2tTsAd6LVAQHI6aCNX41WZSeY16iDg29Io
YM0gNvWV9+vsUnVDrxVhqzBFcFUUxatpg8ftEjWShCp2PhybjGcq4Ku89Q+Cw4Z7
uJXBLBTCUf3KRc25AJaIRA0lEW8P314lU/SROoyt2GCvst1DWJinQmkb3N7RuQd0
v182IxwKGQav5dYSJNk8/wU5bF/ziK4GZXCcXC5j2qQIWH78Jp6nhfcqefhHYq/P
UOH9Yte/HiODuf2blhPSOHiYXNIweuU+TDKdV/CCt3EDrgJEhNMpwHZqvEO51FI5
/CCC7AvQt2P7I8Wumn8ow83uUAoh/+07w4hwiBc5+fHLt+CJDoHpSvcFIc50MExh
V4VqeR+A63o88B6SdLLc8KquB7q8599ISEznOBmQR2EhXvc/pYFo4ObgP75DGrm5
cm6CCdWSaMSQB3R8WdBSzz5EuSXcEl/ODkQ7g4lNYctEpOlKTk6lt7Y3Jgw3vcOA
okErD/hyGdLQDK/a4jswnys3K3Y7wcWTrLEjmB9jEGbpjIkEPx0Xp0MAvhrk0zGG
vhB7uWZBGLLG2PEKZlmilOsYGnVOs7KbzEZj/Tbe+QmKcUA3AQbTtyvJF1TTtsBy
bjbR0BBypQm5QqiUzZTAIlVEU6JhZgrb52tEfnDNYyI=
`protect END_PROTECTED
