`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wD/E1CkgoQR3YtnjyF4GYexIkvhE3TMUqze6EkesVOx4oI9aRE6UwUZs9tnvdWGb
hN1n7rOOVat2FdRi/qd2Is+XX0mK4FP90yxJkSSUahkBpz7blbncSirS/IuknU+9
bI+rupHSD9o4oGvnGApSQKCaL9ncTapGWQjY4o0pTX1rul4kGT73V1pBVK/ILs9H
d3t8/tJy2u8928amBBi15yT/yW4sftaO3ImEC9lNb/bRDHBLWtozHK+w+14rfjPR
Fb7dr53iAEelz8Ocya1kgbZlhTP2Z6xcEJsP5Qq+abg71UWG7m1Up1HX+rHju4gh
tWgkmXYSrLes5Zmu4FlKPJb1FclcSd5eY0MypCxOG3yV2oxqOhavH2E0J71rTtpG
IGY3MhVB6Nom++yRIZ3lcwwvAtv9jetfTiHqaqP49LFbmvBElMkzJI4q2IdxSdNa
2jAN03EE7NIGIjA1+u1zq50pBQu8j0BPTUYS7MH6Thmnee284Ka0eLVGCmiOnEfv
SMsv/ileKZl0ZZGfLTthcdhVGQ8B0hXd4hB7BqHwzzlzT9uzgzG4tOgREhh5GtUh
A3XQvzvK+T875z9Mc0QWiYa7z9JuWfDUpgdImV3aP4GUVPenhh/5S2AZlO6NxLG1
CX1R00Gm9jnENhR4QUzeGBZu+RbCEvmYQWMWx1EPSoZlVos9uVTSyuEYR8duGpr7
OynBgSRdvcP1FAKrmBp4pispxdCu8+0PBY6rXm7Ietj5xv5iGUc7i1t7LxXLtZmq
GGgm5+e7ngkqW+AtNKMZA6tPoot/z22DoX2UMGJAQPFUnsaArTjGVC0yjQzH9hqY
7LZoQDFhqbMaix9uewoSaBa22UDkMT3/DRSSE6PYNFxefUKFwSi3/iEKHGVGkvgh
FQ8vZAYjLGm5T9y8f2g2ON9SPBVTtPK4WA8YjGNbq8gUnTftwLx6VqRZHyEppIAF
NZzX7PnVsNATPBASI4r9JmD/JLs8EtCf7hMLLBlbw2w5hFXNSKZipOSYAEXCOb5n
E0hzcrLUS42TKlXslJbV+BA8Ic5F0iQUkTHd8+XUvNRaVDoq7ql5ZqfwZUo6T8Sz
pY8IQvnzx8pkt5y1oZBsnzsgYhMWNoUhtlsmAM1IoVskQeciKJZLnUVcSO2cFklE
HWC7loAIhFJLlkdHuswlo256Z0vWJdz1ZiKHKMpcEmcUvSIITGo2DlHtxReMeppi
CU6pRtw7tdOyjsbKZWLIQAxubBEGibZYV+j3a4hva9SRvUkXiN3th+EcGsndjmSz
c53fsHjJ1nvkpkILpeMWAxJPJQQvAYK8nkS0d3HTzU+k+Fwyt9QGaSgOT5qHrt1y
3T4t5ngddMgaeEKOwy1LIByC4y4HofENl+hMfrK099ESy79Ko1wz1ACI9I07d0iD
yC20UCnBRKqjmmy1S7J84MPCAqoiiRhODbICm8yq4+GXU4/LQbLg6k9H/Nj5pqDd
L6dc4JpMjQj/NSJKBgCrS2MqVfS2QJ/x3HMiU0SHXsKI9hCzULxqrT/ma7iXxKsu
AuyReF8st3bdD8Dg5udr9t9VzK1C4xtag70GMnHGY/a31v7BPqXFeh7YAY3aDyQE
7yRcqm8IUcGi3Xd9jzqzWkl/WJFsRLp/fiMwJE6AnyRZf393RrY0Ul3ExyEQRNUt
V10u6TugRRk1b5vN5JN0CitNOMhjOpBfJh09iWc9MrHL05B97m7MliNSdKvuKiau
SAGGudMQYGa6ZM0s2ecTDudP36DEE5QvaWr1aC1r1PurDD7tFaYocvtKmN8j4LJo
A1JMcqen7uTgfbTtp6Zp8lgS+yTUBLheuByoWhqEe88pAFVtSIX0xORVb2H36eQX
cx8Bc0vhlbuhscUgs2MIUm5+zELU6sn8tMlvTsaxNb3UCKoVFJgh4mEtF9BFwp5O
HWq6KsVp3s4x9bKRwF0fnpq61LdCvd6LQ0yFhaTa4pR0g7NzmkLf9sB6iwjDW0wV
wvRbWAuIzdcH7e3JRCPZoI2hlp1ivYlUfKTaPYPuFrouHoiQ6RtbYxNOkb5V1G95
jMh3tLxLIz0N/we74XGOombruv7jK0f5zCXWzdf+Q1Q6vsc4yS1YKcXOO5IYK2Ub
waNoSC7uZEeWghPsFYJxVVdOtSw5De3hwVyxg4IFKAwoU6rmNy51ZntGwJXhVUwh
VEPDkXJCOZWaypGfHNePDar8KmLLqnZOLo91OP+EsjfdpQzdmFacJirTr9RYPxFS
s2b6SKK/inyqN3ONnJSZo7/L5wIQJT3cWL0yUjjs8E0riRMlukGVaI8kM46fanWy
5lvoENwXgaO8qSBj+57oIIAAbhI8Kr9rR2J9Umio008w565d8IT3TDCiFjqonqNg
wVLlLJRtJvjH8nMTgvVxLf6rnBhWVAdnfIxObdTY/Sssno8CZ0zQ3F9uTpg2Wlu2
oyvtNGv55tpLzVbOCafd6xKN7BMh8p/eQtuUJ5JRYs3xRu2IHUbEG4w1O0bw1sfZ
Z/KOqbJTN0vF34zKlEu1maiB4ModmThnXBsQkBeBeElVtURSVJU5YDchLiLeG1yW
GeJVRhDrhxIiY9/H5B8J81UOpB3t1g8/J3YYAk+qf85kfQKvSAbNbY0NdKs4j3np
zYWOZrg1p9tIVy4bLWnQ8wjmFZ6dblGg0NshRKhhwAr3HrByCWjwt85h4l4xk5mF
tsTHHqoVemvllpXAfrdLPKFMtPCtTFpPpBPPo3ttOcZrAnk4ygKsyzIGZnILfg9P
v27COn+s/+214PGh3a6WYiX0uNu6eeuJ7KAnaci2Iqf2XdT0kB3OKsOmMsIGhjrA
A2A3y0fY5xVX/QAcg+vhk1yrpPBHX2ny/SES24mSeg4OSzhxE7Vmz53RWwo0eTrY
OJKp9Qaz5V8H75cbmgg0tn1+NJBxom68+333djkP8O3MsJ4CfA52qUEEofkoyGQ5
wFqIGVF06DzZUKrXKucIf9Tp7QCtBMfvL2fA4nuNEhHDqUJbFO5TfapcACpyGMmr
qfW/cG2z/QWtZeqecyYK+yNIp0aJ9Y25vx0k70oZIjnXi8oDgsQ7O0VOBiralQxP
S2X/HQ1+/8JhKIIg+RI9D2YoVBFpaoqV6UXVACCF0RxmUIj3lngxx26QEU7+zQzg
y4XL2x0gO2xxx6JLnnnKC+eUMx7lQ87SbORV+rvNcPZ2HkQlHMjHE8lL2h3o3VPZ
dGwtPAh9FJ/T3L5zLjqB3ZN7m/eHvSIYv7e9c3tiQpuQp2xx5FIryZxDI4XeC6ob
Ihp4uEH0ZzijTSjWD0zJ5Yjs91kSJajMkKtA8Dx/DqRXrj9hEuQ+IbfaPezz4t2z
/lkZsAhoOr3LoEfazoMzHi2Y3lV+hMzPAX1ZQrtr68K3NRmJ1qElIEX1EULPMy/X
tXqplz7qvwLdcX+0b/XkNx6v1sEZ05LfBcTpiyaZyeSXr8IfAjDvorJe9VvfQ+HC
9Jup5Epr80vfSly94V9570CD1bCT4AFOuBduXIIGVlmahdGub+M66SVn3HiOY58e
L079/Gtxukjj0DxunstHtMBpqc/5aKGn8bFDuA5gqWxO6Fr3gVFWGR7EVWmAjpDO
QbVXtrIGIRIYIiVFbNag0tLVb9qrE80PXMitwJcnKpgd1kNIQ6+2biJWGUu3cIWI
atgDtDCM6U3D5OiSSW7IQgwEqxkWjV7p+ngjIBxD6JASpQRicvi5JDCpG+j+EXJY
TS4/hh92wUopHYKAgHVVh4Ia3FiEf98622rKYGMjpMl9w4I+16c7ra21F8piY7D7
ZoE7XBsP+qYAHKyuvnAq6oDXop4FGBV2bq5b+PhT3ifg04sZNX2LZdaDk4PDEBck
iUXDflvMVDilfL/pgK17bsixIWqdv/cNVSfjel6X3v4=
`protect END_PROTECTED
