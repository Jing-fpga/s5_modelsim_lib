`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hMD6y1Z0X1FTQkp+Ip4eBnGZM2sDizKco031xZoNf6wVlxDxaRXBXc7TvsXbx3Jp
od70lC/FE+vto7RcLyT1BHGzo7FCdrGOvDmP7uYYBPoPK+dalZZn28/NH51fmdS9
b9t4T+TTOhxlY9iRPwwOrg6LZ9N0Eh5fzN9fNaSWdqyUb0XnMOKREQfiaghmIBQK
Ta5cSceL51y0Xf6GyIfbbiXItUGWyyyC4tBeYGP/iH270BHrOzTu4GaBQJ5Nm8KV
KZulYliTcIigFmWtxn3Skr7n60z8H011n3EbF0UjpzuPtbUSI5pLwFJ7ZEhrZVb9
bPADqewSfxkwlC9Dv7jaR7ZoAcDEKfrVM87EC5g28uGe1HnQoVU/qXNNLJMIW7LZ
0R//2HFwg88lmONIOcKXLhdHvfta1lb+0WTVJunYAn+COQccECdrdsALvtddEaM+
I3wbRBTWZigvQiKRQG6ZU/DXp+Y5y6AtvPDqkufzdLo=
`protect END_PROTECTED
