`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gFKgg/l3oIwG7ZsTzOLEbhOUWD69P7vqfUGoZtYaZMG35OUIp+gL95BVxpTENaZ5
Wjw8W6duZA9zYLexkMbtEUf3gk4qFXgHgimC7ydiFvIpnoqv7HtCe24UDF7Kk3bq
STD+4z4E4gY7ivnIWGoI2wHrN9k2cLuSnBdSR03GPPCyJhRHlFsRgKMO1r0i5W64
DbmX1ubVGk5AJcV2bPV4wMnQQYhWMNttbVGTuUGsxs4JCEhDbfcWQZJGUFWV6LMS
CAQRAhJ2tQZHo+55plPrXa+iro+uthVtR0d1C7HOgiU1QjQY4uxItjHr4/rw1s8F
+D/6KDoFydJstR4I014+4DUBzqGxiaHuFlxL62Wp8UGpDTUAZsL+uJsb9srZ3mW4
LOrMrAibYQncV8PobxQTUTIigJEp0WGG4xLKXHAuXYYZebZdhYDBhbalJc8MLlZE
0vj8ygJCAos/DJuEl67V2Z1jS815uYWmsmO7qps7dnl0Mv5UbC+sHe55CihHX4CP
05acWb68doTZZw8f/og1ZefCYzF7Me9q1qz7XEboeO5F3l+wznftUVjLNmSV8WPi
9xvyHZwKACeWPWHXFxmKUSV87TladmO9iMYINMHAw0o4VHj6PU2VxriVRpaSZ4ZI
FC9SpnIKbzantVMdv0LXwSBFt2LQahDIesum3/WkFf+bl/cLWO06ivlo70yhFtjA
JWsRyM4BjKO70oK2swKyMKcpgVcCQSFWi4+3p7PgoHgV7hZlFTd3B20/roRQiiys
ujKh8YT6G5mNZf3oOYUF94o5+BIdhjus/BQoESC9QXbBQO5ZppuSZhnVkZQJzYHa
6dE0Sns5yGQjwasrswbg4SQxmBLfxRibmYSdYPUf2rmd230xN9oI4tYp1m1qTj5X
`protect END_PROTECTED
