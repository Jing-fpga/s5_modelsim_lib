`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LgkfSd1mwN1xZKX9njB1mc/BMo1dL2bK4sWABYMD9AcefacYkxcE99wM+Brl0jg/
iYgCsKMBbmE+1RL+ufyYxjp/7bXyrVo8npGSZPVqg0ZNXymQwMjyC5ChDr0Ad1HB
hnxu/pk0ZhPzcPfeCo3aQc9+SBPADWSjWZK8mBjBkNYy9MrpgoB17RwhbwJcg4yS
IUaFH6cyPz7ch0StO46OY58JO3woVbRoO6asy3jJmFB2eNwfJBVxMyGZCvnE5PTs
rER0b6MANrI+hI7WMvBUM5TOk9kpzMIL/SUmVTS2DYNb9YVOJhLkSFNbe1/Kny96
/uFSWo7q5ILXDrWauOGT/+7XVtD46LPfFsTiouw7yCiGoqpR/5thZ17Ij/DmS6hA
2fOW966LKVDyvW7BhMzgppTQrvTsonGs8hjRZQZz12OTk5lh2RJX0qb5aXVegERF
1cW6rVC5Sq/xoR5hZED4C8rfIQFoh62f31+zqdLfrf0QX9P53ukX1i8Zn/HpDTJ8
4kVBi3ihS/c/3vNnO4Uf2Kf3UEdpBd9eCF1yk+09q3NOqYW2aKuDZ97X2DBPdEQS
kMpwryV17wbnql2GDi5bZPTY9NXxjSgbubRb5Uq2r4TQC3AE+627/jZEv6KXNzXp
FpPZEooRLOyvrl9nMB40ykmSp35DWlyuldvuRQ13CncKnJXvtU2T8Qk6VpNGCRgy
F1ouOAM7sPUHVtUNacAUr9BZ7cMK2bR9hKdLDLx3rI+jGVp50NqnqbY5OSGpeS+B
BthmbUIyZQLPPWHfbcQprATw+eTB74Umn3KVav/YLi1Qw2u5oCctuzg7nXpuGbeS
UItARMJnI04cRRhS7H8vrDDZWlBAc88NqmZS2XNkx1vY678WEj1ltkQF2ZV0+Mt+
3hhM6cVW1YwmuoiBVIUP5+W2ocNnIfyo8tcqM8ebwwWyZWdoQQB4XVp7uZ74q93V
cY40Xc0lNNH5AEnjI0KzALbziNHCyY+nuEcEZW0A4RScEJ6reVOeOEuUHBK1lWfi
XfYED3lE4Vw4cO1ytvwG4c6m/6UPmPznkclFSB1mxe8w0JRKyixjOBGmnoWWr8ng
lm1rc5PdChMxS23tVwAoguOKOQTzWV61/TQyywup7uAMFcxhLPxUokBHHjiNLbAE
H4TpFswUtzdsUo8KIhv6s5nTDGSEgKwaXPZytLqQSPmTi4ukCWKPCFy2GAp3vq+Q
Ehu/3S0euyRzB7q32tWr3L02AxArhfH3hnrtR1kwCoEnzEww58BP+OE6X8lJlEml
JGjtshIPJZk5A2M7XhXrmdEXDiEe38tKj1T4OsHan4CW8dTxUhnR2fNTJXL3kJUg
ua2HQzNChrTOP35q/mtqQRbuggzcaAw2LxiL/u1c0m+qWKyLphVUbjQF7bANzQAt
fjF+GAec8jPWAcUIFKY6HGuAaI61h/MGOuvn0iErQkIEBTc/Eg2YPvSAqJsvLjKF
gNi6PCoxwuL6pR23PDduj/9S0ymZdHR9mfZBYt+bNdZJKhtgYUsaatNu+wqURIxA
65bJVphQr9qwXezEiUP6Ujo9tpq9pIrBx1+cOi3y5Ojv5lz8XbcDbQYhWDCWH5km
LuDjdKdDMLZ2HnmxbZkk690PMAJ2arDyt9J3sJ8fyW3f7Ivc2domL6L0lf9AqeN7
9ACcVSvFUdflWIluM56pk4BCwKBK7HcGHtYDwead+YNFQqgOsQoKZQSfOSpc5Iyf
jv9oRThn5gMDrw8qWbt44OYYgf/PNI3GE1k/DD5lh0g1s2hvI1eo0p/8btQbuGzw
pQEerbhIJpe9PyMYhrpdnOivaLSGm3U3LWz1q/aZgXgaads5FvON3ZtpNUImCRZS
PY1JNAiUZTUxvCDjr8jpXXPvPMxtV7rK9BTnX2BHjLAhmgP4gCWqTyKSJqXndLum
V1aMcgCZM99vIjtGgo/T9CaQykao0F0xJHZCZGzAmqVqVsqYwIVP2uBPQkwuci4P
y4q4ZrrGiRR7BscBmP8H4th/U8rGkFjPz7yILvgiaGiKTRIhXeQaMngHYVemg7YV
gZjzLDN5Xx5DI9NoFxA8EDuZIb6Lp1PeFQY7znKgSaPtBsupAo82rNnrBri1FTb0
XvnZQDQZ1UNR+hfD1kU3aLoAFoCxZCSgxrWdRArCiLkJ5Q4eozBRGIuR7hlBuDa2
fSSX/Lsc7qrbpQfy26X6G9YwMxmKV7hFJH0GI55jRielSHIrB1t9qDVsKnIggeaT
z3UXL38Z9a/KCCj49pQ2ZAfSZOq/BNkkaX31T9frRP5sXapO/kHVaEUOiVD8/amt
WNui7B+7BGwIwwpIm9u7f335dPL4oBWpW3DH7+1YClDSbF2pgj1zeafwX+WM0U+7
cNDakZIpBso31vXb6rZ+hjZvPawI/rTZClA8oh4HtavMOwKr72wh71QEUjRBg6D7
RD4/10vL82LJSASharWBIxuAJ7bhLnJVxCf/eMy/WXQaAWuO2yoT4UBO3reFyBLe
mUSjPYrzHOZpI99bWlocjRHAuIzHe2itv653QGwnVHEMyLSknP8e3WI1r8hRAf2m
HsIlDQMAVVYeiBvzgZUmFyDf2PS5mzlytdkD0g+b8DuDDsda6mfxGCKHRzCcBsTz
pDkLXsJaZJKNarVf5/8GSXGq/zkXwccYSCs1sF3VjLlzVF+ZtLvPI1fneG4qeFZ1
EBqOMp8mnR+95j8DalFIrIBr9sToCVSA4pzv/NccBFsEZTLU0G5I6JZT5Ejxt8s2
NhPE/kg+MRnRCn5AMomUcBCyMcPNiQ0wtENAe89Vjabpr8QHyjinnm+bTwcHQKH2
cnS46+jOL2TD+uEJKOxGGeSU7uJKsYrsvGyB1PurACIkg1E7pMD4SqEVOEk+PhP8
qoT1f29DOO26Wr7XqR6XaUSv9YR3WeUDr46o9cj+vdXKNrRhzSJ0fOMkTbn9rXlj
3AmSix6pAXQ5aeNDD0cvaEmHZ1CxuMgK3rJzjgGcu59upfTRv4zTx250kj6ldRbu
ur1+GUQz0Zf2j0nxqqakZeINCkvs9HT4TwEbbYl96/lHFggXhI+l4l2AIyDVxRZA
jSdIlfkPdY7UT4CILh2vUsESmt8HwBP1pIKjiHw87YxV9kRVaG3RKRqoen/C9jHn
/ZcWiAKj9+0V4PyVUKroOYhZ99DaVbjucWJu3R6RWSv7UinyDVtYrtUeTzBk/8SJ
udd1gietTJtdTuGJqriXSPWG40NfwnfyA0DV+2rhuLg=
`protect END_PROTECTED
