`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MH+7QLArTiwSaFQ9Q8dQC13Eou55OTDyPX5kOJYZsfM6BZxYM4xzdKWQ29Gqa1Tj
ua2U8n2OGrQA54mhh5QG7wK/pGnJzURdxxjGd0R1Z5mwpjO+TausY7TPlEVzgmPG
+VwHArWJl5ZTEizaX2lX+uQct5RvoyVTUlgPlHl364gjf3R2ANcS7n9VaVS+MfWc
C0a/qTWZDfRBDEKEIhqN41XBkzuXxwUVC/YuggVxI2jNZRRRojAav6I4iAbkXJ0b
h+Hjb7yACDshLvpUz/5mXY30rBlf2d8rlHu9Am1tPstyHuFJHz8WJrg/+iweVRxA
WF6RmFXDrokgCQr1R6faEgZHB8ZTbMug9JXrpBsWgoBveo8sDgkpZdh0CAIvBCLP
PYGzXAHkqW7L8kk3iIgnV251pbW9RjLHNgszNMtu5Z2Q171bc79Y4INALTXzGVpH
iASsLTWqWJhCaALqTtYBqD/v3ByDfmGil1G1tvyOl1ArJK0C1QVqEkSFnWbL+KEU
bx9rjk9cCjVLzBUeQkTokzi9MbrhcXxDW8rjen6QpRgP98nDStqyAGROK4k26Mr9
wzO1AW3JQYOhInEE+N5axTgL0Bcu1cFNQUCfzTOIQoU=
`protect END_PROTECTED
