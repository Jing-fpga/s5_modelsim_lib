`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ex0pSY7EZZYyNMwa3+2nImEXLugO8q8/Q1vAR8+xyXGTQZVPZT+/KKD+yc7X+FM
sMby+KnTH4E7yIraiHx4wt3huqhXehiBFCqWI9wZ23Z6kyDCs+Pp/UIXaDCj6ai6
5a1qBJa//uqsnONckKlythX0KPrhFF+ldh57NWKEyLyhaEFG7P2+c74tQxggORIZ
Zn8yTQwE6YyXdcA0ziZqi/VXQq/rH4g+xPtBDVgw4SZkU5AayZ92y3MB6DE4POIp
UqWYxMMDzXk5iaUjYpITNavl0S/bkIWEP+d0+0RUlys7wAFYR4sEG4l9R8Lbe1gn
VhGODZuJG41Ku0b4PTZ9be2s5ed78KUusco7f1bhTfMeRZY5Ws7BVYJho/YNBaXs
Z0ckTtNscbwHDrnMtEiMr+sZiFHp5Hrq3S+sov7/8oPbQ3xzgDXLstSni9MVba8Q
SPkBB8tvSgyScKrH7Qrqg/1Uw9RGaZi/i9ARc4y8FcF0xUoRAL1HTexHsDMYF7fW
Pzsc/l+6UBo544Cs22wONDhKfUawT51nEuJsc10ZLVkv7JNUWSzKbCgNubSDXrT7
Fs8JaFl5YOxOAIEMxiD3JYx7D7wtrsGcUrYLqsSccKMyFUVFFnLUlVe+KdS88ljb
k2Au/5YncMZxOBgA/i6rabq+Y7XnVUVtl54tgINiP3uqdMM8SkmNbFGuLaBvRAy5
y++KBuqNmFH7zdNx+Bx/un/erYUDRQm2j2SXKJnKQVic0fgrqIvShkaDBL6M2Iyv
90dAlyYDNPeu/X8zvQeYGqGmi4+GPT2GanPmehOqvBuozFiOlbSHuAuLK5cqo6Et
X14q/vVaUqnXfOjc8SXm364ACR8yO1u5PSDTCA03B7egHgAAocgZ+D/44FdmmbL3
W1eZ1iDE8rWy54TLuhKFKgDSxeM3YliucE10v30IBRpqX9fckTvxofsOSw92tdTL
yqXRy4uQdQTkewFDvTnDKEUK3li3DqrinFVKnWjvnXJ8LtErMn6gV7hvMro9J+BN
uHgZVbS9mDRbm9KYpoJkHsigjQkWAEg5m2OIRo72R+NG+jphWwSENZZkHwSf7CzM
StGHIXiC5Ia42Vk/VTi0b57JPTRSO1+pQhucdwv4FqXwhRPI8TFu+PWvpWOGmz5a
w6do8/pesEGWlaLKyn194k7BHJZH/6CVkd2ToEQ9XtXtrxOEKkc9qHbrVh+RGQnf
nMGNIADC+BcJnv8KttrVyJRnA3jGqKCgKIWcHpj4s+MOMfUm5/bjNRJMo9AQEyzy
NZNd8bNWm7BFzrIeWJfwozPmcdpH/R55gQMqt9Eis42OSNRfmW+7YRNX5NI2vbX+
5orPOiaiC9fE8x+si3WIiwdGj1UTtaCFzFKo3H4D4FRh6auXocvvFdjFK939aBar
mH8ihuG8sy5lf74demhuxlTF49cbu/yh9Iym+HA3JcxcmTIARCPSW/7vVobYwUBV
Z6AT3OCF54UEVcJwSe0wBNTF/4fcp8UKXAa9oKwSquu5FTQXB5N3mOSf6S/gWOKG
51hlbcTr4edZvmYrJK4wh6DtpALLH2MM9Nmch8Tigl7cqHmnXJ5dYD6lDWFhRhnH
OWi1jGLzdrrMmX4D5CDCvhnzTdU5cfGs92jGWc7iagCePbgTEefgagEw94hPsO36
QEpc9+EK9hTob4WaDRqJ0l9RFabx8bJmlav5SRprJaAphldKk0ZKjKAmP5wpYoFe
9eDVGuczZNOjclJiVQpUjcZSU4F+YWHoJsi5ruJsDkh/qQTgpLS1yN5fBLIF00dq
tUV8ElbvnLOW+em+3ACQGivIEEwNm++9TvySz+w0Z+hk5G4qKhki+pJiD7D04EmM
w1MJ86vXMHoi7mxp8yBpUSHJueQ42jb66FyI22d4YRKnes+h2vfytY36+nq8feHj
jm9Gq581dgeuGsDbeDS3zbkuBAFtMbi0BaITJtBZ3Gekc5jln4hHoSREaVPgBn7w
n9FXdwmfc6kkVKAjzR5w4NLH+Jicg6/RHY0aQzr9rJnAt4STM+S1bS42f+wnSqnz
YVcMb5E4AvSSOzFody8dPQ/DFjeyQqlQ/Y5i3YJaaMqPUG/ucTJcY5wzqDFer8eP
gKmKqL3PZig63YFxQ7P/liGkSxGU8SsyZf8/xhgDNaWdFy6GUStFbkVRiWs1gxns
ZURjMVCT/oAhRQ0ml5FoR0Ntq4tisi4INJafGEpyIFTl1OJKnMNMTdlen59le+HM
jf8sSuS0JOgzYo+hwNiLLTdLMIibNqbDlMXG03xUllucmOlWHqkaQmINnRM/C4RS
4MrDLrjtdgq2eKFGZdYXA2SBgRL9Ur81YG/qls1m2fIKe+DT7lHm9ninq2K+byA4
c8hyRSeLO4GljyInFkY9WVITmMsP/pJULOCCpxghBMXck97A5vyDWo7eIzEJ7mMc
webTBxn7etX/ZGRMPl8sRrRzLNk6ldheL5EcZf9r0nt59nKhntEF2i3/OPM3s0Q2
OeWyxAqlytTjS/BMKI8b8zv+gR9iZSeCVlUP/MGQHB51T5LoAAVL1odajO4XJ3LR
W5KKAEpMTP/IvIzHmy8AR2UxIEDJqlFop+l2Zlj85orVb2BUHqeJTysPAiFlFb00
7/7onMX68TNX8XTifcKAbHTh9fZ6LCxgnkfY1IojrnqlA7bK1c9t2w2ZRjXE/Boj
dQOK3GNM5i2ce8q3IR4hhHvExrM0yTj04eu5dnYQdIg6oC8ArYIfX/JRYDkVmFAF
e6HSBHCVTkfTlrVyuc1fnjuadvSCs08lNNTGMsNAndCYe7HhFAvA6QZ1WQJKXmoh
BuBqi8sSKOMEHExdiiOsuNcOXO8IO1+yjNGD2PGXcJ+XPPNo2mDOX59+O4345QdC
KsJT/xP4dsMGc3HASkhzPOncVCeonO+5poSGVdXugNkBTl1SrG+1xRhjrVCeSq1U
4lEXcHU3JcslJEoo6rNwL8Zw604g2bI+MdamM4NOpdq9K6CRl6EMxaBoLjCyRVfj
Af+umg39bG+jGwerSttqyBwBPhkxAF63IPXpZh5yiuwflwK9xt+rMeGz4LM2gCN2
BWQEq6FKOx2PfBuINNN4ivkCZUjRm+klq8pPLm5wmMLa2R3jkwPjQ4PbEbAaFbNc
XVqMzHUC5m5R4yJUwMu2oNhEKBxyJ8EIYW677QJ4kpzr3/xqobeUfaHrZUgXJihw
ZGMmcvwWd9ny30lCFZiuVKn6qpGIol9xvqjk6ogV+Ww=
`protect END_PROTECTED
