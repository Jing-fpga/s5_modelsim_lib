`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Hz/cZixq3+4LO7mG4CYwj0o8GDL9K7bR8XHsxjIndVrwgSpx8tDPAvf6rTkAt1h
WAco9/bNhDMr0EfSsvF/lVlHlDfpUWDhLXofKZqFvHEoCmB/tbQPyMLXWlyIp0AZ
QGlSUJmqyAYlN1rreXK6B+YIjd4VnUpWk6UtoqMNPFxDtcmduuePG4Wm/VfU3qZp
TKL7DB2Qf4pcMrTFVPf1yLxyeY9MN3N5aeIIFp7zECz35OhhRivJppJ4QeU887B7
FOA3OkeL0yR5ww3kmCNXgvPVY/QLdCTjJus2VxnpVXVWR8BtauRzpR47GI9mp8dU
mQ5Tk9l1Z1W4H7U7rQfkkY2Qa9tD0nYqfW1Zr1TU5eVVWNrMj+9JE2c3GcG870O+
jdQBY3P8UmsWp5tRetJ8F1j6Nfld7Fq96y9Ck9PH5nlogtIV6xHksO9kg+prC+LK
scsrCuqdJ5ZOkbPkQX1ji4u9/5n3oKYJiuR4jplxZ+oWymM/QJVzSChv3mxlwVta
8zji7Lbb5gN+pNfnDnQxDZ3B0r7L5gW7/ZvjXeejm11SDsVAmOwkqH0rFkeHmp55
cq1YC++5vyv1S8kmy3lDyq15PHLRdzaez/b4Pqmfs3uRfStrCNr7yBBWDM96WBVz
7vVgiG9oUYeYd5ydAFc/9SApAuMDFWecJ01Dm34fSrlDkh/e9aDq46/Y3ep1hrMF
959J7ej8pyVbPdq6kC5Fu7bTIYVrn2I3a9nEhRXIEM3S16ib3uRPg7YcLVYqRxQp
dnGXt5mUItF7PZdZYqKdHgCQfpKvFG414YkSvb0lRp+3TDhDFPGQCJEK+S5HZ2ts
NagQG5xrL6cJyDi8P1HDIQL/pMW0vktF2ZaPdUbVWlzhyerNR44G0tqo5YaOZxhp
jxkweaTXpOTl0+YslUwZ4O379kijNTF0GxzSE9NPdhB84uSSSyo2r0s5cAAqDNAt
XUrwu5iVtFx+GFdVC6DWc6InSJHuVmiW6PRcxfpH2iW3Kz5iAGf04teW07w+4bpP
tW/ih3ngQ75Tc/0L/e59V25IUi1SixVVxgIHu1mb+BRONl8As90CLRKk2aAZdZSU
5TGb22lIsnU2xesy405B40PKLiQ7uiEsAv3TzTjOO/P/9IyEvAPflWaCGx6Vktki
hpIwCCemwDWLmwWegkBx66jz0XQTf8QvKBKfNSv+q84nz/zmjSg0WGemW5RhiQGg
DIiBJODA5zpk6IZvrZjzkRFLSgHvSkoU1StsjvCIt5RHo5HdXItcZX1F2WBFT460
ZPpTxABSfwDYywdG7GEHRhxhcSLXrzU/9/DiZ/NTYJ37B3hJIpEbQpPvYv3IGaul
Fw9hb8iivAKAHJBQVJA+CEbUpSVKxrzZPhHcVRuf5JBX7dKgOL/QjB9KG55M6W9N
ZB6q01/wErFoRv15ZsuFVnA1jRrk3YmujMYol8J7r/RTmeu7yYyCGWCiUD0EvXjf
4M4Knmt2YHPaXGlAzP+C39uHuaV6kqPMExHX6EXGONzrxf04o32wz5skyl5gWQgG
SORoWO94tGN427uCZ2zcd79HINMfqzfLK7tduR6hDlq/AnYGJW/gcm1RtwsPSULd
tG/vhFWtg9XUa92C67fOByESPQ+sUBOXMRUgBx2kRayBWm6Ae7Ynx4uSD/B+Ab85
uexSd3fAdX+ep4EYDcRt8KFsC8N0XfUvurNpYGWterxsFfTxmw6DB0f9Ksp2Beru
/lGgMfkT6Ka7m1pMVhwGVZM5ozpYlYJJUshsRhv/1N/Ab4EcpcaQ7JgYKusaQyau
0Fvs8bj3GlLI16C+SzR0KAkozmFAQJ1XdEkt+ZsN7kHlAhezNG7VkenNSm+eHt7Q
LX1lPzyGgxbUEKEJnR78HMncFEUCAQVRMizRsUDQQz5+MsYLQlhefttiAJI1WYrt
EWd7Ai2GGKcglhxeT17yBJuep0AfMLoQqCApRyJTQO7LuHkCIOku0+oglz4rzBoz
F4z75VnFnzXWmA5lef7pRUAovBcm0PWGOPAX0kzKgPQwGKS/OwwhzreyAatVGu9T
qMYz67Af55S4LguEDixLeg==
`protect END_PROTECTED
