`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aosOJkVCELRj10lKl+KN8KRx1oV+20TfrWSbt09bSjhtxx6oS1S83GxjAhPn24Ox
z060pVV48/lJcHc8t9EFMlet9039xT2/5gqi4nleYfypaTFLAWtOweOgS2gRpWPF
MfhqmmPXJESgnX9xnvBTGHmfwW793aEBkn0x8+3TaYoFoTx6HY/18jOYbOw6Nezf
+og3puSehgB2yRye1a6Idt+RH6Lmlg+5oxj4Peqyk2hn6lru277oh5O2J/xHrhEf
xmdd1bS+OUukwdU2EdeDIehtwDrgwlu28lDd0y2qF7vycx9O4j01c3QlcONM5+jI
O/OFlKDDhU/fndW1OY+UkN7OuDTZRk4c8nfvBYkPCyYZRqJJK0wuWmHSNttEEgua
MKKGiw86vfr8EViDwZzEUsaM934eCkUlaZmSAOYOE/iyoeVwDrkKNOSDLLq+PcFh
McEOLC7RiJXV7RidjsJe8WrezUWaPT95ICtQ2cDxclOCUsySs0x95T2VBABYAypc
b2yqu12jsgqNiQKuJPylePZkloBE5W5E6IhjlX/x1lld3lZhREg1mdbs3UaDem2a
B1O9TvRZZ2Sc+pL86Xl7y8bwZ5AIfxI+NRL+VWudSiPy6ntP28jWRBJAfIT0Vm15
e3rHMoD4evHx7dFlFi0d6S0PBqZjKTysU5wIV7MqRZLuv7aZXDit/kW+vS3HLvUK
SZD7jY0tfBpo0Tfkh+Pt6eoh5Sns47m5D3h1Ed/jh4ytK7BBNibQQMqE4U3HgM5O
xzmqAXt7Y52d8k5FHHEbk+Z5CvKWgdjoloGsS2SVeEWCZ9udiDyrNYLAmiJzlESF
HyH88Uq6UZ+nKzFppGHgLmVY9LemMHaZOp7s5EeWHaqHA0Cf5VmSwZezejOX0TD1
qE7/k1oqZcmsu742ZqKSa+zIY1AYgmzW6ah4uza3VTLU/EE84iXPYy3rG1tV4oqx
aV6hxm7pY/yyjHhHw53nnKgNy8/tzfK5yfuDTCkEq/TgKVEx78rK0VKS4C0t9kZb
UI5KTZsFGG6I3oDkCK5kAT3A1KZYchB5ew4ECwmk5F1qIDwJEoV/8fsZ3LI25JpL
NIDVD2Iga9f2cdqjyMMdeJDX7Aqfrbsn1dBBKuyWLK2HyG2WUvNSQ4LbtmGity6W
18u9GRYXgvoUg4w6b3HsxXdxQlwWzhavfI4jZMCpQLEDSf9q6S7xpxW/6oFHVIp9
dcKHphuBu7dY9DOE+LF1EFouqy2aldvEaD6XcLUljkGxrXtskQ6tTDdM4i6DS7rV
TZET+Z3EwfaFjya4D6yOtFuUcs30xgbxyfMaW1eT2CkCtAYBSyD43N8MOzyPO7AU
WlRa0skUvNiqTuhEU7gsqa+XH++HDI0f57vvWBBK5KyiY9xbp7zizHtv2Vqbod0I
mVYfxjhQC8/QW1aDpwroqXGVVRQe57e5xO+/g30WfXKeHkoEQuh4AzAECqlPGhkb
SZ7hZw2udPOGo+LxlUzUdPqrjCnncBfczUGCf9JTE45MWmqZERYC/qEKAi79ZZ7d
zZgtwVPHUP2pf9RVfWF3Lo2UotC0rOyVEhTREz2h30+y+WbtddBx3AhDjnQ55vZs
5FgiGO6clIoW/lAHrnQHyiii92e27J5h873Fffxa9IVKiwQUPDC0FjM+Wsrb/bBT
6wnNKb23qmW8TiHqfzrrBpSaPvg2xze0Yfe0+DKajdlyO7Vmusw+Jjxh4jAGW6/p
j48OvRrAqjZIZmBcPdPGYnGy4E7eQphNtAXX15ZYGhzJa4B7k3rQJK3XNPlb9XWl
4FhZjIGRJjBmBvi65F2jaE4Dl5MpS7Mpb+FgUSPiTI/ZJ4so66KfbdzM054U1RMt
04Vk/WuBYpsjScaYlvaTnq0YDOUQRywgQoOV7WCE0zTN2dcdWKOD/FXAcVKvrjAE
TwVarJYdz+dJyFZ02RMFAz17qdVHzk3Ta1PRfQDPtEBdcAqmAAzf2rBNrsqpE1fr
SNdjrk+5nGeeQ7CvmqrtxILQqgmnk8sOEHWQg4FaHxkWHU5XPD90oawf5qcdKEx3
8xSHkkX3EdqEOp3zTEJU8QgLZ1IcjlIBdNveZYQq2l3uTxKMxq7FI5p2n4tGdJii
EWbhYD9nzI91r8ouWHKQj/fbG02MkK4SFilzPF2bDW2YoeCeXn4amczW9RZIEbpm
cbm2dqlwjB4F3xTXgZHn/pJ+gO2Q8g3PL5zxl+rbeMLkYrshjSMhqXdHe6YXMZ9O
S8wswiXDD7EiBqLDCzewZKXShsTv1V9XHwc2N8Hg8EYtr1es2UunhwrZ8izFvdPt
4xwzz97Dnesh7mu+xDL50m6RslCyMLGElmyHB87vGMf2h+F0lWOqNHCKJd1+HGrs
emDQgDgwENrxJgxCFkjQ839R4VFSwkhUCXXTaGUV+CVLxLLyBCOJtM61u4V5mcNx
4tOxyk8bscPLHrXw3rAl4OesA2j82ovhI66ar8kdtv/NZ/ijTjBk75QnVjPTJn8j
lpgFUhOd/+n3JJk0Nbi4g2g2xxeRXWQ5ks3JIK0qaRZz7ncueZiRMHMBNlXhKe8M
6AJIOrrIMa2m3vtXqawsazWUJPp0sLfjiGClyrAuZY4e6q1qN4yiVgo/oSW/z7q5
LPMA1R2iQk7ubMdsI0u01Qfw9Mrh9xaqSOTRgJ/k3ZL5dSL03m7zaH1VfCkHV0A5
iuv5UEGCFd+XPskkBD7qQga79XPb3t4wWfzuYweHkrvtDL0b13Od2H44xv+ljV0Y
LpWVV+nSSNvk5AWs2N83SbuPvi0a+tsPHTZDHJhN99lY+RF3IlPO9TQZS1MBpAhb
jhkkmPvLLht9PpZ7fWgB7nhDtT89x9pnpKSzz6iHbifBsVP0L+XLM+W9liktl9FO
bZEFS/HddZP33xfMfgT1TgwPXp+w88INwW5SBlpRrxMRvOOwRpmyxOmID3z0mrRy
v+LlVJ80hxMbGhgMk0+wuEPcyoY3zgI5ZHgd2LFD9LWRLwyxV/JlGMf0gtXzfNRF
v2vCjh/7rki0OOFUtwHsXPQWcey9vy3VS/uJfg41UGNGzJXSWbUyj66mJi0O7G+1
raWmHDBveEHNtv7ePNJyNs1lF5b5qttlPivlTY3AXbs0XnLA7bKpXBhFRxK+Axha
bEMCl0J7EOV80DQE0bfAfyKENu9yGurkILylhs1iKglukXrCTwHt02GBdkutwPl8
iIsx+Wg9sFVvOytL9QEUa+GURUP/r+dY/pVRyC/F358g88QjfgTo7zCfX3mb63nh
NhRxAqwAOIL+uMZiihX7YFWWyixWAqSIpKB9hizOdDtdNP+jMOvDg4Nm01vQqEpJ
3F2fqdmD0DTiJLG70baMqb6DBcEQrOegkbp7dvbioSO+huqJN47ajCrOdloU2P0K
nTw+O//gae4plG4QFQlqbcnzZuH7CYw3/5QZa5VGrbUohVI/dJ31Gsm7JmbWBOhb
xcihXYzAUz4CwqvcWUYPHEyV0aRmKvf8z3fukIKWToB8zkJbegYym5Rt2TCtVeQh
821E2pfB5jEoDzqRx+ri8LptJkm0gCcoAVP505pYQgY18IGIOzsFfRf+OsWN1XH6
76GAo3VsoHW1vKwiLIpuVNGY4cg5+azvyvTAmSGsgivCuLyZnkRyCrYZGwFzlMZp
mCI+Z/IAwWO5f0KrccVtN6bVTciKAtzRTLxjXX+chNgFEaGyeSae0feEfIWVn8lG
B9ewhCcACt7dX6lg6MahO6Mh44SsRVDzzixb5b26OT4CZ5m7cCP9GwtnssmJYC1m
1n9HJ4McvFK+Zh8Ye0oGNoaBZi4cMMu4o2lNwoVnAIKNQVjJUxOVCoHa1QEhTfZA
MzTCMybdXjgelXD0IxPnICPlFaeUCaYm7L2yvoM722DLn5olStOHwUB8Nj9FifaX
QTPU2AKeMy+ndgYsp5oDaulwZRKRtJl1GLMJ2NyKxIfWWnxQxNptFTNklUZL/XHa
nEqBeauAKLVa43f8oVfjNF4tB+9lA+qjClO0sp6/T6uPmwtyoNKScp7TFCCrIGG/
PHMwHm6t56RUXt2ldLSiC8WyJ1O38cAkGyYgsCSB2emOgaoZ3lc6OhNcVFWZsD3z
BMvoL7UXoxcL8WQoj0aph5akCD2QobYMZHk5H2A2izIdrTWSRljHkloSZjO0ybdT
sOvmgyo26nLzUDBUoIU19dAFbEGmegq8uIKQeLeIF8lHGamRHIjL7ZKXc+WBDLun
kIPyq9m+RdrDm3EF+Nql3e8jp+NESHJkwqolOOTej69szZHe7o76cADWpZuJ0EtQ
Vq5PoX9bA+QtU+khHKuTCMQoroHoSWqvpA714KmW6COdcZa+LZ+NhdumI8cQLGK4
UKtbv2JVaXXBTV7ZQSSZURcyRmFDaVbzYOW+/kUUTPa1/fJ37u02X6el3PEQypS+
ucRAHBeGfm1+NFLD7Ji0a2+bre4PUtGcP5rCzHsSBMVPRwes8ZBkF/Il5XODOE67
VSS4aIMV5AOgEATJ7j4Fwqi05Q/A+QbE3n3NOKZqXX2eOnGk9w3oFIbLEu3sysn9
0KDzVzbSlJy9UWMizR8UtDRt/vPSZ3niwG/mxnGXfsCb5wM8sAF1v6/BpEI+uCxo
0qDKCgRZIyxA8yrP7ctDv+6rNNY6qDCPFmLyFmv6uqv1Mlmi0eF8fmwvNLKnWHPK
dGl+80ng5oLFhfInvZfEnHnIgJFMyM5hY5b7FivwC3nmWaiFdQSjebsHwOeJULAw
GQ917TtQWGOG8NwTccYYMtV9iKh8IznnHRv7rrMYL8eQ1jrP55xRioJUgitRqLws
emyJ6c6wknCTk7Mi73C/95Vl7Mjn91dN3N2qIEsrIwaRYOXYXRR4BZjlArb9o6HN
1Nh69VUevMSJo2wtJtvWROcrkoW+pMcP9jtkevYsZS9OoWQFB5v36VgLC0qlufQ/
O0DueSd+pyhl0RQk7CBQl5SVsAWAmmJ7v1GVU6bm2B8i25EzOdjVhxSpSknQiYqP
60093OKXrq3Pgyy6kjyjBaTB20XLi/MOJVk84N6JFuNGwezpsZcGcR6vjaozi1Iq
NccrVkdiVGBKmwcc2Z+YvHQYjHR7cyDvO7OE04W/K4liRx3vwoEHivmN0TIp+m6r
+LNlM2jHQauthyyi81c9HojY4vE3p4aOndKG/t2NlEFb9GGYwZZdQQP1fFiYcPSh
V7xQ0ALYPpTYsFcwOM+fcvTjO85L2IpiAhpJB614BYIBpvtM+wUSDst7BZLY4oFr
qDjPVUDkw6ke4aVOwHzR0qAWbPrAlnpb3+yxIK4Gg6QYws1QL0IMBzUmwRsDBC47
Q1CFQV6xi1ODV4OS0fiPfgLjSVroM3+kWFLQxS8RPUBS6VnikiBjAWxzgO0s0hFM
mE9eQDdmIia+OZSx9oiwOdM69IuNM4Oj1lGnMb+49MMPB48Ndtb5gX+CM/ZWV6Sx
gVaDvyASgZ1iO1qe/LvV1/Jb3GaXdNg93DpZ8r0ILxFNFh3dMydikRAqFdiHmko3
HrcfdUSmTZTwhurToNPly6IrJOebPEZsOdp/JkBCvLfJ5I4yDSEubXmGwC1JBu+P
+u96Bl/t32zqozY93P9HfFP5mCfMv+EBe3FQGerPJwN3d56a2fklLHafwuvd8uJ+
VKSwDL57hD3AsAQfxfON+ENAnToe8uFr8qlyXRx1YRDXP1bEqPEgFNRJCtHUjdcE
n54mQy+LVmsh6BCiyASp6R9y2U8/FXjFxwPDvBDuaDvHC5gheWdWwu0tORa3j+7t
R70Nrv93udn16LPMS/OT7/1DgRk6IAyTxurCK1MIsJ/JG3EUkIioJkuMbt5CtnZm
PQD/z8oOirQ876VRI6CLl5k9c3ypK/sgWVdbtzm+A4q2kLfhNO4UgQ+0EP6PAVjU
BDGVxc3MfbDgDqu9AcQv3DeV1pgzEfMR/KdCWnk2a2RvmOpeDcQXwfR+m9N1ZSiA
0XbMLtYRPenYUtUe2+QFF2KxCa+btN9/Ke+kyPWFysKSsbzN9ZZaLcLRtwRpRtiQ
RMURLEYi4jjN6+3NeggFuspDfYIgE/GA5QVc5C/uwcJIeFRmrjyVGj2twQEnDRke
kFhQfkvgywZ7xYiXWBsWDOy1BwkHmwqtpiTFoR5u7IV2U5Gj6TYlxJpTYUvHEnER
sqO/LbEmVJXaXiGp6QGoyXdXM3T80KTGjkImjjqg8A3Z8GEAS4Fv7VSjq/cxYD9H
0yvTF+srUboLkHPVGwc0Dftt4ozyC/25ntFYUVBRsMxN+zTW4jkKB4UEqHvppNwI
ryQA1+6BM+xdqaXp6QWZzZY4ujET/5IGVlVIlIymCFD6WIFx222PaPwp5z482ZhE
+bOqNZ/MpC5yV7UzLO1sgv4NMw+H6N2TB2bWKnwykcX/RUDn0eT7tm+5NAI9hPUU
dmwQvtMdss8/0RjRqzh9Aw/KNIhWWeJEGMZpyZsvfZbfq2L+VcO09xPwohxHnPoB
y44ft7hNlxU6ur80YS9Z7foQVc3zMUSBugqfIabtFe48pohaT+hAKyMq7bFDmr/5
F1D5spZf46GLXKWNW+twCDsGIesMECzjtaxuQPvUgi45xpA0XzN/HmIM7Ir0Up5a
2LIQuv/1r9azX2rArJLOAT2F9yWblG5ye2jKgUNZEzJTnXqcv/Es9Xm65dQGhN/N
IQryddwQj+i8Bea2MgVuDc3YNAhhSqh5ao56zqFeRktszO84wLsWkYfZp4w3bvBd
sGMYYDa2DqQN7zsFyW03XMj4KcXeSn4LRJaKB5nmaxdfbF74lgmNy/36kzcAhNCn
zbbJRjDpMBSkvwb3jt7by0RX7Cjrk7ZJ28FEfPMY13ccBmwQMiPo6h1XdaX63Cvn
d82E7RjTtaXirYS+PshEEfM6rUX/yD2WpDk38AINOuEfcsOrnZQDaISLN+cnWlt7
NJdDWgNYL6rsFWe+U433+g==
`protect END_PROTECTED
