`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JMTnf40TV9Ckm34CgZFaeB3rOgqMpD5BogQaFl8IXbATmlBNjULi3MlmO9mcUOHc
woN/g2ht2KSXjWZAk8DX639XafW25EBdl6mOhKZmuI1eWpaqVcOBdpYvGcwz5q/p
GJyFhNglQh4/NQKYafNNhVzguA40NSgJGc8+07Za0gMTfWvKgh+8DXi6ANrhfeeB
sHU69rtNs/grWzcg/QJ8L43oZbzQQG54MSuF5TOdS5KihtSi/6DPNhh47CZvOF2z
IGZQLv5yshi2eSN8FquQTDbRRW7Q7YhIdAHXzbbqZgYJr5jrNT91nF5E3h2/C11A
FS2JxFNsHh9OJjpowSUvwutaNW9DulDKdH16qSrxG8ZTQASawCLcVtcwEyynnLNZ
jHJOQ+0yVX7keMDDFquUpqPvGYSsaN3AQvlzz5xQtMU7tYWGFVFvghL78niZ8J3w
/BC7YViIlcEOT1tlOPQO2jAOi10ybgxGopYDJ+c4Rzw=
`protect END_PROTECTED
