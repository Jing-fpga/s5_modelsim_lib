`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m4i0T51EKBYhvfRoEHjUkv5SsNzFXhoODNoEFC5od4u9I24Ml3FsoNonLT9jjpna
IAvBxUig53sXHcxD5g5Zf7RM3s/fDgEcM77W5yaYnp/3tEX/3kqZx+trcGCmX78U
x8Lj561uZz/wOlm4WObRFUj8/V+xvs88XDFlqhXIDxshoxlo+sTLf0xMqzOXIGsJ
ZbJqVXj7ojLDGtgcvSe78PF08ivm1nYKWpQTXEYcEjTJHEy5CIUe2dglbhgu9DcZ
e1teqniG1c6a6KuU3WzQRHl9lf5ycFbVg7jzDyYGXSyLHw+MMkAGNfuhfDlfEbvd
iq4t0Xh6xRnJPU1h+IaGc0xq1mXItHzBhYRO9czmYYpEpwqRUgQSyaZro9F6AvmV
TYBpcM37h8SyBfg7RfVyDN3qmhSusGcKh1pVtdFW9dXqupBOkpg3fJDvPEWVtXen
7GX0RITZgAL2hcVVSyBI4YIeVCMijQv/72PobmvY3/H7BbUCqLV7FOP4Yza9F1mb
FSfmLE3+nTEyofMjrWNX4A7zL+xDog6Z3gteL1YpZm6B9WSpbgDLCEYAtVDgjNS4
n+RY00RdNIN+73DVfI/vYrNomMX0OekhmV3oW8T0yO3w3VBWZdVuZiNw2xsgpkSc
dE0UpYRqkmf5h5XeXox2ypuEWE9jpn1dHBezo0mk9MBYwg45oC1FVRVcGLLAOqrO
pZAt0dGA+NowApXB8dKf2mZ/D8C0h8RVuRNYGtYiOgK1JFOS+59KbrjO8vwNxtQb
cH42+C0UO+DfhGYqh5MOH0+3c5o1He5lJWff9Hwr24Sh+Ka2EX8G83qPv+axke6c
x4MKiNNffuR16gjeqNeUl+Nur1ROq+w8qxnky/ywcQZBb9jphEW18X7fDaWNYTOY
yFCs0Bpon6rOk7iBI6OfVgnZfWp6YJT1V4XX5tNGR07IR2gMI0PxASZe1Vtj1xYe
TNtGcZyI01genvmzgYqVkq9DkivYjTWu4Wd3AYM0LF3693uN/kMYKUAJh+S3Vf+w
1HhEnRl0QuOF63X4KHXwK2Ghpbj5eT/XYjJvhVHeX47XPsR2JhDNVom++l1DzrvL
YBecDomYro29hd+h1aLvfyP43dPYZv6icedxgVG1pvFCuoSXfkgMlkcdEslDQAVz
y8mF0+irc6BdBIIq+YiZiE5YIrHIMVvIXPmOXAaNt5DtRCgd3bbdrBiEKICxBE9n
mEUxYWKTqZKfeMBX6TKSXI/T7M0pyA4RG2OeFGaYADCaJHCxRjYdI6rpGfmiZFHW
NuFiv5opw2DuODSZihvfdn8ZVyW1Y+G7mr7pgzL9IO7uv4ITyZ/tpM/7rU2dADW/
UoQVmGfrc4tmcgAp6XZ4zDIfFZTvgdk0rDIKzu6UiTyXgupZHaxSWAvjDTweMc7s
zuq8w/Bo2utsGpOQnLPuf382zITsPahaNzfCc3oq4fZ/wfmpTSiJ/eboqwEIfOUN
pxHAgopTw0RxjbWw8Z5pnB35s6hQcp4Xy0uMneCMf6wZAe3jd+3Lzc7yoviRMfXO
f0ZGAJEZuFuQY0a1PjEc6OvPqyBIqEEjKEj0GtSyylkuPFXjCclnklmVaKIWmX4/
TSe6/MXsXpVsbdcYfew9M5BU7yUxopuIjrxQaiiip/rwxBN/61ZgeA9uZGN81e7R
CsO5rDRzc4LOWwjiZc29mDotR356DAYK9ZLdvfwgkzbiG807sqPTfuo4hbxfvxrx
mPGXZ2ZRcRw0LClvdDYLvE+qEWwz4oJpnSDrJjvMR0fvJK/WykavOy55ku8ECcUb
a0Nrecelr6qBnyMhDhFV0ZiS+xnSdrfdqhsmSgVG409qhCq3Zh0agiBHo9RBDzvR
xM4DRZXEz/Jy299ddENUYoY3hwHDmGV3PVtWp/BmMpFnUXtEnDl/kuITE+CmuBS3
lAcOrx62h9MNCNmhDdo4jWFo/vCnaOSXmcWU2/+VUwEbISKNFnnN2PTlhMh+8GtO
aTydmk7WwNWYRsvCPhIwfuxerWT9676anFDUfzPR1xK6R3BtaR7lUO6O6JmDMoDn
hsKBHCbV/WBVSEPALuy37/66Z2JNOVgZRUU+khsLdy6fgeNDPk+tWZV68JIsAlml
3qHaOsO1Agnez1kKkYJIY0PcnJ7RQEA5jGwvAOB/Y8rKX16b/GBmYlmvz1eGKisi
DuIPngP2acrl5jXzi+hgr99PocRAkBAm5+NNbhBbU+H0MSmpgMXUG7V2yVimcWGr
uWA5DQ/lvLarC7RCLFPVXe1Qkn7aSa1snY7cTQIVDShGg9FK4lKEEFgunfYy9404
Z4EScp60Lopfg8wHQ8DY0au0C8XlM9pFbHR5pUxINKPACt78WqHdL2gSZTikOrMH
L+U7aVTbF2qqf4Vwwz4D9W4SUKscsToVZA3onAlt+89yMGBe8LmJXAqUzzUU+fdh
iIxAmQSdG9l+Lr+gr8iN8kVFUoyxEUFnbles/UPaTmdBqVy6I+9Qb/MVDB66V8u7
NHhp1xt4W0o/iTuQtxZtNl2we1mtrMRMpf4WqWscWZEAvVmd1YTc6DVeLh8aTC8U
Hb4GkwkuyBXnegOvS2WOjxEvxXpi4fBRWif1YmPLzXG3N+SHfpFIUArF1AJeOezJ
wjIKrD/rZZ4hHrrRCZP+Zp3ta8eu2Fj+cSvZ7nWoeMx/PK4+6U7PyRi5mbHideSs
0cZN4sQE3zOzl+JVKbQDOBjbjm/k4BFo05S+nagXhqpS9xpevmuOps/xJ9ym92Yc
GbZhMlxP8FtcQppmodTShQXE07scaVrZdOotMcLc9/y4BlOY6Mug3Cv/y5ma+zpw
QMsh/JeXyWx7jlqQw9p6k+O7utpu6GulUGIvklwFGSHk4+4jcRyKAnRLYw8k5X0I
H3GZmnCRtg1+OSOGdRsf7R64vGVozHKuOadhs0VMLP0f7/MLjTexnMbe3NnBKTyZ
kzqSceHLdoG3SJ/ATA+ZhJH3acz3GuEVhPU/8V1L8X5zlBEsNLXchZ0S8qWrIJwy
+NLvBH5VPHCpCC7XfI6FvDkVWkIUsK9FnMpco9pIkec2X3PvHlg/5FzWWjoSdP2P
9NEtrytKjGF8GZYAXmlGe8MAffQaYYKfX2ZCD1j4InH4iSsZmK6eXnKqenEqpqrl
udhJMMLzQ8ipMGbABEotYUYvhGcNT+tJzkBcKXiXV2xw0d4qNO69PZVdfXPK0Lo1
yC7vXA4jKalje8RO7w/C510k5C+leHhfTnHgdAB6uaM3aeJqsvS0GsmdmJE1h42O
1/LnpwFa561uYb12byNYKjNioqqdv3xDOmzuAN8xIvNbH4bQDqA2wXpoFA+3qD2a
ud3O0hY/TF9OtbG3kT7rsQxFhM3bISM9d6/UMZijTA9rNAfTe55Z8HnlqXbXj72+
plad2XlK3V90pMrQ58Zan/pK01jvamCvPQ53zEtyqNmcpAZFjr7G7pyl/RZpBDGr
Xb7vBFhX7HKO0FLzuTVpSebSiYO+FJ0dGKnB/GXkYuL0AeZjleECr2Xxy/W/RgNu
qQa9NXzg7bhImw4x7kPYcW8iSMt8pqE05XCNb0ZKC1i78F/MBcFzpywQGlwaRjcW
uIoTQICexgPFu9D74rBgiXQyPv+oeTtg8Y5ZGu+suS9ZhvwvmI1daGQaryjg74Uu
Xjjg+RcxLSADT0v07yh2FMrx1TQdYdIRzWwqEkehHTZLfRRiKaoa22DVpSKRwd/T
oQiaUFp/7KXAUYzIgsWkom3HMiwNtBxtOJfPBAe8kntOBCfP5WFwHo3D9Gjj+fbH
Y3+f++vfyE1AkDUeHMlMtz0KiHYFMw62iAvelyNtRgxqu80OfhV+ue/CSXsev4j4
GvKQSJ7H/fqB+Ih/bgjOTaB66REHtna98nKjSfWlLCRdBR+2BoBtfIBoh+SqPxoW
6nqvyM5xYKzabS9xvaralTM9fhX8CpW3IPpM3K9p0xiUEUD9Q7TimFFvEHrzduNc
ZrV903VHLvRvwTIRTYjRXngyreb5m9a4tp+Hm7pPST0J+v1nCJa59YoXTn8aEdbU
Qj0r2ffwDEJ3dNTCUovGdac/6XR6OgRQ1GC5lZVEjDvMSO2mLp7a7H930iODsM5C
MM6uOhP37KrKe3VEiM4mjUq6IkQNUSIW0yoIuV4Xj1lcFI/jqfzCNsmyDwpPoDDA
BKnUMjyMk8JIrJ3FVeQ7CuZ2bQ4iLu39acgxurqhuN785udEZ/6YpNPfis3sNuzg
ZewdBhZdQTgxN0qpEz/hbel47962Z7cYL8Q/1wwzP91lEExTuCOueoFAcomL6Qtx
xmRU/l4k/ddcRrwQ72lwJv6JAFZspNyxRYOU6xH/CYo3tZQtA6OOd20S0mAh33tH
OzS7s1hRRcUzgUgRSumPK9C1YlzcBZTRwF6zWZAGKDWbSGaN23NxGKhAKPVvpB1w
n2RmlgwvBqTzp2Fv3bKWy3oQSyVPTd3P/A3bZ71XXO/QDJIO0ZwxHo0K6wKR0/gE
7OthmbwYnNedbPohWWfnOSP9vIYPKJ3YMopS1zgN+DqM5qfZ7M/BRfwUfpcR+3U5
9PesulwIeHRkxUbQEatwYOBYGwepJx7Sh7DYFXVI4WVkaXcxyaf/Rhgvm7qV4c1g
6Kin6yWkPt60fvg8il/ack3/2x1/tUaXTwZqOhMG05IMUeNDNQziVt4+PUzYIwwy
MTvm6bWuEg/p2yD3uKFxg1xONY477mtTf0iilj6ctuxDtlYsghqtucJwdtETnNDb
dE2QjthfbibYbehSzpkzxFU9fnGRPQOJ3kLul0itvVq1AKG4Yn3mB4YzBIZBwGzu
bE3V1oIeux1TN5RiRiCQixDVq6ZTkeXz97Oa6zIJkC+fLlX49gqhek3zx4/8pn5b
QjbDFuRg8QY5SAk2WTt+lasFvj1GBNoEDtRQtaQMSbglek3WS90Q35sWKqmBdna5
Qdqgtj+mp+0r6Nry0JIi7sHjgHSqbW8d8wetVO7DQ0vXQccziSGYiXoI5Hk3ukPH
Xf/F4zTMIC1CW7yH2GscNzNeGk/oTvI4ak6qJ2GKg076YV6VS0SJmm9Jp1JBfdVk
6pLDtrrecItbSu3Cpy2EKvclSBZ+c/PnwK6GtggFRhXrDGNwH/yv/ePEyFsyeidz
ahxjUchU6Sfj4bm5qXOQoYrCqzUuP7t3uzbfTCrcz5ulFEBWESLZtXJsR/Bu6irE
Nb0qsJ9Mm2h5nMYFq0UB0EpXaPFsJoPsaL0iIzDyufd2AHFbPDjmReubkO2c2/jy
+zLGR/1Onnp5tXKXPCAT4TBTzMTeEYCAxM77iQQUjciRb3ArhhoFpQpWsKgD0BCE
y4rc31OvSS4tNbwsc64dJ8iTWKJ9uUfHGjEixYktW+D+RK0wbuGr9BUv/968mncM
VnbOMqs53tnIM5/CXRcCEUmVYv3R1gOqiECM9uDysvPJ2qYpMeXkWAf5Fgx/PzhB
LY52ER/rSi8Kl500hEqolXAKvA5kHKHd++sux6K6rWqUTFcuAOaeBR1t8VcAeH6m
yUOI7McdQw9/JL3n7Z30bP2np4hSnNcQUUlyk+ChNHEh9RIj848xXO7pl4C3pyn8
TbRZIqYmmUEY/TxZDpOpVcBrnSr6cZ3dqO/1xEPRqHutCv2eXz3g+UMq6Wu8CJF1
O2IZOLK3tHaGy3i6912Y6C7s9sPBxm1VssaFx5fPdJyaGUM73+Gj1UhrZNzSCPEE
6zfKqW0Q2O3AfL24SHSO8/QM/QlcjsZ88ObhGZRX+L85TDGcpROq92eAFQdfm7mn
8WaIPa1CGrVquO7reeKnsXt0MfrHkRXyJhBexr5Ze5TFcjEuyc68fUjrD/StEq9W
TioAWk1cN4AzQ5nG7W6WLHSTKj5ftMznJIKWLxEdOHz8QDttBd6tx5kMuFmMpI0i
S9XJ1pK7HZEgPkMXeEOrrGK2oy0iA9ENGkmlauzIOO062FY4NgOseKvWSzGWjBiA
rkhKJp/RiFynFroins1wcoUThoQEowkrgjfVwyJFlhnQOILNTcxgpUtwYMADoLSJ
Ovypzwstlht7bf+WMTWbLFoQcetDADv8IbkOSCBCW2vIeqjmq9QBOs43U5jGpBnR
I5/dHq3mPQx0xcwFTz8DfsQi2Nq3sFwL7ex3ICRa13v23KeTaRoGJIHXEe6KXrsL
GdrfTGlOTumCDvK02sqSATZY61bU/uryRlQU+OmPfYdOPzmwJ+sIvXXUlJoSHpnK
5RapofyClF5NjKUnlDSdVVpHqiCsBYfJp9IzIoMNuDt8yR/7tMbjtcui2V+3T9II
Nuu+pQ6FODvDCvLma5VxdRcx3brA8DbccXftfy/4cEpsfS8mEzqvZAEMpreg2qVK
oNqdyW0iEWnDGixLCRWN8dYsongITXYtFyM+aayMHDKxXZMuNkhx5YgQUJzsEwQ6
W0PPLdFU9QDUH1jNII1xkvEB+3BvsVEuA+JsxcpqspcKPd6PGIjgOOVKqvOkdf4q
CjSLKTX2kh+Y/ZkGAHsVBzaXj+UxdxffgFyK2FToghlkH7yQ2rBo3Z4t2uUFu2pl
1oRB502acqL/DfVdj8pq0b04sOlRhlXPkc/5mtfabDCg3XK6vJuLzQrA3r0ua0Wa
2QxziDT0ECKUl3SK/g2YuZKMNWQajbN0wMsqMlnJfkMdKfrbwa9YF7clxibDZnzI
HNh9v0cFDGKE/UtYjvjYVuUIMkK91drYP3MoJCC1MknqkSN/YQJm4qW98Zx5lLHS
N2+GbjUnIP8+BEqI5UDm/mBvDrwz6Ykdf3NfhAbeVlZPAFuOcq5cmEY90fE9ler6
3pFl2C9NcJcUgK4VwDXRjpEecAMq3+Na22GSjFTGEEDNzYibPo621SxV9mb6heol
4GKV3Xg88yceJPcZJg7krzWJzgnBnI2gHVh2YVu7syjx5Zp6pefGw1RiiRHUKEqO
O2xMxx/3fR76BDdvVVasw3bKoWMYdoV5trNAZPV+VrXzrkbt7jGD1D4O4iCQP7ug
OHfFh4gHGL66UymGwH18Rol/yT/0wsWZklo57vOgQAiVS3sX+6VNIx8+nOwiIoUB
fTOTFycrt2oT+6DFsU0WHWEhszjTZmsMjbTd/Bs3An1GZYpjbyCLKL2nqLCwSYSO
RDKUnle6tayG02Er93jqlX8ht0N4G6nA3RzlHR5vRss/XwG+e7FDutIxtfzsnyon
L7zafwdomWd1qc+1EPModABbAV48quNQPPnO4XnL2M0WE2U0qtaedYtl2HQ+IQca
XFEVE2L0n1XJ7oLBrpV1krUHXyswuljSsWYyOC712qcqoRL4uOMvmivoqF7wO/dq
4T599YHKaRU6rmX0SG2aNHkcvT9zLBXw+c/LBAwvHl8REFeuXfC8wc66gWFaB/BS
G7lJv5sgpakO18f55/XFRfGcH3Sn4hdYjCfGE+0+NyH1rRQDCaESwJubJG0ccCOu
jsJ2l6wDPlBNdIRm6d3hCXMInUJf1utwsJHsyNgv+nXw0q6hbJff4iJ0hAdqXnct
xB8TkIYJfX6av0rKuVQ3h11YJSQShtVLLHdecfD1RhY1fZVVL6eFS32Kaer690aD
k5TFVwfrBsLwkn4ozJ3lX8wmpSpz5dSqk+rRVwNT/gVq0EKtpF/PID270yxNSamk
BT5zUgkoHVHh++JXh/5grFzz/LT3S5ycqs5qLFULHKRpSlE9x1pAKX3YcRHtHA4W
ry4Ga3d5L6uuOfbVS1hEXsXhoP+tuVSNDNzjM+VaZVm5sMZdnRNI9d6X8iABnvDL
OtGsvlqoCKBAS+pPCXwg9gzXPaAwNASCjqH0Eohui3UGbS8fU9dEqOCRjyH44q2B
cI39r0W5ZyJ7vTiYTsaM+itDzwcVcu3+rlwXzzuD/gUvlVaoiC54CoSRBIk77m+0
9HVgicvy0zqYilWDsseFbm6Y/9NKgXLG24/Q8etEwGSU3LPuqDM0jzOYFdZjTEHX
fdO4yHbnlw5sOrDN106c9csqPU5ZSmALdlqYPtAsWxBwN0HrsnVUmJ7BknuQY0GZ
9tr6rtXE82C0NqUhgL528UaL7vjhIRDQVUmAPqFytD6Mkk9MxHB9r8evn/8wDoRZ
oEeKinqCSEC7vKh+Fa3k4iZZsq+0Yvc5N9RNEtZ47TIl+kHDVV5EAcLClIWne1qJ
k9rbqSGdj5RqnhHFXGDzYoC3EKiTRyBOFit0+onODaeMxyovkXmvEjgp6kwYkeWo
lOtD0tddAZOhxjZ4w8urgAmmrZ1+vSCMQyzDzd1JRLxQ0+iunen5cPRQDISt890A
DYDHkwxO4OyYGzhHBBj6dvIYqQQ1glAKNblpIovjkHgc3iAiwIdL5jLIR7L3d+VY
xh1+Y2NVAn6lZHHkILU6JJick0lN0djVaWvwKCVyHeOkhKS+6k6w51bHbpmpbaKK
ohEI2ZRSKjB4XMHrPUIlUwdIHyV76kF22SiPhyxv309rBLZjajIaQxfJmLMY9Bbk
X/6wwf/ZMns4FovVtpWaPu5CEBu2Sm7lvFDvoWSKenJwEjVwtdhtY5KjnCj+Hrkc
APIg4Ki34jsooIeLxfOfDRc1pygJfqu28ZRwL98zbRvz8B+Bz3dzXnnsM5FALFIH
iwrk1z3QWv0qjLD/dx6qtO3e0cEbtAqsdIK0LquqhD3kjddorDim/bZxwh9V2l2o
bwSUjnHb8kYKVRGLQv0N5WQ7Lovyld6J3NrV4p7Wjpt6viDvn8AbCz2IaLi5GWpM
J4eDseJxRU9/ClQpsE38v1P4Ep45hkUMByxhrKdftt6d/fVZG98/NdxLCj+SAYB+
AeviSq/8PmMGRqeLsuwvoIIlRBVGfNFEBiVed4Smm5p+OH1gWD8+sm2PSDhiHPAW
sELQDUIKSFQo6y6O43fC5YyXOZJlPmOq2GqzLr4qFlvYYabN4xiETAF5+gNUIdyG
YConvFdaKIs2escuBWig33bJcWtPfinOZCiSEeOVz7gMRJGBfPzEHG10Pcq2AJh4
UMLHWeL6Il2hDulQSH7EOBs2ntT33ZLZsF36FXhJxGWfG8Q0pZy2/kFSRdMkqjoc
fncfzsHFwoGHA4MNUqd/VH8dFyR6r6OU0eN5VaqxEYNY1GcpsYje/teoXM0DwWkK
04GPKJLRIP+vcJs1BHLByoAsIXchi96BWwjLQ8F/dFcaXxWJWay/sb7AEvxScnQ9
uuBNFDNUtUv14X3iLOIPek00d8lXU0e4MB1GM0/payEtkfW8iLtQRHx01/epU6oC
m5mn92YMTTWEXTVo/IH2jlagZ95tXum3rowd2tKppsIAme/HXc+QSiF74ZWHgvru
LM+C+kuuSo16Wyq44hinagKDNnIGhWyKoPKlScEkBoY4lYCdmu0bRNeAQhzLTSEc
mi4mz5lGaVjrzPBXNWvtrEnrmflsoYi0gJ6KCLXqwIeIXk7dut5pms0avwUPsh3m
bnrzdgx/e4wznNfB+nRKukalUpDpu3N30JoOxf1UBzIjDoHYnxlqwBnQg53Akrrl
s6krmtJIAgkiwn2i1+NqLirwI2s/RZQ3el0mreeuVvz3REJCe3w8RT6+H/z9x0qP
AOW8nphLnOSCUiK5SbZb3rTN+pcZv/GRCoIfvSANwT5TPGUz0o+YtrJI9e9xWYEh
Isxv+13jJgp7Dyc6NKwWo3bwvpRgohiurQk1S3UZKv6pG8XgdxnEAch/XTDKwu8S
2SuTBs6qsOy7bIuOsp8rk1B5swCyImarOt8siFrbU8F+YiauZVD6doEyD7gjzRcK
0ih3/Mq8onKmYDbAa1Rz2AI8S3EDPAmTy6ir3m58URRKOMsLBUZW/C1+x6XDF1j4
EtxGjdQzr/PRqUxWA2FspzyXuONHnlT1PTX1kS1p5hnYVsLSQepEramJufjkEhP2
duHuBAv3M/z2rEKDQOhioQyEnf5vizlGI0/51tmx9hdj3s5lL9HfbPrgg16UmaTt
9G/ourOTYoGeuaapg2J7GpdbVwrc/d9KrysRi5AuJ+7FlomiD727rzPTeB6Ui5pZ
1crlj+Ovupya3EAS7sEDSsIDiD7kLYWXSfz280dCexOWtps6kxSt3t2Ivc3taaVu
ebtl7H5JeuRSs+ihqgc8fynu23CJZLclaBelKBwcKxDHmJUyMgi8MjWfOcUCcgFq
2zFA0QzVR79CdUcp7B/9D7uSiOwCYdv5N7n1bDHH8xewJY4Xp+7ZT/c4SMqNpH/p
7AY4PiYHdZieU8yQpYKySkXWU45tNTWBEV6iWGuXB29ep6K0rmu9jfvKEoeBAKrU
MRhYoZcgcC0ZKtPCdzD5GEcpBNA9ZLXTfHW8Kr3YUrsZV2af4+5ePV0gO+UZ9Yll
kLGTL7Z6uAzAtqpnFLoB9O0IpTkD3Y5/ghbOLkeqJROKMqJNZBlTr2nTK3aOPhpi
0fEmZ/PsPJv+MJmPsAI8c9Jd+wNJdVCBXKDsmPIsGZYL+sh6t2RHN+J5Q4iBYbEW
U1nSw8YP0JFF4UaYZp2E2qNDA/8FiraPW1A6pf1X5jHt8SwAkgZXxpjwaWsY6jrp
YhaNjPWRq0Bkgc2NMTtqMPa2B1XX2LoS3aQy5kukw05ZRNQIKShxZaFmTj9aR7Kp
zkHv96B2S12lSmOS2RWnGW2aj4iXoH9loBVt+KoNbOo37ZZoxUH7+rLLk1NTDMVA
T5+XZzDiZeHsTI8OaUylQpRpH1MdtYq8QDDriCdmcypa8eIh3q+96ezq425CJCqu
aXZR90brrclbvfzTl9acfVMQh8iRMzbGiki8/LT7z4i56foCzmo/DTf6RVt2CmmQ
aFhRseDWVV15RAwx1zYNJT6cPpVxD32lqhvROR1W6ZwYNTdwu0inC7A6sHqACazZ
j++c4ttNUlWnCcNjTaw6CYIWNW1SR8rKmnbRC/HJLcGAIB2dpyOwqfsX3D546PrV
GiQYGNIlgOSvxxaNXNY3YC9lFoSPMWRT48xijHl+5aVE2RQazfIPxqHWH+uDvgJ5
Sc16TtHcLL6P1F6hcQqtOlV4oWVwQqCRSn0vvDZjXK2ZeeZvT8yx3fEseFOs21g+
kBNCIZ4wwT5GUd767M6yaXXYNjcn6kFEmXQh+78KyMSCG4lGI35a3ZQ60aLJg3ER
S2fjpkKlUPhFfAwhCBVqH3zvr2BgiqhtqDC0gZWYTiHy7BTrp4ZaedGPQmrdgHwJ
2SgCU/ptZ90qx09SUObGZeYX3qesB/XKYAwrtqTMWXmJqfqKeCgVbCKzwfy16n2/
a6AVvc5UMUtaM0KmbxZFANCW5DITIrrrTUX19Bo8XNOHx3/E6Wj0lIvAZjfmSxTB
ZE4xMhcH/2CxhEJVLEjmDw69tulnVj8gkNvoNXbJPXHKBVhejARKByHlsr3Y9UAT
ZFnQQNdvxM/xAOZ53o7sfB/soc/WK/+TkjAUl373isLA7VaI16lGqYjbr+UUiZ7h
/Qt3W2biT+DmAWBZV3NapZDTAl/ZQvgwbJFE9b8OjOjjAgn0Gh/tCoDiMCeIIqda
Yl2Ums1JZmClF3j4VSXgg7Oa/I4zu+pBcbbg8LQJ4YQJNzXRqUBZgUrsAvhtwEyv
tkWwqG9+HhgUJNICUIZJOyLjoXUwOXwsq79hXcFPWn9MUPXqg0U8l5eunvSd9MPu
uKyaTM9E2ZA9fYSMDLMeQ6wx1VHiGgdvH6s23SGYNGT00G6VZxf0aKYVeFNtlu6O
y5wm1TFxP5dvdCWJ1WV/BzPDxpzdU86cpiOMElvvwcc+3OnVO5vRWwwkqFQ8WmLT
HDZI1BR2BqgTeh1ZZCX4NtdbAPGT1wssM5xIgimqRrcTMZ7UIYGsR6gx3cY+MdgD
AKVW2x0nuFC9Y9SjcM6X6r5SG6Xdsa9Q6E3GfeG1YNX/uhR9aXbou251Wn8vXuQe
mYuN6f9kk/iKS4Jj8RwJnNhU25IyjkBsEGS+IPc2iAB+akvHm7iDwVjLr/nNEpwu
l3fZxn2sNTv0yItqBDoyBDl4wJB5SH7jz1J9HVagATxVohlslisza7dxn8VfisZ3
dc6lzQZnm+m7C6lghoc/vcy2R0qF27LbH0sECuU1QfQ/lb5jjg9mywJhrc+DzZGh
YyI6Vsguuj1eTlki942jglxoyy66a+LOnxK/uDFcgcJJqZimbznpHYmMhEz/NXXX
IK2H3ZcRexYNZoNFWFaTjWIOQ5vVq4612MZaWFaGPcM85C/ND7lGzxkRwDnOltQK
4tw8QE8AukdTOwlirpmAoOBgPXjG8u5FUNfkT6Wprmf+9qt6X3WTwg+rMCJteSMn
vzPX5T/JXaxgMbW4fEyrDNyUoFCCOXryV2XFquDofLrG8FIrY00ZtD1+Q+w64VOY
CLMnYjb2SjX9p5nuoMQ1q9WakIRTU77/rMoWdKti72DYr5+VAOfCYf2QWtJXZBtd
yD+QIA/t4IwtQQ/J1BGUb/x2rG/mzcgIAqLn1cWJSUeOL8aF3D+5eiSbrA4dGA99
Lm129kI2HkayOolr+3600hd8ebbwrNI/e1G2p7WPJPo9lrT/BSJZ0cXfspMnR9ba
APKlqtX+JpnMuU3ugr8ZHyuDJLarQoqBCLVX0MXlIZPSaQH4tW444nMywTUHQ1xf
2Ct7XQSUym6AntYaPmgqGdHxq57vMLBSJEyrCOCtuepu2B+Yn+b8ArpPOoooKsD+
MiSKe17nxAA6aXyB6omhDlMbou82SWUTs6UzxXymfGZRX4ZRhT4ZjXd/Se74zgbD
oEdr1f8Tq5tLJcVNCFNjGamr7EfImAy/LFnErAjPX6OoQbeY0oYv9GkQ3poyameo
LINl1kt1j5xY1XpA6trrsjfVUHIt6FDStykuy0H9FLPx5vuwbL/lZ6Art8f82YTj
CG8rWlbzbdnUZ19+9BjpxRI8k970OImgwZX7I3O1VGfGEM6e5hIW+qyyeZY2BsBN
9CLr5o9v4vHmVSvT7nAh87njHjiSfW29PN1FDHMggQUf/7lxRSikL2WH0eJXgxqZ
qmAzRLhiZme9X0JG+UHd9ww4Lwc/S/6IzZF5vwEUdmKRpd9S1y2oKL0Fcnz9FldY
6GR8rh8398rVVPOpy/xEnbCtFBpzXuZR5au9MdqGcNa7KNuERws+JSe8oXk/+l3Z
NOwy9EY+/GptuhCuDNrncUJYD1jr/miLLprPmipSNLMwdHJz8uomD7+Mf80QTw8s
QCaHoIwqRkchk8MlnFZbxrnJbB8Z1r9JZqhoF6CrTD3L601qpGK3xt+y5pGVXgis
UJxXoMdwnuK5wDIqmAKERbP78+zxSuHbNvJjn1aT0MUany43uQmn5YzrJG6f4yzR
D+gb47myWRxtZEDWlSJBmvkAgfINcdzcAHTXFmvNkd/BHNMk96JyULVEG3W8itS4
u0tMZckLRKN7RCODDxIGAmU4BCZete966fDLi+befPqKDt8YYczu0pzosVA+0MyC
XtrYfjwwIriOIGuUdR6veA1xjgRjZR1j4bj2/Bym+NIaeorfRP35lRSy00YFPKiE
7Mg89LLLtVSl9XCzJUOm96HGaxIwk0+u7UZHsgTDheG9q9rpIHMGRGT3e87EMs+U
SiQF1+pKsNZtbbb/nfoqEhzYqCjjQCN3sVoSNPbvSG8ppDqjAx496l5rp/KWsQeK
+3SzMgtAXNNMaNt5bHKFZLZ3wcCuLwoBejrBiPaww+jlvUM9m7jhf3Ypgn8QVUNM
+g1rCVMdk8ylUden05x0MSfogEbHoRK0L1aScXe9YXficeh+EO6g27qcJkunr+qL
dHXDZfE2PnemvQOpa4khhk82m/yMEh6JG35mnnEZ1WWfm3SyR1L+r4RHkOXItjrI
Jd2d+rtvEQvbzRq9kzPScwM+tpBN97zX0mkGCtlQqIHdpyxvpB0+r1M8mLfsFu+w
pFlOajA+cdROfv63rivHDuhkCJWzbzBz6zqPNfQyltA4zg203JnmcLHeIsJeGOUQ
K9l04hzgNUrWCkQ836MlDGLPdILujYeOGphq2s/uxS+GvWXmX3APeJCUZqWeVIr5
82W2bXqwZwy063epkjVXHUhI4pY+q6aWYcD0CLGZIncUFgRUiCRtpaz5WDQoVyCy
HakQmDwbm0J9K4aOQeQBDSuwyjeSBf4ZY6Ty6zsbaqQ3NqemK1h/8PqNZSoN2WfG
9EOcvevGLVzmr+UX26Y1GiKDBpuAbNudwLJIgDC4aE8RHNmSsSS+T19yX9Rs6kQl
2j+Pqo8CucPaU+kajvaNJbwwfMADMx+NoKvMobTqnwv+WDmAGuYHRa9AmyfKNcLP
jSbQS1AhO8tvSd3bYNQVnXN3xWum6j86WKDEfyq+PRzXasNo4dctjjrwvL1KC+U1
5Uc/ISMZjsffZ/yOqz5sg2Ky9OK1CkuNd+GFXqLd1tEBMkaS/3m/d1654drguxZn
HZbeAG3F+1O5FNHrbOGRJeB1CRXMN2hMQRvicAhHZveeg5YfKxIKhhkIQj1PSCvD
eAAoIPsZBBe4/Febntb2L6S9Y6kiLMVc1cl7N3+IdAvPWX/137JwUyOn00RGNeG9
UavPm8SdubKf12pgvLIYftiDIlYWR7n03yTFYcDPBMa7VvCAwgjJ9cvUV5sqcZDI
Qbo4OBofg6N0VYRvue700mNfsW+h+J5m4EqZnJPg5cbmgQdmISN2TOQ1RAE3SYPP
I4da4afXRCnnzVUYXYl6lJL7xo0UfMQXkkxskYew7MAs9s6FloD4iKztU7uBkX2S
VJIzwrb6tq9OCcjxmG7MJIu8P/zxX/y/AYujF6hN1Qt76EC0K9OY8gqJ9na4Jszi
rPgf2dyNNA2dYWqJ1FrJeIFeAjqDY87wCTxwh20N9Ag59BxIUanEOX986iuinqeK
K9nygxN5WV6VnaTYTwTlj9SmAxcfyO0Ur+/IV2rQ8gi8aewFqLjqTQqcmLJFn9/f
m0qat20C+Gb9TbvRd0h6qi248P+02hYhggQMLz2VHBYn9dWkUc70Jr275RFBlYcF
rV+zrjM/O/+xRYOlgkWuo77udy2aq1bGee7eyRRRhj8Ox/xVb0panlkOqL64+6Vz
jeXfEj8aRMmPmCvCgIqRRp2TqEvxiE2pqe6u241HOTDyYgQ504Tv5UmqAYUteKIj
HceWXuIADjkwqJSq1gk59VGC+KHcUfuMtotSKNWfrlYLRidK+QQg0DNAHYDfJDw3
dQMTgA+iqWwa4bPGK1RLVdqsZsCHClxEeEJomiMzFNmOc80HnG/HKZk6+pfNdp7Y
yCH95Inc9JB2DcDGRmr1jkFGa4r3DgOnNHzStz77ScyRmt6cb/fwrLDZone3zosT
rnMyzr5gS2qr8PzTVjUlcKCzAjIHHCVIPsPI3kHON2lvudhFGWovjkZyPcxjYTB2
NH27BNJsVy5N7QECsKF0niWZPATtG0XnuRExsuV2dNgU50hryzzShizb9vsjjGOi
C3/I4tKMfuXViHGzgRocHVL699hYeTRs4wQCKkRI8dfAfcBRypcnKXfSa6WveQTw
Zk/KHSYIoGeEtdEynxKVHdq40ynxlhV/qcZKdLwhJIbI7kNwxZDr/p8BYLzGmw8E
mwYE2HJgkqcZZGbe2j0g6+hMy1WLAKJw7CCU39DSCmoD8KMYUS+sJeFnFrHRnElX
AwFGOKrvFTTeVZLh9iZ7nErvDz2To1iqYwYoH/bH8GvDcS55sgE33kzEbi3B4Wau
qrwzkiI5DTbaN7S9pslo+ntZ9s7sJvwuYARt2H30esxq7nAUmiVWXjzhMfPdxJXy
CgGxqHE4LvwVB1oWb33yzOvB7CnLmjieMrNWwvN3PwuBu41H9f874rjIE+q5gz6j
2souLHSRUOXKQqAAjqfDhhXhzcl01f/upSyb8CFh9nBXxS11FpT5sp2o6bpVnVDh
W7gTR/W7KeDAOy2oeONlCyCH5dFldFAl+V1WqrcEwW9nU5tSAQsh9lGdiMfKFpsp
Pir/ho21PCqrpSFJ44//UcP28+S8rx34tEjg4FdzWYSF9z7N4SSBlyd/MamQZn3I
ScucWr+pCDpZCL+DRE/5i5dUpfYFCY6Pw3RryFycKn13clZ7ZXiANKtgU+2xjb3I
G7f4Lh8P0vKlIdrz9MYCpROBnE/9d+reAsj3jah8kceczB8Q3IL/HErNC4UVaXtr
8jsIGmlOvJQMtL6XzwATUZUqPdR4NWnkjQ+digyTVeekEc/w5O6rZDyS/XAotDvS
ZCFnu/JpuamTp4GtXvyYQXnGi2YOLX1PvLVFnLnmymHk2RfrLarmglT+hmHJwXWo
qq99qAc0ib3/6Kj2zWOHXGmHhxIP2wOeGlgHzeWrb+Ufj8X4iYKE+mzekkBnPZuP
E1uvid8gaD7t9TUa6tnnzfs2YmGbdT1C4CIVy3xjYShfv6lnGyGpWI7rJEW2fjNo
GFICRy5VSKBuKsp6aPfHNeAV7N3YEQCKx3MNLN6T8cJbG1i8vB5WkLvi9Iq+VjJT
TAEuGXSt2niyeh9rdJd9cWG0RKoT5Hsw/Vyqhu4HPRgxh1ATNYB+IBWYvfwlxjDY
dnsv3R7MLvF8CruTQwJbkjHZNixg7cozr4MSQdrPXBomBt5DuhtlLRRbBfTOz/U+
kUWIv569XWzXvcwBUOUWfRl/Leg984UpS3ipfdFIdXLtcXja1WBRn+qXf1k8qc6U
KLPRG6ifQNWSksn5F5ekQQLiOr6klLBnCf0jzu6n44+/B0D8Y4P9K/MGwyqXusGY
qBosRxBkwjVx3kdfCoXagk79Q6Zss0pxIV7FtXbGOeDbFcBdNUGkaUiK4i8sJHUT
04vN264yX4qEsljqXn6sHiJnh09jWvnYO1bQzhGd17IETAbPF7J4UKWZ2pu0ZJPI
SX4EhKnt3sqgc0305Gw5ynF9PfQGEQE1NYXcHbnl36MEFoNkTBE2Mp2VPlw2CQex
mbOCoABLjkiESGqo0swvPjSULDbPFUOIxPvwKiMFhwjYYss2eETJrCJpbegCc9ZH
uFWVL9iQUHwd5kE67OkynZmiMS44mBJVExeSuQfWNfwmXELCMTmnSaNLTq/sSajr
4iFuT4Csyt1y+nn+/jywp2vTEmi+5sVm7lMkEM1FShEoNRqrzkrzo8OHw6EXAjXK
+p95ay/WQR8ozlwdeR4D6HAgkEVA0tnmkBAMnVqB3yeYettKv9JH0+qkYXLiHAb9
acuB0VRetShLJTHwQjOVZB4lnJiAOk36aSZ1W7r6LcoK0B4bI9zwY+VB54PkcOTD
04B2cN9MOKnLrg54pcyluNidBLU8Yqc0b3XpGfydx8M7QZrzTjuGQOBoZx54ABms
hIDRJSbzhOh+GLZ+XOlppwiEbYIPf/U6eSGw4Qn6TgWpt8di29khD34YRruKt12k
tzs48JQpdiJUHpRAxFUmr1Qz1Bag3F322RSMasCBL2yHKzfE2kjpfIwHVSTPY8i9
xCksYHv0RMLoajWmHrao8dA2lGfqgYZI+jt1oVQNGCimD1QRw8Hm7Dc0JyOmsHqj
nig5akdA+WWw4qogCkpmQV7LuNOfALBzDUYb1czYta4TilbHJCXYqcRvHv/YaVwN
JNPuFzgoN2OfHeeXJl0H0CXr6CZDd9mzu2bAoB0Zc7a9qd2uhcOWKA8Ty9DXWj9p
H0STTL4EwBNranOsN1hRmzN5IhoW0qlId1KPkvO9UiHqXVHhI06tZDJ+M522DDbR
Iu35LjF2o+JKMsGsxW3Hvrd77Ty1Xk+6SEzGfy547Vux5t9EcyZtFn+kr553U/1D
TuRrHJvBzez6yNEi+JuZs6qn+ieGd6w2P0OkRfFxabv4n13FfNcc7EnUwbqd6U0z
AtwdlgydcNQsWUIWy66tQiCMKTIuAYqFpsLkjv3LOrTUkKxVmZoLqEGaHpt6tYIC
1VXHgPYUFW1YDqUFLymovrWzCWiZUNkZWRiof55bf/NL63brE+EJWNrLKv2AL7d+
7GIIUbUBEaID72q9+/Vl0y8U3+sUtKpQVju984/nOuRfapTsutZZ0aztrZNXxKIc
XS04l9cuTnvHrw311hJq0CUlEcGqcjrsb+nKuDP64AqNRvVFPez8/tj+ArytP/Zc
7fE5Jjxwk7lrAikTP8ujdsjVYLMSdO/aGcqwkzGnfRgCyBp+SyWzEyf84XaQC1qV
u5hvvs7rcQyq6S2COYHj3aTBrF0Nc6+rCs3MfzmeYIyg7gEV88DOh4AOT6550zv1
C1BxJI40OwhP8XXQScIf9MxXmZ/c14z1Kex8u97YrVN3OuLwYkeutf2Jcn0cVZZC
NmKxcjKvNPAbTMbPQ3o1cbqr7h60dVFYMYnwN9BRp1G/ZUW2+yoUaSLYsnFyJOUU
Kn7vonZcx/p1xu5nxe3Jjw==
`protect END_PROTECTED
