`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sn0cm7rjiiOeZaOLK7rDjAeb/Rkmb1n/qFyFkImSCDKAe9QKs/GTQdz5sQdEDh7M
Q1vPHbMcRDqDp5TcLC8yD0JUBAqseoY92TSGFmdyynWap+8G5Hl4v3xZLV/PH9BR
hYGot9oum+eTa2cAvGQWQadmMhYgPvAGg4xgIy4ekYvdelwtUlcpO9dAU2iTSPLZ
ud8AQTdobVdHVh37wzOS7ZIhYgL5jJUkbM3yOIA24c2Fuvn5QV7ZhdAbi0zMrGfh
alqkJxy46wJUJPPG5nLMHpzLu+B2lxMtS9s3nAxNkUVWl7HL+woQ30bBpP7wlVUE
W4m7DZ3ZIMHasxTcIz9gcdio31EqFWB8rMHWYzLvb6nbCeDJSFS78GS9WoEquNue
5w/TD+1gSo1iqb5k1cBjmLBHONeyp8DD4hUP+pMcO2nvaSqaliLSgJeX4/By3Etf
PWz9w+67BBQeVyqHi8ARWa9Z+fI8rMhuE3kRI5g4LVSqLaRafSiWlGsd1maXxfog
mseccI3EMaOV6PUmUYZDbFACFbOptp/u8ZqJo3Mn9kYvUvTl4JJXwDZdNbxRzkqj
oDvgWcxfhP8x2IZSndGoAJFjivn/FmHwZJJAIE64hj8rpPzWtT5nXdS9iLj+N0+J
RVX0jllw7GHWSNFEAR6mxW2TgwtUg5FImqW3AGCz1CZyyLORqMy2XZJd79GlNPhK
Hx1t/zgKie/0ZB0zbtdSjPYzOX+C20V39wPVCe9C+TgEXQDv/vyyUi+Yjctg0NC+
qcXL5xvTGkb5wPYzJ4sv7eIe9RDNQwarBmvkTHf6kk2K+Wy738/VmE/mvaPcIpHY
AUJkBuQsyPl0OBvDh2qvoXHx6nDylYkggDMa4qVAi5zfN6wphWATUpTVDNe6V2EL
YX+haYlvs6S0yZgmd7V8JeykkllaHu5HxiCVNK8CUujnEIusRJUdzrOcsOz+a8jG
MDb3yzySiw2pAkCutFB02Bz5VcUfnBQvwOOKmDJcrAT415u0papU4uOrzi4Z/6Vt
AwbzHlvyr+bOxPprQQMDdHR/bUa+sgEhGGi2chJlzrvi5LdTRAbLoVR/hdb2OwGX
O4U5/CKGN7q4UKG7OetXfqNl5UkwSTbIhxhgDMd9bMBjDtUPetJGC47twqq19Xyp
kYMabYJ7/ODxAl5g4s/TSeDjIRwlqFFqmLaqjUTBzJ4D6RSEraA5ddhkBbEJdNtG
+uyB8rG73iXLNuidlRGcz27X2Q+uvBpA1g6ebbSTyHNqXt8KjNtEdyr9db32idk+
9kOS6f5W0iVxkR5DQfacP9po+/IBDy/rk0+4nFQmfKVTvIW2MXrOKupfrj/fJxvd
CvijQanD9foxyVC7FjnkyKJn47Uq6a4c7RNMhCsObjEeWi2n/XjX0rRux5mL6VK1
z/ZOUoMWgaLho4m4ucNXxeGqZrJfyWXp4NLFw9YRjlrgiTJIcE1XcLicixZdgd4N
ax9tlGuOGFmvghihmBe5JIbrFVRk6mlmxN1rbBDjZeGQ/eMre+yk1gSvCS8zWBe7
4fzBTZxV6bS/CAPeBVN+bASJPDfjutjKEJR/cXl/O6CK8PWY/+dGzRmz57Npd6ZF
lLEW/w12efIkjhDnyXKyiiVagenf0ZbfBX0Yy0vZfkhRein85Gi9hCrH3Upmk6Ij
+Gy1QurOcgRb00Viz5T0/mAlHODtJnnCH3UwHB8YwPL9JzDq/t2M0cTgr/Fr3MaK
QFm9C0jn99Ku68f1FIOHcO3a0yh1ZmpCjfSkP0SKoYq+hQWZhrgNMAfoNrd4dvjz
zTfY2xvmzrXr51ujfYnB8T+5KCKcPRmSYW4s858JmKIkFmHNN3DvDpEt71FLUk18
QOtFicGj/S8aOaXC49IBOcMh+BU8Yzxz8oQiDVxVJYLMnPOHqfy6ECjkwYRAanX6
`protect END_PROTECTED
