`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eRJtiaT1ocnpQN9+s1y4gDu5oZjgj2hi9C14wya4ja3mroRJtPohWFVnQ9cLldZJ
P24sK9Q6ldNn7uo8xiD7shczxZ5498pEcNFLYmTYXGWE+/AEDBayRRGoy9c3hUSh
s6a5Q3zCmSvjtdL9922/qpvFt1TmyEiVzNJ4tt2pmw5YgaOhNhglJfzFYKiLkzk5
6E+HR+qKoznyYUlZG4tN9jYJRLUP5FkgyZQLQ78o4tuyMZM4m8tq6Yf3J1Cjio3Q
pWPvnoO28Qx4U2xWEabSZ4F/zcILM45Nnpoo/3wZTkwEf2J9ubp8ul884LJSNi2P
V2aS3Snq7LBEVylu+QGXOgjxSesqd0fw+cA7VTOLPvNscQ7l3q1gI00/vrcuWX/A
fuK3rx+vfIXnJ4J8A2AQWgEX/7jrPVvrmIIpUB9wn0NPSt+UbKIsEjBUB561q7Eu
45yndgal1DXDmHUczqUMjoJ/gapOmkZUdYbCM0QhwE8Zdhq0uU0YcRK2U7OV9sCb
5dScl2zCOedCzbH48SxaxtgsHYMnj34tJsrA8Xui8uMUjJwozRAfSXmHREZGyV8I
/E4sjIiXvAzo56W3DLDPgmq4iOLqAH8qUyiTzzUZ/Wlx6HIqy46nqIiY3Gm0gKMq
Bm1hfnwiXh46DQzDxtpbCN9584h1kvU/Gn1oJG9QIOvKJ6GL85uQZtd42gSHMQkX
9e+GZmEvktRYjZ6mc3pEQfLkas+PGnmiHzAtO1EOYYntW9cqBd3RyG3br3WBzxMl
qyhGfAm9o9pChDS4GYwFZwRxk84rnsU6i9oAch9aRyo++fy46OPNCNnNNtiZ99lM
eEnViiXszhWewr+YO8L2Mu05k9aC6y6RqqSl8OxEiYgnV9tudpA38ZE+htmnh6Jw
FJXyLm+DBCwkFIwxZzig6GV2dta+Pox+trrYVTZcMsfM+YNnl5Hll2WE3ua0MPKB
nXcprDkEPZ4NF3+st1ECfOcgNHJA4La6yUYMbTDnwEblFOFf0SXit6DDQ00g7DEn
kKj4+anAQYO688YnrnnlldapIVj6YY8Z/SzkP1dHTTxog0168TsAqtt9kH/QFrpF
Dxm7hwebjYidkkoABKcXsbsVazNSHshBPnayoRndI712YB3xpQgVDCjWuUdpWMLn
kMWJfDWk1DKZcp4PkXcE+R7RFtKinEyT2EXZloDWKTkPSQvASc92B3j4jZfmGuW4
z1p0c/D5isslIRb+oCa/W+YwzMumLLJLmgrAf5MVEyXviPI8yZPyYj2U6KCHUsJM
s6J1oQvrtdDqM6/z/ZzWbuPvTpVRNDjxGvWN3H1B0hNn1tdlozzkTO2/XAdl1mf3
7C//+Jfj7KYis7RA2JMSEe22uOBKzy6jgF8O1stY1yj9MlpFxqo9zD8XduAabrkm
0eEGJDd5CLR6kWA9F0cjCKS3V9+YLNv0l1kOO4u1F54MdXW+hUo+n7R+nAsu1/R1
DHH7JYIsTQZ/6Xei0DOEEq2rcQ35XV8c+qPSDJMpUuX6nSyCQfhoNEBqOdEm2613
AcjXsp34gah6AvFTvnXLkcOx03qJGcxx1n3gPwv00X+gbh1snJ9MDEIk9duHK/+b
21taEZsUva9jPVBqV522+erDJAiROuLbSD+jqL8WhkoC17aK6cqbvERES8t8BB+B
GXHSklcns8euIGtQgR1CME5eSnhPUS1ClKm8guK9J6e0OLviyHH7IALufxMgVH6T
CxdlBeKfjkDxVZXeiHK2NAVYWWf6RtXGQxlYZwqasai1xW23Yo1DY6Yk56j+2dyZ
I9eRrk3R9RX1Es7fl9vM6bG1vV/3iqdOYeh8+SnLMinkyg62C5TMRIRoNrmQDfcZ
3L7IMTyxXyhq4c4jYt/V6wxxX0kI0WWG8WwBoefLH85t41YuHqXC6dF8P+dD4NvK
2zzov2nzpeAhsKmX5mC8v8ZZ+XUX6Bk7XRe8P10elBQhzRVcxLe039btPHb8a4EX
ENaP3uBX7bOLyziFMmTPK9eWAp9kCQerE1XhWlW5x7mjaeIWqo7spSF8oEZw/VZ4
LS2lMsSU+a0wZvh4ta1XNyzySTiWudz/8LFFBSDfVLstcw0Sa4yUY8ofdTthfiuR
zwZJ/ycXYYnumPp18RACS69dAlf13KHMtrS2CEJxvXOtKw2HAakXTm/xrR4zjXrN
eIhfAgCFL6flo6kYySHorfWlR0juWBzXUaJwK2XM3cDQF3YdvirAeYGEkf+S7XQu
n/+45u911y4v2JhubzCjBc9ciUxxjCZwN5Qb3B+dHzG89x7mEnr0erCFDpHwA9y7
wN6bVk1yoLHMvJ7DtgpT6z8f1NysXUqZ9cTIkZrtwLrg9AS+kpaZvcxu0K7nZMFc
ntdO3cXSBilKWn5FE0cPU4fMflMTuaStJ3iOoo984zrb5XR8dnUL5I6CCa4N20K0
2a+lC+Vdhp2VLdjWsD2lvaI1hTaWeevahi73XZ0eyqFiBr/NjPXbBfl7pbh4w9sv
IxFxUlQLAOTJsrWRBurj/wJkClbkHwYg8xrnEayyrfUlavoI2g2/yfJ99jIPUGQ0
ldv7TMps7x0sr8PRGSUwlOCDwHbmyWVSgtf4vtBcxBIggvO5snStcz/ImHfn0cry
g1m5UbeP+yOmWLUZBS4CkFE/9o8jCqfM5akAY4p4CY4W2blzV89tNCRSr0xZagJR
A8cHiUfxdf1I3q/iUbVxe6aioOoPRWzJaMi8orVTrFbxo+X2InOPUhU6eDWEYSuL
SAbLRqFiHS8Fkr89GNyBFb/76q7mrl2vFIBsPsa1MEKnjS45I2Jdc5XojP714fxT
p6ZHaXA7B0fWgWtg5iRnSHiNjQk27DvwJJg1ertGN5W9gPnksjx5i8SOpxxJtF/p
nAncyXmkzw8mRMJR7en1X8VxZOrAHVO8y/5szw2fUB3HSVDIw4yZb12eHlCcqAZP
z8hWop22d+EKAtK4ABTZEwNQ/HP36u8cVlFU0eRxHrCDNEAhIawXQ9s3QUuMABuJ
m9TZLBTkvOKuNLN898vNo/XXMKaTvBjpnosayLevLGKvXL6pREDKoWgZrvVcnSOd
5D6p9Msp1bxOlpXMkc+A98Q0ZVgLFk25BEgi0LGahX68RXHVdNc7G2yXTTD+7Uma
DkoV0tHE7Y/qpccTRId+aODK02tBdW9CKKxU6a+417xL+9aTAbP7PJxfJfO1JcyW
SXNxyt2b//up/qxxRxzD9dq2evNbwLg//jnC/TFAqUan+pC5EiNDUiRdWQOfnHK/
J9e6eqF/Eh2iG0bqqi9p2oEJal5yMdSV6+fTLkMyjkf12Ui8kw5wiHiRdRYMbQqI
bA8OXYipNIhN0Rm6U8T9HddhQlv4Hydco4rm2h6r889k0tBQnXQPAjNU6NhqpLhr
ZU4z2hTxbNEHFU0UeCgtHEh0OV+aNu0M1/lt9dhNYbuaO0KGyMy+cgAMEBB/w04A
ZYrdKKk9DhpWzWk7aH3LKvydWTl0kWfoKm0J16ModrlhNjvuOuZqO4Duber3/Bya
zhe6rJigA5JmWsAkFEEz7G95osfFuHB9YUaBSDJvQTRHCCgbFVd+DLTKNuuBPVur
7jN83t7qMd/asM+eVWzgC3Rc8niOjdb4ZFIAlxpah4Vv113eE4XwC23Rs2jiCFwk
IO8iVaNDG0scaR3wG0dBcORs+0u6SBtA8qLtpo/8ERa9aSL8qd1oLyw0NKn8cWoy
vU9jvRramI/2tooX8H9rk89QgNW2+8L5lxsR75Y8SYXV2Gud/0rEkN+ByQdyPtEj
b/s1FzBlk6jGNO1OmFxWeBnBAsbSI/9v9apWpwmF3F6hHTlJAWBbRwicohHRrd8O
m3YGARE7W9x1PJci7nr/9yXVOpeaQ7Gsst9UNtz7vYUAXYdREPX983CJC5NXxLSr
3/CpvBsAVYdZjESJiN6kO+x3oAulKohr7jtoJw4XYqE8nhPCQj/cxs66t3aEdwV0
5xdufrApjw6t0B6JpyjEgEvvN+QRiInkEmQVmOL1DKvvBkuglm+Ng/JX86k5eq2d
ztqCqJMoEPGAAi82IjRCi9NSyV8LcJVbA2TUb6otCQ7nln91UbHgVz5x5XJp69TQ
reCYwS2SmO3AYOACbRN9EdBdWRhoUUZwpDqY+5zpK9B+OK1rhrroT+4b5YFL2U+L
XuzQgi3jl9J0tjlV8G1poek3uwgxGl/frmDDXOP7aseHIrwBhPqYbJU65VUlbuI0
w+5o59wsr+FCSCtKtK3pDWp5QGjkEdLqtgGq2aAxeohhOfGrZWJS+Z2hR2mWfv5g
yOv7T1SztMs1eH7rrXHMxYVCzh5MhveqU187xQ79Tqj5945xWl+wBHIfPiT2okhN
o9/NTQQqIdj0J5ja9tSWuEStzBZf9GGqL6WztD5OUpj0K+hjOhnWQuLf1YzP4N5A
ovLdmFgod4QqdYFKK81/sjrMhqtoFY/seLide+vbIx0QEbteYqhP8sugPTxSizd1
EjSteXZi1sSKjLvsKYLWRF7ey+HYpT8DgbfKdKsMLS6SFMZCDvFs+3Dj5plvlWIo
WI7BVXrOd3wm+ahb95N9sz4cCXCXUQ7tTcq4azcTCBxADD7Wjl5hyStM9SLaLyB5
Ku49u0zZDzK64nZjQo9BaAVKfR8ewvt+J0kFbZQoWxbfrRwlnuxYIgjqDN24YCg8
DK22zT1uisRwQlx+qtntG7HJLCAVjIShXxr1JU/7OjyWw2WOpvLYFyKDsOk1ToCd
T4wFaLQC0DJDlrDGUO0tuiGtnrxyE5pHIy0XMRAr+joA7xDZSPCdoOAGbWv3KICq
XLGxRbR9Im/u2M3T0RwsyWZ8berrejMg0KXcg3pxRCoCqzf/jbNoxrip9CLGoDjl
sVpn2OVKaKhY4KBoH7QuE7+3SThT5ngqzNEp3TGoPvwDO45G8KKRPv/KjLkgGpgt
tnncTfy6YkMEgMW5hHhTSC4N2QLIvNExFjyQfDKy4acouLjqku5yoYCWUty15xd9
Stn096BHzYuRSuTrGEnrEW5gQz9BN6cIfWcyFx0ZftRz4wABsFtRs50fkhr2W+g0
871I8X8B7M5M6VAwgg+wc2lFakWTl8rFqd8lKvSef3rpBHPOFc8zH6X0QtKRqzAO
LvhigDi/en9uFdQz4VIes5zSpLk2UzEmFbkMmZLY0dZppBfeZd4zGOFPmsLpLenq
Bna8Vxqre7LmG2K/Gc0PVcczE1xIpYoeKRzqMoVfXazrIcP9SAm3XR7h6kbUaQ78
twU7aWvO5Gd8abG1VxC+oYBgNjM4VXJBwk9Q1JGtHxWCH8PMzzdy/eWnFXckqexY
Vr2B9Fv9/tDZuYQsJ2z7gfPNP9bA/QSxeIUbevaorac124Lf9+/AunRGzDhCQdly
WLD1f+GVpYurAf6lrvg7PzyZh5dAhxI0qzRXIqx1D58=
`protect END_PROTECTED
