`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VS5xEwpkZ8xdUjSxbZ9nqbDV5IlHCJI3iwXtcDr/rh69AAaooSmTZZBifdtRSUHS
icfc3ZKj3OrL+7oF+Bhla5eXrPRabpmf72fdGTNJRRRCDMC/0rwogO3RyliNp59y
t398T9yeCxpjPGWEdMRcjI/U2sSwmRvU8HmDGw+HWWo3MrokcrHNeRptRSEmq7ML
PRUylfHiC1WwtikDiiW5jFjM9j1GEYiXTU8N8QN44Dfsj6yW9nKef41FB17x6wdT
hj8d5BC5PfN+lkRdW18ZN/T/55iEY2JRk6km56xNutSYE2wHyzLvjtMPkQO1j+Ae
FhoqreWveg7vPqDJ4IgIrYv54cddwPkVSKV+4kG9khAIC3Y+mvjorCAfIxx41HG1
R3lslqPTMWKREe/hAHX9ZqBv6fhI+Zt3Cf5V2T+ZVZReoEJaXobNk0/xbxJx4PxM
ua4Tun5Hw3YqSbAcyRoYrZw/AILrBlxHRXwUtWjMYzMgvySu5udt6drcOflD//P3
0GrzAZd7inm8ow2rJs4y9IPvaHqQjJHqWxWE8HGZ+W7CJGtk9PN3WdSn8G2YXwPP
NaKDwz/vs4XG+s5k+9SXeFZuglw3cYPMcj/uwV26wM7W93QTckmHxeWJsSb/Rhn3
jOn5a4iDhjzpU52o10de+tIhfarp0gGh0pS6FnOFaZAUTpA0HkBOBVIVP11cosvp
zpO9kdu1pieYmw9WcrKvp9XmyTccDxZfWf9k953/kifCqZXvmPkdMdoZ0I/qEAtK
+e1NxB1Zg30HVAFyqR39XCMKW7O6PhE/EacbBAGeDMTMerNtbVGBD/EFDGPGz8vR
RWIlMkvuCEcmBrpfaaYLrR5iOWb1akX9NgCuAdVZ/aGX+CnHgBICMirfSHSULKWL
XQw+cTqY6W9XsQgv3vaGwZ+WrxUyKaPSganhSVGlH8KnTtC0gtComHeDm3b1Hso+
OstOyWVH2W9lhN430kaBBN6OKyWfeH05iJT93MG/rkeoN2QvHE/R5DR0DSAWAnd5
bHu9vlzrcTr0F5mnhsxmghrDUqxUKJegBrzu9F+o6ZGAWRkL8aKe2MId41y7zZUU
zfUnZsSgSQFu5wqO9a6IhDE2p36gNqcVDL0sgelSZo0aTvYVq8CONEjdAfDB0K0V
`protect END_PROTECTED
