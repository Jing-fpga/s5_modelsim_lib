`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jqQIXgQPCHHTbVcD3DTPQ6AaRtZ0wF8L4yUuhAbF1BS/Rva7aO/DQiUCXNFSKRog
o/3fVVwlRyCKxz1UPKYzaV42mNE6QmequQgO+kf8lLNB73vdi7ihvAK5VUZfEujh
QtXH8FoClb7YZ+xmyhwyZgcdeUYigz+J1F8GIVSloWnjc9IgO7ZRRSVZFE8Ykm2Q
y00Ns/cD6yMJvsOiH51vBX5Qsz7RAsVHvxoC+T0/0kDsx7/ZfVeKa9lFSL8Bm8ZZ
/f4+ZG3WavvYENwXP8Iw1qjRaENOP+cAeuz3XD0/LI9rAx954M9rtuKzjQwP6mXl
UBsxDBdAT2s20iu9BNQdRRtO+38AvZD2+ftNSEv/nKYcGGgcrJvRxRkD4E/qxbK1
FDvi3zExwda5E99IeEPQGx90laMmJI5h/VFJX0++ICU5zvN9ocpMYcd07cm15VGu
JO1Lh8PPHEjvG7oRLB09kyaXLVIsek+A1YXdw/GThlY0ZS2BbyRApcBQQLu7W8DM
lFB94ZZTbYkxD8/oHLnpkjIyqqnz3RaZQy/iqyGf3E7JonRLdHR+0XFmoIsNuLdE
Wf0A/MCI9RYjFcF8cDcMv4Ecm9BC1m7woS/6sTpljQaDxH6d6HFbv/BDKHNNUjTI
Vh8K03/zOhRaZWck0LPBQvijqWappPFzQoTS/t2pDNXgReZ1wFw1nxbTOy0ZcBH7
gYHFKI2wM8Tb7U8ZkHDyAL0LiwsU6Id4DRyA55rYa0mlkOxDox4PgorzEcajYett
EO7P0cpBD/ZnaUtoYxzc4+T50E+Mow+iYfQpAcH2UrNcHOPlOeg7UuS3MXWi06jc
BQtsP14624GGBPksL/lGXBsJeDqiIfGitgZP8JC0JEbe8wc9tZBWw8zSCfxTKt7V
VJLElFumc67EfnygZ0+IhTq1ibKVXK6zt43on7eXNICvZj+A3sAVb1H+yDFLlPe7
LILMJggx5i2LsIvcVnBJ7QxtK+JEqn+sdTyooeAVS5ZG9yOG34h+DkBwpQ5t1+wj
SqaJtnYb/M/8NK9BRskNhjlXlJ0U+DCmVZw7VtLxXLE=
`protect END_PROTECTED
