`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZAUOA4hi5RNux7FSsqjeR5A8nfP7TF8Jh6+Jw6wXG6i/WkWrBTGB+4wfRfu9PXX3
UTqz4l8YPs9aORIgwAr21Q2EIg9FGtign6oVprUYy8D6Rior0WH7WsvIdn5xPAA8
dnBDLPvfn3Fof+lyKB2CfPxrWn0bEaN2yODEbk82IkXuKB4fICub5kVxWtd56Pz6
q/kLI/NzniKI5lhgLDpKyG6XzvJJCIDWXNr8t77w1DejQWXA+JMCr30eWxIYR3HF
GUqztMeI814rqgqoK1CSb7GNvH5DXgvsdweZ4zb6Bex8SoOkUpa/1eNuzelXNRXZ
IkPe5MzD0VSOPxAMfQnDQhPwBbdYTIhtsAa8OSdHJr6zk9MHNKY9U6s/NPzRAStz
1EmQRnmM3qp1e4oimH6SsCsXLBIHA7Ias57Mw1HDVQfaOHDl4Cw8ujCNtCAKG9hp
/YAiIssQc5+tRv9Use3W4pjhh9x66hO4Mc5xFY3pPkEb06OePRAv8lDXwLPO8cRj
Wq0f0ed/8AFJSznL/QHXfPq6Q9QnT4/Y0qL4+kXPzyVO7Wvc+QvR2h4th85pyhUt
m+kMzER3PsTV4Xza6qLn1FfgCo5zG7vIuyCEPONWa4WUga7jyfryMCXlB3Pq+nNT
dFOJw5kly5XKVgkIbHuULXXWAchbvMUsr/iOWv7uuq1O+uu6C9dS+bn4rmz1H0ih
uVmnWK2ZZeRdT92eqU/TVC+ROA5dOxatAEwQb2xKf9b59bUyR8I925NsU+XHzA6e
db+hgDRqH3gL2PWjzYv8/GiduJ2kqVkBSeL0OCTGRh1BVgI9WNSKh9KcJ7xLretr
/kytGe/9TkHS/O7lYhoUdPtB0atMmib+EgHAN3txX7Iss7wzjiZ5G5F1IzfXoLKd
Prei30O/pu7ES4u3GWBrNMykCYuUMvwlIy3JD/hy1Okb3PuUWE/2NPtZlI00Su6/
wvUPaPzUzs06RThLA5xq8oAvqvjWJQ/2p8IBZE2haSdLQCfBu63kS/OPf3OhLOP4
HFvoys6I2WsRTD0CSuai17zC5Tu8Xj/oXSOd7BPjt38Z7qLUikB3+jl69LgKH0R2
sWC2/m1cEW6YDRQ1FMz6KBppqr/gQFlMCqfsvBEvfEquAJOe5jFE2LSxkL0FVHEo
OJhrz2yus/ftBJmrUguskiOcddrEKjqvCyenSigHQH0sgvLAWUsNRDHg3nw7ZiQ8
8KLtEaocyrjRaO6fk2xrecFjlluBnGyNXpXyQvAiXfHGw1aZF/Ntkc/8BcaAj1OW
sGhGtFPWi4VUYCCZP5Fc5B1P4AxwZxJT4QrLqbP9lSnVdnPcIVaeTGf8h6A3WBXR
jXP5H9tP+bU8V5Yo7updTLamtTnjM25nT9wG8ENqnpHFEqlc6JfJJKXUnkKH1oBz
Y+QQrIil8DWxgnqnFo8i4qTTC9DwFWagbsF34XONi2Ywpxy+atol4Xl7yRFeaLtW
goH2MbOKii3zOSHQqYUniOFj77wCF/LLJdVhlsxJ7E7nBbTvahLYfALSpt1IUcDp
Urq1EaIQ34xBjhB7ZXZpaoaZVPJuYVvPIQTtrmUYb1NCkeaHwcSSzIWpQ1zbYwJ3
IzDxJL48K+EDlk9ZbzsdoB3aZmKP15yn3hIXXY3AIr5C6bsPTkidX++M71Sy1180
ccaRD+A5GJ+qXhR9Hi+iw93mDjaKySdrAvKyK5QYEpQ1jgFPNdCBXKZy7ShPWvkE
i3PKhFnbwOGWS32XlV0Zi7UvnlWNg/FGQVgLrm9b7S4lCYzRIPKVCoQB/91S3P/z
`protect END_PROTECTED
