`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pY3dBF6cAj7bJVSQx3qEBgKtrP+i557O7ieAvxHk1EgItMT3FQYQiVsk1HLhCoky
0zh0K6O/lENQODLOV6QcZMtk/2kwDUwB9EGcTu/b9ub6FkMgO66H608nFJxmXCj/
upWBSO2aMY2sUBh3sNSWilEB5p6xxpfSya5/XjNG4BeItIrZ5XVXVQ2wZtjjQHa/
RRrJbbPUDV/nWw2O7UHRcW2wNacoPrAjoDa/RS5LzwJhOshGDY1pxWtHJjZ9nqNb
w9UeDDr0yQKkv4Wiq9tth+h1vu74jv43y7SOrxxSUHohCeOXwF7O64tagEiMp3Wj
8IegSGx6yPuLLthSLTjiinmCFaZkDIoQHa3T/pET8GBNTCMSbnwFCvhTNA47nfm6
FEzuQDcfJa30AhHkeccHjSMsZ/DbwGXwK0jWnxjI86VrCT6aqbLmlLWaojseJnAc
nMQ7rDLM7ZNgfF0OYbp//UK7GN+eTpLZE/1VUxDj+EGRGoOEl/F0tx1lUhlk0PXR
40I0aRSsIvCPbbPNKxKD1hBjQFpavfM6xk4D5LLvIpAydekzB37HcqFw1iLxHvBY
STr2wQXKe7YNIl+4MLrE0wBDNfgH+veBSmezT7fSVw9J/IBzgf8Nh00LuESjJ8OW
ltkW9doEae2vqXmCGgXE5De6P0buwOM5lEwwnk1jQwMsG2Da/XM9WO6NysMw56zC
uIp4vN05wOOtWnlP66bB2YuqaBqsH/MOERcbFMWFIopIVgAT6buZR387shcqGWiN
zGUzhipcbzh9GmMRvea+jdBvAeAuacb6+4Tp1NQ2vPTk1+b96oAtiVnzu0ny8ggw
dHzjBzYV2RbbCiMaZZCgzbAoqkKdP0mRJZ/Z87rGVDzpz5g0JRekeZdjjKUjS9uV
jyAADr6jSzvRqAe93P38pNfE5H/1gSip/QiDd11qad4=
`protect END_PROTECTED
