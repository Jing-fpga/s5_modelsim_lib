`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3KugR925hHnykdXhLmj/qkBofiyXRtmazFFlV2dkwQDcwpgcnG/AixZFyn7teoov
CZXDuTfla7Fq7kdDpIY5EQLWI954OIuButhpsLTWOJutp4dj3eNDEiNBNw6fOCUX
lkjKvO5S2Te/7W7CklHLRfbfUIC3ZWoRr65ytapBPwdlw1ExV9dWjNNc5/Eo6Da7
o7cCmxfeCVRgyVo4snuXNWHVbtHK/NYqiCeuvXgUSdT3NXWGF1V5hy41YJQjK5Yz
PoE5EqIkcRrf6WMBbxcGZOQtL87tW2omQhLp0rN8p64KbP+xXLmFPl+EQGrW+MbB
uIZn+jW/sPSdCPSa5Uzgn9OBjZygNzUbxS3taJFUU3hEY+u+Xei4KnJs0ASxZ1xM
qZ52ZNhDzEjJ3SOkpmB/lC6y+jmeeyAHXBlcVY6y63pnmCiE42yPNIxGNVrhEiGf
8aM/kETKU3mOhdPaZmobOrw2Ieb0jreGRUZnLKlZA71NBDhdbfSnxzQw6xra6YMa
ktfIsuH/Qc7uOFt/yQCO7iEY+zXC9GdIiCi71kdExNV2p4ZYjsgCGeUWiydbjEzQ
3QlgMVRzNNqYpxE23c6IQh/AezZfsfEN58cf40CKWrL+Vk81m4i6tLN5v/tWZSwB
OnX9JEAnLwOsR+tWw9vB9D3EtAlkxBxlzpLni0KIXVsHIObB7QjA1qN+giOBv6VI
iiGXpiLkwu+CGu7DfVP5bdfYMvqU00XOzFJfOW2IwMbJs3xtIZ0wre5QTFFMeQ/B
Vw5EQqiK2lDC8QvOlogq7fYX/SJBwwKedFujHBLgGZPoeucUI0Ajktceu+Ix7Od4
oz9lH4J/bH7nT+ZxH3dqbAmJRBIhXoplEd6FfIhq4AX3K06pTy7Gg9sBiTQQ9nTW
9/Xsk/gwmWFKzvcoztuq+oiNxPxTrLHYao7CaY0zTKGeB9GdAK5eX7cDZnhiU1Dh
W7ZREGbA8hsgwxUYU1lNl69Nn4fqTD6Zn7n3SUwtb9V4Kn+IItAGFG2h2GdMzVC1
zaCfDzwAFjvF/PV+mSG7F03I4sMqQmGezCr8z8jeruBfZnnBd7R9mBtQyaR8WGwz
UHi5CpVbf6PvEfYKlXVaeWemHWqdNUpnumY+94OyqrqCTHkemxLMmyl1m5otvZRB
v56tT/Q7e+zI2IazW+VJCIW2RCBhVFeQMNou8zmiPQ+HSFcNaesy0LzX2+kyVDJ9
wbwY1ML7O1OcNswyzK5G+M/YXVc7JhpP+TeSvycKpa0qKmmgEp2VTjzWclJw8boi
6VA/QaILhWSynkxCnBkALoo4F7XtOaiZmTNzF8fxgMPsr/X/j8HD2ibtHLqDDgmB
iqQ4CorGgLxCqNPyH11meWFdON69reUaCP4UTqRSc8X+eY97xWe0tGxa6Uj7KDlN
5JyHfmT5CQu1MINrPWEFoEEHf8lAu+tOllZ7/VXRzoOe01Mob+sNdQTQKxLv0fv2
xa1Ku5ioOzbqc6VPisiRU+Rj6/4PtrXqBPpRAw76MEdND+gamWwzzhZCAzjlVXLo
MHSGuQ2s3eHAR32qqJ0KOKfetxFEbX3uSlt9PdjHIAjMIast6r8huzqn7E9rFpZJ
gnzdTsUb+OjBhhCdqfYvEBKOBgXNkkeSGRON7n3gZXUqMWwdbK1dq8LZiGaWJryS
Vhp2qEgBbjy0yXYZzBtPDGaoi9wTU0sjUbyJDIb7CGfQvWZpelRXWUskGDPVKMw8
UmOLr5qIaSolnFBNskQHylMBDwer1W5WqyeQRmYrApVimwUMQR1qRBWw7ev7Y5f+
Ugl50MDhWBabySwhgGCzHllNEuCG1fcMEfIIXRHs6+wwoadxvIrAVvyzjtnqryo0
TBaQBexwgp4UjH9bGY7H6+2eAhSncXXVXxOZ9ZqFEyjLQkFq7OYIvoQa6BHKO8D2
W4C7/MEEf3i3bbQBB5/5WBEGFKtL5Ua8kIslrXlnGUD72ErFlZbS7YxMEI3E0buD
DT8FtuqeCO4DJ0wmtAaTeJ2NJxZykd54GVzWjfOqZEISYSru+E0ggzz2x8hCrpeB
ptdXBuhNOQ+5dRSuOmALFDDB8PQGTOqCqa15M0Fk/F8ciPC0QCWCDfCUvI3e8O2k
ipKynV8pUT4jS3sB9klMQ0YBztvlGkZtny5s4qBQxDb39USAAhcPT1lV9GLzw2rb
r+zCIwIV4VtHS83tQ9caLCa9FK50XRE9qfFMhtlbrA34Ll37AZxazZtpox8F/IjO
hVW8M30DgqvauiNnHEeLD9Tgy+blRnjxiVwdJmevQ0iMAv8wonLXfolBn4E0Kfzh
lOXoAngU4UtRGC0dFg/rhaB7cT8IVPr6qnN1JFNuDqSgfotJX2a+MDnvs6Bt634k
QcwyqofdCRdC2SERZlBISDSfv4TQ6fbd3XUe/Q6iYxy2ltL0W9KjvLf4HZkOQyEs
HaKExIdSfA4IkA93fMRGwDrjhWv+MtiTWHxiI7iNdwOO3Qep2eXXdlk7k/vIQqKN
7aqzb3xBMUxHfXfGrI3m04Y75u/q/Q+Fz82baxjxIreRf+06Fjhec3OtIS6yUK83
iqQz2tntV/PitOcjVjQEWXzr9RUowuvyEFPk2CjH4CHP0hgZM5fkk0ynDkto903P
EYH6+n3fJkv/xSbN3bD7P3T+dOtCV8/UMRecKS3JU2R0TZ+oWB/7NNs1K4v0VU3K
OXQDBVAj7gYqOCC2dF2mWmziOLGQL7kMisbQGfOXZmEHwAwEzar5dDyj1OtHLxXO
dq8KNODtrpVI4uKkMMa1N45UXyt21x09JTGr0d9kAPBKW+oE2bSHYLQcV9SQm1JP
Yi+/f8ZxgissEqE7k7tCFLjoIwgNciwVmS6bD7SnmkXLai4K1byZ6UK6FdsF6y9M
qqqdwFzhWs6E482jFrldluxh0fNwttipoJnbsTngFxmoqkvaVbl+BrefmFfxrkkH
qYFNMyar2sGT8nZ0AEdNZ5Dsn4enrLgXCYeWXxx/DbkSZIpB2OectDsK6SLQKA8I
6d1rBbpB2ySnZ13QazjjytqxvJQfSx+JdJSIcG8ZydmPv1N17tNzy1yLliizzXEu
vsdHahFgZhSpjx5cfp7/nMt4XvtNHBTQX6sNGlaNE+3aObSQfNuPle3FQJZR17F8
TQFF4iGTdFFftJx9IK8Tid9EeTFFu7cHdziEUW3RT6INRELgCRiL3OUzdF0p9U1b
HpvEKzGtTTYm3YI/q8BzM4/ABpBVGJAClkRlOBMm9/MU8YolkNYdayzHe1JiXV54
5VNnLvmC+dn9irrktVfcAOsoHapa6kos96xU6h63FtDcpRI/zsFHwTtIHYMYQc5C
6JDuDXEGbmI61BPpptJ6AJOJQ4ZLYiQq15RnbddXt72ZNaFOL/Ve8zyaXm7nFD/b
KRx++TDSnSbkcDBZcb6bF9ghe/2Jbu8pZWw5jryOpv0qNL7WrKs+MHjg7KAlE6OF
6w/8Ke2GWYN0uOI74nxExr50Qt/kX9A80CJaC3Cp11fvOwQxIQZEAIEhvzUPyyLZ
b4xm/t54oGhLgudp5Wur22LSk2uXM2LTGs6Qli9SKOsEiK2L89mrMtriOeqAvA8J
mSQrlOPh0/P0fKOQKBDJd+R1HAQilbDJ8DDwpbwZLXIIjs7arCyM8INBiKNss2AJ
iwYN8PuYofEjQreLKbzoriB4WWPntz4HnaoVb4MmC58JvYF2QMog0rD/1Ltpypxb
cuoN09Uh3yyS75V3FJs7ag3ZG6TLHmaWLrfAGD8O3/wti1+g3njJTHUnTMXjxVBK
P/ec7Z+0qBfQmBwMQcDRXjMDFTzO8my4roHxDmY+3Y+a/DKj4ToqsNY3bp/kKNQW
VaGuXqY1uVYck4s78l/JSsKBuha8miLn0Wfpau0QXjHqdTmXZRv21GEQUjB3vJ6m
rVFZS0yDC4v3Auu+N++UgdRaXvEOamaZYF8e6XbiKinkEoEXykprpPdVwM80nA6k
x9qmog7Bso0XxuwPWBKuSKG2SCKnWemJBIoFF52nt0IMnNniJ/HUHwhLjPNw5E+S
9KpSB4U5sO1LT/OQ44qGN3rsQZbZHl33xUCkmloj9Vk7WyZgYYiYtB1enRh7ygCM
lG0xXFlV3EIYr5z31K+YLC1t4iRDdLxTZSyoYq/zcCG2uAJDXDutLn1VAk85JazB
AU4Zmwc5j7IOanBPmkSL4KnXhSxdWUBZ5hSz5OjeuKfHVNu0Fq1haPjl+28lod8A
0ndDPCCniRB2LYZjTGugsQC2ZQD27ZG1e6Jg+yXR0k205mjEI3MKu9MAE8hlDQZG
sg+hCochCGJGZ9Y5MP+I4B0GBzx+27wZrJUChkl3CEmMSeMjXYgfCZjpQzUwou0W
+Jmxnh2+VdGvAiMa+HNjEuPx40VezQ5ilFm+VrH9KaYjNb835TjdfHMzySBz60I+
KQX//e1UtSK6k/1cQA5j2K3M7lgAP0E2OoTeabXdmYEsHUXt4GRa0OORTqYMXPvq
CHIMHheZEQaEhnf/N6guOdmSFX/YNLIDf9aiR23sJR4omxFPVk4rLEGpB23xtCYp
bZ6YxOZx9FSgbvt/xM92HM2iA30WXtvqA5R1P0zQgM+WjunwA+w8Hh2aiAAb4cVP
OvNiIyVJF1ZrQCasgRZ3alB7Dj28QtHfzTPRZmdm/KEpei7Ivf0NR8M05jqplMbd
Pw3vxavdSoMPOyPoFLs9gGuWSzyVj1duUjz1eH+7fZSeblWPUN5ZzF6W8/EfzwCi
`protect END_PROTECTED
