`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mFLeaBQNXv0U+85mX894hQxYb/8lCL9C8Wjb2pmWA6lOSMDbDSvGWVY7F9PTlQRR
lzeXJ+M9r2kslO+gG30w+D7/E/STL1pP8bZTG0a/i0nHF/coJsaVoTvxXYeMpSrL
h6G+jCV3zB5gp0xRGeRsprmwgA4iZxHygQe27saTNPaUckPo0QQYJBnj87HBZDM4
tMXcbZ/yyi0A8aB+xbAwOD61ngOFq1d+vAJwaovs14KTpJWJv3UZxkTqOEJ78eXc
sas/mYdW4jxCOSAJe2ASUg+NwmiLAIsyJWOtyUgkKDRGf4VSkUGCq/S7k3V/AQzC
VNWv+kBJyxD8XKo99LQSTSAO5kq/lvhRx44yv9rsax9IWX8gOHZ8kpV8TlDsCXKH
IpOClGkjKaYECO+cBcvOrHCusLQAUzFMV2/oxfsO53xlAeP7MhhO3zoACpUOWnse
9carR3ZdbAbdJ4Dy3Gs3dR0U5XqC32z4MAxvCuT8JIzKLvtw5Hc6bm/ogNSjkESh
CyQjn/BmFIo1gq6KDa5oc1btb/L4FG2SXAo6ZK/3uQc7Ib49Dmz/LhPvvsIr+EnO
Lg+3SKynQxnVQ8L3wxjEnlyfXGVbt+u8p2gvMy0hUTrMst8lUKo19GrDAvnJnzPv
kKwi6k8lw6XeIKKDWbFAq6TzR59BDlqZEsKYlRpUsSR6jcINATVIgVKGL7DEFS7n
qPAMfY3HwK5hwvrhPmB3A9Ou4uagb2Er0zZ/Os3xwOhBs6bS1bLy1i0byjS/UBZD
ohlF2VGdSVPQPoVSO0885O32bMl3tWY1P+R4Z2K8GLRfBxJdLpBB0+ZRyY/hHYQp
YROC5dgVWBdn/yyBA/NcrPyGNFQWtcz+lG/HzKTbt9YJhEMPI7r189Dwe9aHG8mv
m+zDc3gj/mur77UibZ/fAOcTQHH06qV4VLCzbp2CC52DuWjTmkgY/LY7Brk2qQ84
hCVlXfFjhugP2XR06hCdrBx8SgYOE9qik38tVkZn/j7uBWqjbTpmQIvMUwamivKB
8BiMLQmmT6X02VS5+QcmLAqQ0GtuQvokSsIQSzo65qvQF0nl2/xuio6JW0P+X2sT
Df8XroqpF26IC5ELznQ6dkCeV+o2Wz8VIIFf0FDnHbThO8mkJKr36oBQ734klKIS
QeQKlrO4hv8fEixo+Y/13Gm3+k4OlFokBigMVjADnFWBHLOkAgQBEEp4w0T+fpgG
Ewok9cGJtuldt4M4CCs222P303eh7mfL3/JjUEeAQvId0O9LyYYbUVH6O85VELa2
Kpm+PFQSrzJ0QAWuzy43Sk1QnyPQrdf2ustRAmyQK/4tcPGJqg5dDhgAHvwNZ48e
3NXVp8Nlm6ObFA5kN8AYMFwMemlhz4pfNFeTFP7CFPV5gGb2EsUDDbD4/AHTcG7s
RItULPNWcGreTXzTj7VAreLpU/usmkcjGyx2pb4ubSMstbbb1js20cjfD0H76ynw
ZANxHa9njbziu+UXQ1M/C3h7mQsBzLgKeNajwHUjUHZXnI9kb/fVU0TicpPPTzUO
gc///g4IDL7SyjJMO/oTLpU8vUHOGkLnQLIytCK1XbMJ9+8/cm/lTID8nK99Qpwe
kgQpwsNu66wMEST6XRkkVtcDAbiDtdRV+JRLIH+wqMcewwlLu/10dTERbvJ2/0NH
mEuz2mbMQp02460bpLkfFEvQ/U5K6oDVaspfJxvhm5ipRstdmyA+Uq8nvzTOGsDg
VFJDy3sdSIyWFcd3J5fkK5d2UKnPLw/MAPYrmWf9ei9vk0AbGKeVasKUuJ0YC90j
VchuDklTBCOfQ+cF+hFj6SDCTJf8Cxi3NnDKFSA91ooL1N8WWtM7D77UrvDcMVat
RmOFZoLRiR63QIi3MGrp/j2PB7mL7bVSpHee+KoxGswtniSqGXepJltei4WOpNmt
8XIyClpCJlEvhOim6MCopzITn0jAfbzjEGv1w3LpbEDRWXoviODQ/5zFSGV4XUYU
lgZnZRWLuUl7hoihm5nGVooWvGXrZz+h3/l29MEy/jfgY0YLoMN/e2LdD6Nolf3x
cDcKfMi0mlAzRlnxXxByeJ0wT9FaISMDdhCddkk2XKkiNPiB3vyx0zmyUCXNhTBD
i01a+7wrhfESOru0BumktjQpXHEG8VPzq3vAlJ3dHu2LTtn2/ciBaEQtJ0AbHdkL
xhrn+3px+DZ1Ant0D/Ierx0YP34eEcSPSBdS3At5mK+0nk0PlL1qwAH6ku6FO7bW
lYAkk+f+wswKrcY/ydkrBYNUfJsbdTexFSylQF2k+zUTWwQCtqPkoKx9WK5nzQK1
g/D2UCNk3G/rYNAdC9Z4uYZFcMMGcCn/u3jiYRcbzr+ETCBEA+7oYMDpRIGYHVxI
JoPLORzQSkVm6t4xtCBphoJEK7l50B7amPRsWD85zpLsIIEbt2N8bVXvAu4FU1LR
fAVnfGg6QFY9lnh5llJWFwVzWWYgeKMxWQqi3aA/bcfdZTjHTrEZywIPfBvIT2zi
PsLF51lRZB4d7AHkKf+0QJRSwztesLMlbKeuafiK4v3CMkoMRzioEYaK7YF+MYq3
HNQdFanaZ22KTpWFcIviedY36tw9hejCH080mrs8uE8=
`protect END_PROTECTED
