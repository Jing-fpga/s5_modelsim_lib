`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hUEAd/f5iTQXpi5k3vbDrU+5VJn2Jk+jgrVulyfbtcZsqApKJYskWR3dJkrDb9uZ
Myq0eGuzmey4XUPn7wpE6z7Mvhga2xCIlFU3/G5Pr07J726T7jWhlCBMdUJ2gEEB
uIFl1qIrfZy6hgsApFBxyyuUkZqR2RCM/aEm1YkoGAqD/BcMAxkw/38jYEA7WEKs
3masBIe7K5M3+c3c1hc2OtlPwtCnGatVBvKJYHxA/z1KUffeRmeVg8Eqhcn/3mMy
MvmyilcH8G42hfPOyYTpx8kqk4z2cRcwQyXZvoA658bxqmqrERPt2yCuaog06sqm
otoKnObo9lWGHsxCkLQy941EIR8mOD5ufY/v2r5xZQWvQ9oUpHTs+4Fp73wGY3sO
vpsZwDY82Pvl6vxbmppzUi0aFVAQ3XrkPvQilpLThbJXYzpfrtLRxzBZhd00NBcc
SLBLZqGRvB0CwQ5kc8iK6F9nYUr8Gk13MR1zShG7uQ1mNGKsdAc4wonyLpFjGQ5p
ExCTzRv6jcy5ahmAzwuyjGkbW11U5JOghSUXYAwv/CYFO6ePIw5ThnpEcb/c1POI
AwfKuTf7bGqzFt0/N+7hn9PMUNZb6KXjbu0NMwmhxPwLyvdy+U2dPbFx2ZFJ8c89
lSwvv2pSERjZCi6kYcP8Sr4+5eEnUqSbqfdphbQHwqP1WYcUcOx/DVkEdghwCR5t
cUpEf7gzirDd4kumr0maMOvlcppMzAbom3ZT5ERxn68SVbSIs31FqEehrZGlw/Q4
56eeAecoDsBosIyHE3GKh5T4hkDxInVydRjnui94FWvtVNpT/r3MC0AuXoX5IVau
Isbj90KqeXuh281N72eIs7I1nZIm91Z80dJkByzIm+HanHiSD1p0jSSeaE76RVf5
oqVbwJ3PDSCTN9zQdUej2EXSl59wOxskJ7bmoJqRhFR3PBe4GQ4MVYwtVv4GagJg
2AhyYtWvDf9VJbT5vUdkDK4HftipY9xox/xpKM9Dm/yEqYHRwx6HLg2s0LCmS4Kr
9Somli3DLrrxHiMHtfIg0J153hyCpRPWPRK9QTOX86wlzgBYGiJYj490MHLYhlKs
EKvCiJqUOKdEYK3sFnK2tHWj6BIIfx/PqdWxKrFgBosSC8DEAS/Me7uBusIdGee0
OYVa/c6aBfkq9IXoy8xDlJTeVAqqLBqb+jJRrA3RssLtUN9nV6GAHr37J47CBiEA
gGAnDtFoi95nOnxJ/24/p6tdne8yh+RDHLYWoK2nEzhBjTN3y4Kj0MHhmXLXbyYx
SHUgNOJbWnhswoG3BuvtMvpdAf8OMYhR+NFOIO6yX3VxRK3tjMNMsCmfN8eqWC2p
3BxunmeHlr9NU7vtx7dv+3un8Fu14TlfK98nIPNrpZIZWKszQxRZVd1Z6DDOJQD6
3eWVZd1jciiIQyP54gGcmNTjQxCLOR/5l6t66omhG9rCzHiIhU1b3LSWeG2KyOMd
zDBVBWDg9HkTtXfjhEHWiAa7QUcFXdg1MzL5hDjAjcky8Kji/hRGeNVG7UWpuN0k
Z0iZx3bUZXNXOxDLerzP+vLLLBDSIulLZgFQT+IOXhduADpL9vjwfE5WYiY4gBax
Y2oxGuhJjedqjZ39VZYY9hHTMe4HT2tMP0gT94sbaXWABDvT8QLJS9J7qWCIM/lb
NkPEFoIotoJ83TCxTcK+rGcX+W8EMylvRCbWDdH8XTvvSby7m/t/Z63kkko5cMn8
bDmhJTP44ZRqDjgnyfisiBp98KG36i0QGRpoBRoSYwoaJZSckPbaew7KFmmiK96Z
yYSocnwXZyBbOp4gqsPi2ZZURovUVQJlbbFotwIQS6potJX5enHTfYt4fif9GmSz
p+0AeGpST19UmqQ37dyvjrsMPtV+n4tSW5JePOa8H6X2b+etsT6o0DXkQqjs3bGl
OP8N5KY9gfviHRTQgCcA0V9JRqpvMDAamYtTxkpLdTNNNrdrfCG+HluwSsM3JXOn
HDeLMW8uJOy024qwybrwHGy6aAYXZs77qgrnakJQe2IBprCh4n7+AXMF9PPESRRM
jnvX8RMCOIa6BU5ExQ2BPprg9KZfnH8LsBpt4xUQexhzlWg3s7EOaByLbFMCjiu2
OqjX9BBWSW7BkwKLGNcVCrV1jSjCcdtmiscd/FRGEusN/ekpQSUr2aERwZ8IF8LE
V2gUGF8u41Rg4EsQays04IJQu5mMAkajgKl7bo85oSDwM16h+tevREVJQuabexT8
sScdumXcrm8+xaQuNK+XoAL+dKUKSW+cPUjOxBUUtBBCwi1Fw3oeomFUh6h2ui5i
uohISbhOdFKnff4j3XYarLmkRjU1W8Gb/Y0TPWRUlQQ5EdxHzA1+tcvReqRT9ol/
LOPTm5oCllLlXiWQvcuyLDvCnZBoJby6IDtloz18ddyiUpcMIPmfQpeWC+WkSdsN
KujnMd69L526Ik/oZvST1wR2LlvfprbXS0SHiGpxYYkX1i/PbwjzJHfMXEGxAmnn
03XtRCusrpud8qkM+RpNDbM6YnhdVuohd+8FyYGhlWmwo2dbC4LwXhAZ3AR1m9AO
4k71wyJWkgIqq6UbEFBgGx8gn+yUc+LsSfFvAn4lmgVadLeQqRpgxL87AXp7S23U
SpYKENnmmwG0bDBlJOdZMxUpsDixUF2+xnz4uPGO+PvlkpQGyM1wcQtfn1jjuuuY
5013iIO71F7BkhBuVez5xlD+/dO7uAiCv+BDILf8SsGu4f5hwkbJ38tHIvNjmmXx
ubb27ezeF0G9cbN3fvilebc8n2bbt8iWdaI3/BtY/v9qEd/o91+AP8YtHDRBcZpG
egPyQ2mdvNqBI34/e8GRRh0JMSA58CNGXDVoFz9i5pRfcVApiZ6QpQN9ycLg8GGf
cBQ8VzU8HzgzVJUGohdVgDHjzGA4I1ItM3r0Di8EFyx6vyQfzIc77d0/ogMio09z
cTejtlZIu7x6MjQ/gaBrgjxcVGvi5tve8t6FqDOj0Rhbyvwx+C753VvkA4d1L6NA
lXlUIXO7YjWxxo9CFRuZEPLpZmHbEaEc1k3DvyuPbrhncKpVfot3flfgSPiBpPEB
wa7LhgYdBEQ8vNiUEcPvHYS8aDuJXde6ErTo7n3c1tJG+5BcVtsOa+P0hFWByOtS
aqnVkjnlVRVnjsFokqERsic+pbGUfHilUQM8a7s/qeBeTjAFtjfsfXRpRw2Pge50
j4ciaWVfYVb7B8g7KfLsdPDK3tDz0gEDbYwNQV3TwScelxS1eim6LiArt8b1r2dh
edlmrc/eMBEyJc30rDlvA3+7tPlCT/1OXAhRXF4WYE2sxt7zzgu+3rzWpWBkL+/b
0csA5O90ylttFuyfa8tnGNch32g7EWnNpjka/rjabKStfDYwrBFJ3xwpxSzR079/
SEf9hp7UmLGZtSOE8a40KN8YYiPKVqhSHGQ5MNdzbW2BlyvI5KoXmphM42+YgvA3
WtPVlzd5pR2mSw6wSLIMh7ddovl70uMI3rxi4520PhiL9YeMURODSjzpLgM8o+VW
gC4XFvdGxnG33q8GczCLPZCi6X6xtxiyGS+uetCeIYLTv1vPfnWdJTJvKOKBZKqt
fkNtFqaFquwDb8d5tw2iVEkZHjfh6GlYhn6OsmcnXBpLF40WZW6YSIwDbUGDCXE+
VBxKbaTPc1ZoeNVOsKRQU5dLbOpYom6TRFlqrflhTS3+agLnuDZORfJqJAFQG9iB
IDLJxyTXOuVkutKtsci1erUtxcc1bHIt+t5JtD5hw0V6jOejxRAyVY2c6DUfwMW4
711N9xbdxGMUSwrAQPeY+w3+/aIIAaXwnIYOyHKj/a1N8lyivPOx3Ll7Gon4Krzm
JdaKweXX22JTxmRi8yVyRhcL7/D/eM3zkOPuIt2yxJgMoSM32JrTOpw7eIzuk3Qu
+XWJ59VGr1HlGpx6GnMGxPlbkhzU0Xifo9OYB79TYEtZMPgLfzfWhVTETXIbCytU
GTqfEYVKt3aCXuqVMey6xhzanoubZSyIlvE/9bKJuCdjOLL9IwDkjtOmVFpi+TCD
pkoEu0CNEzRzzTFxmAKMVINlWEL8mAIBJFlmMGZJoIm1szcMp3g5BslLUhbNMeDh
OoB91OgSy1bo40bbo9PqB/ZjU6Pn4jCMWkdgt5tuUiPXIt4AUqaDUu3W7zXDDGHA
tewZb3lE+7iijAVtve+eEc1brNNLd+G2AqTrmymCjMPmRZusNmBA+76aUqvvq/KP
Ej1QF4s0Dr5HdYmyl3lC1D61bMFkeu2Itb1I8VLBL+G15TWGFKGVhhWYmPB+vdpE
a8YDoUa2t+QigsflhYHUDsiruniCSKpZM6mo5IIL2tQn/YM1KgtNPxZ//RcXcyU3
ArVJTX4cZbXXUtj3NvCfGIlYyyrYVlH0Mf0gxwjQUToue7Op4TPrzrExyrkgMeCs
6+l5OAF3Pn3lt6P3cVsOwLNtLryyU0vRuNPHdS4yFORYh56FMkNmBhyAFGi8rLjd
pWLVztPLffxDEDKX+5zj12iGqooa9k1a3wVlwmOmXPDinDEzAq8WaCrfn+JjVcFT
sG+Zj7b+Uyu7w4Jg4xLY/yYxuszL0omCp3v/loD3qlor1KhvJtGkS31zfU7aOn5N
xjbhHZdaMbgxy2PWbAXPYhucOaoyc81zY9D38JBzowY=
`protect END_PROTECTED
