`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ox2C43Vd/N2tKFriwml6NtQOCUeHlsRgTnm+3Y4GbUeFMsBzNvAQn7EWMewNqEes
3bV07Jbcw6CQTWjJjbM9gZLzawyX1JHH9ibyyjMwyhGK2y3bZKtNrewFaiWmTcfP
s/EicqVzYZJoRI5V81q3o6yC69rL8JCdmhpvVFdex+BC41xPVFsvHmzo6DA1Uy0L
Xujh7PxfFkbGdlhY7kibX1JE7gjUljmWMPlOaaCMMijKzQPrmRyfz92fF84f3rnp
Kk4cqDT/ulMp+YHWyCpn6PltshwsxOUpbT2Fmypm00K0kbTIFMyG8CT1Sa9MQHIu
e1SMbcm6Kjtomx3sDqiKtDTd7Iqx0QKE1sWu+oR4aQpY07hG40oglY4LSwxjItB/
LoANpzKIUkpxWe9e46Yal119jj47dnxShClh0ZwCEmKP7wsbmi0L04OIEN4s7kwZ
ode2sRyYD7ulO3V/Py1T6Ie85B9jFTIUYbBiwcyQ8Wri2MLM4nqOS9n6E8AyiqEJ
IEbjz/R/rXkQC5DM27Q91oajjtOeW1cxftYSBbHAhUyPDWKL2b5aXeF891vqGTTL
DtT1z5+Fn0C4iV00z/QKnKV0JcMx1ZeZ9JN40HhE81fpyyy4C+LeDmkG1Gg9vGdL
yA7bBRDmDFDi+yyaEFKVDi3sE/C0CHowIty+wI43Q2iYiUE8eQJsHPhStpt3AZbs
uvZTUZuzd0xDvCjc7KfSinaXbmRDMMsCJIV+DNdUJPDvtNbU7qqt14TakZS/RpFL
a8EHq32s46BWqIoVtiY++tZULng7iOsLPyw5XfKB526MMWmgPUKOxDlwb/KBQRk1
/nIHuY+HDdGTpRVKS3I4xUkNKfIR0w2zZxibu8RYrE9TxkvIr65gl+Ab3Q4khHqe
`protect END_PROTECTED
