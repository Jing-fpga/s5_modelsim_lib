`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r3YanAhAQZlfQvnlrz1kUj0WX71aYmF1AO10v2AIJJ81C9w2CuEaAP5hu4ojW1CT
wJ2uLdY1jHZSb2UFE3dyv92JROzXUntcFH2Sr6zcdcLPkXffv7RQR0s3bzLqWxEc
JPj3EKhCY65YPLXjDIn7Uc1OeJANZyTWgcKQoGf2XojBnjvn/oO4h8CuUzuAqxU0
BqE9TkDeFoesWrIIBOyNjdiBw86IpmVNFNFDeGRbrMBp8TGoPwOfMjLR4RwjbRlu
7S+DIkcvPlG4xCKkor2o3by0k7avWo0f8AnHm+AClIP/KdjSXHxaLtxEqG0eDDak
/+E7U9T0vR8L9QH+c99pe+QC1CMsLEq+NjgIsRN3gJ1uw9i694n/KPs/Am6hyZRb
k3Ll09jowck/8jlM3QbNa/ioJqZPywo+x0aO/Tug+vXvAmyY3tB+1tkFqS8oRVEn
MniQ4C5PX13nSNYX36FLy/vUhMz80S9EBUlGP2ynEp8+2ApfSezQUMJV5A/N7eGm
6nu2OfaCJpNtA4Yj4Weu6FlItpo1oQIjrzDNglAPwoyZcKKh7yuBCGqYN6iQvXkC
jS2GaQlwpdcjtzmJnR7U28GKJ+uskOrwN3ucXtubS59Cf6jQhbs7yI1wJZdbTBYt
BtcFPahLBNxlUGNsFwtFRfvzGCcJai+Fxa0Go95uLm2Q+lo55xJERxsqcrypCbzo
TWAo3b/fBLeu5glBQd5PjNeMRJ3bNphapx64q0ZJ0UlFofk/eO81vzDCeWwpHwCg
RugJfi5IxCn4ONq4tpYzwGYkpAMsceOyNhwdyiu6kzp759wxgBxBYwBQoj7E3zhq
su0p7AZln41oUNCXrRYYNv35Ji4MX+ewEZgEG6Qf7A3UCxa3qNsWHm9AQzoQosC4
pEPTLpv1HIKJaa76t7JLEgL/6+ucr0EevhjzD1nFxAYhgyLW3/VbW56WYxm8ICAo
oaq7i3xEnebpf/f5zuhhORi6rHoM2Dm2HQJpcWwc5eF1xWYfva3mWukSgJ8EIdgV
MmOVgH3IP7rxFzq2RBy880nACocmgd/A0SfA8BbpFzKC9QxNYh9arjXY3406tTtG
U88doc/t79PS9qWeNVP543WSyMxC7oHJ2htzgBEW3yI+06x3DH2V5eEKRxVbTwDK
UKrax3G2b8nXZAan0N9xr9el2/jU4AByaaNVYEuLXQuyCVoRyo+SLC/IovCJpEAf
52+7eBlGHnEUlu7POuO6sb8NLQHQvPygUUMgP2Poa26cx0g6lO0ouOtyYQgQkmOe
tmUa2HiBF2PZWfNP/rnu/rzcRTKA6DbfDgVYnbi9cdccLJp+Z6QFuyUs5B+/CV2N
mGf0MVWMdOfMqW/CsTESH2vmIabWFsGc0aNPFPEe1Yju1+5JKNn8cJEvu8mEIw5P
GcxTW+J+EDaX/WykaVLjt2s0LoWUc9kYfLb5t3+OuhvLIngoih4i/5PwrsPW9os/
KaSr/Dw9YyVply4LthwoTZM+ImM+HpAKqxuVmbdBWfmTuEHwYRc110MS6Zv8wZRj
fWugJYkxGme/KzKD23O1n9r3Q5S4S7WeR+A72wYx0kllM/e8aj97uOMZ8bXmJR7O
tySNQaCQccNexN07+1lJ/2Ej1qVIuRw9AushIVtQd3Ra7eHAl8ZLMB6XQ10B2se5
ltDduGDs4GbY56DWPpfGjQ49tlXOhYavf6tHoIXQE8DeFl+hq+7dkbpGXPmgw3q5
GKTMaQSn3grTTLb497wdoWH++WG8URMIIl06ACEsdPM5r/OhIr9Z7pFafnBfKYwN
p0y5huLcf+5fPQeLHzJ7bh9nJTbecLhTOwvBCSvgSPdaTqQ5UU/ftWb+yMyfKpOm
TA6OJLrBKygTi/7J99oBPO21mPJ0uD++tVicEDGUUAcqpiP3fu1fHu03KXiIZetL
j8V6a6YGQSH52Kc6eEwmo375oIJStg6jdZEs1VVNoXuSMYF3EuXjOCvmMDu9QYgp
ynA4/djlvDv8aPdc3w21jZ7O7zlOeZNjcaYXz5NXgCy7N5Y7TOIG6CiY6Wa7ywEr
GrCs13dIq7r/mb6k5xhEZzt92pFLQFPq8urtwAHxRvqGInhgyvo0elX4uKU7Da/Q
t/bIik9bnSvBiNnjmyAolj2SeY3Y9orPBz2SZcnO51FzS5hSvcazVEJVrd6R+/Pn
d6hjB1itagt3F3xMH0vhpVOXz0wx1Inqv9Zjj4cx/93FEshfEn1pSNxmTSTa9KDA
LxRd85niBjc0PWNIarQ6qj6ZJCs4FXg+45qrUvYnZztbwxB9ELDkuzI0tciPpPgo
W8CJOzC9HmWtcdypc6dGJaMRpwYgo4ey7rSk76LA+m4thD7qq+IQOQZw8B8wUI4L
9Fb/Ubzn5iCf/MHIOTC/0is+2y7FR9YSdjYUa/OUuG8HGH5PQQhxXX95CaGG2+jb
7SKAiqdfTE3PFWo/erEBjwPn03bolo+W6IXFqJ7jBmORF7XXvOjTuFfE9BAQZc9K
R6/qDkRWyJP7liMXsXSn25T4ahft3JDvRLO+dtQxiuCJ3MPEn8JUDkffsNefH/IL
j/3oa4SiPLnv3UNmib2WcrluI3K5RiP/mqlMM4B1fM7q9nUCJnQwAL2UqUg6uy/l
9OD/VnE9/eK1dLGym5L0ixhr1e1HFKTV7lxF8f5Ek79g8rKzxu1doEHYeKbNFjwn
zv3Rhh5L1Eib6PqOGlLpWj98tL2lMcs2HBj1Bjtjg5a1nLxxkECGcUcfUlH9c9pU
EVZqXVW/1cd9qP2Gpc9fR2xNlDUMIh/YIjNnwcVzfQDKdufw6tOb3P1Kj00yiFfF
dBVfJoqAojLB5oIseE1PSsvrDb4m7T3N5daG7na9aKjMOU49kOTAkkAw8KoC13xo
ddvIyY4hsAdDIUOwe0sKX0aC3TFbJ580RqytkQoLfvFtbALcLLn28S5RHZw4DU4R
4hk5x9si8FnDSJkrn2vOXFZAZNgy/Yx8Fpb47OV7GUAvPUQkHMRAJZItFZfFLfG3
jGoigr5bq0fVIyYifPCljmFY6MR/lj9Cfg/mp3FeoB9ffvKD8ErSotpGQMgydstM
TzRHrd1xgLG9ia+CBvGon7sUQcfFii8sxDgQJ9/ihI7B80UDYpdGSYyLk/vX6DZn
WnLSaARAz6VXnIk7CpyPmOai+kTLbteVshqIark/v/PqqG31zWXPB17lDxGz3fK2
FMhpcZJOvsu97BoBuC169xBrDbDB0O1C0XKiUz7SXeZ3AOJDhtBSXqn7/r2joPho
lcCUhom7LOtCn8uAWz33yrsTtdy67CqlvTiTGoWXMrSO6ulDHPczFAXC/EVb/KBH
vqlAvazS6j3IIoQTmzJBR0igP0Y6UMULXHFVbE4dOOZo6ATQNwfsUlEcW9xhCPVz
F2mcj7Ou2o9Bw4HNmELBPIIEqisacBiAxy2b/YzRdHh9wlLYHAn7+cHAMv8q4pAu
lgWDySZLGzHL6SPQ/BrTHMmTd3SXPxao3PUdKnoN89EfjAaD6HR43sd76AzkOkKR
NRomT4Prbzqu5FPs1SOaPeiD9mAxNCs3kN7cLMHKuz+ly4e6js3yJRW3eZO9O90C
cNTgtLZEotdW7xytRNkulTzlnkZ1aO2lyf158UC+xkcxAGqPa3oa5kAZT0ByYeqm
X2bRRFNRn2dagu0srPyJFsr5jEhG5MwhNMTU1IyhW2getX/wGf1g7Qg/UQKzknUO
3Sk0XZEoAUgt6SxjYosXSKhaK3QSL6ogujf34ZOB94EXOMJ0vXVIMqFzX5/1mnsu
VLqT0nGuNr0UvR9iTWXbfpqrO3t0OMUwtZmyNArWDwt4VTPOESnvQiO79e0ZCJvg
TaB1JPKFMhjWf5weqHttUf/0c+jMK9Ntxk5FTn+3swxbu9vj8hzKYZcVf4nFEDbM
gkQxfj08uyG45sa4xATj2sys2DpslAUqwsAWHLOeEqzUyPZaVmaKIGu1AUoQA2TH
ZGt2zCigj3SVnjJm8I8Z9XEvIbGsYCNbzUfONhcQTJ3CbR/nEKksuHSBm/7fBuJS
2k187EdGJVfIyMQPZfhFqdvPh3oyF6hhWMREBAMNNgp+ycWjU7MjL1315LU1yULx
KsmqHgiQjrlF4HTvK0b5x1uDXqagUSmfkBc922dP7DUtMilE4txudYs+6+pY1+PR
gHFi/jDAMuZ6rzoD2mKFxK/3SNReNB8IEOPT6zJ8CrkJZKMyVsc+gI/GG8Lf9UHI
o4fTYOkh8Yj1mGZgQCV9tZfjTQDioxzI++MSODdxajFDcyur1dC+8ZzzdYGRZkht
I0hRBhW36yGwIqyQIhHJ2b3qcDeHM37iG0f1HoPFTj3HNaS2QWhFY+dag1eC4LuF
iIcqpkXjVxK/Ffy0Hw5fFuFeMHNX8S25tdGnhQY9WZTw78PF5lpnTtKDWlIgoEVA
B6BRDnR54HOl0m3m92l23Mry6YlBqzW/B877DlehzCnpvP5uin8xPEAyQ4v8Ic7J
V0P8bsJHmY4H/zbEey5HYydqxpfNh9xX7rehC752i4S6tZgIvP93amEAukAIRow9
IXkT972pZ4VeeKqHCCxISGE9Y0B9s7IhemJaY5rMBZx3Vq/hmm3HfMgbnrPIOVjF
pbpv/p87CmYiqyMXC8T5N8F7P8Jh3gZ0nFflgx/9WhFtq4CWnBVUVqU0sDaDhzCz
m2NjB9sJzIb9hXwIhvwqY0yu/GjSGcQhZ06F/IipI9cf2RNdHhaJWus1ptATfd+r
5f4gnMdTsXN/s5f6XBluqg04mDzbdFN5XqER7D4bOsFpNKiysKJT0HqkJM77nG23
0fW5+kXjzEvFV8Ulxvn0mb6tM8ChuwNxEt8nBIYFrrFopFUZg6HAeBGWG5ayxJOR
GIgfLexZfRa8re5Qe2k2O04qOZoIfC03Anc0oyyJTqB49VQd619GJzYl/J4cx/+M
sSYLz33J/fMIbUsYnM35gAkOt4je1E6FjDaBdhfdztEAjZdPSUzvTxzHHMja3/qD
K/5yIpqLR3++Sx8x5nNnyWOv0n9JHSipaYmk/nao9B1H1suCqDSj/HWIBF1gJa3b
UPyovxf48q3fG1L67uzpDVaHZ/ahX5I/qog60pEsUnk/TcqXjhwFIjN65VTw0m2p
ePlFJtxocY3P5o9+rwf/3P9krxik/lX6KRtrwvehzPdCsDPZ2kgIC6NIB0z9DjxN
ddKcQ9T1/UnY/IVhrvopz7tx8gEwAcigqkc+zhVZN/itwnQN529dCrQpD2mS/9vW
X1O2+5at/WBRMU1GnaqH3hMnBR0zxAoEJVXGhfjMJETmwP3ZFxDPtYgpVRwlmtOl
ZOo+sfZDQIxxYKdgtZR7xnmYdXob8WVSBBmLEYI+sfdnPAuk3mInq7hrC6LuEq6+
nJrF26ulOjH2PLUiRgWNtXtkI8X6S9gmTfXqpdoTVxTeUpXdm5ykrNv0uHNiUZUg
gGN7rNHNbaJEgUJbh9Coz+h0GN+SA1+dRCYxvKV4L0P+aZk0zBZHVEarQn61oqd4
4S7gj8eTlQyM7WM8Urab+qvNy+BsvbzwWPiUtL/2atUDj7noujUtHmiJ3C9yVu/D
FRmomWZbz5hvD9tRw5026K4MlKZVOM3iVhdcilDLfCKi90YJOfQ6jPmNeWjfwUD1
EzKS0VLGxH9r4hlIEbDSCTIaF3p5C5F/rIX/YTDZWYfVXmDCfcNDltGd5CCbSsI2
8uc1ODCxNCwHo5IWdsBRggsSaiqz7bi4m99i3N5g+yggGQ8pOJyxZnI0iVKHteiO
w8HoDHVQpm0/ZPBIG5pS+rh27+yjim1xAdBhOiJ1tWfsWNHdoTOaZmxRxt6QF8+/
Wmv5t2UJ6GfyGvxUJ/f9X5zZP46SHpCKQuJ2dk8XDO0EZIDipgsH0K9RECsEieU4
6cTuFO1zYiKJMKLC1XQGzRSGKTLs0LG9PxR7lK8Jndl1Cw90e5AHpIt+gAs+N8SD
VIvzukWzpCKX3xXQoYFjCAJtZvOzPE6XvQlGyCfly5ipqFY71P/DwOwwV67n6g+Y
`protect END_PROTECTED
