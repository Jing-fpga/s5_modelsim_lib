library verilog;
use verilog.vl_types.all;
entity sh_reg is
    generic(
        SH_CFG          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SH_RESTART      : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        SH_XML_WDATA    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        SH_XML_WADDR    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        SH_XML_WDONE    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        SH_XML_NOBIT0   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        SH_XML_NOBIT1   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        SH_XML_RDREQ    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        SH_XML_RADDR    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        SH_XML_RDATA    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        SH_XML_NOBIT2   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0);
        SH_XML_NOBIT3   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        SH_XML_NOBIT4   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        SH_XML_NOBIT5   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0);
        SH_XML_NOBIT6   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0);
        SH_XML_NOBIT7   : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SH_XML_NOBIT8   : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        SH_XML_NOBIT9   : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        \VIR_BASE_ADDR\ : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        \MKT_BASE_ADDR\ : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        \IDX_BASE_ADDR\ : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        \TOTL_BASE_ADDR\: vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        \ONE_BASE_ADDR\ : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        \NO_BID_LEVEL_BASE_ADDR\: vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        \BID_NO_ORDERS_BASE_ADDR\: vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        \NO_OFFER_LEVEL_BASE_ADDR\: vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        \OFFER_NO_ORDERS_BASE_ADDR\: vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0);
        \MSG_TYPE\      : vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        \FAST_FSM_STATE\: vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        \STOP_DECODE_ERR_CNT\: vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        TOTL_FAST_SOP_CNT0: vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        TOTL_FAST_EOP_CNT0: vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0);
        TOTL_FAST_SOP_CNT1: vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        TOTL_FAST_EOP_CNT1: vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        \MKT_SOP_CNT\   : vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0);
        \MKT_EOP_CNT\   : vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0);
        \IDX_SOP_CNT\   : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        \IDX_EOP_CNT\   : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        \VIR_SOP_CNT\   : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        \VIR_EOP_CNT\   : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        \ONE_SOP_CNT\   : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        \ONE_EOP_CNT\   : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        \TOTL_SOP_CNT\  : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        \TOTL_EOP_CNT\  : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        \STEP_SOP_CNT\  : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        \STEP_EOP_CNT\  : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        \FAST_3202_CNT\ : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        \FAST_3107_CNT\ : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0);
        \FAST_3113_CNT\ : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        \FAST_3115_CNT\ : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        \FAST_3201_CNT\ : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0);
        \HOST_PKT_CNT\  : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0)
    );
    port(
        clk             : in     vl_logic;
        rstn            : in     vl_logic;
        cpu_wr          : in     vl_logic;
        cpu_vld         : in     vl_logic;
        cpu_addr        : in     vl_logic_vector(7 downto 0);
        cpu_wdata       : in     vl_logic_vector(31 downto 0);
        err_cnt         : in     vl_logic_vector(7 downto 0);
        step_sop_cnt    : in     vl_logic_vector(31 downto 0);
        step_eop_cnt    : in     vl_logic_vector(31 downto 0);
        fast_3202_cnt   : in     vl_logic_vector(31 downto 0);
        fast_3107_cnt   : in     vl_logic_vector(31 downto 0);
        fast_3113_cnt   : in     vl_logic_vector(31 downto 0);
        fast_3115_cnt   : in     vl_logic_vector(31 downto 0);
        fast_3201_cnt   : in     vl_logic_vector(31 downto 0);
        host_pkt_cnt    : in     vl_logic_vector(31 downto 0);
        cpu_xml_rdata   : in     vl_logic_vector(31 downto 0);
        fast_fsm_state  : in     vl_logic_vector(31 downto 0);
        stop_decode_err_cnt: in     vl_logic_vector(7 downto 0);
        totl_fast_sop_cnt: in     vl_logic_vector(63 downto 0);
        totl_fast_eop_cnt: in     vl_logic_vector(63 downto 0);
        mkt_sop_cnt     : in     vl_logic_vector(31 downto 0);
        mkt_eop_cnt     : in     vl_logic_vector(31 downto 0);
        idx_sop_cnt     : in     vl_logic_vector(31 downto 0);
        idx_eop_cnt     : in     vl_logic_vector(31 downto 0);
        vir_sop_cnt     : in     vl_logic_vector(31 downto 0);
        vir_eop_cnt     : in     vl_logic_vector(31 downto 0);
        one_sop_cnt     : in     vl_logic_vector(31 downto 0);
        one_eop_cnt     : in     vl_logic_vector(31 downto 0);
        totl_sop_cnt    : in     vl_logic_vector(31 downto 0);
        totl_eop_cnt    : in     vl_logic_vector(31 downto 0);
        msg_type        : in     vl_logic_vector(2 downto 0);
        cpu_rd_ram_req  : out    vl_logic;
        cpu_xml_raddr   : out    vl_logic_vector(8 downto 0);
        cpu_xml_rden    : out    vl_logic;
        cpu_rdata       : out    vl_logic_vector(31 downto 0);
        cpu_done        : out    vl_logic;
        csr_cnt_clr     : out    vl_logic;
        csr_shmkt_cid   : out    vl_logic_vector(7 downto 0);
        csr_shmkt_fifo_th: out    vl_logic_vector(11 downto 0);
        csr_fsm_restart : out    vl_logic;
        mkt_none_bit    : out    vl_logic_vector(63 downto 0);
        vir_none_bit    : out    vl_logic_vector(63 downto 0);
        index_none_bit  : out    vl_logic_vector(63 downto 0);
        totl_none_bit   : out    vl_logic_vector(63 downto 0);
        one_none_bit    : out    vl_logic_vector(63 downto 0);
        mkt_base_addr   : out    vl_logic_vector(8 downto 0);
        idx_base_addr   : out    vl_logic_vector(8 downto 0);
        vir_base_addr   : out    vl_logic_vector(8 downto 0);
        totl_base_addr  : out    vl_logic_vector(8 downto 0);
        one_base_addr   : out    vl_logic_vector(8 downto 0);
        no_bid_level_base_addr: out    vl_logic_vector(8 downto 0);
        bid_no_orders_base_addr: out    vl_logic_vector(8 downto 0);
        no_offer_level_base_addr: out    vl_logic_vector(8 downto 0);
        offer_no_orders_base_addr: out    vl_logic_vector(8 downto 0);
        cpu_xml_waddr   : out    vl_logic_vector(8 downto 0);
        cpu_xml_wren    : out    vl_logic;
        cpu_xml_wdata   : out    vl_logic_vector(31 downto 0);
        cpu_xml_wr_done : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of SH_CFG : constant is 1;
    attribute mti_svvh_generic_type of SH_RESTART : constant is 1;
    attribute mti_svvh_generic_type of SH_XML_WDATA : constant is 1;
    attribute mti_svvh_generic_type of SH_XML_WADDR : constant is 1;
    attribute mti_svvh_generic_type of SH_XML_WDONE : constant is 1;
    attribute mti_svvh_generic_type of SH_XML_NOBIT0 : constant is 1;
    attribute mti_svvh_generic_type of SH_XML_NOBIT1 : constant is 1;
    attribute mti_svvh_generic_type of SH_XML_RDREQ : constant is 1;
    attribute mti_svvh_generic_type of SH_XML_RADDR : constant is 1;
    attribute mti_svvh_generic_type of SH_XML_RDATA : constant is 1;
    attribute mti_svvh_generic_type of SH_XML_NOBIT2 : constant is 1;
    attribute mti_svvh_generic_type of SH_XML_NOBIT3 : constant is 1;
    attribute mti_svvh_generic_type of SH_XML_NOBIT4 : constant is 1;
    attribute mti_svvh_generic_type of SH_XML_NOBIT5 : constant is 1;
    attribute mti_svvh_generic_type of SH_XML_NOBIT6 : constant is 1;
    attribute mti_svvh_generic_type of SH_XML_NOBIT7 : constant is 1;
    attribute mti_svvh_generic_type of SH_XML_NOBIT8 : constant is 1;
    attribute mti_svvh_generic_type of SH_XML_NOBIT9 : constant is 1;
    attribute mti_svvh_generic_type of \VIR_BASE_ADDR\ : constant is 1;
    attribute mti_svvh_generic_type of \MKT_BASE_ADDR\ : constant is 1;
    attribute mti_svvh_generic_type of \IDX_BASE_ADDR\ : constant is 1;
    attribute mti_svvh_generic_type of \TOTL_BASE_ADDR\ : constant is 1;
    attribute mti_svvh_generic_type of \ONE_BASE_ADDR\ : constant is 1;
    attribute mti_svvh_generic_type of \NO_BID_LEVEL_BASE_ADDR\ : constant is 1;
    attribute mti_svvh_generic_type of \BID_NO_ORDERS_BASE_ADDR\ : constant is 1;
    attribute mti_svvh_generic_type of \NO_OFFER_LEVEL_BASE_ADDR\ : constant is 1;
    attribute mti_svvh_generic_type of \OFFER_NO_ORDERS_BASE_ADDR\ : constant is 1;
    attribute mti_svvh_generic_type of \MSG_TYPE\ : constant is 1;
    attribute mti_svvh_generic_type of \FAST_FSM_STATE\ : constant is 1;
    attribute mti_svvh_generic_type of \STOP_DECODE_ERR_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of TOTL_FAST_SOP_CNT0 : constant is 1;
    attribute mti_svvh_generic_type of TOTL_FAST_EOP_CNT0 : constant is 1;
    attribute mti_svvh_generic_type of TOTL_FAST_SOP_CNT1 : constant is 1;
    attribute mti_svvh_generic_type of TOTL_FAST_EOP_CNT1 : constant is 1;
    attribute mti_svvh_generic_type of \MKT_SOP_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \MKT_EOP_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \IDX_SOP_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \IDX_EOP_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \VIR_SOP_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \VIR_EOP_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \ONE_SOP_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \ONE_EOP_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \TOTL_SOP_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \TOTL_EOP_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \STEP_SOP_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \STEP_EOP_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \FAST_3202_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \FAST_3107_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \FAST_3113_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \FAST_3115_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \FAST_3201_CNT\ : constant is 1;
    attribute mti_svvh_generic_type of \HOST_PKT_CNT\ : constant is 1;
end sh_reg;
