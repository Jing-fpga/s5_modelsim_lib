`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tcJFSaa20MC3uPRNQsFaIp7df1/Yua2OL++8r1Kj4N4hqYK+4GzR/WIMbU4jVDFb
pA8XMG0Rjle2GZ6nIrnM+G0AEsW+e4W+Vx59OujyaKGPH5yK6Z/vZy056EursQC3
VdVjtkFYLWNNkTlDGWNJQ4mQLt5uAcMgx5llfvFYav7o7SrJTxa3DpUuTMg+ijO4
6Tq/a41SR8Pp9xWkZpzbTacBMUx/f5pkJ+/5uraNBAXE3lZjzGNY1Pex8BAxB6Ea
nYGXgB4XE/DGoGmJIFvw5IkS/nzUUJBDemhQEX0uwwwl9HfMXlDc8/lWTjAjwuH7
y1PbRo/xOHSeTjNYxOJTReTMvZyGxhkAqcym6fWRFVgL46q3uyhuySvb8Num5+R1
Bd8Dj+HL7DkVDWHpYZgAX19FGCmLYs4KRoptCyvMD/b1mUJ3ZdOSl3c4FsbGgZH0
WFZzVIXm1zEfbs6U3XYIO+RRjFUIpcIjt7ch9jDM7U04Un0QFKAh0Jk7uix3oFdY
o5e+1b3aJPvMswnfmSp39Q44KPmTDOXG1ti9UlWSrg0/73fKHLytl7mnJLfotwVt
mvdiZLln/8/eDyc7mqCB1udlCi+/BS+PYGYbBAzvyNr4JWx/z+eCJ9VKOd9KUGah
QCsOUJHsYohWw3gb1KtNSFIp5eYKCTf5BgqPxMPsKuBa3lbLuHGQgOQj8IZZDbW8
a0Z/n9jwqIENzzbajs8z8cK9wAqknMEOIJo+coc8Z2M5dcAFOaXf3Jk0uD00t2nO
U3ljJd0ewDR2ppRxsysZRpKpqmxWYLJr03ZMwFPMPEo/BdECQqLfH86YApZrTAB0
ILuSoTEo33KDOISvo4/LS4X46PFbVXKiDa80z1Q6afoAcwtLl1nbyPH4Ma4TVWW2
QjRFlZdexPGFkZqfLCFqtA2YFxeTF+xLfOZvyal7kSEO6Y0V1Vyw46ykevjuyGd2
h8Ufdbsp4XKMLsjW7m4P/nmULx8z+3Z5Ue8xMHuqS8a5mr7QShcOJGchBKVmgwWJ
+FcWH9WrBe/xx3pfjfV7OWRnTbZxdNlCVDqzyF6i6UX+7GpIeEnxTFtjJrtAl+Hx
qszl20y50it4en4cod5+P1W5SpAiHidVisrGPndYMy3m+r4BPgkOcrTNvdGmorce
90+Njzjj2d2rUr7HV0Zj/mJlZJmc6VHhp4qCrSbGl103k/2FgMkdC4FfwKR71dZj
`protect END_PROTECTED
