`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
74OsjKMlgcf6j7Kjm1HFTMoe2/iT3UfYxH7apEKD7RcbFemcbg6biJFBM6OWa62j
TRygpA0E8W0xlaJk6+rxgyJDyedN9LGeSdd/aWetQMgrhgE6FoGVFFnVZfipykd5
2Xia93oB1/T6erhaiTi6jVPKAug9zWs6whUu5uih0SpnfqdpEo2mkaa5++ZeWJiP
7Br2mYzcufb35oA9MtUiKHHKlawpYZrF92tRcKvzff21ykWbPpdRAz6XGZerA2tf
9bzEqyQalimqB01SmvMsq1R+Z/EIJhv1xWbysnZ7NLitfriNRmPBkcjmq/g7symP
yISVQCbH+PbowXS8auBmyse4iEizfYiCXt/BgWBvOMar+JciTsIj+D9fMKfzzkEr
nnP3ynCDp+dCOenDWiEcaAJyiveuH4CVuNkRS13ztFgkwtsDvGS6+dNjK1svPIP1
mTXV+PwB7A1BlKf3s3pu/a70IKjj6YLcaSBUNiZ4lXs37/PCAOGXENtPq0BNbuFw
Hi5Fz6SbVxlaLWq83jBF74Kuy+Vl2IylQsZ0XUKFvP6B3nA/8kbcyASXevEmetHK
5CDpODvSID5kc7gbeGz3jyyx+in5lKui0StLa6JgcGzFoSkWOFk4VqDnCYRFgmwV
gnNxZ7hmIz1bjU2U4ebeHxhz5M26ZnZnANDmTrdy7dTmMq3/jPD+P7Osx9Xo1AxF
uovhPDj7fEmlGFPTECYscwE+rlF8Vngr8UTuTuiL95r1V+fAZsZPhTGw2WaAdhSw
d1MDxdgEMmylL+8tAxje0rPrTbAkAyeohoRQaAdvSJqYVEftAcqPE+fu8w99hInC
YOj52ly/MAuPqe3NfYTEYE3NMvmSlwlqNiHVn3ZY5N2RjqR4G2MOKWUuKcwu/LEH
6oYkE0KNYt1UZS1ut3j6sUGTVuGzkG0P7dR7G3SW3dffskmGx8S2hg58D+heFqnx
mSO55BNVjuDr4ODF17lnYQNAbwPr39z/rvCDiW7tuSEYntIK9WeJgGjREvBtyx1V
WK2Q8TkxRG5P/XwOqsszK0xdnEDvohabsRIJHKK+M6IxpjcrT9zUL4Mesl2yBWif
lz3rc6B+/wI/Fi457vBOycWFoW9IVc4F4OLh7rLn60ObE7udnONg4P3AA7D5Fcyz
Q3mUcS7zjjeWmdEZyaJ7VP5RaxCs+XpaIOvrxPWtUL0ak+fjYqe13ABtgr4wYnFD
QLVqOgLsryVBtJ5LyKwv30Ef9tUikOFhJWOPAn8Q6W2J8RsAesYhX5IKdJ3IuQTB
MrAWDHPqMk9ASJ9XV18eDJ76kPsHd3gpufqcYaIVuklV8y9a9qfE3D69/fbl0PBL
R0/ew6VcvrMx8CfcBHiiDIlmHGMYWm553GtIUk8d49+sXJix5NHbhqSCBYGq3pSn
TQlepl8XJEFmjPO3688qrfKuIlSSq30OSA+XnXsMyIpSGl2SlW85QNYQhDzny3ds
DMW4LHJZMMB3p/dR6fTDhShqOBTNl4rt70xbKLQw6G176PvRyHhmSRuAtSsY3gd+
P7GgIuuPck57TC+LxnzPvuNDvFTtX7zRt9oy+Oo6h0Ia8TWusK1pJt03d546wK3P
OycSvH2OfRcD2ZJLgpZrwRxlyZdgXXJqNaPYSo/AMymsZO559cosKGWOliXEQJM8
fJS5VperfiW4Rd9CylR5sanp1Alub3spT29Y/7nAz3yRUUsjRu5HcEQYrex9wXkr
mGQmaL2bq2qau309LagXMBlUnnijQ+XXqe7FRqZhmjJzICBUASrVtqTn2SXdSpkc
S0BJpv/eopq0WDm49AFxuWlNe66Wnu3OF6Key2sor7pV6xbvi/Ch/xHCT0P+wSIt
TpqAmlSJbCcXxvLzMGzDJ35lJJLd/jVpviDTCOwt6wH4i6rWGtM9CW6w0AAb+mym
MYAoRbypyGCC49gSe0moc98T6SvvtuQZJdo0UxaN8ztPsRo6xfV349of7rDb7KQJ
f70c2kBUIeNZjuz8oYhLSf6pXtcAnhs5c+I524AvBA6JOe11chdZqd2NtVTov3T8
HzMtWbETErHE7C4DmJ/O94Bf6544uB1g64izvdJaHvvU9YKglYeEXWRuqQk4VPuE
7ujIyApId3ua8/3lKi46UteaONfCIi7ii/hviQnxu2/8GU+D1KlKhIUK+CVu4mi1
Vn3CypXxeoJ4PfmXC23fEh8JhPl1GEjTVWncgsELmmF2/AINLqca0l8QZOEEn4I0
jax2Fq3IWBlOr3UCcpiTDVKskT1YqW10o2MxmPt0i8fA4VFol7OGlhh5ZEvrkLxw
bClj/dqrpjxtVaZLx+oAd8iSFS5ZpT7VIa7ZrdDXQv6RrkPJWF7utv+gsxYjK42O
4on7+tMGgiD/lt/10hSbLuj+SfSQYsFip0bGSCaeHHqdHcJ/c1Wy3HGMY0YEKAJ0
3rwvHyDZiffo0JRp4mk9FgjREZ79mtO4ljOrcRerqK/+92IS+w0EAsp5ZVa1wLkE
6HWvil3Y1i+DyvL87l+pNDMxKzcMveQr77zNsY5DEzM22ePxljc4WJpRrCllfKmB
a4KsfozbplpOyhaiD86WFmWS9PpLrX+wR0CHnQRjt8n5KYLUoGW5VV3/7EPoZ3nM
dpWqnSVimjOqupmrvA/vwzWzGRVOzCu5Uuy2IuAJrWtu29Dfd8gBa03ueaSr+g3a
s2rHXxyYk4XjUgQMSQkec3WuGkCu0DqMsbHgDpz1EI3bz2hcaHhFqIruFFCH+Orw
jaI+6hOjVlfdohXOcIC9evWjkehkZrqkQdeN3FkIs2Y/UgsZmW74GdSjZLhLg+ks
eLDGjcO/3Lz+jC5hxeUDeY5fx30k2rQFFmAnSNdG7b5gJyT2lT0l0nlhFqE0jaP5
+VAcCtcWtdsOKwobcCKWxrdSvA3eiUBTSA4YEROd93hPSGAfWFKFEP29roI9lgrn
ToFpJhEFeIpnARvQy0NCBheh5eg/NQrfYhr73TQIM1/lVpkVDyrSSm12fCIB4oAa
dzIyRYAJkd3aq7oTSRsR6K4mwKwSyNL9b7030pCQPeEru2Y4GF7K3i5AkMQwb5WJ
6aLN3OYVCYhVgNXn1OVvWTYbs0xCo77U+sIXyFaV5V0kq3l+9G5YMNmQBsew0YuS
hUAwQlepcwmLAH2JgxCrajjgVmNFVDPisiwCyuIb+CPCZr+YZMhAzkKYswOr2he7
4AYl9oQSwugSSnsSClbW3c+UjMdMmIgubZIR4fCnxpcM26QhdVv9OwfIxlQImFhi
5jLBj4sVrK8I4TQSUaCLopnRv2jtmttLKjdUzHPKtb1UPI0Fo7pIA3OtPk3pD3p9
OvDR8x2vbia18G83DIgrxqlfAztI9x4thcDBzl1aIST/eAW9Q2X7P2VIT/JRCFoc
yupEc9nx0TMFFNqRsnk+ioKzQujfgXfaDfLx8YDf7wYX+N9TRdCmtuI8V1fbUaDW
MYxhNJZBnWDbnIm4c//S/U2rVOXJUoEgPLIv+oebtankcamVs+Kvt+m7GlNXoYRm
CQ1By3HivWwLvEYm/mMCm6EhThNuR7IMfAu2E86SBd62hYOR0uzVGGgO4juFsoaa
xc9LANswt0XvnsyTdiMOKm+MHugVw0f+agK/+nfTBpjSRo3CQIcRr/qZLYZNAeXo
lmbtFU8XkWuDc5vKhqMFuiRjH9Rx86JV+NcKvZrXI2sRLgQ8B6WMk7tErGX8L0XJ
Mv1MQelH+g/xTq0tRPZJVSn9o/ZYihF7VcFiaRj8xGTLVdbwkA1996YwfRigOzGq
uNNyY9EZReKlX/2j08OYXs7tJcumpyOogFU5aRpK6Tv4c8OAJoL4PjKEgL95p5OO
eiZoaoBQC5rmd9viIw46S84XzxLK1BsXvaHXUzJLIHwcuN3Pjs73YGAYTTYfLBBz
dbmL6Rn50MBuTVDQO39pZ7hgXZIMM7sDi2xD3qjkI9OAw1/DQ7LrZdIM6o/x/Hg/
vsdW70EsUfsAzH8noxp9oaAlgsIjt/SeBuzIytzlhu7qapXtwLFAdwCOB3gr+3GT
kjhkZoTdk0WqGEfrQpFkr+ED9w8DvRI8ZKhqmoXPWlQt1O+L4HW7L5TfzAmaIGHu
n9SGngCJ2QwFqmwoIShU8ys4kPzv9WIUst/D2vSUb1+r+SFfVMLMlcXSwDYNnxhI
/vM0VCZy96a6XjapCCdX6A4SKrDjQU4+116Wa5uDfQN7+gZQFbJIIp0kHeVhULAK
TF8QPEAX92UcTxVAn0dujtVWb2kJXyEV02VQ4mxCBzkJbQEz7BhzYGTrnlZHMKHh
HmSDIJhjq2Xg5MrM/Eg6NgbSy1V2A1JtcNvmBEvwoiosilHXCOy7hOBmK3xa6mlj
CcOZuXKgB1qs5HzEnio5KEbVlSym3zZfRE/OrCyjTo9e+rcUT42dxpBuE6VH18MH
RIn4MYnl2LDZO0WbaE4wAvVhJkO6KuANbpuvxoXg9tK3JaPkxE612X/3yx3fUqCt
M9FSiWQYjc6mj2CRxdMvIxWrEwEGByzeuPU0Tr/1YwTNb/PF0DNCJujgZ5SzdHG8
1BGNZr2fHSyU7gsqg8PRADFKgzshJa0vfVjHD3EFHtJXy/qN/HV2lbTe9+yn38zZ
iOykwoNEt9EQ2XVXRYSZT7urXjHHB9sb8r+8kh7Tsw9FIZJfBVnRBnbi4+TmqbXQ
mlwFzSFpswEnTZLZArqy9GZlMjVVIxXMbGhvXhVw8wyH4Tk+y4Bi/AieIy6f9Vat
SA/T11cSIF085QtbppsWzseRVMKEtLm3tc8XTCbef60CLOBj8ojkuLXlmExt3VeW
NVOu8Z9Ioxi1ETQUgdfbT3naqCDvRsgwlJfNAh+bUQVuTSrrzqXvCC7NkNZvOJdb
N0awW8UivkKfkzSDPw9qd7dgD/Njj3pK7ZnKEZFf8ybug2lKyMJUs1YTHOEv7BAZ
hICiKGhBQeSiiT8lovzmTdQ5fxBNmY0jMtccAol7LAhirexqK9+FMsf/362hQsu3
a0dRXHPadfSrZXFcVByb1iQJ6aAI0rbLbyZIyz4dySJB13RgK6MkRbgjD9fnexoO
CuTp3JQbKltEpPHqu3RHkiE/rUDR9j5QUSjBebNC/6U+xOX1am1Sr89+An0L6Zra
gH3t7QDl9E1GyGtYD5BTWpNQYGWXad6s20zT5NAmebd3j5eT6vMhlXP1vSKw/WY7
jTz9i6zYrFQNXwYHPPgrmxHK7ZcyhqIHCLaFWlEaXAncWLHDIW+O9Nuw+ivkYP26
UyI8vr1fo3LjGsYCfJRZifwjFJG3OrVuNQRK/XA0g3SfSrjdtlc6CUMkASd0bRuF
+PBr9OalS2GSdkiksq2PEIBsxNEQb/E5W/NeyloD2LyvSTanEXKXKh/I7TeXH7QO
AgmUSP3X/cv9loxJGrhqC1qjMk2D42D6ruwgsDrs5xXbtCxxMMpiVfcJLquzF/ww
EVIXdue5TVYW7Mdc+fXQTqpnS+yYtYZD3x/imMidV2TbKjJUaVcb/75L9kNlIVMI
YTOVNdMFEFIfJoqWi/Man3yrSU0IzyySLFsREmTJS1r0d6G0soMP1d1PZcmVT5R5
iRus9Rbgw5oYSjg0XmdAl+RurMnTPvmYUUnizG+AydTyjKMkKGB+FHC42xrhiMzj
CmiEgJ78CRvjPIvQj7NZ9QeLeVSjkdsjgaRep9HO09Pf2HTgOl8QAZ8hA9griLMC
KgzN0TeyiFBMoZfEurxBdb4Hk5KTJaNZFlOQ2ifw+WSKEMPE9yOtp9i9GhrzZmRK
Dc+2mlJR1AqAFPRxNtmQ/5ncJzgwib96M0RMirNdb/Ng3lOHTnZpC5u2L6xeH2RP
UXfC2auFGnDeloictDrG8NXo4e9ad7Oeuoz1UOiE/zFkJjMELycPRrPgfGa/JG/5
/z5tjjSsK7jLu1qsBF01uILWnx2eQsDkmqsTxbtnXHAiMV/rW2UtrLK70A+jUYEp
RaXneWo7v9oowuwrCtUGVeWkQ29k/qHjknKT+LcrUKcAouUZjlDpLnBFs3QF90t0
cwDs+g8qbyHZvwz9R6mKUdnEyRm1sURZZzE/S6CYkb5AF2jrv6jk4+vY9ZGpFeXU
GBzS8J8CZlluXHEPMqjNnzoduUYK2/qd57a8d2O8Vw6onUyE2lrw2AimSnH+HJyz
MZ5PApvE3RPXrtADRyRxStwNNPJcW6Xec6O4kw5b4NHLNpwNmG1bIU8jxH7OCYLK
qpXgcZ0KRK7HEMDK5uDKorH8+kuCnkz7vsgwhy+jXLmSFIIfY8T/BpiHBqUiDc0+
obKjAdJ65No4EL0fBpx/XdINy1Jjxdva/PEt1AF7ES5SuNuMeC3u4nd2PpGCQPZa
phtTHqJdft5XwLXocKZHRg28ujROLDh9LQfSzF8goSvZXcy7rGXqsQh62YhY4ymQ
5tjGFV7icrcqd8/QfZLhPlKehBnMDc1zgBqSebA0doQhJOpUCflMATQusOwTltIi
CunKaEpWufHEILk1jcsVpXO93US5u2a0IIsCnJ+r0Rxel2+fOhlybZZIh53jw0xs
mQgVuTYC3kpzshna0A7ewWH0wwVdAbOEmrh65zx1xdkpZdnEpWcPIWMN5YkE00dr
qUm0lyXxdEt4gEV+ZePa+XxVpgrSzweOGh/NjmPmSinflgrS7kmBk92UeLAbRcsx
u93ZGvSGSTnUbzwZrXqZjbGNUBQHIxxYWkSMDiTkfY8s+amXmVW38nPl4INHoFwj
z7JLvVUE1m+fG9eQAltG7jd5dfXNn/2Wys+7lLTf6OafMi0MaScc9vMP8YiLshGn
L/2hhCU/5HgKhQGZOPQlPAosFhA3OObAJ6qagNwpmWIDaFg7L+D4iDagska2bc4i
m9ES6609jb7RBaRkKbEoGkZjRIQCKRRTgqd2LUfTf53v4GY/zD1MzeHkvic/GKOd
BB8CqA1nZf0DMHw9vcbmPqzd8mQhxz/lDQumtVyuvNbV25CmqFGQ6NZ3N93CLfQq
yU4jEdFQzCn87pPQPNpnphBorFJ2lYPQFiE4ZtrJ22asMd6bFWFbt5Ai2rD0Erk5
+Cs+y/yyxyOLSjq52nlLql1VVTpkh736w35KjW/UmzDzVf6mLg8pyO98rSaUBByF
QWu/EuCHP+mHxu0C4/Y61E+DHwMf4yGfb2pUKYlCI26fZJA34aUZ2KgtLboqFfcm
fX6Nr13Z3aPoW753hr0mjcDba5Xh2yDLralckWMHapQ1AuTxstFRhlkvmRcjMtFL
B8zlmmnHEHwqCdd6Veno/SdnU+08Ed3+SDBk/nPZ0dq33YUR8Q7lA3dgxqrFTh4M
GIBwJJqLU/qdgxkGySh0nAo+8oZFW2lCns4pODF2ZKS1/MExTyvheO1BIIY9YnJj
rfStQ9mOd17oo8aO7Pwa/7yd4kt5IQ6jWw8k4sWeLbutp6TlB65bTajEOYabqFFf
75W8tKx8/AP0dShnxAHNf0Iy6nsJwyGgdauHNBdp4+EFuRzgNYdgtFexwv3vJFcF
MGvEGtK2xb5eRk2UJx52JQUy/9Kg8ZHOEh3iHK5ZLaQdoH9tNOeuIiAts0URXjN1
MJy5K2sMuVSIkgoCbKBIL4wunDJfPr7G8I3slXJPErPksXk5YAtZbKWzJ3HhbylL
RIbe+pAVqEDHsxaz7om0qk+bA2CVr1PCBpBaVvQV+4VmsRNvQnZ9nDF6TeLJ1NpJ
uTjZF48Lz2hpBFvXxhLYINOk+XTGwRbx/eyRNEPHx+LcXLEEJt0wUMjB337EGBhv
DZ/R4Qgo8zNS71wIxJdtlxcoaWV8fn4Yr6nn4z8nYH294hmuuDaXGA2gO6yoUtAP
JvPiIGEsDkXw6BPfZBxjhsbOEoXAzbNp9EqO2WlrnwvAdxuxSe2wP9WuOOz0zNR+
NzXqJHl0AgdjntAk7ab48nrSWMBkunMGRyc40uGPWWvjwUkbKSHKmlI2AnpERyDL
ix84Gzo06+Rfn1mo7C56ghUmJeTQ9QRJl9kPepPDZ/R9tCfzclePQBBxcf3AkkNk
2yc3wnWUlJEWZpH9eXSt+p4sAKrIF7/CEaAA2LEpwwBjjMTZx3u/3CZ4ctJ9xQIj
th9pYMWjmWw38j6qTmcd/v5ljS7RCzgVqM3p8miPOWs5vLIziOMWwp20Ho/3GWmO
6dQ26y4t1jScat1SGZHWmKEXZ750eeeoWa8kNWYiYOeTeAHdwFo6ycb33+63j0Sm
e6vCVs3ieEzfPXIUW6ObV9YnAq28m3fAh6qIczWfqW2RhwnDrPVVS5lOuSptKkfV
i4jXrlSF8Cc5a+VLjT2fBIlQj2Di1Cq5dQyrNTCIjBh+jTz1+vl6Txdz3I9wCdrt
m/GE442NEIjLlVqpWe6UnvozbmvcYAsCheO03wq03OLWWSjl/Kts2MVYePaCOQi3
JLrR3GXI9XY8FTnstjT4K2wRWdl9Tt7/14iJLf+MfI/+wq408XXfO0+japTpNtuQ
Fe4ZZCEgVeT3cka75jgZGcYxQjoee/Q7DIHbtQNiNYAL/iJgcMhrfSS3Iw6NVdq/
YHsWagdt7yK0toyo8MkEgE84CcJYUArSYC6O4aXk7uJ9ok0uHOTixgs3e+OBzQtj
GDnUHAZuHukoGzeLY4FsGfXwqdWFpSPZ75lBjNibTw0bDkaXiS1Ca7jAFNQ6JXFD
mR7IPEkRMm17ZNnkXu1HuWQQgRk8toTLcSnPHVMWZJ1jMJHuiNV9jx6KHMKeL1QS
Df3p3rKw2oo2BHzItNmY6wEJY9esPKhx6uQACS+Tb460YEbwv+iah7m+m4t82DBH
57X9BfL/0JPxzQz6Ia5qOS6C8zxSEdv9oG5T0Bar318mv7T4Mbh5eV60A+dyZA7x
tqr9YRSAXKVFSWGqlajKMpdl/MbsjJxBgQKsi2Rq7ebxu/77bFQ9dhYXQm9mOegP
182Burqkz4wnAbarH92kXVgQVF7Srkg90qUeMiTrgF1wuBDE2i9ewHqH2eGuCgVy
gTvh8ez/LKIHSwVsCGBVa2ZJg8Hy0dbbuEniWh6pi7VY9DT3gygSHO90yHI6xW2Z
NpNo5ZQFoVFY+mRIVEw9uBlP8QEn//ZnmBrDg43BFkGWy0GKD7THtyOpc3pIsVHf
hjdCJEe8q2GAB5nsGjuPzZo7o9YdQLM0toauSSqs3XhU9UqkrtH6VTKcWxH6s4Je
4HP6cl4kBPMPftiUqj3XXTh7qEG8OKTpAmhbqwNaZI94NjHeOpPEfZngZv2oFCm/
m4eAg/yrvMlhCHLxRRyZMCjLq/9gAJswtj6pBduOlGnvbWiYHd4PbJ0Y/l/KXHOY
yBcXSI1pCvgTyDa7WdvLjkotJNiI8igjjcXHohkqH0M2iLf6mrAKNqvL510WZJGK
NmEOQtMqWoDuvLbC1L+aykkpkXCWEATbmNnlrYHtNK9qrWzRRplyPKrof0i0mQRu
g06Nv+h7V/73ST9ufmZakBegI4n0iZpr/51hhXL4PooWpx0CvVd42Ufh+iDAg9w0
IT4akyKz6MlRde3ZAkFCyBr72kSs3qtI2/5zMK0SKxHOlpapAdF9/XeHgRVJBb56
zDtktQGpxXSTDt0BdpyuAM3kcUevmv01xt2lQT4nCkA3MYTmUJ5Q1yDvUjXvHA1P
kzwHBXzUzKAt5kJkqdoKzDWYOt7Wz7SIsEqz04RlX/TcqI7aOJbQtjttmOHzScGx
Nn1KCOPcdDYGuMRnM9uH38nDOs7/YY77OxG7zZm6ZE+Ud9jltKUjQ0nqSItCIvsP
uAJAoREdo7ZINSgnfwrrbIndFTTAdFsCkS4fjbHA9wgRcSOXTn8tMqXKfNRz6uyf
KyWQWPhm6fUnn/FJqWzAbWQiiYK4kekGYIFc1A4asEg3jmnbcmKtX1iD/UdyOide
w6IDWTz+MEVTg53oW6W8pyY/0iEGlPI676IMia+yprCIp80aEO8EQtqjB0Anjzs/
29oTRUHQ4kPtvQqGE5Fnj8WHHnifeT/lxmXvodxpVuICN3t1KEOE6RILE8g+cksb
LXHrpugmZ/bOAi6VXN32cRnz4VIS/Cc4+SO41oJotR60l91MO8PoNElP68sjNbqm
tntkQ4vIgassrFlCHky8XpNz0M5b/sDRe/9MjVEa4EH2u70Oump2tYGZe8foJzJL
+MRlfK1Tq7sRfgyNiO8vxG3pZNy9ybNrTomUFCaX0rLR3Y7YYebC29OxE6vFvcrk
uYhytEiGmDazRRr1sYdUn/erDMDkXc5MFC0fL3TDjiVzC61myaizugi0OVr/vdxX
CBsUCi4k+H3WUB2EQVnU+cKVvU1OQyeG0okyfDwdshNWj+S1iW+osX+GcthRFZqC
7XBGEADZq1EvVIDCj5idPciuA8MSXkit6obbXKMLCmd+8xwB2FP52GAGOZSrO/gR
7HGBCHc3nw2d/sxKt2expJ1ua6pSpoW3rRstpiMr/Lk74rv9Kf0ILZz+PaVrLbTs
4VMJT2oeLV0c7Y5j3bdNpnKvMiiVfZNf1t7srmJ+TixRcSGeAlK6mT9SBxMhj2an
MCsB6hJ6mD6cziEH01GAL1FvdZ/BmUS2hR0jvO25AXd2xtKu5088CVhaAqupx3Ln
JREJPaAjbgfoMdzZsFVKLEOV6j2aDTRuHyWJ+/SOas2T+VbVo8Bt4ICwh1Mekf/U
qeMmcfLGZg3UNA/DaqmhwIS5rvCuuozENTYZwuikjJ676BVVGsme00B9txaoW8aj
b1tyTZVHgEYLjjoicbP6CTCZyCTndXYxlo9gxeOCaiE4LUmPHahdn8X0/v0/xx7o
IWUA1yqtdyzwuACESX4SDmsLoeVfERPpoU53EktMyIlEIhxAxAKYdn+qIryqUvA9
DJFKeBl9NFoc5yKmi32LJYCl8kOuoPnMy8ca1amYsGaErMz7nj5vbFKeW+5WTspD
Xs7pwcTvwSXx/lextp1auiC0VDPMluBLt7XLtH93k8aYMC5E3k2VPGeE91/o0C9l
gsiE6YBS3N28VN3AlFwSLC0kXeeQJw1OTyUkNYqTOhfbOSHvdcrHc1bLWajpLxph
+Tgn9C2BWs9AOgQKbWxl2sdyh7D15wQq/OUcIYNfOCgfRKrJfocOYlgfAuK/lJ5y
HrzgGm3qCJTGscGvbrXP6VvU0V5F1B8fXf5Rj4gGrNpkz8M9ZbCIjt87IPel9fBr
ECYlTcNHKVvBeL24B8XJdlfedK/p+FhiTmbvB7y2phPi+aWC0lgKSchmHwoc2hgg
XCLvx8+j8Y/RfFeVhzHE0svFdB5R//NN5uyfZWf7hgOIXVdKsWnhkbKKRvUVWpYP
N+ALIn9v1LvhVDlSP9HOvSPy9CSLRf84iZOP/rkGxs0gEe/zToyFpoIlUg3CcT3B
4zsywVe1CVB/Pt2Tgn5FJbV7xiAUQIz5KjIiM0g3S8DNfNXBjpPrkmne9D0Pmad9
9+GiBum7BOvxFdTL6nsCLbsZMA2jCZMqy4t0SzujB3eiG82HwIk9iaDUrp7Ne8X9
/dhJjhkkuCbRtIlPSPnHtjgp4knnKWezCa2WcDE/c9chzsJcHtS8zQ/PGyU6itAe
YDqDHZhu545iwlNikv9UNzVF+L0cRmFRWWF529zUJiWy71gZwnxfUdeefn4ozUTB
JhklG1uRqhN9ZGABmTZlHLYUQMCdPXjqNnyArScWm+inJQ+WNxuoN4aRhx5uGWQ4
kZItcJN4uxDN08rxspp1hA8PHumzYj6PXGPlILI3JuX6AMOELyvzQYmzqPFUQdfe
cXd42vPdyBDf4UVaZos+U4bPCTvbbJFRB5A1j4PjNOEGcbH2jpI3yL6xWEX40XEE
l6xuTr52gTYdPnZtizJcLtXDgC2Ce7Ws/UpFBTS1YFtezV51ZHUKJidA327vxDYl
3clHLOvEe29ZVf73YkB30i59ZGhhbrkGukmMFVOMSOd6hFQv+n3iHDAF7oGr8tSZ
CFLFGwt726TnPrvLG4jjr5hBldpwa980OEe9e6sj/gnCtA9n6AYG45akRf7BP4Yf
aIMx/ktJOiysATqmcxcScpJnmt8MXUlEGouMtRQyy0RZC6uAVayCn3QxIO5Mr2OJ
Bid/q1N26bBP3jx0foUZximK1rLDL7GBshtrYgpn40aHk9toqi1Hfd54B+SHrvCV
ATwxrGFxryTV4RdtWoZvYVcphFn44+bRAyo6qUTmyYGNn+SDZ9pvI4PvQMYFS/7L
peTWpAZ5a8dRujf6CUf4dtR1YHAYn5eEJqpKJlz6Rvm/7DGFfsOtJzjIyZ7bFOqj
IIwEpc6uBb/bKAn2WUV6l5r5LrTBPpIHyp2gzRubg83XhL1D2SvqEoZNKUrSxT5K
aHE4apAB8QeKp6EYH08XNuJZ6k4vZkWaypMduAZ2Xp0Hu1LQf/8iQRpXmtOWaMWf
vr/RzPBMWsZJKTeFvqYje7Q/sytWoVWKePQSSfzf1i0DFntpSVSKby+SDrSywGdy
TjNn/thVw5K43bffImfxcXbDRARahH1EQDzbyKt2HDwi9mwZJcG8TVYC8tUK7UZ5
QDv2LIKcqk142iyb1USsv+XGpU6LTDwL3D4QlVwb4cwn80XbPUUzwtp84zrF/MiH
nEuadxQCCF8Ls3wUCM8ODnoQuR1wb7m4ZPI3t95Uh/mOWrSvYIH16Y8xUisapbrG
hLJb1Ix22ToQTJiaISeXJwEiORWzt3RNmG5doAXYE13hItyvAvZR9s0PPNjgj0dj
mhfDsGHhS6gGcMTd6sFK9sBZzwNxOdP2Sf6sjIm9TaQZyaOXVb+zmJehGd/Yw8D1
rnx8J2/2W03VXuGH3nMysiAq789LkE6mrJi90uYTHIWZItl2pZkXbwHynLlrnNnG
G1Pn3fWgXK1kiErDKqIaqm4CpUANibuOIHTkVjEx69cHtneM6UDZGz7YO+nv5REw
PzrGvj66pidGP01JpGUA+vJE7pzEfpSAJBR/t7sL7n7b9lDA87PSrz2m1EIW1DYG
lwag5hnzkZHv4qfWgcL5a2I8Eh4vRnY/pMbjRUqeUsEi0cy6sdqjZOuKJyqFCIyC
PxeEMRhzznja2Q+0tOIRgJbMHxWVW2Vtc1paoUG4G15RT8n+gGlszSZ3cTDIIcrU
FQc0vM5asZc8eqdbqMLlFBuvlP2F0uIXSRqVVmZceGIBFYUiwBg04mVyWl//aq2P
niMf6hccpyUSotXs3QHw43q9v9SaNKEQ5DDiQJnRoJYntUI4O/veCeSmolEiKOKv
ZRgOg1dPQrjn9f7PXdok8GV1ksU0KdwSLf3JZwb31tl4iTJnbsqT2MCLll9tjLnR
NPtn0JVNdtRj8lAndHntZJMOuBva7nqmeeP04amLfbSOkaWmHIMjTNRWjNZtXUe8
kNotNewB3Wf/qOvzAOLtl7X+BFcKDv4nrtxprBAO1xabqO50EdTFqIO/kqG7WL/b
HPfPPgpCWGgU0BCnEkKiab46htRRmYEfdOMyp0mkUO7rxBi6GEVpG3EB/49Cij4y
0etXVxSkubqKyiqzdqBGs+YucrksLT8I+SagvKw/u3YkeUJlP8WIp/DWo2VdcTq5
ZKjHqa88pECNPZ7IFYIeOuVPWUmj9kGytWnGtDxsTfjxrhIwM8V33k+KjZ3wi3Tz
l4iYpw9gAD5nlzgV4c2G1hGcEzvyHb9sZNrTrSXpQFgYl2O78/IUw1ep/XpET6kb
F0F8Ck/G3M3X+ggJ3B0G2Vo++w2RA9nNWCNt0lWj7DYk3ulIq7yzWWM5F4xKfAbQ
za/i9ts9nVv2sAm5VujqiRuEybgqj3oB9N5jc4iMVKj4aFkF3EN2EzUsETIPTJdy
vmkifM3Mew3Bxyu6RYc0LA08YZMH0VYkvMmqETygNH1FOylHDYpH/WTvl6zYwXFE
KwfeLWI90To6ddCDj9wryQOjIs2r/Y7UkTqK+6gyYmghAkmNhZtzs+emeScieV+Q
L6LwamnitHCUYE7GHwSekTxj6HYcUP9NCqFW1MRZyiZbRYR6hh4FH9/chfuqQuW9
kAABoL7RNfurYP1N/xgj8zkICGqhYvRb18RQBwn6iOAcS5QeOEl0bfZmvTq30Wm3
/IPxHvV6IMWxrhgUe7qph8M1VBEZZmpVz4WJjQJlAAON4vZVk9U3hXzsOqH3gTXT
LVGiklSat4ep7GfZHwQy5oQnp1X6sru7nn0pTJ7Y+Btl2tfwpJehYwL9yYmvBwos
+oTsjL8NBibghFB99t8b4/ZBJq1OHADuJTT9PTIfOjczM1lVbuDwZRXT2jRHiTsx
yzDqyKsli4WqLWbiIZjX718xlY5Jp6XMwVHq+h27Ko30Kj1vRfdlzgr0uVWQ8LWO
UP8PBSjuKgPSiFTj3S/UJc/rY/U0tY/1MseUTlVe5RLtEPsigFn64GowYSEoc27N
QikN+3Ba6on3aHtOfAQgAV7jP/hOm9VmF43PZNK9j0gd4GNC9feXOcIA9Z+lU4zU
Y+4nkn331P1kmrxxpUiaVmbBktuiux581O07gSTAY6Y11qFhPxSfgnvGA/IXXe3o
DazT5rBz31CV3ui0vzO/0qpjQfcxxA6fKeVlTa1ZOwgaFpV7/ukfMNi0WGBlS6vL
MQ9JpUhR8TABUzkHspNUjm8nyZtnBWH+LbM2e161Y+M0n98qm02ewQt4znffWuPf
w0E3Lt/vf8GJJtPbC4/Z0eCoKwpeywkQOqD1UdXOkWmsQLExwNEI50I2BTbxyIrV
0btMB3Y6CP7+V2tUhR/zA9UuejaxLlBAfgZr6nk6c2jmEdo/VyUXdVUqdyfwjMD3
uzMdPh/HoQkJa9TMBlKgyFn5t5KYEUMAfvNR0ghSTki/j9TRDzDFAWTyAtE7t0qh
VSfBBO+nc5cI7O/UxIMB66LHo4NpXkBBXo5axrRQn0fv19hXmje9JZSICoZcrjJy
S1O2/oe0PZYWEDzHI37Ueay0f6ar41AyqsuIHEp/1etQeYz6m5FPj9d8jHI1lgUW
5HcOvDHDSm2V06+K78gwbM2AgZb4qOcA2EiUO5tbvwKoihV6gjinpBzDqQ/YgVVF
SD3jHt02qcMes9wTYQnA7Gip66wPnt6uf5mxhWz7pZksJ9WHegcU5WhLaj4sjMG/
7D8DHbqY3JN2gnY/L+F1Rv8enYQ8aTD+jqCe0sjUjyMM5oWkwsfRgYhnp5Aza0JP
DUELmtpwObHERnIBk2+7Om8BO9HDCmRgQavkTVDeWz4MoL9l/o8JQbRVzsDeH1L8
XeBkeHvFwbY8ghBLw5K+alYJ9pwxSb50BHnZ8jweBt8w19YIt/mKRXeE7V1R+Vlp
HtHxd2hWKs7gt0OcOELjO6Nw/GOuSG91qSbgGWUiEvhPpORBcBQTaBNWjISZHB9B
axVO8O21DMO7lz7gy/36Nt6vV8/5BDpNahJsl2qJcKL3DmC0wMWQv+uCmFfdnlci
OjljgDYm5MpU3kuyrgKxZBnfQDdwAtEzoAAV2JsWBNc9UKmoY4hrjRZ5KKlR4WKn
vykEi5sSkqxtI3JFSsciKZEzqGKVO6HWqQ7P3IKV7yRm7avJpKbHFgQzO6w68EeL
3b1vH62L1CgjU/o8fwtPwoKbLU89S3E7tHFUEl5CeBK2segMSS4ljC6hCFfemEhf
+F9umonXF78xWxaq+NhSloySTtc7BFv9UtzAKyie8akGxk+vTI1zpS3Z+76d0u+A
hK7MPHpKP5ECPfHx5rS0LrgEew/ojaD3iXxcQcru+3Ou07s/1Ws5oMM3I+GYWibd
zUxLWd7OWuY6wbVugIVA9P8D6Ww+viOFZku+z8LBVpkKhIJUOQvKG6SWU8pmOmQH
RS0x5mjZjjkWV0ixUfrIfKPDl0arU2kqh0nhKqUP5CszO6CgNgc72ackgE31BsH5
CjrSwQNAAeeu3seHyyzRxCUvegG+/zRqrTWEfh7bGZbpX416GlPe2yeXIFqTfbEq
1Mq8F7LQVXXR749yqMsKwQToB0QhtfU63wcDocufaOoR4pWKj34jX7zgufTSMcIE
/MZLxJejlA0Y0pB4A9q4bisPPsnO4hAHGFtHRmwjZ/74T329gQqTLBqsiVTBkFrq
M0SrXeBmp31TIs0v/R3bPms88diE8SayJr0Hw6KW+lea1nCfQsAaBOZksxavrpFZ
fH/BYAHcRpWCHK/M2NUqtFYtdt9P627Z6zlorIzxruQLixj1C95MEdpGMZ937Z4h
iUOQ4MX7F+nmcOud1D1PR/3NWyBUAV60x9PScoAj00/lmajrWHdPcmhgQjiVDmgW
CQllEn+jTw9DFaCzvFwmGZ5vo/IMkkUWX3UGPQinzWG3NQw78g0BEdexVbwKpwI9
sO8Odc7gfsW7XAADFUeyMK0AcpE9wlNfcVMlvMwYbmdUDlLZkorJ8uCZoJSSOTpx
tDKocsOdVntK3bS8KpEKkkPGM9Pep01eoBxuiLGZWy8b6lCsB5fKTD3b3/FDB3KC
uZBS0VKCZB4lRFZxMlrBa9xQXA32SvjEQbAQ29MZElsdgTyzDINNkuutaUf/HdR0
Aq7P9n2UBIGls1BR+NVtx5TXnkoR/CLJ5Wvvvm+9hHa5Re1EuiUQunxecj1gSx+2
dDeiewyz6VGw7ydMaZGQ7yh/Jt4nPrbXZFBo+m1x/BdWtddZHD6J0Uejl0wdK95B
LIB/mcpZuApjXw1CEpDwcbwG9dcctwL6D3w2mr9ZLfwKBmcp7okiVB5KTCQNmXpd
05FwINNqJHmI8jCPySXrA9BZJ6y2r4k+iJQwi6ayJnIvhSGM0dRH/rflLbFCcbq0
RNIC1nbZd3QjNQmr6qGV4ffLN+GBmeaNdDhyeg1ogW2bnTm7UNm8k/sHs7NJl6/b
pMZz9Pwt6osqwROoxVNnCxH7lTNnHrz7fpPgHye+bEI+JnElyiisWLQYJZ4ths11
UG4mwhDEYxLw4P45ruPqS1dvRCtpIyz0tAQ4Hfje1ziRRHt1zGJTK/5SEKf2tRO5
hNF3pKu00WoreGv2Nfm7/0SLgU2BjJYYbnpq6lTQ3hSj/1JFCZHOJdSu8L3ofq5U
L93lxSNewZAK8IoKWQH1ocOBHWI65U84Gsr/HQBjp2H4QXyAt3q/ychPRvWAMBOS
3YugdalaVY7ocKBoI2YcSvXpkmjCSwziTI2ELEbkkB1kL0ZFiYpfuYUqv0TsMT6b
mpldiLU8/a1XQUZ+nG6YPoVeUrrjhBLELua731Q1Zs8hNqRIIYnQSl89YPSvuKYd
9tdrQVhzFnE/z0wAOjJUCS23Qx4n4eezpqeA2006lrWYhb64ogI8DMEJ2JePRAfW
CmoR0rBqBslFZktsSk3zikH6WkvcJodrCCJOwSZmEIBkIZjziboD0cRbbgEgMNVf
Ba9EC8RtxcmsdRZoGKx/fnoWOTQgJYGQEgrSwQIybz5Tz1FFNKIMEGUHJrTVRZMI
ln+iX90apdFwxn6sEHOATJzwPa45DNGwPS7vvURU1Go3Y6QdgQyFPVkI2KFQLr5b
6pN3/DDEq+Tjr7FKuDxtNibB1ngciaIEkcGi1SbmBd8jZYRWuAh24NYIfT33y04a
K4qNPSLQz2f5uEcRrTSh2rgifGVJyAeLAMGhMBI/S1RNo7KYmXd8s76NGAoDovAm
hYhlxHsHF2eZePwCXWHSmOejd+/BtsKlsNQOH78NUUb3RTfuX7hY4/peD0MrxQ7b
9QGFzLCmSjEavGog1UaqcQDCBMBJXw1X+vXzqkXuWop/wUhCuicc/KWsqufApru8
3xjPN0KRhhmc8rzCECbwVY3gx1014ugLLia7ua8qjwYGno+C3zD9fDtbB2YF/Ewz
GGkULi+dNPz9ygiIYZQ3XJk4cz0g2B54Nnb8Hwt4K7qgLFUF5SjKsktAItKpIC3h
tjoXvr4RFKAUDJRrc0l3c0Sip2fA030/f230ge47anTJNPdo2+HYdLUBd4k7Y/2U
SaP96p2ivZnqW5QvEqohCmVmzn1xMHNakIX0IfkNO+UwrUy3PS47pKkcTh9jlAZb
gGm7CB6LwXHedJ1sDbR+1sQ0JfXWsV6U908+S8Q7lIyuEo5xejC5bVipeYFpMTRy
r8y6mxdkbTJNmmSvhB3HIINyWSSg8oJR5M6PQOwQlQip7gqqn4AQx3gRsrjlLu2z
1HrePNWjvlvVXw/dq5xYDc1qTBaCp8H7PS91NFxITIeK/dvnHDSWSRUsur5rV/wX
IpPUdQXaXKHhs0B0FN/WInDxjkhXl4+vVXetT0rLjQ0FgLadnxBN/oVamUax0Dxb
ldzHkyIzk2D6w34s5T+SfqTnzwj9s2+7sgTXmFnPYC2gY1p8H2w8S9VqTAS6mQIr
W1XAXxte9GC0A7vb4vQDAIpHX6sUebkbrH3UXEoLrpyR8+BoVEm34DvzUyD1/yLL
O9HjQGZZmE1pQdvdBfWLjVq8jNuLQW2JCQ/RfZ81eghP8ip/GgKlpgqXIgxNqbNX
nnSVujiB1mNxSSEh67TW6uNuS+rBNt8iJUTer5KnmXlQN+6OJx2svrWHsZOiWWUv
f+xTXELoJ6L9KcaWB5SoJl8GxkFStKSi0iQIlw26yQo3g9z6/9wdncR6QnrzcZui
jVIn1Sgqj1wCFq/70u4r3FsFRXMZa9WpPPYQSdjUm4rzPjCTEfK6AEdfdrNGmWdO
FLv1BVftySEYEwUQHzi9xCo3lkLoD1NQ3yaXpznGwhW9P7ym0a6/iDrL3ufWFypD
Y4w83M3GdcxssndsKz2TOxNEX+R1SOky5dXtThtqOjZHUA9Q0xmaZfNLWX8nRUWH
mNrjH06xA0HDsNxpWOzx5Y5jaOJqUqwiMEgATAcG5YCy687Y9zedF4dukq3nr7qc
9uJQAw/9V2JHs2fmV9sB9pE5e6kDzZrrRuKisFw1ctd3Fsk5yMiMhqqTFWELtuXX
uVNEJQJy/vQFfsGO3H2rTvPE+ZKS26AWkES1XAbTLcvjSuUcL5PB+3pd85IpAZLr
2kVWC+0yYCF8BW9qfggDseCnC4MBfjYPxvkuEnn0yTqERI037oB9GbmMH7gTGFVd
BFrSI8jzdCjzVPkC4tW2I0VN4Y+52qSNlK1TH3rpDWee5Rga2OZGYa+2Im2XMMCJ
XJcdlX8qIy64r0MAqwxoNjMrO8PCcdqwCkIgeZ+h4bMd4XAKxI5o/3zHhv+C4M5O
2hBQY4ngKuQzPHjUjYit5xHMRfwxqrF6GZYKpcsodP1hzcVGvD2HQ1VziPA6Fnwq
q7nFwwrm6wV3GwvYjejEW8XJRYiVuoVCPnxLqoW/R4B8OXdM1+sXOLZMM0zSKv49
74hjwmIPyX9eBa1q/NwOxhBN4nMNLoJAqhxB1ioJxpGgT3+J439U3StWAREo+cMT
5QC+wZgMBJlxSxJ0wy9s+TxXvfwAoHmRF8/ZvSEDrW4BGjw7j6cCl2Gz9Lc9c51L
UWey+CFgFVWJda/s+SqfE3PYXEHaOFC6mjcNCbm12sOXuYZZ1VvTJruWtwxboNsD
5tmffOR8kc1GQuq1179lF79QHJZmygZ12ev9CwCRmHqiSiPCT9n3a0u6wmWI+Hm1
GZ4aKvomzdBhhbHznXY/VG+fUEXRkJIKUIDT9XC1bssZKN2geNnMzAeSrN6l6s+q
R78w3owZ9Zo3xdZ+bpWMoFHHVJQcoUsz0lF/jgBAq8e9saXiCuCDl/hRLcI28ZHX
Hl/ychErjLrwYSEs/nDMBiXZ/BEDDs5KBaC6O4yGcnqHihuqbfeF12rmd1z+4bHR
kbbkizx+U+UYUk9pWuh4y9N8+PPQNziF3/4sItjESVsASRqFvYVDKABDLMqeQIiq
2AW9XZT+R//Jwq+hXM6WxGhKNas6ScMHNsFUBgSuoK/Ndc8EpTzK99FWW5BIkqdL
qvwe0dSUHGtINmhHuGAOVXRitJ3+C2w8kJvpaeHtKNImxz4W41fbe1p4sa3mdcoj
8/xUWtjD03eSQse5gJSsXw==
`protect END_PROTECTED
