`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wU5I9BlpvDHZlCjageLBrjuAwsyWbsgnyQNnHdZKD2542aqRRv2JUDTY4pzfsuFR
ZiUvks0IHCl3CPLYsNMeikWdi+KQvp6/T6kDKFBYPjqXLfac3mtiAuN/od4WyYIa
RZ3cIDAaTws4b+p3FkYM2+OHuKJWX+WCQGMf/zEHCfYjjNOGk2Cfv6GvEr/fiaij
bn3tItOpdcGCT1l86JnuoB51OGhZeplYkAMcizLYIXBR0GF13TXhZ0fRlD4rHuIu
DOx0jM00fWIgXZ2ok+zG7wHbWhcDHMCzpUZMVVfOeStVsVz2R6x+xpZkGEeDJhQx
sbfF0N9jdlvygY/16pDm8HTvqcEXhg97vB+Ze5eYH+H7ywTAr/dmrd9OS1YLMIxx
NRZrtoOszxPy9gTKD1/O8tP9q/A9DHcIp2RLoHEzBDeXDWk2Uqhm7CX0/jVF6Xi5
+bqFwP4vwmE7PGC/x06QcIP3J0/uzAT67EMSGIc6FzREU1ColWK55/vErv1KEfmc
bo7WhQ458tYdJhZgRLvTaPRsel7mWOT9pcyyj0GgEwhEeOIVta08jjGUFsFS6txB
BZI8z2S6jfeTdJfL8oniII5IZnjsqslMO7w54+PsmGsVVp/scnUpuUw7lHxQDEd4
dGFcjwOhnS5CexCiKXf99Yw7kBQe2pcASB2Ixv5/jFHA+bKqiIGuXgv3yLGSlN4w
CpewagxnlwLqVh6vdvoI49c9yLCl4NyBc1GCKhhzuTvhWLM7jxkeAssxLBf6wWXF
0mApUEwEOlAaYWsK6D4tjoU7P/w25gshV3gTUUdzHnclxWydrBCarp0FOsuawBL8
CNvJAzDP2tA6abw3/Q1tm/Qen2duLW3DhTdGVr8BObrf71HJbE5zRLjdHyIr75Rk
TcvPQ1nMPA3qNSty99lbNpdr00zGNFBMVuLMvpkfzpwUcQ5k//JcQWO/hr5/l1Fk
TunnGNK6/hvmJi8j9Nir2JRi7hhMuOV3e3nxciug4v+1mNpiGrhsyQhNp2wT5D0J
vcz9Ou/u60wz5ckqZJE7uBc5tlwDhumoR+JafI8rZDFSgyLtyuyhroIjkFLaOSt7
Wiu8EC+Ryyow11iZ81I33hajoWsP+3t+sMTJYpugHe6+yzmFtmHRbtcvgSGCNvuo
q38GQ34oJAIo6Nbksnp6ynoXn4mKYPIB35JOL4DXc7skKtzDZ5uWDWPYG87zhdWp
4xGiDEFK0EkDu6PfWbxbj+cRvgfC0YPyjb6YZGzK6pedLFpFhRtp41+zwzGKBs2l
ECkzz9KjgmSBaO32M5ABGgaRcRD+behzuULecjZPOpPeW/iQIRluRarMbPGWiQMr
9OtzVWVEo6qlW3xifV9MKaTushtbl6Z9RTC0OH+guxyh59WwnWY3FJjXtEe/fdvi
FBiHY0KElEj+6G2OMteIoJm23B51l+xFLX4Xlm0NdwB7Mp1i+9X8t9xiL+afPUsY
SlCGIZTnRrn+l5IlIZfp8mFEyks41VviqsA5IGgOWv/daKA4V7YiqD/nfWZwyjy8
N5nJlln9LFghDbHCkwE7xL9xkg/L6ySVBcAQlnVY4Zwug9XkwKWPrYswFCwUHxeI
UPKTp8Xbv+ijyhoc0N+RFjnlZCVSBqjX+FZi3+KzlSYoKNhD0iXk5QFw4PLtfMw/
Xe0N1P4SLBy73kaIAKBnhleZM7d6gUNPKOlSQwj4sMshsbhQ3ixDyHc6p0H8zlY3
fUgiN3YR5ioan8JcSNhBHEPLjqxatNSUxPLT94u9BFBpPwTubBU2jTZYV18ZzWMJ
3fmX4ncrycgMUavT36nc9HwLh6ybh3dYFR0bvnbVrPCcvgC7UUz/NdqTsJuCGNT7
4pGO2evXVq0SNdMxnnp+VMiD2nID+Vnr5Bf8QDX9pB3cE6hgzETJ4eJOpEYOPnkO
VnU9YpbKCTwoEosl1k150stIQbvsPaNwqED8zcKmw9fh3V8lglVTESBWL34H84hC
3AsXkwIa8s3rYjne6eMtWFjgxXcBSAfcOr3yghgiGM9kDbTBP8zN3Ep5RneS4Jm6
yrd6GghvmXjDW4N1oM2dOi+vlsfYTorN3Gr2VWe3BhNjIrTM0Meii5Z5oNX6Fify
XN9RPrH1QKYI/tvkij5Fkl6t52gqwd7zNSZ0BheWWmfpAzKZkkKlrxWD9fJ7ZRSZ
6QUN4vbL2JpMBi7MOBNuVDqAtdqIkJfIfi1OZg5WJxwJvAidDT0Dt5Twm2YCGC1q
J45dJweiR2fo6qjw7Ae26Wv5FhaQNnUnCRmysFJ529vnW7hqxzHBB0OnPjTw3/X3
2b/7SCBUI7fwFN81wd8Y5IfGSgYyElaI7gFODbEzNmo8t0edQ8txpQIRufmbV00b
Qcmzi785Dq+RlwLHz1aXZ9dlBmPxWqC+njRp0teeTfEHo84AIQV7IrqNqgCiqi9p
a3PByb0kB4dSa9waRO/o8hkNf5GalmS/hYY6EDyyr0Dkx6Sh+/ToYMYM563b6zDG
J8CFzV1QqKxuXRDMcK1ZRboONK+9CwIkUFsGGQ1yHmTw7VQinD6kJAs3l74a++Wo
bFPlmeUd78GeM8B86pQS2Rf1I1lfKe7IWrVp7EwqC0Tse2T56NLg2kDZJejTC95R
+y4/iXiejEvtHO27oK433JEOkJRPinEIQV9h8JKvhkHtw2Iy2/v8qTX9sqyK7TbL
7203hBD4MQVanN8SFRTFUUKX3oTTfVDhmGg5MCthlGUPPYb/RKilL32K6eiTHhhv
5E11UQRXFC1aT04Hiuh4TxRaXE9BD7NdLasMO7SWBgFf+BBryEmPgu0cXhmIacco
lhcvm6LVK4G6JQYGqtKiLS55f896rKuta0i424FiK51RtcRVi+bmrq/ENNKeyDcN
x7GgYUR2HiiytDlaLg9c3DAv7orM7TdwRG2s+SrwtdxwSGv8PGlFoDkMZJvRAtQY
jGEIISEYdK3n3JOHZkO7rpVQjW0Tbfz0ANJ/lhvuOD4ARvZw2WeBLq02rXMqQ1ll
HblsZswWAGQW6Ymm47FftvKSUCKr+knZ12QYqHipdjMsGMcOOftavn8bbSGRxtCo
g9R065NFaa57OAUbFn7D+zpYh+GLSszkW58GmSJTiI565ybJTShv3p+aXZEAJNQ+
NG0BdTzVUXJUTAekGTVBt8PMvf2UiH8HXujeWA0z3rCEnOL4J37lTTU6oRuJ4oiM
BHEcrSRv45ctd4Tqd4PNFT8i8B4AFvDwwkT60YHgRjgCX2pjUerz6Tug3tEeFLxH
5/Yixp/saQGge/fDh+u+GFuYwi7SYeTvtdQ0w++JnvJ2Bkv+0ZWBrXNIoGU5KTKg
ySEpd3azA/6dttjA+09iC3IVYccIoovFHnhOvA3ia3v0m9vCRvt3IOYVjz57OFps
pCeyIM8aXwfqpCwhtc4AERZn3f7I0dSrWzHTt0SohiThwxj8cnm/EL29GF4vbuJK
p11tsKtb+Wxyj+qGC1GsrDdIqmRQDhTo+77nJuMuRqDv89jjCcV9hck2SkUm7vN+
d9G1AfJ/lDBNj9p45KfQ0cw7wpWcNpSQhO65IoTZTRt3tQsn/CUWRJb4+3zRRwfO
8iiTmhFxMQ0lvkluciD+fP9/SqLBSLSO3VJMf4OkZ8iJoZmX3d4asUhUqJh76eji
G7FmF0iKjlC/oT/XTUVXJ7pM9nzmjsR4ErAk3Sf77VxbNW6TjQxVwaL0zYyBQUP0
mVCD2KgE0Gb8nCllCQraq5d3DOjSlunrzXSpXpwFJyZ2TorawiHM+aUuVeSFeuV9
ryeFjKcfDEB/IfQwruz7kpuKlsoVPyfjMch8wa8u3Qg=
`protect END_PROTECTED
