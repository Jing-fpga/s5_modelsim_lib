`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vd1wEWM91XvC6pgODX7izWFJ8lRftMliBkCkYGi2KRAFpxOTSUboJKDUKvsFNkP/
OSDLYQqn0fBrKrICYpvqF/ufG8fntTYyFoufj+qndBDl1WQ15tsv8LAaL/8qCpW5
wpZHDDXC7HcPvdEFRhzu9ZxmdMG8yQ/KpyW6owehYIeeOgImhnyNHvayikARzavU
ssP6HSSsFk209i6VqVhP4A8gR0HO646UBjmmyMzBkTXi9ARYWSMAAlb59LhJMDGu
NhAoIgsw5bDtLApnektwWKDvHlQgMQQWLDZdnbqoyGRN4s3yQ3u9I5iiBV7qVP9G
4EksVSUMIjmMqVHGvBbP5ZrTQFQ+7yIZVS8KEmux7ES4Qg7oCOUq0Pt7pEFQ91e8
XziNDMgxU65KVSUqxS5pLQF6jf27ekekSHofNU1gRvWCx/88ilSlagiiMCoXYf7g
LfIROWUl5HCb+qTNLV2nMXi9UTm1zmPLx+VKLflYS5STQ/Npfs/C+Nun5QcscqgZ
EkifbpBKikstsdCXgRHv9ZX9SifWaqreITuAt0dbCzeORYlBI4r2Y5wQTkD23qd9
7ilyhEh/H0j7HLASEaZa59dZhOxtolAMs6ujK/5bisgRG6eVfQXbQeaoFSR8zW7M
wTwRrrALt9oueW5Tw5bcHcne3fRaecWTYDJkcDQY9Tk0pcWozokq2ynfHwU7deLa
/4C7MQ5RwYsNcNY0rSwEWEIDXsoYoW183lMfVbaJ1Yqt+guo91muO7qzgkYymOx4
`protect END_PROTECTED
