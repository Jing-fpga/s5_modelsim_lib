`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nZY64KhmguOTfmrwNe5Hvh5iNI8aI74qDA0zH4fmgGKegzuuNZ7+XsxnaHVCti27
kaYTKKXpr0aFXHBpVrxd2K1wvcGLPU+2l7FfzM+/l9VdnpCp1nYXfuVelKaKk3L6
diyRQibBPHbBSOOI4EuBwS0cWoYjcIH5M/m/qiYfQEj3QKhe0cOENr4hAqkRdilO
NzL/mEKyeTazJnkbO9HDH0HhqiLRi+f3VidsL/7EaNAI/C8IdJbbcetWGHnIttQF
81fMK8sr5xlKOC5lsJRsSFF4sbyfbMWkDcpvAyUlacX6rrhD/YD+7D6QgB6c/R3v
AOfs0JpJ7wgXWfnhkzns8y737OD2I/mYRhKtS3AF2WJd2fOvgqitm90L0Xl2iDt8
CDjhnwA1SdyzX4yERq3aubdlA5/nnsNsceeqXVdzk+27DLM+NZa3DmpcNkVYTiqr
yr37qgPT1he2hyq0X8xSn7ZaV/kqZCR3wyr0qftJVZhpzGYeoCNX+eBLPxxNokWO
3GM378kyeDJNUYd5FVWTvvhItsAq7copQYFspn4Sb3NLaw8E2kVaZmUQFYVszhUY
y5VPImAxUggyBgJKy9IXY8q9h6/55BIcNK66Yn08k5MP/nu97yoBmTBNYznylI3P
J7WFaIwuKoy7xciHcZSbwR80IRg2+dzAxxzY24B+f2F9zkSD1Uvuqt91B/qrVCkU
n8I0aAXsy97AeEWy1GOnjp/CR1vDQze/j3d+S2y5e6mbDrahEy8wjWeiDFBLH3se
8QsBTARMTbdsTAIaxFBdWQBusOu4qqjM/1Cgmbe3WGY4Iab2Lc7xwEw6f6wJARpi
0KoIDbfinDvE6qO/dIJ3t1023E4TBpxhe5aNCCcjuf9PG+92DRTE5l3ai8fEM7ZD
CqhbIZjYKE1q77d+Ey1JDzClBl9uydlfOj7DEh/d3r0qAzZKLc7m162VgxLLvqIx
sdFcsYFb/RrccrD0NYIFFNdJCh+sEEpTfms4pMQkQgBF071i2QbXasqVtmjpQHkD
M0dqpD47Sv7P2kpXIrFgylJr9qqPH8MjMYIqzWn8eq6igiLkmeChSXxjtzM9tNcw
4GfY2PfDkPaXLnO/of2Xc8XcixMcgib+sHlYhAFtLXcEgvHx2cIchJfx3jM4Vlnw
GRjlYML4sQ+ncsJ1rriDstsiZUPIelH681mhkah7NoFV2yp3mpAxpDYeyVK3e/Cn
BvMp/jBmMKZ0lN8sQpgGPcPb1QbnBjuZRFjopByCdiUuXSt60hX6Kczig3vqpwTC
BiIbcYGDXVQMFb4Keotbv5KxLmgWoo3rcDMdddId/7XdrMj3uDZAHrE5G64e2pg0
6qdA/GPponA2Z1GTdRwJlA8H/Fml9wGjU9wAB3SEv6wo9oqLqnK75+lDPKD1DAjY
ujRPHA/Ng7Wd74a34MrBI9HV/o1RIA31n6Y9rj/flj9pXYxjRRzWZvYyphgtAjQ/
Q5Zc4m/1ozj9FoC4Ok9Zl0LIE/zO8MnMfNra+jbIhObXFickuHreKViq7oGHi5Hl
7STxSAsVICyZRgi/RlCuFlVt5s8s9FR2x3k+T3DVRwIheH9Zrx8nOWsFea8z/Esd
dY9pa0f3bCUHvas0FCRkXQRyleF2Fh2MVzInPH1qx5pkNrWA9DTeF5O8UdqBnpDb
vNpme+q8CB8QUuAl1rhb/JDz5Qat/3t5ELYOGYapGen8sUQqhV2vWmDFWxQiaNbD
uNELsnCnyAngeygSAiE+rfBHZ2jMmSu8oJEtpbkR0vnSxCDYOT+1VYo3ATU2GFYw
trfahYuPEfstn6Fw7QWY4cCPzQ6FP5NeBiOsyKJcrchf5u2FbdV+hLB6fwBDSq4Q
YMklm/994qwVsqW1uNJuV5kww4paWriw0LrQmkMpuzQnZVh74+gjRcJcs6fpxQ1n
61aqkOl+1OlobSlBBquO/v6tmc9EtKMCla/srwufJtZ9AbsvZnLrRi37Z9ROD+Yy
GbMoxxF70MIjT9zIF5avfwbsrQbWuvRroxoDpr2KnuYbfEkS41XeUdytfcwzR4qr
6WuawsBLGH/hTAo+CGz1LLB/s7iz9dBX02Qyv6EOkk6GKHc458vtZTWvHdcUPqGy
ZKrvTXyi7DPsYJQ+D+tlVTQC4VAQxI2IVmdjWjTvnpLYXJDqD9bx7JOE2jGl1Ckq
BPOk6AIM8c/Wa2VJB2jmBhTxcSQbIx+N2UES9gB67Kz/gJ3DaLyExDDP9pmiiY7j
fJSscWDijWp0epizbu6F+b7bqbi93CO2awRZlTe0bB+Lyc/TQCMFesuq/e3DVYMH
TtOvs+7JiMXOw4klzx5nVbKBD7QQ9vPTZbsMGbW97I1S3WINHg+tx4zCpQpsKXIg
tx/2KB4cqngFKhGF9yQA5iV3sowzuXnBh340b2X79Ci4VaZOR+obHGdTI0/SsUlK
ebSDFgmULB7vo41b8TwP+d1sDhP4+b6EEocoNDD5FW/zWLB5AZxuUaUyf8pU1xe6
C71SkzH8BbdaE35BBC/7fOe3K6xYKODWFOyY+S5X8Pc7AGnlSOAV8rkUVJ5XkOyk
+sgOj4/U/iDaEqCeb0qhPULxRdal68d4Wvn2FhIxf8O4IN9vOP42tXlop7R3wbZu
QjaLctD5+J42rmOLRFrMh+OHcTtPoVJ9RHkhrf7uIVero2wqIkALh/z5TU1TAKiq
VI09Md1jL5lDH0eL74/w76cTUxemI59mA99PIbhW6IBQUeDLLzHskezS4L3y9lrm
fG6Q8OquYmNYJDZpORU9vQGnwUZFUbfW+1OhmTzQ2ScgB90LHp6lK2g/CqFMZaxI
mp1oR+tG5s+NgQ80hPU4jy7n/2r0ki6kn03bFrSqgFu0Q7/zlOCwSMG/sf/KGYOh
7+dL2dRdw+73I9hK+Il0orxtln9r53Qryp7QLLeyRpFgp6EFTDN+ghaqrRSRVVQc
jTwEdK55u4UbkhzdzJq16rcSiZOSLQLHFhxY8ceLWlD1onqOGRZWHmPolwG4RSJd
oeRypKzffnrb+CWXIMFNAWmMoI6Z7yHnY4jy0c8La3FhsU7MUvBVqGjJD5LwHcHr
krel8GeUBN2MRSPM1s7n6I+2Vv2bJkNhRqpfVPuD+ylmt33SloA5p35a4OflZwhe
lo6nHqEOP1rE5U0lQgBcEgH2g4acpqX5CKxUHo40cCkI7P1aen/BCPIPatxI557E
SdZrX8y4R+tBgsIvcwMitjWnefxH9vYfJbB+2HFHXOqQjW8t09uXSfs1IBBnJT0a
t/lv60F6LWvCJW2DwYd37CtQazPE7+T0gMfZOaGKEDwl9gdhG9Ak5Z0rQTJHJ8/j
O2ZvXyWkr8TwflvlverFqDMxw6q3MDSBaaB/rW2z0YrLLoVeeGdWnRo8uMaU1beA
5IblBEQdsIsF/nRT05xGBcKSRuOfTCnHIrvIq+C2z8F8R+5sqfmXSjhsKeVykdUl
iJ7HPRK42z8B3PIdI7SDK0aTWOA7rsyqvRsINBBojO2zPd3pF9o8LAZV98ePimFh
71AFfW7PpyXfUj2/ZqMBt+Y4fp2uEJf2IUagb2bUuDMkKPtI9sghaHPrka0V+2ly
vg5rrD3N9kXk5TDVi57Qjgi0UKDTdpS0BLz9amDApbgR893aTA0uwPPVltr4FyeA
zjpBW7yv7FrOXLBeER+Y0oF5eHhkwbiR01Jaw6uZh4o1VWVooS25gQT/6tqh00m0
gymgD/ft0keL09ZveWoGMDgNVB94+lIbJ9MmwnmhnNPvdXhrhR8yUJfjuRou9OTq
XOtcfMu56vxGZwlWHH6CSa9KfXhCdgiX0b+v1gu/+iKmrixP0EibWte3tDVn5LUH
zesYuDxbIYUmxfHdRWhw9fw+BHmiYTL11vX+sTehklboOD9VXMIxewbV+AsGV+Af
Pq+bjz+SpxDF54p6CiaAfmd9qdNB8JQ7Rx6KIICQkx9lZvNFYGr4JVe5bfA3A0qj
pjjOFwJBotbAjo3t/lqVvELDo2zjc6WhoC65jfwo5x0Us3eSNOA8aZcvWrR4ugK9
Z7r0UBKsZLLlU2j+3rXjY3HdKxtgrNp1ER3xViO8Gml33NLx3zM9r25JLhp9BGMY
15fNG/u/hsO+yfCDQ63HEzRNoGXFpIfTfrclolO+k9O5pvjTAcoJowJMr1umXKqy
jEXuXwGiZLhMxitW4ojHJ8JvHHm5uB9/CDKY+73f545r3sNdYBw7TjKtkPZE2Z/Y
KJiMxfZ0eae/d297YKB0mcosqYg3EucRuoYoeEJOvK21VT52KsvznBqcSOv2S9y9
Sl78SXet33Oc2aW6JWFplkT0T6v2smkpbKpG7mEzfsJk+NE1DzXbS3nQdcM+cWvZ
tQgw7uh7qqoqNHJG4k6xGnyoLt3PT1+5z2XkNA+zdt8HWIjuTUbNELyvV1T76vRa
xQVXhOV+LZodXV7mp4dt2V9EKJY0ef8y0+vYZ28lfAkADWrEs0ofYsj/oF6qhc0C
lGz6wu1Fs3BiXmAT3YIjit/Vk+ov62WYm+qbY5FgoqKQz+f3MahBmgUhfqLPV6Ta
yxFdb+HosOFzFMYDYEGvKwZZvwPkJhRxF2LvCIRzWV5JMFoCqU8R1i9OgswLpBrj
TjeJ+w/8NV0YAor5vqXfaNwqP0egS8mzgublPRm/54BnAWBpYACL9bcs3uYAFXls
tQKz8q1RWJLxqi+K8Oxho6J2mhTLLucT6sOPWaNWAt/fppixLsXEmlolKHd3vc17
M5wgMRneoGbiXb8srFckZky4Sg/rS+t3/xY2LDVImW93eKIC1X4PwD0kRQEjYLBS
YHkjGUz+c6coMrFARaNqniSnZ3sO+SKnjrb8WULvCr37RM5TaJB0RZ28DKD5RMxH
IOYiHjLBZVf7Lth+DGcLeuHJ6vbPw3AbuQtd5Nbj6gNn1WeQPAyfgruZfrWO0msZ
ZXkVXNVDLjkzWXYH3pVU82UQOvlC898/aXCvqCAvTk2HtcUhuzjito7bdQInHSzN
lsHFykB+X3NSRieLhvA0YDqNJa1yekHop136T4btBNvJe3G2C6tPWrwrQepPHlvt
y4PenasJyXX9FOQhGm67yKEmpbFDgKFwa3G/dqKFPTn7LaIy2BAiWhZP9tZFgun/
T1G2zpyeDcGiAy8GgCbOBt6/odS2d+BStSWQcwStGPpK/Bap0fIq9vtyW5ARHwMU
+baxiSlN9Jl5ATE+n1M+bkoLNXKLIIC613tX3fJmkycVtQ9Z59kIuCXEAJRs9xsG
+c3FQaiI3ZDvZbDpb4xI0AiIHd62tO1OkX8Q9L4CP5xHe2einfDslTogzMMScQfU
Tg0xg7OWffJwcaW2lM0rq5ZE5UFy+23cmHunIDPhnhXiHbVluV60AiN8NwLXet84
VhKEuGk7kEULDj0yNKV7mKWSHLAFijqbVYBo5fiRbSe1MaxHhoL7E+osE+QrN0I7
x/u/aTSPpbOuWnWrICn3EgOjTbh3/IaUcCa+86Xp7HLXENLlfKiu25rZQtmSKANd
MYsgnaP0bBEJaQciQhm8CkpKQNx9ZgaErJEl4aMIGwtzUDuojqe346NzgMdcHVCg
b+slg1zheRchyA6bNXwJSvaV3iUB8vwQzkbTAvCpwyB67UGEHURAqNm3dPkTClOm
2ehnS55nG9NLyscENoXpY3J4j/8+Um+LWl8jGepwWYwT60G95lhWrZ00CBvDh+3o
bduOtZayOItvlmMSzbXOeMTRGjO67gU8FDBgFCYuldQOdmfEwsRwvFXXkDUuh6TG
uem9jywJEcDTzVBTQbxmifusZ4HNY/7Ltw4tHpcyhD5XfLKlMKVZzNXIbIfF2bGE
r9bzhJx8sCgpBUxG8a5edcniFILv/Y/mtzLPOOA0QFCbiJNiaDWQvGq0gBo8DM8p
Ok7SnGy9iVAGbCIzQNhO7Lh9EN/2HpaSRWd4O+RyYOLXw2T/YSGVvwRYMLlnf1NX
zMeFP5bupT2MXKP76AeASHs9NNz/tU+4Bph4B+2FmZWQra6jYio2foaEfdIrHc6M
bBS1kQbioiv263cUUKz6d+/ybFzqsnir6zZip8xN+U0vnDOOB5YlMQbCf/D8Fecw
l8eW+6QR0oDvroWJJFUEXTnzj/Kz4SujZSDVPrIdfLV/u8YMGYJnJwGcfmIs9/DB
uEpfwMPdvxJ2ugC5DU7uORHELc+4EVcadQBAz/O40KOjPiyzIaJH7bUajuKAbWRJ
hi+3iaPN10rmMRlRYG/zmx/acJ9/t6ROWiKGXamOkfFk7I6ceRNgO3nTDP368G3X
AoWbnj1Bh3iSJbOwBbAJEmp4OcZVzEgCuphVSVep649KALpl86L2LCXxpwzw58M7
kasLTUGUNU5/z6x23Vqrprgpsuamb17IYiaDMEpZUSqUu11thOqkM/ag74IdaeEX
NyWzYs5jd0QOSJDFkEFYgGc+nEhHOu5VDOMFQaFVWh5zpKv7/ZNOk1MG173SJNJ2
19SfqddYtkz6FRJ/hT/02Chsh1FNwoDalYcT/X3VMTwl37P+WfAqgz+5VUUyM4sT
3msRRyvDx9UD1kyD7D2k1XKH/ibpiD3APkV3DFHArSm8NEqHN46/d1QMseLD+8GS
RrSzrNO8vDHHtgsG+fGhKeywnRXY4uJtqajLcysfanyweMQCykR1TvzscriSIyUU
CwUPNibY61SEo8CPjOXRId6U932443DLWGuRS4u5R1v34K6DlKiDUu3w5PetlgtF
YPE8OZCPMCSL9Q+hr9G61oyupO7a26/KnodGoyTqLgYGzPCkfmksaNQRrEn+lE/I
Wpk1uyflg4uqC68BRiNLB3ttSlbo4kPcIjZdhpSom0dC+gcyNmlHsmmuwxebmPUG
x+P/2LM5J672lCoH6GT0C86i5xp7ryj5jUJp2QvHIOwt0cEg9qOHbLiHAkEkiUGe
wCZTfvpsj7dVhkr7ZCbvaqNvI81vjjpIF4i7y4bhQknfZeymrWl8gMs9Q/tZr/+F
WrtINyGS7Wdmy+FatMnOqN/rCXhf9to5Sw02vRW5bWtSakHdDud6xVfi0m4ZWfxG
gwTA/uPXt5TPKhtFszFJTFijATf8nVRrawMyLHmlMkwuy54ukIAzjWia/0+6HU2j
4t2xqVGLxnnNvmNNiKJQXyY0TjjSNffhpeAtDqy3IWgFvZqhoqebiWfeLBo6wSSY
y4bKF2yROhgUEs1wjxMs8h3jDexrCwmpEPHQVMCoHaYrbsMNH21O5kcxTokX/0qx
fLDvj1L9aEXyeMe66Ee8VRI4aPk960enZDMU+saIX1JeCDU02XQthuMstUlrZWZL
SJtAiTD77p3C7O/m2suNMujbgbu3hw1vB7VyykS7Zm68NDdhmcLGZ2lj3ghSR33e
gnb/Y4ryzDhKfWtlZykm981S2Ob576gzBtDmf5f3M1jjR6d+gSNPPu9SdNqvg80F
T8WSHb4Afb5yWMC+nw3OOM9uInST3jAK3PvWUaIXQlppIwn0UDNtH6VJEi74kByk
/rGHHgpNq5jrI9YJNvqPeS2sNJ/KXj/c6GWcq3bdPuZ4wvDtVqTXl+6SlB0SmZDL
ef7pnM+iBzILBcnPExKOZ4GMw10KW4wv4HiNvLLCZrHBIk1iOh2btARy0A4JkQxs
jq3Ffl7OKh1QdhlWTfnYvtmQefVmmGwKTOi3Q6LrtlK2K9OJmkCAoZHRDkGpQ80D
ULIxVbS6bCC5HPS/0+ZNwLnrSKA0Y3DZ0vkhqtmKWhxASn4C1hZ0gJeV0Tv10kMl
EOmvqmougl/IbOtFOMqrQBWlk1IUlPkO3G6xJi8LkNyEdesm9rNS/KPdpRf+D7s0
VwW+DWExcIpeDrZKE72s3b1CxDLHTRnI1Vp6ALbh80DiCLq81FnLi2T5bQfMU6R1
13a/daey/rRQGgLXJCYhFHoDctwclaBBU8DwNnykAbsh5Z83qxNlJ9gIhrCAHoa8
0KR9G5FxQZoeiAwsD70EAMljLOGb2fD1QlZ6fuTyGJnzxl+pKiH+iNnaX9/ccu4m
FIHvUfFN/7ZfF+V2T5flOgQKngzqxPxsoxNLBCB6HkDbjmQtInt3BtO53UlYI2Wt
iARe+eWR8iBrivjIFgLt0DQbKkUYDLnJuVowH4zyfYa55KiLXiiCFalZtwnRs3/1
x4ffTp/gg7+eSHpRkxQrEOjSRWnYueesmRUibwAE1eo1Pc2WbQ/0qDC5REUK1OTU
Fk74I7s67FoVUFd8FOwk67BfiPGjbFaLh33QoOKSZTfJDzRSFNtH35ZSZo5PG7x9
N4QdeEy9iXUohFvXyS7Lmq5Y+5d/z/6dpJXHaRT7etsDR2FDdimFdU4mG8JqgcHp
WSNjdn1o6U5eML5GjvhGqxm6RKaMzaXNLqAAT+Z0DTSP4YAY9oujWFIkjpNitLIo
YQGtKRLrbI6EWtRDhEkWoOlYy5y7sJ2ikD0oQIxoRZZdThIfn+VgHGOzNI7+Esab
P00Qu/8XRcNMxigk1UPY0kjGqHBSLTacNiofM2MMCH9WWF+s+CANqDo0Q9DOd+UK
NCRCk9nhD7LmvE09sFJEhYLjy8XYxlgQ9BcT9kG8G8L0cijFOPkxBHw3CP0iFv2C
unM8odGugxPtAP8mf496NcmKljPVnK0NsWbYVmYXQfvzuv7JVHuqvL/x+rLP4SR8
OCcFMQ2FvmItRluV8d8j+BoD+XXZkQ0iloUKpooj9Wfn7piEiCBqIb5MZZRvOZwZ
/P28xoqpHzxw19E/A1qWEIpwV9pmCtJRaeo1zf8o7E9ROxYTwViKpH/ii2gOoFsU
WnmwDGwQa/BKQTuqbxAx52NGQ6UCO+B1WPIG7JVwKEz5D2xJrEJlkQ5sIoQ4RUVG
Uh+5rohbehbKLw+xR639qQFSXpffoK64EDw1edxjsEFVXHfEePOig79yvXJL250R
6PiAB3HU/xNifU65o1byMFP7d9E2tk7AWn+ok0U4NDpAkgCk3ShIGa4PXkyBG1Vs
9RW24sjZcCgo6k5co4iFF+SZgkyzVbTWUKSFe6d7zfbcicQWEhoBgzkuY65xEc4Z
DHnp9ltbaacdqYLmA8NDwo2oMlOfjZ6P8J/fs2jqqgF4viWvF8yfOpA31YAkGz5z
uPYzcgNQShdzpPoqKHCEluwX5uw2v2ysXTLwiguao0mvQfraGYVVfLRtnchQoyWK
iLLRQ3LFVkiOFNmDg7j/q67wpGmTRxmN4vbu/vQdPSPUHDhb6hvY7z1tKF3Dbt/P
rUm78BQT2YOq2kAtKxHElIC4R0/MHq7YMBoiqlJ1gTMycsBqAH7oSkgDY339oNHh
zE49tzuWZNs/k3UlATs0Tqv1/Oi/qE45hcBWrK2aWPGas3ahv4VjX6tfgcExKpXR
/sdIHyac/3lXw4hWjNH+Pu+93RNX7L7DOT9ifqQ2WPfKSqWsqoRMfTvIok2xY8IR
MIzafhZ9V7BdgrhFTWWAVZmNvvle+XaE9MwJV/fsHmgeIPyVRw1/BX95jo9KtNLG
DIhTRfX/G9KsbC7vJYgv0HuVKd2X5OSIUIgk69jp/6P76BC4bPQUg+Jm3eyX75J/
tLwVvargqsk/LrdezAbz6VutBrdyf1FlMbSuWa6cWrijZsYtHer0GBYbGpSfDmML
X88vqNpg37ycmKradIKBLGuko8IsMt5Ht6H10TieLNCrZJXDaQbFKRt29WDRz8fU
POX+PzdQnCSbFtPSYqlQ3/aWlzh/FytUQjhhmJafBF3gwsu6fDJYUpBRGNwopcK7
rZh1KWx5OXiRaIS/zs0kOvSeDx7IO4Qb3p2qScNpAqFfKArSRj1breq5GaTKMiXr
KpWXDpqwcWswDJ7zsz45zikc5UAgSMNtSgkEhBWFWz4gKTMDCyJ6VaKccc7ACuRK
tiZwt6VK8UQ+apKgfodgl7ng6JrXSR8hlGNrWn8RrYM3Wu0HPmVuqMHKp/wmC6yQ
BPmgCQI9s9IP8SYUF5yY9s1jvfupu5V8fpvtWUGxsuZjjYpyigrx0BHahhnBSeIh
gbQewwqvrFYM6U1+uJ0RptS0YupwSmCBARhty0d194FNfHbqiz85/kv+FBKEBDQ6
DVAtlecGJxxMO56qka3u5zr1gz1Z8TGM89WGfxumfuj5ISX6pVVhk0zmC5uS34Ev
QrsMOTSdY1IrLbeES8Mmse8EVkVVGFnqGgSiSVRbidYUn4XYN6BP2txUfQDkOqRV
0R+j8GsV1iAyNtKMKTPIVkXLvIjacXNNdKeqt4irK4pnLSncGwLdHh2n6j9W7irJ
jN+w++Zwkm43xSb3g1d08Wvx7UkuT+vhgf83Iurj2De+sC2hlDevuwIBryHKcPB0
+Ijkyfjg9fvRscLHGvZZiwSflV2UznqKKeYzPpSwDOFxy2kHcdU+tMalcKTyxVkc
gm1z2QFo/KV6qsP1ISBfVmydXaPVx1rzl905fF5Y6fIpYYFI64ZVTwBPk/+zNl7E
jaI4fdPfVklv2OzdFdYsKO45sR0HGlGtOC06NZF0nS3BKfy0vwU2FSugMbi6KGMS
4MLb97IBhhwqqeaYSyZXVFolNlULDtK2zi7H7ZDhuRuqZ6B1mvBLB5VqjGMjWrMi
23PaNRY33ltWRy0PVDmgzyyq4NCYw0cEV2UpPp5v2blXrZrtepTRqffeES1urYcm
pDB+KtgJ0tHEUwc777EPKVQbbEZGWihyl5e/uSDt9tzg1Uqa/s4wfrtp6Z5j0l+l
x47HNcgXrXr7LwUkSMVzj7G2hLNSjovjdhOTWmsxZ1DcLyVbBFeaUzISV2W9dDbM
YyIJA3AwJQp0yorjqrGWcSCgq67/xeFfMjbNrFLKacNwge9G9SFG59xPZACyesLI
J5Boam/MSDphASq9O8yKtTBkefg/MZEGVDdSvPxSD9GD9JomgEU3XE0H79xNyQqv
GZzA9IvSPMXZ2R8Xe+RLDQbUPPlEmNiNDdqoUmkZHmn6fiwgfW6aDJp6h/EDCVN+
iuquZ6sR9Lfsy6qS0zz5h+uUUPLJBDCAGiiGPv23UfAynYyw+lFLuKpBUwB6fnJv
97IUCylBb6MGlBTvYWMhOxEx3VDcO4rRYA9QA24lYdrFHHe3qcfG6hXrH8fSH2qy
bZAop8NhH1nP6TTQj7SDOpKtk9AbPTamcyLS5Ly5oABhxnGdn7zHOn4JiphNsp4e
orScC/OZ+YEPhuZI0HqL4iCx9BQl/uAhkoRLsmNDmdq0GDJ34ByGdsYnfUPqYq57
TFreKUQ6GBA6YwhXv78dHYiYQk+KAT1H40DuE/M6AS6yfhi5Q4dDs1sNSd2eX8Lz
Ss7lCXI3SAd5PNAIa4OeKhHu7HBDIieCmAhwPuFbIPf/RcelKmnJQjlEkncDUCMR
w2SM6nIThBOqLeTn7xv8b9tFon8uAq8EC0RMshW7Q5+yASZBFOjJxGcISIflTArB
0g9juulJXSFIGVY+j9Vm6sf93rZH51e3ub5eEPYXhmDZN8cKoVvbPg6djiOAGtO8
ujk+XXspqXyWuoG9+51hPCRvfdNnBWS0yFcRdLUteWHKwApa4zYpSfynwI+pBQpl
XvWeK7IE/WFv0J9xXmmMthELPoFBRp0blrBu1uNqVNwux0tuONh9UEeHGimuZ0Uc
/w4nj1KDAkI2kjkDIO6QZXGKPCET2+JzecnWTV56F27NLhXoxIgNbYCfD64jwsnh
1L7NQJ+MLPuJ+CSl2M4ftu+wa/yCnc1EKA+DUYEPdH3XzJsH+ECkPSGc1lBPjzdU
bBrZIni98+Hevlkuh4qb+JMhUqVEoMYZtD+L9d3Hvza2FloXpLOJj4ZT0cVLpfud
kUOvDWSeRywVmWfmBArxHpR3O5RbWoRnuDg/jvpwkJNTasLRED1nd0SGHTe2oV3c
ZZVDKcqv1RvOzgKNIZZPlgaHw9Ha6/uipPYs7DcylSUQJ6FjVifrj1SH+6HyNez6
8UfecWIbfXnG9xRma1EoR1uWVwMzUByZc3cs49aBeSDGERy3/W+jSMfJOOPMkmDE
tcvT/+m+bzr8DWGpD4iFUs5WZxE1nRlH8xxQEDntDT6bkocD2ihxvhjomQsVVa76
HCoH8Dp1oXaKpV10FZMkN3a72ukZd99r7pRKN2YN6qUEpiYS6wGBsxmSt3iqRIi7
ek9vFNE4zixerqc1q5/mZLEQoRr61t0moxR2+5jUew493V3YcNeuehNFmH/9B08D
+eQUqxNS4+1krs9tG2QakgxEOgbZw6wpNnOM2GWAsUuCXgB7fkc/nA4SBU+ew2d8
Wk7g/swG4eM3hK990oc/CA+65egekIqjzwfaJmcZ5J+QnDJwaFiZjKWZ1a45JaDi
2WQqO2vSGdhs0Du5mXTLl5UF60w0BkFQFGcACA2rpTmlfbltV45+QHv+VyQCdQLy
KZRFEXLDhgFYAPZAz0mdJHRJb/zh2aK0l49dMlfIt9s6efDHa8XAZ1ylZX7hmNyI
56PHdFwnoEZyI8wsUXYS77PTP3RkK9SKMnBs7csRgugX1wj0AVsCymD3RR3IRvZs
eiTkcrZnt47ai2COPXtGgYospoIHD9RUNNRn4Q/1MKRMEGW/4P0j7EIxJHvDukl5
ABeyQBxa+VGDgd+KUOOJoksJIc3oxTW7VPt+Eq7m1vvaehL5SQSqrH/fIQWkBGvE
JFC9SzUi87EkblBR0KeANl3e/CVb630UTU6MzKqmP6xB0VFF2Ihv46j0ZoqbkXKa
DzPE2WzF2+Vdaw4kh104WtkJGuOQacwryjLaCxwJyFVHZRfLXgDe0iyK19abTh/x
eYoT5qmEEQlH2kWzY7QbZePGeJabawqJIEtSVDEqBusVIat+SO364842IUCd0IT3
P+zLZnCW7CljVhz32ahmXIFdODvdx+SQgO9md+F4iRboqGodm4rwI27n6EEuqw1k
3xUiyIv7OBNXpiVyzlG4yaSd6l6GpNcWx4XzaBBkqcLdfTGH7qRdD0GQ/xPqj0wy
dr4sQL7qjx2M391mhJLYRjFebsm1NwyiAJC+PUMothhucqmC0VnqzAH+/IHkTobL
wz3e8VdkVGO6Y6WjzYoUxxO9WsNC6J0uTEFT0ifglTI111nw3GlV0ZeofTWiwkzB
Y+YSxqR71hrRa4YLKe5LJRFYrB2hxw87sdVP5Lxnq1f2jmhKXILR7rrbKRPkzf/6
G4YOlsr72XUuuQun+HOEpSycF/4lWKPQq76qSqES2M9TBhVt/Cf85OVY00evo2nN
275Qll75eoAPErY+JSf4eoKI9aI+nc3JPnudmL1FBW5NXk2hVwVTZ5sXD3GV1pjp
FT/tZbXqPoZgUNiy4tQEgJRBO63pXOj4JERQzlM6LfFNfTexPHKWu+8m0+x4rbc6
cjQ6am5nzOHl3bx4SmIsOacYEu6bQ5xePYSGs+sGthfOOna1uCrv254J1ju6av47
nhO1sKG7roSTRSKA9BRZLrAfJ+Wxq+yJ16TeSA3XuxYZiiefwDZUFZGgMTre1agN
lOpB9hrlbsdXTuBa9paIiVasgM9SZb/BeX4mjue6uVjbN/Px5pHfj1OeoUFxINyB
nYKmSU6HJ9D3b3fPsIcbF4CeMS6UFU71WYmDL3EpGLK1FpKd64/sq0faQGnbaX+q
6XB55ESDGCVm4jn+oYbl3+mzGh94DuhF4tiF4t+sPQpPi6QcKFROJZsEDIO33AzE
hlPgBz6j+JlsZ+T5vQIFWFcuxUc8Ida2W7xPMKF3ErBhhVhmz1PN3b3Yn8DR5W9w
0f7AhScvLeUzSTx7eQ9S8VgLUGq5z3oUFJPXiByRobwIW+aNn01SWsDMvW40JClz
Vr/25IGicz+pdJBNTGV0B2FBOa4IqttDZGA+1wQxvbPkN2M+RLF8ho7UqgsvaCNC
uin92iCP5Vj6UEDpQapUoiqLDjLKxaOaZYv7cdvMbpIBKLCCcw1VSb2f1LOrlhC9
Km92GDQdhCcKQYf+5OlHncMzQGVuXui4k0ZWhWO/Gj/WP0Q2cWSUNc86E8MHVRnv
2ll/Iw20kusOTH7yzAynyYaioYt/VVtpVkUYYlRh3/2jaghqKZe0VnmAO7dhAYsl
XLV1W7BZqGVeEJLNWwFQWWNnPAgTLSHuUvXKgit5uLf42JK2o2yU0+jR1D1DSqFM
yXhZDBsr0Pdb6U40clIQZggn6365NgrztSRA2hSjshdUACtyoj2Eh6MdECbDtV8C
4II7IE0uVOiMwy6mCoZg4xNMDtvF4XPnmwXxdOtFSumaBsI02w6KZeN/ATn3Hzr6
N/zx0VDNBejiwlkk6rOMsj38BuW9ntqshCer9S3EJ4q+97Pf+HVbiICzx87ns+cz
1p/cMzQOBevbXsaFfbecoJhjwucBP5diYmznhlngg39kQKDcke5L7q4INplneDJA
cUcJn5Iu4tm4juWtNBGsXIwqy6tcf10o1CqDTA3I052WVyUUUwtGF+oOtIe0vDtZ
Ue6ekDd29DOrMwoGCql0Tp0ZDY+ky6MDnJwVEyhzNF21AaHkS5P60SkFiBofmZp0
CsGixThiYGjOpakK3rlkCPAdq6N/LeL/+X4VUvA1FPJjcboidYZJd0jhrsw/t5um
OPXrzaGQNYZRZP36Eco3GthAOQz8ZJhQlYRVEK3IcaIIxiswu4NBQ3YyzmvDKh+r
tk0h+86IjGn+xnCRfeSsjkB6iAFprLfKKdJ/YvZt5VR96wmKRHVTj5YWgJPeXgxq
2TrkLjpd7m65LYFzGkVSF8yh274/rIyH4GDpbHz7LFUYdc8RVIXs+fV36gCAZm09
2Vq1FIXWzJNgqNT6b0okqlqGSB85D2ryAcb5lGoh+KTW4UKtP0S7RW0OgN5ksVlY
zQQlhDpW8N8vyflu05E08Wtx6WA77+KK9JO5Em3JlrXVjSFndvQlNjs/P0SeNt0s
PQo2QOKuGyMk2xnGSx2gsUKqc0zQIfG6RngzS4gSbOAiInVOnYMJq+lT5SvcUfIT
aQWRSHlVBBqQ6DaixOl7b/w/b9GJamMZqXTVAfpb3RnAHqjKGulpSoBRFgdgEd+L
uvWrFYBRVrTjTYqaGmeW1hqM9IVK5UWeL95Tb1nDY0nZqiTLLbAdPc5XguBwAHms
BoSTMVBbBDLUDWx6aFgw8Bu9RAECH9Hny2B+j35tnzQLpP0AFnbmKw2RozezRqDi
FBVajI/k0noGGLrNnG8POWFJpzuRmpsRhHGI/2Ul9Ym2f1nnLq9pBguoQo8pn3pp
DxS/uKlPDVZR1KLFQMFbutQ0+JnxHZeVE3W3SFpQ7EQ6enDXpcqnUfrh8wPusono
W8JgL0nHkBNTq7sBIWIzJBKzGKZJYFaw0fT57GJ4fVhCz6f49HnJBba9LBx33rDz
YsHwhMpiiEq3MNc5rvs3HxT+chxt8aqq+IhIjh1dNk6uclN44N6gjY7ASPjjOChI
UDk4gfox7AFQuHczphv2LDybyoRYSP166pGfnz3urBa3ffnpy93Tq62UQIrDKd2k
2XXf/nZFQZJKQNLS4dxP+2Zfpe/qeWiM6+I1qrXJtftMs32octMaKqja0ZlwJLks
ppFSJxDDPBJHNwUu7LHHmKZgQ9B6KXtlvX4CponxeORD1ribto06FAupbVEAhpyO
xs17OjwM+kRHnUugyuPWzy2QhLTZRlj9pMBT7g7l2M5eVbWmmR6pB2tXL7Bjuf7w
w9mq0lK9oCYpdXySWVVBzDGHbc2Qa+uqgQWWamXVxPIX9RejqiR4oaCGpwI/oiUT
beJMaJCADo1dLqXHoXgrgox/o7J2tucdbPO/v2SY3OwgELr7QtMNHlPHxruGDTx1
UBs1mvlAY7bPuHTf0MGNqXLxbaSm/jOf0LumpTHHIxeYkh/Z96YEu7sid+euf0Ue
Q2XmHu/V1p5ar7ujKXxnZ9w/OWHo65JekE/8m8jpt+rdV/fm3o+NlzphhdWjCvkb
wrdINXUaWVgsfbp8nqDpCrRsvNfvM1ZxWcADBU7MV8276UuSnC1g2fqrLGqlrt2s
Cshg5CkN3eHGjmKKH47B4lz3qEQr3384eg+N5/ONGWCH9LG3idj2EeiNIWSEWr1a
zXpQCYFu7i2KOmMZxm9gIjGRc8I7efhB73cVSgehNfrhPpmRFtRoSaVUfzVp/CAO
QFeiReqtXKp9SQgq5v1TMUP0S4hhsENktaaDQeifmlO8jxuaPWIn3OQxMsubmujI
BWSRCYyyoSNzqhVrBA82aw0t9fye2MbnRcO+YkAElgIUgTe/heg5D1GqF6nj3Kld
BGFSqhFgmkUgbUXyDWMdXCn55abU/MNwM/YMfcYcYgOIC+G/DyIs+SPoAbExWMTU
UpIP096cPnfEffUv1f7nGA8I/igVp4bgKJW1QcdhzShabDIvaf+2Pt2jB/6QNg+Q
14DY7svGtrn9c0y3F8RUIAAO5ZYoq5PkepqhbsUg5UCrVnKziHkCdxhlj7Sob+ZE
uSyqCd3Nc++uC7eDc0FMH0dLSC3D/fm4KOopeGek6boxCEIlcvhbPjaPj5WwtvFB
aIPzw4qlGHaeQ2NXIaCNrqpf8A1y80RJV7J2Fra8xZ/ySXlL3KoF9BZ0pHkbrOam
+rH5sZSKyS84D9yBysHu7oIBaFnl3PdonQMkb9nsE/r60RxzICUtGeZaM9hp0HaG
n4bLUVw6PBRm0YZKCIpg9XHpd3BPunQ4Ric/NN70IFQJO+EaFvTIv7eJt5kuS429
3IdRiu4fBm7b9TQqGo89ydhT8a2jPx9RHOeSVUPPcjrcXeQIq8J5Wkdwsl8wt2Nv
IXFsAyVXrqshOUmJNDspDdokVNCjclYjDI5IE2nZQm4gQREdIkDp12LKqgUb1zPS
piAUp9Tjbz7mRwt1zIZGkgDKzjtx4Rt7I7nDDpF31K7JFkWV5jVHwdKnVj9G8k9k
JE97O7I7Qk8pUL/fuNkQFxeKqj0Jc0fGYWze9CB6CwEa9nDeXo38XLaptWfziqnz
ObbHbZfAJmjoGuJ/7IOQU6fRDMpgItdnf+GG4NZ0OzL0e3OuIsOwprkvqiDInsV4
/MQtdBJzgDrNgJ4Lgh4IQ1X7kCAINpVtxoEQ1ByJPSrDHIMG4PiJXHrg2H700LQw
fCIMQMEHq9OoqItH5HKXzOClONoFJCnx/hxnDkGMfipPWHsMP/yVF8gWFNhS4Gp7
ZNa+W5q7FLsit5kdMlxRIbNpEcB9VN+jN1lu6x7YD7u4lwO5lfPhu8Nw1LxYtN0L
D1acQ1+fn/yE351QQiisw59D5e0STP5RLPkk66INH32+TUAnCu+fk8/RcT8ZXArT
3oeoxW75M+J96yGDm922iK2dz5kEwbSqemFqDFfSR2H5U3spaTDNPjtVHQyhqGV5
3fp5zlUjvvBtdg8Q8lKfkTqEpYAWPlMG/1iMRiW9cO73qJ/FAybYUopVTZ3hkQwu
P6lSaUNr02aa7jbtOlkXeob2cHU8CAuoXOaPEHIJumFjZkGlX68gA1FzlFuUR7hP
NOVQguJ8BtTCIWTTHD+jynl3hcnujLrNspXjoe5Wr57OWvp7k5Vc1ZnLOB7zoD+p
yiwsvB685EcXEgkMVa6KrlOxkd+1K5hVqlJzTV6gp3q0p+CELB0zHgkPwHVGp9F2
ojZViB1ZVnTHL3kQCsZscTQHcHV3eRqPLmVmHKFwfbYigBzhYFsjmR6lOxeaawMi
aTE1/i8C3PvwNGfDmrNSCMsqcTA86ALx3mWFd53Xd6p4PIRC5THRtzjp3mAvHAiX
RrNY2yLtdX54k/QXjAnYem07WPIBnD9SsuNT0i9svu67hu+VS2tfUJoe+m+/AJ+V
AhEmh8H2m2O86mD86wUKRkodvcsQlmQa9loBg2BblhU4XolTs5LLVjGAj7kANHYC
yg/5Igw5bVELmqwWc287GwkodtZpWhXZ0XM0Q7QFuRmUvA3RzL2TmYuANXr+DGO+
pAT7xa5nbsTKnw10mQXmWjYdCu3nD51Xf5zYfGLGg5Y6U/iqyrKZgTBQ+B/5zpt2
ADz83upn1u17OKu/13H8M6VjDdT26KEMZg/co5ixEjiN/rCxnCtI1fAeK3Xi/OlN
3yM+YohLE+yQvNewPPBVSBXA32QsS6rMTcKQRIfXABA/tXtNPZlL6L74WIREyssx
qQMBMQbEo7FhZizCY5J6LjnRrJyKelHvpth+vG5sowbAL/Ce9Buf2Edpo3ZzHQiP
I7Xc/zMdhNB8mHkrQNehfHZWI7BDfGiq7ySQ90rmv5MpP6JD7XscM8bg+10AwaiP
FJH3iCOTOG7BaOQ9fgv2hP4GN1qCcshhxkdhTjeP8bS2KH9fbYNdpQPve47XMSxn
xIAoBOsiLm/Ocn6hIp+m5EpiCD2tAyj5U1vdhVld1V+fWF6CuCWXQsM9ePb3b/qB
Re+aYiFe9X98egXEfREJrT6jc41CiorJQVQZY8qBImXlqk0hqk1mbEhsEPrGi2va
nPES/3SeloiK5mlo+CIf4GR3mZPL7YWWTD5zg9MpEUzW5TQLo3t2xUfGArA803ak
Ar8qr9K/fKPPjM4gc3/1Roeb4FhdWy6/ZklmDGj8FRGC7Nxxgd8k+51MK01ST3PQ
Ceqsag+syfCI7DntiwQLUbKSUgDvg50bf2EBm0CX594ZpBjEYVa11myfqOzHPQO1
t585f180vrG9IRrDZ3icYgbLzwKliZp3G9/I32qvUj5v2tkstH0HEcjdGhGueBTF
cXpklAKP/Hsto1WZZiYFTuXMuXhh8xVoJd8mdTpSC0WrIB2VJ3cACa80tcX3sK0E
EIvqOh1Lx9zxhnS29PSXrpnLXgZjgBblYprl30pHoATDazjHqk7B12ldffQUb+Cn
XB4IQJdhORUolGEpg7epUOrD2PUUm269bZelhWmY1D+abmT4RCSYdOX9bNy5rFxl
z4Z4dAhuU5hlkILmqV2eDrMJOmOyK7HI6vipvFrBTIi5/wgYQfzG8Wg/oge5uxNZ
gmFR7K+CkvaHfJm6MFdVtNNXJq50xW1xNdHfxRQUzCpq7PtYxwNx+FclO09dlCYy
ZLkXXGyKkLsGLrVw4lApJLBogIfoz80N4EWlAhQl1nxcMk/cib+cgvKS40JnKZif
tnDppvmdgaBgztIVfe10Ny8Qm7BX44HK/UFSTf9QbSAEgjhv0df3+G4SzEvN7Gbi
Q3H/hDrb6SBgfSK8pEyWRuhapiuev72OBwk0NjbxkfvGuvzVtF9EbQ/aAU5v0nDA
taw40J+NGR33aNR2RAdk2Vxujrft0IAVfou364D4DGJ6+mdz5fnyDQ6y9p6cxi0D
2GaXmrlE07sjpnfHIP9NG8UDnuRL0JEN0ILZLRBF4hvLSk66YCnxrHDK9z5HNolc
8pC2c/F0IUDZ1EcUQY1dw95foTLrkggQTvV4eSFLHE8QFR5K8tevbN1cA6jc+nMq
ic/wnawdOSjA1k4FqqxsX1ywEP8NZ+CiIXHfnLkT92gO/+NQK1LfyvRpk7dh9lzN
bWWFZ8C4jl8cTYOa7bGJcYVcP7CZPrliTXAzmLBYbOJE+O8KFc86WxYwyOnJ66kA
uDAOwiwFemqrUCmf1rBMxVh15BcddF39/LoDdzqIhmQeadnt6Y8sLhfTgobcmg6L
i3zhdH3W+MEiRH1o9FZUvdQZop5EqMMn1ZNUhffNDseSjETRNdylVjjB9ZhhXExw
Tgw5w+ElX4AG0mut6oN4iMFeUd2orO4rD6+DeZHFhdOod2A4BlI7fOFQoqUZaHIV
cQKZ72qu8Jn+PJpq+P15a34fhoEu227hcvfO10ilr+2XAOBkDOSgCMFe1GjM9q5e
n7D1OFF6GEyTjCsdlyAA/z6uUJNMHwna9V58NAcsdhqctJhsWWC+di/ifUi8PrP5
3+DLo7eefP0c3xeGITB4XZp/3CN5lgIbbjtP/cDayx4Yi6jOXTs1a0RIYhoO8xpQ
HiqGox7xARWL3O9FuhuO+bLjdLRmqyE6liVPOImG9SRuWUw3nJ0WLzhvg6KkUrdA
k18Nksv64mByvvhdmLBnAJrpD2TKX1mZmFZ5tqKV+tFTM8AKdTdZVS5STuKMy/j/
IFt7lTFQ/IJRd3w4rJ2+2kSfg28NTVRbR8yFmcGYV3VdYBEgleCz7RDB0HxrDCnw
HSCEXQFHGFkiLVGDeEYMY+VmLuAZWHS4vTdsjHG0EgZNWbPg08LysZJis7Q7oawp
4zbjI6q7JrIHppF8FL2hbne4qgN7ijDCn+xAZqxETG/aFlUyHDufhH8JUPTtlSfx
32tT0/NYIkYRIRPwndlGCgV12Nbsg+gmscdAssM231OHvUhTxNKksg5Bijs7cxtW
LhzqsPVzDXcsu3VsfIu9MSWc+rEgHzmfflTOcl8bkgN7k2sY5eTgwLnn1kTD43OR
aQHaSRBOfzNFpY52n0VviJHm64I3rr1OuFkoeMqq2H2ckM7OAF2JvjiEyx3xqA4s
sZzNlZxbTQmlIG4RfsVN3e+9cLwak58tWyxDP1k44WjczbwgawXbYu/H/4s+qA9L
Jqi9nWC8OpxZA3tqBPL2bOjsRpjSX7b0U5ijtYHzSrH4Kht7MIfBXBTZTAlLdXoc
YOHrBqOGl3lE3LGWOFC3Nd/n+obWQcL89WYv59/kcJyieV3iyFI76ef4oJ6hh20h
cj65QOO63yrAxark6A1CUq8mrHGvEiTMeBPw854go/RbPXXflB1jJGxTWMs21bzc
o9HHkjQ7+CXfqoYdWuxeLdvIZQTWAg8z4ia2+fILTvr8j4whaNBawJz6VYdm/fy/
flol0/ZTCvAQirtZ4cQyl15MQv/1fu+cOuGGUYha8eM5olu6vLf5YuLEDadrZKXs
/C6ugL2ii49MpxA98s7dKOE5/tbdqVmK8QP3ZSYF/0b3jlD/dL57gFZEgwdHJuq3
ypgQYVOWQ8efnRQnXDFs1q1fxpE20pMNXtG9t9DW7MF2lrgDz0Iaya1dGZ699W8z
JmCtvpkkRoynaa28Y1IsvhQ/RmzbzQ01MRY28Yd/1f/BDwDXm1CiXeLJn2unxl8K
z1B6N4HVVswBT52N4mBS2rgffTtV1WDYsb2ij+ZZLCaRy9ObQSnaguVhAMs4YEU4
IHZIxf0osHUObutS6A+78i6eEPCjt4tMmhp4Osg+4EKpShAejzZxLp1Zdz74BkHS
8n9yaDhL6SCIy81g1PH7tLMRA6GA/Xf99Ugwqo6+6zlkA9gY0ISquLHOHLI+Pvju
Uu5efbU6YI93MiRMyHW5dAzdDw0W6Iawf38I06e/8WetO2WLMPGfxRl8hYtPJfVi
bWM/IS21wYKi5MOSQess1FadMPixBFutmlQvyo5ZB7J1Q8ovMkN4ziqO2PIWwTRN
tPtHQkfeovS+ZcbBIhsjpbwDFLGuQPOdL+HAZxJFPcm+I5LM6OU8gdhRxgaWEbU0
VfEbXfq+npg7zqHfWJVNRyQ9Hkr9rlK2mCjbXfqCSIsvVraDq4yQ5Q9Ivixk7Iv3
nGvBVbess7dCipFXgXE49Twe6jkL9+o7R2bRmQCD46XewTHVQbe0feqeH6JZ6Qaj
a66YnYMzYKYfa05zNGwMckupOdOXG30pV9FjDo17Zmw67m6DiM+jmFAABdJZHKf+
0RMux4Mhp3eViy+4Qd9N9SIslY5COa0Sgcst4mD0ovWySSpYlb+vWAdvtEqU9vZE
ZyR7f7z9LPRwGEM4fHLZLFinbW1s8926VnU/ervdTeYLjbLt0Y3J5swS6bLu408q
tylo8U4g/y5UX3l3/MIf8kUZaEl8zKKlm6+nSAAmra3790dlCRpHXdxC8yHiC9Wa
NTPkzx2is3Hv9++ZzM2Q1P1E4HuuyU593KNIb1zanqSx9f3+EaaObpwsQlvP2RYF
iKIerCHG31OZ4CAc+PNw/e+Y7+u6j6BmlI2VD9KSFBa37CB/Uf+AuQxm156+ufFA
PPVXJE3UDU96gaGfZwmTVHlXPzjqYIZHQWfhrkhMXH79n56scCVK0roe4q7igeJm
ysxsQH5uBTTW+CGkEi08dzi9zc1L9P/U5kqWLAunD9cxYmP6V/o/ItL4//ywma8Y
dIeae6V6jBDl3Py+Ih26EcvbsmTgB/4vu615XjYvL9PPXbgRkuYGTYkYu+FqLt2t
Bm31qgC9EZO4oYXTvCPFkoxUBbRUGTU1nwmic7lK2R27GXUt3Tg92Mu4Q/0Sh/Em
0SaS+CRP7TP0pducBZDpr2R0JxKM8mRQZeYIhWxs2f8mgqKL6TNVqy4M66se5jns
lZRc3pUJUzdVtC+byKZosLCAVcmidnyoihzLh2YAKJeda958MZHT+J4/86hXAmV/
G2W88Am1bz3ctvgOtVzashB0crJyLlYObhKI1liHruDAhtATDptcVENQzsO6nNw0
rLgaFp21xx7a5jmhvlaDMXYO5vP3zOmZMtNSME8Pg/VrUvwxXXBtAbhr2nWT/B2T
BvMl4JD251KCIwkkFbb1kOTfiyMZhUpEbI04Hy42BELyEgHPcUz91COLeaItekrU
V2oOIS8w8NOODoZfzNTEQ5qjhVpAqdVt7m2pQ68q7ltddIrOIR11BhPs4Hp0KQN2
6Vdgz4um4sFh4rwq7R4PmqXhXBhFbu2xqvvxtm3p519TQVeWmc2aztKegVCdqDr0
m8aH+K2g3gWSdmO8ipTSDmZoJo0F6Y40pSV9UHRi3ZjGQRg7e0U63QOV++J8cWye
VZ++9K3X4RYf7fKCSyCpJV6fEr10tSsNpoLhGKgYhP1l1xpwa6MLHunIxKPOR5zj
yHGicJUL31QkzS2gfkI5G0lhoJLupqmbmUMpV9D17761x78QDYctc1eb2LeaHDf0
DGqUPytbeo5zrbvXtYaezUsHHhmoFAR4owvCgLFDhucFohZz1nIDdtMPxbeLc61K
ko43FE4Ur7MIcgJiz226FM9iNGEcJV8cdYif4g5+on4ER2twT9vfXY5i2w/svptG
DRgyVb96uVXxaZvPD8Uv8CauV1poON1IssR1ssr7RPzTtvfyRwbUUKcLEvLbw0WR
6Dn6/KpZJPcU4elHQ6Nb0IsthvQ+1R+vszE3i5TxVQtUQiHcGMiDLjVsDkv8uNwt
pGdh+yNWupZg96MI2x1Jpsi3Ulk+BWDu+M4ZXTOElp0DHooDOK5j4jvE1edkY+k7
g+oTatzZMBrlLqShKoG7vWbGnmsSHeSD+eEJpz3FBg3RvRsEl1reHrpTZm0MA1Rg
8UoT08AcZdBEOIZ3mihjDwLgfjZlQ3OMvH7OLVZT79aZxJIcj6NQT7T2897g/xqo
mAZ09xP6BhdgoLOEWjmZTvwUEGpd2bQFfZDUqsYS6VgObDrVqpqaKFOAJ+ac8n94
0Z6RGqQ4Ld4Mix92nKZhZkd5j1uALrhrBcT1oVEPG0OcYukghRyY2A7EZ5FtXXTt
4/2f86D7fMh4jDP5klCabYAGeHmcgtwhtSgvxoKKKa81h5Wi9w1RPARPRWzcL9AV
YeQ1TOiGvB085jBZ9bKTsgQhlTJcFM4+RGKDvjFBulZd6qiC6iZ4JfFB6ODwoOZN
UPD4P5KJvf/q5YJJuecsUrQ9D4vsosh38R/eqqc+2drBVPdEIPTXYsOMJuhcXAw/
eZiGNnWI7w3a0lkpd+tzTJK7RQeq+5PKhr0UnDIHlke5mN2YPmhjeen1NRvFYmAc
vCd1gHThn5z1ifv3Ls9euV3nV3qTx06mnoo5q11HuKbHk50hbUrvlT4bCXpulhCD
INMTJeRrp2uzJ5BoDDvDeMa2Z08YmFULX7Aa4zG8QZETfvJxMaCB2G1DtFuk0agq
LzNZBUVKvMWEtddsIuOS50smadclj6tWV1BViZKswjrm+amNV5bQO+RsQ5ybIAq7
IRE0dDZg4hBfxjIR/0Sz3mEcs6Fw77Xo7v3oqWOKaGg1sh0mNwRj8Bw4Rqt0aRW9
OPBSHvx/i6wjJzekw9sRDWai5Tbmj8DYrrMR1Qae97a0sbeLR0QDhRUetEE/iwH1
JUVHajlrmmnyaDb4ZyXCVVgOB3WOXSAaGM4GYKAF4COy1vAtIP4ZHBjYpIe7BqIz
ElHpYjZMCp/iUbNVgWRshnCdL/K6pVVF9tGYBWe9HWGzsy5NITS/nwbmCpakZUlM
XiQyWLb8L7gSgmUqRIPUaxl4Pt3FSfSRRYRWXDUexOlz0xcXYN8NJLEzC+yYEOzy
3hQHVr23VIZM5/9oDqWcGSqOgI8egSRCzhwcRlBiCRLkRoL5NPVCoQMPB/nSwc+B
nymGB7lJuD5fn1Dqk2Lp1mwqAxP3SYW2U4M+rk+Tridc7y5v6DlO2UBxx8VAYee9
oYa9bWHlvo+kjIGhbTpPq01EmW+vpeLjxSkCXVFG6wFGuornoi7zoRrJN6EsNimb
oRh3C+tMBQn5xrLnTap8XseP9pcb3P84NRMTImB2dANfoCOxsmHEbQ2ochOVoQL5
aQnyIPcMUKXoXWxtamuofF9pkft0yADKDZ/g2NbpwRp1llAN+5MtJmthyXLkD9VI
YkAoqGEE/KHrzClTCM3pxlZFFU4NUl+11y9jJX7TC1wl+4ZpKuz5NCI2rHeLw/0n
LhJAxuNfptAvOPQvTvEcUzQPZyBag5sLb40EU3Xa04Nl8DKsKERjWUnTqrXtU/50
C4TTxiK8Dk4eECz4mHPRB+kqH4JxULV/xKmSMo+WAzypp3WegM2z6UKHdrhIE3LI
ISDN08QeBXts4ZYckVFOBB1pLMG4Yr54W18gFAqFCPQfFMoElWnXcjVf1aYpqzeV
vCaj0wwQVmUNFUs+hA6Ipe4TmlH3d44/TsWs6AtUD8COJKnVzPIp43Xwg4NGqHdJ
xJlOWdOaz/eUeDIV/ZfxZPpUcZuREN3dnsrUXpanvhyWVLP6iga6301nPeq3oRBs
8X5EZzzadPQmUrjRSLKQfbFUUKSG4Bdjo3QTF/kwqOqLtnMzvCEvqz/HP21onVVV
HfDFCUGI/IKAEsMto+7k3nyKN6wPIMC9lMut4vxmqdk9Yhq6eR6SWzWDBr3H7G4Q
yWcyVKgsIUxR/Up+7V6EhsriJYiVmwwsmxPGvQGZ1uxykdnM2lCLA/ir0r9j6p5w
veTgVBPGmSqfZZ7OVNlkwH/nX8DrCRwDImNZARkoQSQHX5XhA1ivj4zxNq2ope/z
48xGb5aeY9L5ErW7cJMOu/KmthJAeb907azBVN49/ybdNLCUBLZhM283YJIL+1sF
oa6TpCou2FyAZtE//znO/l2VAqrhLZFQp0WRVF9b/HxCeWiKc1cWICjCHWm2/yZx
5nhQb4csDdW6MDNyxI/1r2uHrvfdXhZdqGB3xYOZSH+u0Pcb4ReU99654J3Ozu9U
ramVjcnwbyiVIg1V15pFZioIVoMPnJgg5etvSFlh1gDcrs4ZCQkXLvvcHG8VGZW/
85RWuwN0zHP6EiuWXK8EzcGnQfJ8K29KpBmY69TKiNWwCkgar1PSllWUrIeR3I47
Iu5AT/VWENf2UUnetku9TlZNYJe/3XKtgLwuARaAvFjSey6beHPoSXl7SOS0wGDE
2woxANlZ5MJV+NAbdG1HzcuQjcbRtklwWXfIXIM8Xd5Qd7Q1IaVO4hMpjXBNwogD
s5+5sTY23yysFpTlgXWNtjJn8ttIRpGfmHkK+GlfgDv9zjhrxiiegURvx+RIakSI
V/BNNViUM6Ha4gEU9BQsPm/nrEztTL49Hm97YxTcAh54+IPIVr1AVDxbSwfZH0cK
1OtCwc/KAU8NVSic08UhGU5dtuCfOlVOuw8JU8o5wRUcZWVRvPNb49K7BzwZCdYX
qpPX/WoLrVhTinOxCGjrxUYE5MGy/Zrsf0zW9BxivXXZK66cZ2lmOCJZWJ4r/hpa
4gd6jDXncUqkf9xeI4Ljmki1jagck9XGRpWRXYhRmjJ3as4ecPCf/cUvS+cjRXUC
MVgb3fL/fUesIWCdb/7m8oPX/EawJvhNuCiJj/BbNMklW4CmszjnLBo0XKTPvKN6
Hh18/w9RFGiaOwKoX5Xce28ADACwEJvnw8UonEMvYx0D6jJ1ymxsZw93VWvkTNkx
5UMl8rs/jpsKFdbyzSiSOBRaQ3O+TKH2SoyQJirbLIDqdB55WUSrIvWL/JHhjEhc
guE9KnHbfxKIfGJn3B1Yl+ef8Ceal8pchB7xMJg0N+rj8brJqYHJg7H6FNsBz0yB
SaasFN9HxZOUJA+OmAdX3Mvajyj/8o8yBuQ9o3b8wch5y9KAmXs62cergH5hMorB
t2F40dRgvM6IyGBizwYPyA8uuerr9d87dN/8+WZ5jUaU4DTcW2zk4SCifFxdKNmn
HM/02Ok5sf6Jvlg8vIJO4kN0kpY7XQMXATbFXz9WPcBsDDJ+a7tCpn8MKJDp/dlT
gVDwP0diNbmwfmGXwKy2MtFQBPrThn0QYVEtIk8X8BE3pTNKjvO37KVL1QEKNdH6
CB4BoyK9Ps+rzKDqT0N4Rib+eJ9FeYmli30PUp1A3Jm1ZFUS/P2cRIFybVMbLUoT
yT1dspGmpxDyoI8JHmNGWfJWG4CcE/kLZxwMh5dSSXeHnxDZB6L035jMJc/mXWGJ
/dxX7mJRyzr96PSP7Zgiex445PIWWBOFrj6Cwa4TTzGP27n7anMn+W42g0gaeDRp
rkW3iMePx6QJtIFwrJGk7GJfO/VnTluu10F2FkDS3Nh+YCIilSWpG0i0NNfb+SPn
H5MrYHuMG1Uug47foP9C+GhrcBN69njcBfvNCAaCRLTnWAAn9h4mfllgg482dip7
CDyaSwH/vLuCxSjpCZ9yNy39kfgFvjrGvAecUHizTEIUyU8mweYbzfVjJIAggR7M
l4CBqYyWYvkPrjpgUWKY2h6BIaxQAZ/Qw31BqURgPoq9OSTHE10h8iBMGtWW5S0i
w7HTT8fIBQlrw9gNZMvoC18IhCB+7+bmoB+KNFDPuTxL/P804hMvUo3p1PHwP6Rw
W2Xhy40+rdu7QCO83BjBIQF/KXpDt0tW34x7Ir+eJ3lyNSQyZH/nWnNalAKe1yj1
nhS3U6uGHGb9v9BW/Npl9yEQ2XlDNKhppBhWpz2dl5cQdiNy085xywpup211drn+
DsDbCTRTC6ED3Y0s7wzX318OFS1y1UOnTVe3dWL3dBSR5zTJ2BKp+xbq3KATgA+f
bQbr4YrAjg+rPOgMddK88G9rqNvqXRWo96U6GaFkIEGqZpr32RR+VjWRomaKR898
xwgIEAeRIDtTFDunagxf0Ph7kzNY8dY/UsQ9fnlsSyk2+1M0LY1Y5VsGotclsA9j
PsaUhhXBSKOMbU0MfDTaDRkjHwBH1VmjaqJym+DX/CYDMbOoBTtHvaLuxbPe1ScR
wGBE2hlZC7psloPO7C26quatHG3+QPMXZklSSzwe5VWpCvtuaPRu3aHjOYNqm09l
zkcSBwh/9ktj+P5JCROTgGU9c/1BQbEmCljj8vKIrVPvYXMU+tGfMvw1RKU1Yjy9
lQD9GG65Gfy6kBvOhLZOJl/i/WoUIkZQgUmo4BpurYf/IlZh5y/XdpK5VDEuGDiC
0z0OEQJbanwTwrbpYbIV7SMNDLAFrN8GzCvGsGwe2GfTlZHQtbBwUJU4tpT3jv2b
Z6seGkaEIc0RK79PGGblcd2c2UGxiUS0EJjLfBQDN9s5pPMDQm13A0F/kKutNinR
9WDP1Kq9WDC4gGvfEkPl6QeFgY0rb6I+lGikEyUj+w7ryiyTFL0Pjevn4ekjmyWC
YZ4yJGCMvv7Ncs/A8HAM8nidwgrCb+H3CO2gYY6606cjznTpSBUjyaNbw0EvlOCp
V6b0tT9GhsTcRYgXTuGYJfkiUVQaCOI68PbccTt5//QCYdXwjLH5VmAC3GFur18F
alyV/OPH/bX5HQv5rIskb8BEW/FFbRMKc/hmyjDOV8c3n6L/Bzxxa43SZuCxkiUm
J0hSrh6keCMyjhHyJV9ZUGbkI7wtCxaChkx1FTrL0FMcWN7ZTtvdMVH40lGWg49a
7D6IS/bLwmUF6dxbejmHHMCBWIE08hSEEcGUNf4bHJYqQLRNHdhRXph392BNeh4d
bOZCM2hSGS6+whA8SUPOXJacKHBmGKIS0IBqis5/7AwDWM3nXpVUChaB8O3mAJFZ
oRqCkyHm/UqVfdnwWZIBHQmJGmabVq0nWaIX1slf1YtAgRjvWeaX+XghAKrxx23h
4PC2Q8SAiAOTzE8RiNY7K/0EfayTgRrpWozYTrJQZI3r8rXdca80InGSM8ySJBXR
qw8kKcCB4njtI1vJp4KnXoRFxyNiqgm1my5Sc9OvI3V/r0zCyvw/sSRNqPOziv1+
akwVy2QyWrrQ0CutDHWb5m1x5MD/xkoGJgwO08JBmYz5oqFRQ2866g8Wg/rSIMA1
ncI2tv1VkaSLsdhBWVSIREX0dpmhggmd3KXjV/BEuaF7paZXKXupVYbmj3Y+OJtT
7LZzPn0etM6e3xNMNIzD4iThce//ybYR2X7ORBwCSxcqGSmAg7s7eYgSILY//lAQ
hvJO27of+Ym+LVGUnuKKVcZV40moivWMjY/U5KYU8PlKT2JUuwDSzrX5twSGtEpC
f6ErM6igW7XCUAcREPx0/2hXqYgTONsmCHNXmIK69zLw5VGxHCvBNKN05SO5GVyN
EzFGudXTfZ6RsyBomE7D9VvkDpPPxwxPGB4Lnj8FrmfO/V+ziH3uG3HsnuTPT74t
nABMiUqI0zzkVsh6mJUvyyftY0Bt5ftAh8DN3mqyG3beJpC+0xjMqP6fJ3zvZetg
wSmEniE/9YVku47rsepQ2loLV1hnuaoeoqPdCDa6iL17kGcl4ULu/2gLzGE8cId1
ws1vlnzO1E0a5VECF4jJ0tZgpuRynScmARSdmuZAaGmahlU8oHrhmiN6q4kiyAOZ
nGJxeWZe1MpV6G0uHMymNeHnaO8KSExOol+Jcitd5gaR9ohvhWUeDClzmL9dMNFD
s/6Mp4Idb7YrUY9cg97Pliu8iRpiGEzb6KIQ9/3ozch2TW5CWK7bqNatJHbh/a8n
xbxvNlnnyzAkudNWpWYibmEcpjrJcfhnzTBL6lxC6+77sEORc60KrLpSR28yLx53
tep8nHQkxrkEUlPvdmdZ75UfLVjWcJQWiDRwjJQ2uc6LJhtO0a+mLeGT67pR7oi3
77uXbraY5o6cBBOZwAJRqpWQleMdM8C4tev7CTNCtU5aRx3lCsdD+sPPv0cGlx8i
c6iT1ssXOe1Xfpx1EG5n8CHm+SGs4nLd/GMNk6WhPXOTgM4PcKD1FU+ilsrtLrJZ
SUzXnaLLX+X2sJ9KnRURaxZxirPbEXg5RJOQ4x3aPZrXYgOwidk4PVsWwiCacJbN
qKXQzBl8V7uUHltaaQIS4TKr6JTkuc+FxLT6ItM2j5pVq3lvp61NsIpfXCp2ksJO
eyo9ZvGDDCMAJ/DYKAe9/kkEFYyPTB7WhGrzJMW3RmP0zW6tMSZj0sQzToZLs0jd
VtuxM2VOKT4nlA588yyMJyh7ImwaoFyzlm0oslKUgJEg4bKhAgtkvYPVfg0vv4UU
HpOC7dZdDJgy/E4UhzYwANMC66pJlfMOcS4XDhw7a2Uuw4Gu6EcAC1gHQtmhMGq2
IgorGtd1JkZHzwggHi8IYwP5oc3IGcDwLbNyJ8EleZY9b2EAhXL4X2KuJg4UoZ50
Q7FJZhvKzU56o671e5Q7ESuquln8XnMxhE0vpbxOs0+gtLTCpj5wAoGEFCtp2z7k
+mhf7ITW/B1I3OhOnVP0L/vc9MGYtjob78D+5tKDBGdUWFzHEdg5fix1C+sgmOEF
NDvW28reIkNDlsXR+zDp59Oop8PCSk0b9pwUW7WQoJORSaE4dR7JPaV8hnxIllQ0
pHOk8MbYbqIZObOIOamX2YVspNg+0BzAhRDjdsouvfn/NNLsUTz/WyZijJzysv7H
rxVTN/cJFpCNEXEDZB3msNiPruesrJc1ycngdU86Gp+p8LrrIJmt/JfKZwh9mrZi
7tg7iJEa11BapwZfLDqKewXBgmYJu7cJ+lkuCBgn0TzFWcPvwfyDIHJd7IH95Vtk
cQQ1Lda6ZIf3rdSYt5782764/s5XZeSIvMErFiVN1d0BwIDpH7nO6JK4IhUErsY5
31VbzmJpUXWdd1xiabZYxJn25f7uK9mHaJ+2USfOQO7oqPz1zrkKuOBbmFCWmbya
UnXCbOgJ0PzUB44m79XvtkiUPnl21f9wsR0jb525+V1CuDM+CW+M6dD1d+3v4ek4
nF5/6WLXyu368Oaj7yGAiQcn4THiid3VdIl7mI/nbZrQHg5J/zNfRRar16XzXC3o
ZKHvWxgi9ZuJUoWl413OhlhXTzdX/HzaHMh56HuobgBVvcX8GQbfdR+kea++3iCR
S91LrikMb6WZ/738a5gJE5cpnTXiVQjul/qYEE8JARIzKsWssRIJ5qVf4gR8il31
5a4QXBglBX+FCLBy8Oz/3EkT5ncZd5CXj63g6Ni4u4HaAb62wZFOenEi47dp7r1a
0obA+jcsaxSqx3tQKF47s+bF6gKND4G6maY+1kJRUK6Wk945JhpLWO1x1uNx/swK
GkHLhBEDVEhoaOcIoXDS5Bvfkxjm6PN/9ly4l7GkfzbNbO/BGbc8flnn4wj0T82R
qGSNjJ+4A8nzJ6ALHeSm/Ok0KJosr0w5JSI57bmyihPG2fqhc+EtqTTOuDDe0mxR
Qi3jlhvSxjcpNpZ9W8w8BywBY6BS5Pshi9ZrUxN+0/HTGz2GqBQnef5oDbxJpKaY
TCc16gvQ+H8YLbBWL9ATgcVsSa7yMK+EScUwhVgCUr9wp9HBpYvJTOLFaziWCLYi
Yz11Ttp3Y/5ZyjpvmjE9tiU2aHTamDRDDdJOuETNXlY96EBBLOUbSRqOnyxxBxvw
zOScYZMlNRzVwxadoqeMqkQlNbbnCzc/aRPaYsdNZXuuv5quHy6aKx4N+HoXQhQs
uEvzgLKyTA9tLQPfO4G5QMGH0VEeb+Y01mRC6oenOwgTb8YHvOSLgk8BKi+8SPAD
IyWszJXUNeH1EHAsE9NvdJYqOlxiRupUGdeeKZyvmxQeHGkKk2H1Vm80VM+eOkDZ
z8BFbR2VmAJRZzfDGIjsvxljdYKuhm9fHnAEvKsYg8C8druuyACtEORuF2SSKoo7
Ho7aXq/GMahN9dSZXwbhMLwuiqshtWdewjGniZvQPltOXTYpgv2gx1MJVqz/Glgq
KeiJfmrlsNh8F450lqKI61i5bQiAdpg70vWYoNnSzgjDyshUjneCqxCN181zxEoA
Lq93+ug3ILXPcnGmuS2pWi3xmXMsM6ti94cyZDVqbL22A4dA8QhxMoJoIFJfGjp8
9++dJeJyt+Y5nvTMnQw2HTvHl4dtslzWMxr/knml5ElzXRoVuCOFvx/fSlLJjT7S
zhK/bZYRRuY1ZLTfeh3zO+CriliipiNaMp+rQ96jQqJuDIWDN5qFikx6OUf4CiSe
bU8L/5F23yc2S2GhIkuw5ORea1EuigU2RaSiwRlGzEKMSkq5t4oWqGd3PbA5UhQk
YmVUOUmGnpHObWxGFBF2xbGWGZ87vHs0TIJ6m1awr6v2xOWTwp9YMZ3PTnYx1Cwg
aMdL2vT4J2PIn+ykXJ7tm7xK8bm7sJd8jsCmmJmj+O7/8//N6KU5LvQhSEEyQhAa
+z9w4GK/l0iXmGDEQx59dQFLPvypOQmdjpE+lYEbkkgqEnHRZx2alOK+hp9tphFS
unFt92xRx45IVNOrvIMF2w9okNFwSJWVZFrsLUDXjSY1t+03QFiGM7CTkyeH/qXZ
m+XhduQHy0BFY8lOrMB1WOI/+vRzkY2GmNIBW59qyyiMJl5zrDS9PHgtfeRJLm1o
z1Id9DYbJkkZLMM+n57oo0G0TmrnkA5KShGd2fFiXKjJTfSya0xGi7g7aDTiwIAa
O8jNPJgpoB97oIjzv1FhVlc4AQ7mf0d1RbEFKUqnz/oMHxIzBYX4bKtt9Cjn/SzJ
HD+n/TNDGFrfvKCDFjVZj2WtnS0nV7adbw9I2MtpNM9CThG8n/DpVZuiKq9DCtqf
gvV0esOrCrukerYS/PIF7N4hHGbM3aMD4/APy3NERfMTh7xhn6gZGu9sVMRvKf9E
a27jVmkPZq0FSd0r+7y2c+xQgUv0WfIu3fkxqbAj3nJ3nIz4/6x8jr/1D2KuGV+V
XU/guAP2vuu0YFqidvSsImR/htPehkBDV/B7ay9Nf9MYOswcSdKkc9MWaYDYaD7N
UMYUnjfj7betIk4f37tWWieH3is91GDu20Q1ys8LEojK0heNI/Zuvy2yYCNqECu1
Rj8YDzAw1Ifrufs0q4uC5QWmxHzngBRRbVZen2bVYrmFnAnCc8NpEpIBUynxuctV
GKyhOXLyd81731CGgEKK0g8bySujMlC2DQVf9HXzjgpS79O1ZTIQEACul8cXQYBM
T0N5VGBnYOg8LXjgt3y7CABVxH4nMAxkGA/KWly+mcOv4lJSn1ooXg4Avj8hte0f
CUwAIjXm5GbG/68oujT5doK8zpJGwosnGbi9JtT2N6IrvTpg2Bc/KtVrao6fXdAJ
TfdsbmBMsmqU/oOJUBwKe+upDclf7lFQcaqDKWoqalD7p0Ki6bVoLdMXoxz81MnH
L/IPRC4YVRAyyfQF147ataetu5sOAFMUQPjz6iENFiQpnWM9V2RKskGqkez9lF74
EpD1JPSPehrN2F3CaJtCj/Tlga26RgmEdxzA+C/nUxsoVfdwRFO8NYYPGUaCIaEC
/OEmQaZJqB77XnMLuGWkt3jMps0HxYvLWkzKSoXaMaRMlgoLfjMS141fYUR2JHt3
6r5mKE7m5nU9kp18JjMcY89QafFixcEHdwk6iFa80P5bjkHl46SIIAnb1bNuVr3N
yQOcWtjca4Z72iGKz/YWN/qcb74wGuAsb6Yb68mdTTbBOJr8g5l4///cjztFoUeU
WtRrUl+G7cMC3USRNilNeP95gKt2Ky0WeVhiM8qk7xzTNePRoGurmG0qwr9hEy3B
TZzoso5Il4m0bI1N9J4LF+e5Tf2yzH4tFSJThgWhO2K84upp8zEwrgWceEQRH2nm
w8LZZbbPg+vncLzQe7CW4jhBGlH88K7ZOvNxqg9/0RKw4+OjA4Dz3r1Wp39m+Dyu
EcLbC/A9xuJUEsgoF85hE1PQSL9FF+Xonge2YCf9GPMC1GgKat2BwNEfcBxOP305
mVVf8b6m1UVIHFF4fTr/jW0MhumJ9fYolqnHqMji4B2aP0g1T0/e8xCXVxIBi0AA
ZgM9AUrcxhkDBvrkvWvLwVtle0hmAbcZ4Vyohk1pQaQUFTG4TJpwDrS8+rPJa5eA
tdnoBizWp61LyBBN3+JX6n+Cb+/hjWWzWdvep9xAenk=
`protect END_PROTECTED
