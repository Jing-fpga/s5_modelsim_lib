`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CE4zlk0M3OfREEQxsiHyXW64hRMFGKAt6EsIU6qdBgO4w0yeoM1URbzK5KkUbnFr
etedlweqi3AGA7358TzsYmDLOBDp2GKtOk9I5l0gj7Xl4JzAsY8dyaY7bCnJvekJ
RIaf8BqdQaa7rOyyDTVk26jY65auUkR5nDa14tOor1v8HdXZFoEbl504n/4B6Qwt
bsXKNmuZJEMGOmPn31O3HL5iF1oFZ14GqJ90VvSDMsistxzy1QjFywWcBNsXO5z3
/guU5gealF7urLXFj3sfQyy5+cgJwLM+pjBczorZtwcg1ZNpqtV1AOw2BD8kmTzd
LA2rNPEa9iLQ29MfU63GCzBIyhD1ETeTcBxfZ79grnFkdgedvy9V10tWxNy9h55R
nNSuriR6Twb0i45DzDRN3mmtVMz2F6NZMGON0XvTowsEsypmLKk5JJET4Xbqucze
9VtDzcgLo1zD9KIcuI9r54ohJYLQbaD95cvSXwF6+XsdP/UdkFy9gsa/5ck7qmE3
4JR3CcS5Z7K0tZFIYvzJBZdr1xT3a0q2t048ScEydgpcaajBazgjsXNgLQAAAHQh
guDSoBqgmND+RUSbsFB5wlgHgwuFgViHJ2aV9ktDl62TL/aN18qrt2umiuE2TbGu
pFWyoFD93MEbH+/8u4xao8zXxfNIuhvzBgsH2v/6RHsoN6BEjtImsfC0wqOz/eR1
3vd1ArIg021bifk666NauVlteeY7lwLC4edXDaklLXJsSaBf+oAaljB8GGo8KtLL
KNYtmFOSsK2SU+UFgOP6vv/rp3FMrJiqzi1swB4ySr636avSeZhbi2+OD3gNpygs
JzJS8QxR+5GwbrEttMdC5s3tu6v/BLb73qhuvSRwiPOOV2IQCrPxgpBvGrEWtT07
T+1nNGK8PcujoOM9h+DKcRUVByOxtTHyyPJgaemXo+MOTfmInpKN10RbyFoBj/Fb
Nm5SLw46eLaSTb9HOcP5FO5B5hYmOW85dCiX7KvlLD3LJDeB8Ed9zIPVZ1mnL3P+
rQCSGb/+eQN+Zh5W6t6TTxmvW6d36GeAIsUziIEcC4O+dmGshAteu9um6jrVS0LM
4BoPcPo/y8wSA+KwhsdOlyP6T6tTg+2V1STbMX8gtzUeG9np6ZEjvvg3+N0xq6ju
bFeFyBWXD46ylmA0conN+r/lOjTCSncBn4C1yUIPIYPWJG7oL367cIVNd7Bs63WO
e78XTVEo21IjmNnl+liFZVdkOsJ6wA2z6PAa1SWXw0ZoIdoE9kIwjPZbB7aeaxAa
rNbfQJUXy3nAXt4cwhFY36DMv4oQ1Agyy1cJ64UNzlbhAGgUThlos5aL55oyrgeL
KuHhuzloHgIv4/DFfXKI2sTOvcVo8g7HNgFDJgOygrVM7/Vy8f33AZm1WT3CK65d
oQJu7Q+O31mx9X4F0AJq/zGkxrT6iDWvF20c946HsM0SeM/9dloMQTBacCZ1B0+a
WmtJ0GxnnE6xw3IGHgzLE0YdOfJhvNd7FQNom8FPw2PFGF7a061u9pyI85hR0tbl
kRvu+oZE6tFokKTOb6K78Gc5NcytRyDkYTnHZ5r5P9PUTYWoAVjSNZassfjQVvVF
kilP5kPLUJXcflEW2j5zp3Qsz8q2zsEyt/SXoj1ceJ1knV/Tlbe1alprCd9d+sXG
L6imzJ/cATPcNotKw1Y9cm4GfL+J0KnR0apTtnFPeVhQAaPZNXPH1GBNrivbAS9/
QssloC06MrgLcLMA/3gl7DW5XY6HDVpkp5RxF9u5zuDBrql1ywTYzdMAVXNY9+8u
2m6S2qYXZ7uDyfM5UagSIaZclBnUx6n06VoVJflaJ5bDNcf8zZDC2dlx2FrtfYFh
jPJ98ZLdeUA8Y3z95Tpi/XydXeJY4rncRyvl/9+bmyp3JQ9j2zecK/KxFF/hrKBy
uaX6l+97npUMeWQFcudGgM+o0/ovyos0UwuEcRP+Nh29c5MJRw49lG20vWrQv2/O
UO3jh24Ptn3PkxhdvfqNFGKggxgL9JsloCoedNfXQ0l/6w+haka0vEsXjLG0NOL1
L2qMVDcaUYNipYR3vRzpzBkiVa5cH3f+/I1yJBK7qxDesnLKHVxFGN1l/JZK9slm
L+paRQUYnr7V4ewkHqSuK7sJQikpE+tltzf8e6gDTW7AanJDhiErxAaoXGhMwjQC
HbpX00f6sOec4NQmZVdFu+DSmX6eH5zT8ujxC6oEv6OcyR490urYelaUIioS2lYh
7iwKVC6BDDjvYEXulgiymgZpDt5biSRKVxdzN5AfIJnr0TlNqpmLZH4aY17RMQQr
Ze+WiKDDaAsLXtzb5Efb6j8B6l075oNU0BmPM1xQSyXj49c1YlYZsJ5TC+peYiSa
3BlpYwbiR+1MW6zI6DGLBAQHv229KtiMGZM53vGfaQglg3c3jzA1NmgUdT7q4f23
dM+DME115LnNQZY6KUNJztIkYX2e/rh2JVAwXxfv222Y/INNv1W+YQDQiczXrwg5
rgYr1O6Z7HdM1zB9h0UhfGfYevPSVESQp9aPRRLqnVdCTwZEIFEXpSVwEKqH+OyM
jIha9+lVErWKj1DAUGOqag+5QtJU+0kPY5GNvTt4YNvAEemz2jLfAU8MKv2Eleyr
hy4s4dTwBhXqQpxGDvGeLcoU1BqodKMFOUZYNEL1JfTBzQ1fuleEQxqmkcelYbAd
jGwIHOCyoMSkCwTDH1J8ASwZoOSNl6MAU10tvvu/GSU4JD005MXHT4lq2X/LfjUt
14uu4i7fdKspzTlF3dtZbPVo6P/I5nChnqZSMGvgBsMWemZ205AdSry2Kio0qfRA
dXSwGF0Ld6NVTDnrlnVxYPqngVqemDpS0RaeMkg0L8hBz2Wj+s7a9Zg0x81+4KpS
en6CF2llHQI7+IuCFA97v9t/Eo3lelQ9yLNnMqjCF32mZNYidl+3Ln80ax4s13ot
Q7jcv7EZsG7E3q1Nh1lvTkvvjYD8z2/rReYBeTYrT1yiszxw0Wt6Gp01yzQIP0mq
+uvFhgUi+bdH4HhQ9Zq0QXtVoiRB4Zz4H59rR7YIpL1OYT1QgADOibtjIEkXIXwg
hWzvKaQzaJSxw4LVOdzlSxi5BYPMj6bEvZ7CFXG5LrFqY6/RkxKOLVNcFb1YhbJi
WY/aneeg7A5OHtjvQIbeP2Qto2RJCI3zLsPLf0R72tZOJ7PfGILk+4ZySQ6Rlk1c
4zc4Vw4iMRuhRIpznJjt5zlo/WJoc+I1LFTaPB4WXac=
`protect END_PROTECTED
