`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yZHFqgI0ICz3L6/Bq5gpeG2JuSJBzyupKaFewqDevdtZF6rNnWOISae0y+8J+FCU
kuNcQlhkCLQwTyGV7WF+DtdRVbF22QWmpXTwcTRx+XC0nCrk9rghMkxEcAD/B+Lr
glUx1a91DeyvPTnwQRFgWG9LWq4slM5PNeE/GEToq/Zyjs/YvwowtfZ+14jgse9g
m3DtOcRLBEal8dX6fin/dTT0sFEAdXK6QrfN7IvIWXTOyhHXd7qRk/EJ43VBsAPm
ptXH758xGfvV2UTURDoESNsDftKo9R3en5vaiICRjeJKPocdcC4vLQrGR6wp6xhf
YAqr7rXfGdCr23CGPxAG/pP28ZbWl/fVjV2sAO5zXYyAH/HUJlp+rRGL5p7zZdi1
BKcp6bRyIfaRz2Xpo0x4GKkpyx0G6NC4zyccRbNtaeuL6jrTgp+8AnXnbH8W5m1C
ONc2bI2uPlgKqfOvimCWrAgqrKgqZvaBIypf47BloqO42DuHOT+Fa9uDwUk5iPoZ
6I3opZWMkG8xaKLWecF0eOkt3r6YelALkTb3bSg7YDT9FMPbTzXPlMPgBIAxsJT7
yHN5OOmcpRaeZ5Xb34DjM3jK+FTR5Jdy1Qm/JEeGFnoAOjcjbcCxVX0U4UK5qLMi
fud7ab3Rsj8gPu6JIwCBVTV/IrFaraBRvAcM+Q3sgKiDqGiAHScc8w+6ea2v2Sbb
EPbv1lG/N/b79HIvj3dXOTow7Ky1VXlfNwP8VZRb5gf+3aifZq84/7q7qg4ONXyE
hvFbZTMrTY4HcdaacmHUMFJ1Mqdrp0ys0xqljxUXbpQ5uHHjP/y4PgKQ4XhXbDH4
s4dtTPZjbBSpPdFCS4Mr3+7aLCohIZCgWDgpv4Je6rwoNHoSBt/od4mJ+yYkwqBC
brjQ1rpjS1bK53GCMfMX6guK07W6HEklA6HhjWoHAXnp4GJtbacskezMJVxU2CTF
QwqEZUdSZe9vT23C7mkazDbRwaxbYATfbQlWpora0UTZY1/OWHVEMYlf98xqc6uo
1/Y7jwfDsiQb9hNOFnaFQuSiH+AvP92x8t2EFWwp+WvXDKNRIsCm1gPTE7aQEoAC
279P5XEQveK8M1ciWPRWiH011KtrOVFo04FG6ld2N846CmMX5ALuQthxWpEAvXI1
PMfb7ysFwxUyeo4JB3bZHxJJi6m0fko9ZOi4C73cZxNTat2FnANdFnSkLlaldGb/
KH6kFqjTbLlnyeAAgX3swmUadoXzTvbz+Y/RRG7K1AFiKBjxHdUrKEp3lgLR1PqN
Wy3ymnCd9dc07XaZECDIopYFLYscgcs8zlyI55/EJQwZFY/pjDxNMfboHCMMvzfr
5FqaqaY6QcaBKcd6SvwjLABJifj5xhJinN/gwwO3FJicJUUDTHkYMa4AVGrtJuWW
h9U2zOdjdw+fAZfFs7sYnsXmAjAZ/QReOdkYjGj2BxyB5NInINp2luM43uZoQZL6
z29unHW4+kqsrSkcaTTgJ+kbL2mm5KQiJeoLw6O0Cl5iudr39ae44hWCE34jyfsw
MOoWIr1pKInppxTl0n+4MD6gwmxf296QXcljlg/7QrZf4wmFnejgCO5F5yu6TOdx
qhpfQ8217pXPSZprTvkTjWQs0owaOmz9hsM+UVfPy2r8WZN+hHBuYFfSv7dzCbdh
1v61lEnwCbYa7Hj7umtoz1IFlbFJMgqi5p2y3+Hy45ql+6nkQTIG0LRsDQ+H+EJ4
+mlZR0Mxv4jB4fhzvlsBiZAqYwy1nFYwafb62dT9pz0qrX1TbGKfpL2eVDSEyNAP
RjJy3DzZp7tv0VCg2Aerld1QkiWa6QyIZvSwPVVaJrA6q8SWvhmjrJNUd8V2zzQa
DR3IgYqLkmuS0xLhrV+OCfPoV85h0pjnbrHCw3kM1DDm72PRmoHidJ1bCcXKUPXm
1DHnT8MlPe8UWy5CYYEHfa5iPT9XMIu+uVwkankl2TXkl7LL+rTls6CHM0a5AszS
EkjsCGA1LvtMWNF82rrNQj+hXU/ARMF1bNzAkbR/0USelxyousmkbbauWgwhMXIy
U158db5Qw3Eq9J3wY416kVpVZxIwqElVkEmpsFOgiqgu68ltNW6Yi+rZmbEgnjWg
LiVVDAdj/8c9e6u+bMPGWNcMUyyWhRVR+j9o0lIcbmOjheZIsFIh8UGy78izz7ur
hW44jtBNS74Trg/kgdebRhHlQw1ptOXXRsDEe1sipYsLZ+cgPtTdE5u3/PMGcf2P
9TB1Avk4XeqrfCd7P3LWJwjCigfhcZzqV9W5gCftwiXI2AKP1NyjYAWPDe7jqT7n
zuEkWWgoxX5nHZf0M7Auj5RxBnRwQ6HGUhOwOXX0gB2PK8Yqo10oLBFTWjCYvowb
VKXyoZA8IKtz7sNV5KsmdYWDX0lBFIgOMvnYzLbBWZ0DDFQCJ7TDhOYfaMGf3498
kizfX8Lpk8SdXd9VqASkIUNfgmKjZGE5/GcyxKpJ7dHORqiEUcvwuhmO3794Lu1M
s/y3CVEYj5i03xRfOjFi4APE6Dg4dB+ufsOj3tOk+4Q1Ty8dWcSxFadH2paKQKd8
7VmB95gmSScREfFc45I8nzSloqNem2bLPSQ98MU0+d4yn+1v6DBdPbQfPhzBor7E
avDxZsTCDhSYhCKNO92RmWMP4qSwH7yuJQhzdLN6tVWPKNxgYtODu/3sWbR70eZc
ENs4mW7ggaWnITwMzlV87EFEZ9kTypbMxGOyafwuH+pO3odjWBdw7W72uU1QtE/i
/ohAw/1oI36yeEDYhOC2GmBrJ1OSk2fYVTmT2v/izmye4ftjVy2lQPAnXsG/MyQz
I57SAXvwXJlXOB8bnwO3urqdBYr0oVOGMhj/tY6egNhBx/Xu7iUEsIDPHVAvcAkx
eaHYVlYsrCveMsSxwKOgxys5ksnvsqOE9fJ2cPpPpKIyNtUvtqVHKUIMTPEvnnQZ
kMB8Wtk1pqovnR570Vkg+1/o1cPAKDruz2dm8aaitUw7Vxtxu3cWCQYGg9BJfQpO
BXPN17TShBXAxKMzem3fSaxiqzJFE9o/W7woMj/M5yZ8OfIUTPhcP7eEqHyH7TxN
t7Ue1nv26NnV8xbiFnbV8fkHpPQiLt8gx04QLBEqaIduVwH7s/rbfC2snloX0Bya
M0fodBot15my8BnCAXJ2JQUe9TxePz55iOooJpRw4QA4mbW+JZKKKfpeonmDamCM
Xz2FNXEEFFbj6gvyeQymAkHfdu/rlZP10jidZV255tyQc22eXJ8JRKWdVTfDSEe/
dkrcmxKXoUBHaLyT7WeaRSh4601B7ubGIoBSEj/s4Q2T9gQRtf/MAw44ZXqfGp3A
69OIX32V//waJCb2ProC1MlGqnA3NH5uU/q9RS1f03higbyaz4rOULoYOKe4LpD6
Q2x1qCLbquDqNwFZKY/mYNu+t+8eCIJzah9yiNsQMx0TOH6/M+FmWvwRGb4nKPqW
S+cNaLbJqDG1q+Xmcf8HKPYuBVPDfeVMwFjigc+5kmChnTkW4JOYfNQYlAtJ21tI
sGtDF9Z6D/6OJBGXbj79NQ8eMQ5HiUfyDJ2tkMJxEnDPrbtjoa6a4fQW3Jbv2ilM
i6J/KJYPKdacxkRw2c8BS1cVup5YA3tsdW5qOE3RH90Ghi3VG9uj1jgjRAuE0nit
T3Q+1zDsoGE6D32U5XdI9tF/eOVrCMVoHZCNGwOJPRSWi2nwrdb7htc91gQ7e2IW
zbqoQR/VjLji8UKuN4XKbOccUYWgcNZfD1WRSrvdi/d/cGYS6chxrtxkKhbN+pzw
giIrVv8myMx79OapvgPjxw9BE6xj+vqtumgS3r4kcYURgMQKp7sCHOLBETVUPoRX
zZ4mMdF4yRLh/rlKuE/W16vSUVEVYajJdPg18NG+vdhkV9oAYkWfGmiJ/45HjE6n
rXuEqDp7LRFjK43DZUPZPZNHQ3VH924lbE5Fshx2GHqUpnP1exYe/ZHp5L7/BQ9d
oaBeipj0oOGnRsmdqdhbEEeItfwl+Fdjt1hQ5VCZjcAv3T3onA/rzwbdjCCu39XM
O0yW4dubf28Aujo1pjABMse9mMiBL0o9kWeijlBb7dR8uKGkXsZODt3EsZKYsEia
BK4d3+xp9sJbFkU9wJvOQHHN4Odl5mV7mc7nSZfZ0hRqZ5k1HDbt0EuYZ7Yv9xCj
snqI5P0vVZjelrTG+qDqAZswuw2UmPW6R5eaQUEKgtQFHtrbpe0n2Ct/0MJLyH5h
gmw3Xh7ZENMZU1tiJiP8xGohWuo9gZ/+1oPFcBML/vIuVpPi4+ayz7Zn6PyT9Jjy
oLaSP410QvJKjLkFUQ2uGFmbcYXtKc76aPKml0gQUeBjcuJ0bEAI0ryU1AvRWSeS
hG+J5lJ/q7RiZHGtmnC7P4LUMhvIMnopYM2d84XPt/dlbPtyGsbl6tUYPdHHRnoq
bDCrLSDE988ND8w7UNvV9bHrd4Qjl/dPZGnD1EGx1qHjkHC6buC6APNk/OuGqWkx
c0xs/ANQ8hsiRTtjoG+FgiBWuyP4xg3GMiEt6T0Ai644b5EAMGYtGZC2VmQxKBO3
OSg5m9Y2H9LA7gsWOIZ71ii9mu0KpHDQiNND/7czsSTiZlmuwhZD7y6hB9wkIAaK
TQ6Kxod7Yil2dpnDrpjQk/TNLAZXmWcWMSB5vyC/9uJJS2750rohO1oqCK4BX+lz
9qEloQrV384fnH+UlLtbnMZhj3FoUZVtp8arSlyyU1IaTL1FXzvNcNsqu4XPYmId
wBX+s2g8KRxAlD/pApp/VHIhRqTOmzBLvUTimq/xsOCoBeZiOYGlPN0Z5vIS/jBJ
8z06WKkR/jmxZr5k3JluK2QgSeGywPnxn0GxoCtTtw5jsdlxDCz5qqjxNj9QStSm
vck+qhGQIZBU5jQLqcJO0uTtXwqTvvIb1DNh8OkXIAK77EyuhRpSdIZNEuYVS3ix
V2chciD48RfNWjaxhL7cKceYGx5rSSz2wryiNcF328om4/SQ48rYowsZLqqOq+fT
4r3OhM8X15byLLCbO5n4wdVXWI5XsexapolEY956oDOqajn6Fn1d+uWRXOy3NWPw
QMMaZxZYSVoaN8Ef6Jrd90CoYSoORAFU2ELWwVaORdmTJ8/7HzdQ5mwleq8LkzEw
3Q3ifJ+aBwR3jzXoqBheWmf6AetfwTB0mEqgC72iekiUsnwshXzyp4akYMWx2Jzm
sTVw38IxDBywRn0QkbLrRnS9M7vCgsViXepWZmRM0K55gpneZrhjdb7CsP8+84Bi
nKRVjJBS2IyUShe6sp2jGA+/Kg50fxN9ia32jGBmLhkIHIACipmqTIHALGYWktxz
m4ybRF61QLNmMMpkjgQUWgMd3W45gRGNRt1mWH9BUNgLPY//PqzVygwQIN6BqyuH
5Q72zX9xh5k0KijO54/MpyKaPFFH5LZuPBkErmXDW5OoB2BDj/SnhCdIpd9yIo8M
UOTk3b6+HGChtHrbqOXUBJLjEt5dnpco75SNDB0D9PA2xTc1saW7E1lL7A39lw8p
DAHTZWDJTXssdP0mz5AMZZ6n/fMOeiQdoeNxG/1LDu4LUUr7ny3aqjIT5oFcdmI3
9L4l+s6xI2fqU2oAtxCf2MCFtvW5WTYIudy5JmtyiW1vICBc3wZoYTiKlHsSBvXb
7N1ceVU4Jq1c/6kbyiLJSdfNWmQi7sACxc1eErHK6bKQbWlnbUJu9zfeYtAA13gy
FGS4uKNwB9K6WTIYqsxwo/wDxMv1LQ0fqN64qRdyRViXn3A7treOi6Q+VUOCiZiq
urdsQ+e+g6vK02vLn98lIBU/MGt2cgwmbE88LqcJsYmh2+2JROk+El1C7pGNWM1E
TUbsS6rvreiCUoEtJfPQzCFEB45UnYQWetVd/8XXiWPdoIKTtPlkLXfyKCIU99fm
ob2ey8sb5X4taKd58SHe2ZQyQWA4b9cpgXV78c68GWGBITWW4csn+8cug9ELpAxN
WXuYdELouYlwCPfA4ATn+4RnCI/35zE8otLRPkymq+GKeI6AclNmQAgX3Uguzadm
JQT0O9xfUYHHFa050CRn+vhUERR89FpkhyXFG2tKWW1FzICIBllRxMCJkn8xVBmx
Dy2oDTFJV692wqGVwr5H6Cp7FbNaK4Xn4VN7n09EUN8MSmazqFV2LKsyCm+qBUeH
Czi25oiPfGZZ1mNZk+P7KGJKge/aFZLGVHxWZYXwVOsn0kq3yhhEx6Rv6dlDlIf8
S4ZBkE60ePcV0pdFd/9YTuxrcH5JkTp6k/QSdBg6mpiXbgCLXdga34SJXIkaFGx5
9mjTpxqplpTq1i8OvrhyWcAKj3i7q/EgL22fKjbwtMFKOZ19ArSvax+E2UtAsDLM
kR1KdcnQqBWQXMWLl0hQlW7kS97cRLXmK0xW1zGTY6SEF0b0fI5nemeRJCHHr01U
Pi+bHzEgugB1bVaQNDrM8qeoVajOmbF40ogQTYZ65wx4tSDvBv34Rl0UQUJ0cUWa
G03ZaPlgjs0nd3/cY19hHT8hKgO8rrgU+WLvLU3YkVfgmJ4B1m5tqifY8pea87ud
bZffjzy7fvGtzqozlcI0umG9bZk1F/CFwxf58OF35G0eO7hYmOogDabeiQC9KttB
IW5k8jvvl5JLXLRrzzdu2I1zAfrFjkVXo6PJbpRBlT8viGXKg0eVi+DABzwq9+rW
faHfzHwzwGAionkT6yLA9APQaOzQ73MtfGcrew8eJIW87FMW0WXPNbZGkJMbBUAX
XBvSuTpUO5SU0U494G5jSs602VGs8jReiPgIM94cFDMkTRqxBjbd2DMrBOhmYi87
0I7lLNucDQl2MWZmhozHqKKnEHo3h69YNNBO4cwL7EIkMmQKK3rXaYooualBL7o9
9FVpI5GC1ZquHE9whiaoIVVp5N92Cy7j6GAS7J/9Ag+3A3FDoAcU7D5Vehu9UZAB
Hmw2ZxXPy1kdQZyGMAkpZO+G2bLNPQJ34KTmAOozp1MNZ5DTo3WFOHQXRGn8hywL
uoBE02JXpZKNKyYiNKy18ogWkX80FX5r4sYHrcWgPaEwIARS6B7s7hmdOtfu3a7o
KM2PkiWhLsFFloxfZSSYdg+MvTkGN6s9cpDJtHs0QQZS8DeL7gChr+d0xCKCEqgg
sA1cLPEX/lE9OyyeltPsIzaxjMJE8PwZAgKPzEUqCyAiV47wpNwvMEaa12ljJ1jM
n9RmFihcRRfPvvNo4pPfCOh5BvojXWLXXV8eSAjbenahlxnhRMjHCuTThsikYoqx
Fvr2iQescprfBdeS4meT7TWBI4CVvS493CQX1fPR7AFVrQlxi27/HflK5daoGnxy
uPt9k5NHUOQMLrTPrFu1Zn07Jog/EViaNJKg/frpQ/cjXIlvxQQDO/jDSa0tDwPH
MgtsDz6HRmxYpJTOyvuafU6TSosY/FXkoEQSyLvCON0zjW7dzNXcHpK6zKnHFGOr
fQhBNaqEyA4Vkn2D+rKraYVzCIferDoF4yPe4LW2Lpdmlh6Hukt3qNW2gh5iumYJ
Kqk34u8Nrfj9zraKNOylsh6EnqPYP/oeJ4qsmOeBv5yYwrRr4ogy7+bJz2uUgBnb
T163nyTqghpGalw92A5WiYRl8Pkdz52aA1LfshmyGiK3YBdHjZ0Jq29AwyiJVqMk
1oWFoHgXwVIhCCewZCGPPBOqlEEBjlFxD075OsCr9I0twhbIXOCTroCnoOHXwGzo
6Sm6AHqFNfDCOSMYfSBjE5Mlg/1tl7740v7dLcXXwAkwmZelsafL55FzkQhDHAfR
5fs6x8H7jtYOwpgSPeVj3UHYxr2hab4RJXV59a9nbMBW3NbC6+3YBe8CvlIURoKo
esF1oHrP/TDY0/SnLHteoKUb8a/9WbFUQZ/EgEBTjvYRozdkQ/1wE2O0sgUjC7Hb
JfvB9kNhhBFAw6CRs5e6bwnSQiN+31keD8R5sY+9hZy/1O2SGtL2Mj3RcvcnRYVK
JTRPqLAQkCS7OISROlcV5JLO0ioYdVs2l/fmnbUJQrt2ZfEy3GCYAMg6h1tTqRXx
6xXkLyd3RFRF657EgLFc6RpJO3F5JINS1RCcP3hzabW0Ow7z0iC0s9oaZ9tiSvb5
NMHH/1jSrVcxw3neamCvgNrwVBBSxKMee3FldWAloEyEm3R9sN5mfQNXEzhAM7p4
tgTPOrGmmK/A4UopufU4HPjXzRrvsIFhFCzhUjiVO3i3YIZHBnFHjUWjcBSc8H4+
AhgzKE8D0+LmITYNqwLN2Vci1Enr5h6bxv+8Pgs/bjFoP0tqutJ/EeYy4kpmL5Bj
Cu9ajjESPZa0FM7SAojafjD5RbrnjP74Cmz24pP2R7KXk/nLlVBNBbXs1m0JO7mn
jKyiiW7tfBZbik3kfzpNHHKAVtmVLzVxYFNFvoeaApQqea1WhLrVzyxk0+9ac4/y
f21zV35chF2xM90ezcdUbKxEPBzgDmqOBE1zOArCssf5PnoUdREQSmAqm7M+yvKv
AL7ZofnbMmg3hIk0px8SDhtfSpGMVaGAhpM+fQbBukM3GE/US1/UroS6WJ6LPkWI
moLOtuLKwvFgAUTsm9YFWO6a5SQp40QOPiiDHIpmDMRlqywLVsqjbvl7/NHrga2l
LNCWNH5AsZljn+bvpS+yWgckWWzKnbVra2eV++loYNhI4GJa/3cZcPgIb+I/d4t0
7pNlCEGMdftdJJHHaa7G5jUlQpY1hBb6eoLflC2ai5wK2CMX4T8oFn91jr482fsg
qAdxvnd3aJGPEyJWPBzUxtH3UjUxFVZvgMI+iCjw7Bc95iNYL728N2TQCPGPKW46
b+995AdcTe3U7sJJrRHsHt6WYUkTDLzsCC8HqWlnvgGIYB6Exhzc730ay0ZinuAc
3Rrw8d8rluiMJ5aX5IoQTHPQ17BOMYSBTsIae/VCoMRMuQwh0DdYTZYbjPpfbPoW
KWIaCUno4FUUvh1z04O7UqICX1ZZf8qBQFAxESQCKju0Ke5ON1iQXp3oZaTdlhMA
ErkA59XqZgGG8lIs92145+++MzRRhKk3UhRyuRmmUQlwaWfUydNAboDfP44GyEIE
9iLG9SlMx/EGOQN9AHZqtIM+W0f4KEPm8fUhXuIUapoChchOtURp1EJDOYjrHX4i
n7LsW8/tP4MgmNWY1n1ddYV19Bp2vSyCz1N8HPGyE8AHnTBItzi/O+ABQOqilHGJ
ZgmIlQ2iGKSc+8EoVZtBnZuMBgtfBXyGtr64wnMuBWVkprVKNI6jC2PZdSAOROob
BWs7ovoXaxt//9yd4lLAjceTjQnHjx0J3pDhFHqqKrPlIIEAYpHghVA9Ze2cSPui
tg6qtAKT3KF9bF2wPRhafmebrw/l0L2Mh7jmOn9paao=
`protect END_PROTECTED
