`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i3hQOzKGeozG8TGmMtAliDkyLi/X3Dhv3fjbN89CoXa1584dhKm/Z5jbicR0IkIR
XxUqfSqP47vLelGH6+jywesChelfMFahMzIvNkf0mRJWg2OkdPd0kqZvoEdb5zh1
CwiGI4crdm3fIOGs2P2BEvmG4fYcjG70c3CB1op+8oXuQMBMShsWg8d1XccCdChd
GxPwbMtzTVYiu2jMbIbxOcGuuS55kSCPHEurQ/i/4iByAEagrPzrhAzUsSPwsmXV
WL9qkoT8xqSAg8UsWrf26BJbCKc26m8o3DtHpJTKkK7zdY3DeyEMKDZCap1WPkgk
EpApyaLo+n9xYEfmdF1GgT5TK0vJZsHFV5o9OjX6922ujSEx4b8e/FQ0QyFhGG/P
iYwYX6V0Cel+V5/g0gAOnSZ6aeWJox8ZzFiC8j+WRo9oS+DwSvYmcaC3sTQI1Dcg
4aERvfEXmLHkP+VFYwb7iL5mJ+EZ/Wi52kl5w4Py4Mys3GcxlHXsv6PhKh2qP6m+
/JcZ19FgO7hOcP6gKRJPuBiOCbTJ3Xz4+ywGDSJwpRKt1+Ke3fimi/txIE28YtoK
9v0yt9gcaL56rjUjxMP2btHvxbn8M+Q/N1l7X4Mg7Wjxx5dZENAF7NU8F8mqP077
SnTgzT9LJoizsstU9a7liyZNNK3XC35VdoV2H7ucmmZDIIzcnO7PRQ0S566rVMtp
8KKJElJTXQmiYWMznauVq0XlE0kbFny5zIVcEVt5EiMwTKnktMGkm9x7oPCynFwt
bbqG02+0UsrTNMkj/+uT/GXlDZBlaJOAkk09CyLSEeyH5d6wBuunCvsiJtX3Sngi
1Mmcy4Lc6EeMN+qpwBC42SwaO7SKF1Yq0WZyc3qhhuDvjDuTtEXT4iyItNBTumu6
jAczEWK6s+pD8C8mA4O7nqT21BXl/+5bJ1ugs5RlYHCR5/vf7cDtHLTgZVP68U6G
5zka/NrHrMhIaWRWPsHkuWW2Umf8Hh2nwLI81LiIIqwgsIW2TKbharuxMWnMxPKG
CKj6qntIYkAt4JJHx0zY2fI0EdTQdJsF5l0EHjNT4thOFzfm1+jgbZLyqodYpTOM
ru2CkHU8N2Dy6W5PCjA+Z9er4QyZiMMy1a2LM7e38MpiV/IohkVnhRUFiZAQ/KJV
LESF22Gr2lr1Kt3Sfsvo1sp66f8uaMonqwM/+5lrfFocDr3vN+6H/M0Lz5ZdjHzu
BXaE9vqVHi3TpxIRuonpFOCa7+BTOfSE/fjULlaTH027DeMtk59K4OaaR6Sr0iJ3
Om24lJBopJ3cVKGk4M/sF1uYeuRav7JgTXVbFQqwO5QJ6iwtvgy7JwRe6de7XBQ3
HBecATCeXW0TfKBODADNXIkQHc0/BltAtJ+s6StfJ90LhJ7s5thuBEsPnyx9vJjU
4uy4Ec+LezDGA7Di+oz9B7ogR9bsCRqWbHPnHDpUCMuMNrSv1c4UzWF2udd0IN9C
z+lDZc8tGJ+ROsADE0VYAsguABr1ncQsP4hzKLLSXZ/tn8uASDwJLI6NhWOt5ylI
ITG44Fyp1KQWd1FEGYIRjESSoGeosKEtutTfcjpm/KL0FDwdYpUSdlY9AZqQZmdC
3mWD/IYYS2oB+01zfvZdSqK2j2qUtJhTf61y3wKYLXrIAxmLR88gMV6fcQJeuUTp
WyKBjsistE/W+K7vqSlWIhVvqoKy6ZoF98rP2+YJGeQY/ZO3m1NX1IzQrSxs1r8s
GrtFCq4nmCLLG6WEUyX/JophyyD95us+TqVsyU6QU17DZmIgqnanB98JBF59QRTC
xu2Z3SERS/BpXaXZO+RvbErklL/b0r0EME1pJqVvzrc=
`protect END_PROTECTED
