`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NIOfBRhIH8nGhqhbkZIWvhHDDP+9nF0lD6+xLjNNrOO6CfSotoNykFNcIaw1vjSH
NgXXzDgC8hqqaD9lJ3s58VVINdQ6CtAzB86Wfa1cjSvfK9BFYac0SBhobTo6fq3d
1UAdkWBJb8naFOenxneeL580GF+OH0EUoEuitfwAYuWEs6jvmvlFqNkAFOIjGvUk
CjgpQPw0RfVkVHAGXbWv0UId1MW3Ok0VWmyfx0dNSJfHQkkVf9qtnm8V3IN32Yno
MCVLTmm9FfpnhG/IsR2+XSNURtPuX76ujCKZkugmfm8pfNf809jx3wp4J+whXkxG
CzQuhHvrj9v/nejYLzefQif9xrKzJ1b/myFizmiY7ZahX/kSbhR5fjhibB6BnFTK
Vqex2e6C2N1EK8wgip59wJ1JSv0DkWDn7ZNO9yDI9jBmziLzQUQmf7CNj3YdqkT/
3PMjF7UStOSEd/ByW+TyZ0pfZVfSNLj7U2xIrI/UoThAnA9YxXy44K8zmC4InNmY
bKF4KTSUa7wXXWUlLByEo5+pfN21WzyLsJht+yBp7M43Hjb99/5pQGxTuF07sdtj
o6apc2Y4IwCVvddmpdtQrJh3qZLZSfoGBN7Nzw0Nk/Ets39nUL55X1C5KV725O16
so0Kf5UR2rwWbNPl1Gd3dSbUGHXF9h6S0eteWxdobF/0HDg6KJEm+hsu51IcelHl
5WVzAJhofHZ0zWPqD1Ozk3F90GRFzLqY8Aq8Nt21REVpA9U0tMLScYJ5xQslwD90
PkmRAlnvGaI00S96efE4uFCc9a5tIriEiNOva5K2CnJC80Iua26EFFOsbadzpCKQ
08CE4mni4ZALP9jvlLZLVMyx9WP/NMc7gc4naGeXjWEmcNck9LJFHaAwjHDwfdP5
5ZnqBxdbg0KqLEQu/oUTgFA4WNz/2USG7P2lmu3mnOI6NZW8hkPFH/J4Nj6NR/jD
oXnOSDSaHTiiBt7dJ8HHanvaLFvaDCgcUJCTRhzYvZQdMW2W3nIVwMicY8q2WaIk
8GomKs0ZwVtMyDwwGp1EiU4cxOVAs8djoflz8xkr9Tpfqt+ne2gQmnJhDzLN+Zgn
kZfbAvcCquzkLB+YQHLC7LlcIXWGSmrskPoQfjnGYWhquOPp/Nb2Wqr1T2dJDch6
pUYzuWXaxkAp8p1dPgtOnUQPULPFSvhwohaXkIyOhIsmrYyjfFhDr0CWfE56RUSq
u/m6L2O0B7FJmMzLgR6slAntjMt+GQ8IqJi63xg+jHyrn4U1eDUD+pN7XIxegdnE
MhIaLmr0ZZ5UbheyYT75sKFJrH1ftvUohOKePDZWzK4Gxz4K6sAgmCWZ1jGwPTrN
8yjKCAYZSgs+BMhYiyHszE4JlfMyBly8t4Jn8EvVlHohCrtofXpHKtnO2n+CrMaM
6uBt2p2hU2eB0HIg4OnFqGXakqdjKzFSzFPAsoAoxgL2oWRkJuF/fm/UuRcEE6+i
tfi1m7wQvu7mnNz20fe0KtrX7wHas+FRkNcKk2IeYrsifDNLcKnza7lkjBPZvdeA
JiHWWDac1Gf4j01cb6klZ3x0wluPeI82+AVtH2EFo9Bs3NmViP6JDKyBVgkCg2qM
KP0i1VWS19kVf/c/QUTXWwk93vhQ0iOgBtdjrpaQ82X2fTg8mgmZ2tem8JYildy/
YezTWv7AgW5iUvhz+j2A5PNIdicKo9MRMRgEC3RljjwiWTT4ktt2bq8kTqkq4ZN8
zj+/ORH0X0O1jyrXFjbqZekjFgIV5m5yq2X86Sc+dwuSFH2aNVnVm0YNiH6A2AsW
BGAyV8cCaMihS0STCMteqcyQ1XdMWy1m2YAVB8VfZp7EWZfdxQDSKnbFUybESARD
LLM3QKud7XdROjVdwPfOJ6O685a/SBF9aFh5cW+V0HrjHvgC8xnXhQXR6stRxM8j
HM3NFbb6on6j+Rx2U3zd66xVtwVng/pyGRm2Ne0bSPx3x7B5VQ/12lujXSi3tEJc
H1AelfKLiRT9kdH+Wm0c+VLWoweJoSNSliv0uvO7Z8OFqkDcyBrmHzZWQrBakjcC
zgzzyXtNayzYE0muvw7er93iWki7ZtFtG773xaA4YdGNZSJnLQRcSZPcJRzg/4zw
XATxy3MwqGJhGWcUJ9B8Y/gjPOQOmnA7vTW66GWqbQPzgPZnn4g532TbbhqWKPg4
EjqKimT7ogkwtxhqx6jF7txM39ReDWnYV/791Q1x+I12e/LcVpk/PoGWzvwtD0SX
1VTrfEdjFvzdDPhPl0chilg/6X8KFjBUcflatOhqdvfhtyzCfDa8RglD5Hlrlym1
`protect END_PROTECTED
