`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yrg0jPu8vxpxK3rEtSLtSIFp5y2v5mGMuCvinAJDeprHZ9bAR8Q8QPRomeSfnhoa
ZY0ZA4jY7rZOr3TqvvDcA63KVchQS4EhAWP5XXgUQ0yfIxmYDASBgWP6BsmwgdRC
BUlb5YydyJ6OAlS4k2yskiBoZ+iVSUYf73O48ECFJWbfRoGrwGu9YzFi7MCsaXDM
KaaHQEt2MGuLyPgAEWQ7GMJJ6VF3F5U/6W2ua5t8M4FnbktjehYuq5Uswd+O5ZIE
8x/q00tLnsLWFCp9co4QdC3X+yIwVm+Fglbv0tirtH73pIXIeAhkzRpCXG39rDPd
U2/D43rLz3xI5OkgKUHIsUIA1ZgPSmKKDsQEcpFhJeCxRerPtOPrHT24TU9Fmnwj
zaDsmZxN5dyADO0m56Ult8fgJepJOUAPpRXCdVRvBqquJXEN666dtTLEET/djnFP
CjfzHdROgkfr0foGVzF9EKblSh9UXnr5tKlRNYeyg5vpOD449JeD2Lg3JiUJUQc1
7PPyWeUeXDOP8caWPpzsLsjHM8NMeYLrVfjOgW5enSHDaTWYZ8lIgOaxJLSiESz3
UT2xOdH9K45m4FJzb41xGsJZqQLPvKHJg4o1JnYO6fA6Fkc0tfwBctcBAVgLNELz
wP3QIukD6UfXe+L3kcErfxDCddrmRjL3C1b83jrE6OWkEzlKM6tFURFK3b8b6P11
Q0sp4gcULqFXUsqAsayqV1dcT933+5zao4vt3aXIoflE9dBXBE8qfox9uUmwebDc
UlDyxZAHujrCvS+ExDzlesFTHeEB6Mhb+L++r9+HtHUhfdtRFbkOY66y6i89o7rD
Pkmz7w32q4eFAvjE3+cWDNqEI9reEowKVssjKHYxdr4hmyYEieRWifBYgZWhP/fw
YGhT53/2FTIX4sBQAlcF81jaMvkr6+92y0fLh0FfiKSQOECixF4AbxNS0ajAnsPS
QE3+oDpg6DG277xWMmPfCqdcMUEnzXFrj4fKnZFHbxMZORPnFNeQmXm4lCLK0h+k
1N2URdGi202KmjqjpAU1Jbk2eyA0TC5H4EfeflIUoolN9FUfSBXGWEZzbUIUrDsg
93QVmBaj+nTS8cBz9mwiDKy+YfmavgWlr9zlgqXkD+m0Ot2mXikQ88VfetVjL/7I
+GTzneNOANbouOHcpUeVqpFBp2uUUa38s/qjiK7FrarkJxfT4Nsulbv/DpBMWqEw
cOt5KVNJi8Xs2p+Y7nSNtpzfwTEgwTrRan6f0N7j7EYLnvoxVBSZQwV/pk37Aq/l
Vm2f8N9PMcXZg7Wi51jtkecfXR/WogA68sadHON4YsSMsJJ9Ee9YuIn2eXmdrc1l
QvszuyjIuOMMefZIS/ZMvdCXlYK/UdfgxLIn3GbTD6O4he64HWREqi7E7Xj36Lj5
H3WPHwL0n9jVHwtO4csonFX/3/tjE5chbVeKuRkWBRja2sSmWI4/f3f6qt7Ftf/m
ac8NZQkoAgdtd8p6wNnpVCs4GD6lx8xQGuXx+zHpO1h1H0lzg7rMFpVtvJ8jL4O3
5BynNvZR3FzWtfZ+VfSk4Ym9xQmGzN5qq5SpjlUsEH4SA5pKxAnCemy0bt4f5p0U
rR2BMi/rR434eff4VTb+KhVjoEXp8at2ulAVSt38CQWJtEkzpG5xL5+IwwjxwoA6
c5jUjO3ya7yeVaQH/pGRzTcSVgiHZGsYX5cbiVS2eMPxmRASHRoYVQTjhzoEtdYj
BEFKvGD6b2lKQM8orZtfJh79RalN1ehoQFqmvyJ4yokVwcMoaf8eXqQ9rooJvu1p
3sOoTY5lOOXnMlYGEdVtSdVTG2atb2lNSkvjzOTyTz9MBhmw56oDRGWxsc0KqfCi
VVEn1uQqmQdSofDQlAj0XFWlIo+g4Xp7BXGjIsvuZ5VwIYpHg+oGzcqGoh2W38Js
sxidKEQ5qiqu/5VvsyPLJSy9U9oVCVUmVmDQvFzDa7EYzGCmFYi+xnnc+tYMwjZ1
MmOIw4tBCtLPLW/TbjHiN7NSAEty+bHcdnzNnnypdUGiTVSw7iNctiwT/5BUOTND
PPBRGjBwEshQ0LHRxCKmjKHxpASopcOxDTDj4zzV9bFzszY3FNh9/uXQHgKSAkLv
aUE3KL9pMe6/4Za0FUjK1/Ju2i0Y01v/zwGpl/rmBcF67w+iHfzIDDtMZLkYFKuC
p6fnI4J55jJz4QbEbB1zKmm+1kgATnoKC+kSzOhUB6+FkjCoXkbGaFM0n0l/WCxt
G8P1zgGq9UFK6ZPLoZn+0bNtWBS/N37LVJcq4qYgX/qYchda8+14I7tffbAb+QiW
tBypnET+iIMUHwF6hkxrlI4ncfAxjGC3UtVuhQsV+FcJjxuiHMMwEa3bGLECX/vz
G0Vd+sgkDi9RCcQeZU/hI3kgbqO5nMc5S1/dJLfKl5UOBd5gtZkaMCfA5s24lr9q
nmm6qOday8hT9ym5jitiW9Mslp0VVvVmAuvfOCd+vH0gJITQXJrRphiUbtqRC3er
IqVhoSFjGHY0pRrabClkE0naE0k19fSjVR+96uWrUWwBW6CkpaprtpDPvcuf1ld8
RgyMCG+mFkdd8u2ojukuFQaeWNZpNQ0WK4CY/twxXPgof4jaPQgLhoKNHvswmP4M
wMwHtB/GkiuFDZBzTIi7l/B5mmbOZ3dcFEGS0ePOyazq80eU0AGuzFg3+Vs4wLAl
ElRDAAvxWKgqPaXhAlOomzfJOJZAB1Bj0ebXNMXyzbsl3lVnKOriuJCMsKDxUsEB
x92nIjDLlRA1S7qhTv5u44Eb9bG/DdJqXBMEQEVi3y7DLK0sUdtNnsqBCn7wAtIU
JvM0vFpoKGcVYVwhcXTBQCqTjCVOdUnrZma/EnzJ9TcGEqqv7fImWUOJz6ZKS980
pw9upJ9eR3Zb8JLbdOg1WqIMqQJlc99MlNbfo8wMKTDzk6xuR3LaeAckU+yV5WAs
E53b103PRr3w471ZvsrguNwhpzF32rPke+KvPoc8PA494XNbvUhqkwvBBURlY3El
ot+hT/dO7V7KCT+vfRWHwm6pwCI5IhEHP7QPw/ceJrhsgEUe0Ep5+qmGwByE5O3R
yMXHuhUEQDm/QuOMlA3F7T3r4Yqajd7NgHG8Qzb41cXYplzoWRbQBr0N17MbTp1E
/7b3YJi6czKM0p7E7XbjWg3JUTZaE0lWAKqs9hnAx/brJY7cz7/m3PtDnqWqXT5U
ZJVi5Jpv7i1z7HPfWNhY74oFsFHIlYfhKn4QHni7hlc72nnKNf0lYDSnkfr0AB5E
UoO2TPklFjRnRAg1J0m7GYie9ImITjVYmUrq+sb3pF2AD99ArUzFEnkn75JXYfYx
Q8MpVJ5GlCPSgQYXFddahlHWIGw/OHyAoUEtMKprT65puFQnlvW0vQ8vR7rZsRiz
Bs49PBvp4vBCcTyFO7fcDHiitF1TfiXtAxrmVMK8LVvOtd7rAO6XCtkiqabLygWb
WCb61kRW9WZWnSwlcgOXPCHq6tUVB6D/8h+qAGtIMKnst+ujZEP1BOnSHLdHF1AC
gRJVvWd28uyzgY+3ap8hkEyRxU6iwNYYV+cMMcf2HSqXAccghc2gP0J9pW2z4DMN
PYIZ+6cfGnPUUOD08t6TMg3F5iaFRx9KdPdMHqITD5vzrYBQG2SKAmSkagRHJsDW
AgYkB/rsV98H0l1JTjxCW01+Hh1hbZ3dM0oMs9++YVKE0jzIALGjwkrqx+T940IO
/TeqnkD6D7VJOkcjf24ouowakD7W1e/Lj/WIys+t0pm+t3k0rv0JRmjDMA6uvEMH
ynHdp2a3x4BL4YzcRTi6TS8eXmSCwaEdS73+pFULK9dZrVZYF3oVzdrkIbuuesMe
IHUMBFIhpQKV+NWM7m6emtmA+wEYhCmcks4+QT/yj4b21F9oqmXmznErfGKSLlE9
TnWcvjos+E2TAOuO9TzFIAjUdwkWfohhYahBwuskZMrny9LOddI5GRjdh8IiRw0J
ZhcQ6IIrTGjse1zXolhkUF2WyBxVSBDie3soQsZiJITqtMYSe3liOYCkGPnDKHmK
Vi7FXD/ns/foh14YpFp+rsitXiVvY/YbvI8K7l5u2690mmB6ooleenMc7VbFpE6y
v3ZIdXxWeMKiTbMjFEU4emBk5951+wdBfoOcxmwQMJlYN+nDTNzpCXoagh5r3gKa
O+2J2p+6IytAQ8NgPGChJ+SmZMMnKvLPNLIvViVSKboJy5ZU7H6jhmQ56JArqj+k
JrqfuJcCFrhtUL0E70DmMdalX7QZ+9IUen5Eh9IGw6u4CO9y96i45a7lvtjn0Bt/
9r3M2MCwj3zNc7OYi4CASePZAvZF6VZ9CWk8rGQ692LBKyY52uNlJC3VtP0qRzYH
kD6l3kR2e/1fIwX/tMLMilEsCRlVLugBk4XgshHdd069IxiCMN592uWTkDIvje08
eiGX2UiFxHiVePyLPiIlVuUVCwx4P4Be8vCIJ7s3ZTqZAOWKJYo9E/bK2LU8iaCB
zRQUxzsFBPbTuXlxHEy6yp+xPXk8bOHrRyyBcbePNs94UlXp9kK/A3oNEl9qYyUC
xBxblruqa0qrOn2px3K7o1skxq9znT7vz1mUvV31rF9/DNMIyDDO/A7A31KENPx1
4AENY+nk6/2jynhxR9RvZw==
`protect END_PROTECTED
