`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kg6MG+7UhRlRAeW5fFgTsubd7V6eU8qtIPCbrsxc39LxABndQVkgT7vRAk7AVOJ9
/jxL00M9ZxjQIcaCe68kFwc7T3ERWntslYdbQIUii3MpFmXOh+8w0vrR7BfzuCIY
spIu0F9n8QEUPoPfkyah1726Oaa8zv5MdJ29M/Vw9CQbJmBSsFQF9BwRZXXyk/KW
BC5hr6J4oircZfkNSgAZ9+vc2h461C+EPdxdE4Om6yPSb2fZ+Q53TM6DLCr8zWjB
Av0aG2risrGjleD9RFKNgBCJof50A9nnYwOfnMg0BaCPO8vTKX/P/+De3G0Q7oAX
7MYhii2olRWVudTN3dRAyUkf99FRZzYhAFHjQ2YQk/zsGJW8Do+D9wf3azvAkPK9
lBr5lOTMko+THmCDfjt1548pNjDyViWL4tMx4TdcsG19i2ew73ykIK8exREM/i5E
V5Bex5oCYE/+7vDvofEEJ+KFFpseSGAy1oJvciU3f7OaJt4rruWYUafkj+pUCGQF
fMpHS6MzAG3IzNIyxxmwpfiIGs4dinALn9k1+AAYP1xFU7dAq7G7ksd5kC36c6/m
syKbqUNLjYLc2vLiBKMSg0Rgi/TQumTyl4qjdqDvpI12G6SvGTSv2nP8iEwtUvmo
BVT6S4vGBbYA0oDiWflCV1R5Mb7mWulQXPK/Vgsxa/32QZ0DrCU4UV8vyIEzh1+w
6Frs+0e/JKj0sDJcfyOfEM5XeM29JzZk2V1Zoi30PRzxW5f3XajCYrKck7kyhHK8
U6LzB4CroEe6StBZdOWa4a2eymCmyXOs3nM/qzpkSYLzkC6nDUmZ57nL2Ok3Q5FZ
0skrCqgP/HZo9XIhVNI/wOCBWuUXfuEs6mx/ZeyGZAoyIaqj+FJjidX9owZAsFoa
+HRPNTSI7BC9nFfFj4L/MW4zGuqLHK5+0G1BysyamvkfG455pYGy4gIpnMEOjIuz
7jQL5kq/BDUgwhwDsiNpT7JDOqnHOgltjjb0ApaH4HdJzsKORj8CcLUJxzTdbYsH
kuljNOp/bziQEPWXxNzjyuuXB+xcWcSo5rn1LxByFyGEYrYWUhhotfMfCkrPbbcB
xPjYrZGeyuMAu+FORKhkrffzh3RfAeYUIefPjkJXQCNXXkpq33xbhPd5KHjndmm0
aBk+tngkvKtTOwTfoVoex9rpYO9XSfKAjHQWPCMbfsEH2RkixvTWsSs7GCIwMQ2f
BRvfWW4bYWASqOccJDygXRaaqoko2SGc2MFjfePzDW97aLYox9S0rRlxScj/5Wlh
Vc4G5jlHZV4uhhXm2o/zwykTefbSiiw4FEkkGypqR1JiviBnet0WRUvkzOJtvdbi
ZveWgzCTLQxOAJLvCcW0oSs05G1Rr8Zk9x/SyhUjGp6YWTo/B7DDeeGvly/CmgUV
3CSKNT/fS6EwZAyft7PZKJOteFITxG4lZmIWUOlP6SVh1C7BQwcBN5+eo4RicQxG
JTdoFrahsZfcpJxwAFqQlAcBHYwakY3w1M5B6PAh8EPE7T5xVQQUaWhA6lK+D/O0
NRS0VkeAUP/Taipv2lUDLQiTAjGsXbKF5GXMkdFULrn3MYaO6bqZDKRkP9bkBnVP
pc63lV+rPhtDoNl80O7elvLgHEnYFzLC86Je4giW5dLP2r5TZR5vKda9Kc27wuDf
EvUlqMsM2vSATbZ2JSNdrwF1IHUUMtIOcbK/WUPWPRGdrGA1e0qo7YYUAEwBZ8j0
9pDeMAMVf6BWnB5DlvSQ7qNi6a7ViLv3KfyBaigvI1W68lqFMCVr0AyLbfVAUcFd
+Cg4FlFhwJxlly1l8rRyWcXCJgN2msUCdG1l9Q2ttvr3Y4Xs619QRVqSATYHuOs8
hzQMQYZt141IEwHKPR+5uxIG2URRsxa5mnkUqdiMgSZ32QWDrzzJo3BHDmXbpKiV
ma3sSHLbUX6CrqbPf5acsWLpKcDJewlL3pcHrRjqDJRu2vHEE46vv59RsSsGKLz4
q9nztr2PJ2QMk0FJFvN7//kRIkX4SWESQJ2jf0tbyzaN/aEgKs23n0rMxz9UXR9t
0+a5iXpNKXyR1BlbGHZ8PAu0mCDpDDqnh2THVEEC/k9bbrx+qP/Ye8JYQZPdWQoA
ow5aa9ULd7wR+l4hKGWRd+ocA6N9tfsal94xTUKTepceGx2siL8NKzcyi4STuxxG
50i+dRU1JNfE3rEUh7bw5A/ZfsfziepqQgxEUJXfK88KZhJYT9R5xa9MSagxRqzS
q1c/PfcmN6qPvSGke8W1LzgQI+bvobg8f3+IgyG2YqL6XgMC8seEeVJ/ANilzQcm
t6I1Vbzg8iIkgni5376V7A4HZEd3xhE75xakkAdXC1WCMSJZ90J8xEWcNzO9RYaM
QTM/SjQwyiNI2EpH/zxM8K4NrsHcDYhWtCUhdqcX3FwbLkpAAPt+khCecmVMFWf1
/N0uks4yG2NhtLqc7dpBkKZsjvVI7HWRdFt1xioXPSjHT6VxItBgWh73uabrrjyW
s5Lc594L4MZ0zsQg3CqZaw92Gc5qI1t4mhvCqM+gCprDuE3GvLVsYqJ3FxZVoRz5
KYstyt7eKNVB0eY5M+hroA==
`protect END_PROTECTED
