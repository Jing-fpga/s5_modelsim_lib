`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W8JO/3KN3Z9GkBlqcqe682IFfHOA5qD54IRFs4uBxpg3JDQBLmWGle4Qx9BtBe0j
PoPpPJ95XdUjCuTT3u0StbLk4lzHIW89IHa/DeGTi7berA2dWkLzraE5GRqreY/B
5Etaal2l9NhTcOCv5hbBPHrIUbP036IH12iMKL7bMjZ4ZXq2ayobGe9nNXdky9Yg
hkIpqK24Z/U2J5/CdwjTQB1KA2rPQOfTMLGEyjaptM2/jYY5b82rgmSsn1uopjHt
c6w9XiuUgSyzwTKzgRS6Jz60y+kqZe3UvoRb26z/CYrNg22bO7xcabR36gfXdB14
EPgdeSuc2/zTB8sBK2JW4ZfLnvYR7lkSbaf/bTcAIKl6F2etaQOv2qzqbj+IhR41
6ZDbhVOE9kBs8JaClLs4jqTeBv4ejdY5fi1ZHOFE2/49KVryDdHBfleL3xLIOeOU
9EdVDPvShyBKMh9AnZ/LdQzI78R2r671LqyODlZD7XOcy6DbkbiM3PvH6SSQOfIl
mwuJmr57KD/bSKiZqu2wdUPIoGFTGcs0hsmGaY3EBWmtqOd9ohBe09Tx+0lIeB42
u2aPOeqOunD4QVUjEJ8g+SFKOeC+mXLVGcfsD4DR474xPd25nCL3nsMnT6sKREj4
xpKEr7v8AE0EptCnE83S0VB/kuYOr+88hbrs2YxE6q8DCoxYMkTF1r9gaKAW2CTg
eRZ6OuKubQ2+StSriSxqp5GBPI/AlNIMkrN4D1vZKCjN4K2SMnB5ZD/+55JEJO59
WDKAw6OYuw9V3AoQGcXHiGmML0pDIQKTTa509+RX8s09nwsOSr0MnYpuR3ZmUZgB
bCbvGx8HpoDGfsHG92+eZQhuVcSDydf34qD6W8q/qfORy+B47/4uUtP3pV4nBQap
qXhMa0TLy1yUSmbYKRthZoY29XHqRqqREvNgUrGsDpEsqwEFZti/v8fCBRCmiRTW
eC6hX4NQtfz6x+ixqk9z0NmctQtHTlmko24ERqbXEnou20SDx+9TtCzHIMQLpf4y
F2vXgAvUrgL6vtLVktPxCBBNxG9tXQxlkmwj21+q3mrc9bJEtuNhwN+TVBfzGiYY
yr0RaiEijsNQv5n5qzU7ANu1JxPW7sZzS/Ifq1Ou8ZANEyESX/yvCug0wxD+Ask8
CTzXg2Ly2pyjxB7Ik7RB58L+luc0Ityy51QmXavROvaplp4jH8N48wb+fCxEqZVW
aVQ8HibJW8lnTeS4j9wXcdPykJpW9Mmv7ls70MR1UK/xsKhUejxFV0m3DPh1f3th
Woehpnb9d/87veSUHAbTXsEV933HDUHGKsT+HRwqtRJTZGWJPtd3zBJGxDKFTFL7
NhVe1bonR53SHg2z2Di635qOqa0ANferKFdI2GbHP7NjahY5YSCAFZZ5i15Tz//w
m7xGtPlD4jey3kJ99VzgD7IrYkFfysDQ0gi1rLL/CkFFiq2F0gXASzCr5za566GG
`protect END_PROTECTED
