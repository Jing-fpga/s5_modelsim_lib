`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UlaN06EqV53cXnV/de0+B3Y4XHYnw4M64o0usJ6fv52d0uGgj/5Wf2PsebB1gGdq
KyA8OFNIOfOcPzcZ0GWnAx811T/tJIgnuJozEhROL0NR1nbIpEM9FCtFsUCvzNEl
5Nb3tPxmK3OOYPtlMC2lpE8z0lW37eDxcdo5ngks6e88DhxEo6jqFsqNSI72E3kM
+a7fni3SVX0g2xfvHrAH1PhdFtQxivFjy8rmBIZidobZD82cikW6uELng2kIhl9N
x+mdd0V6JKdEdI+DBdbeQNsZcZCe6ux0Bhya9L1xgnbIgBoiXweKsS9l/pA/mjXj
WsTLQ9mjt/8irDIZUGFfyw1zxtrN8DImD7R3RpEV6s8HV5wErz1htSHQkQ8XjiZL
YRhKrgTiP+G++md4fy/sOvmW3pkyALe6Kkzg7H7+oj3W9n4PSjX6vqMThQ6jOlWo
TdQbzdWXXUdbEuxIxHDSJacjajj2slzdjBQwb3f3NzNz4r/BaAFAqTtfqaDj9+ew
uNhIm/Uj9E9CWfFSThBZ9gjSHDnF2Vc1sLJCSKz+GNfuozY+FKUxtq/qw+pLcznH
WnnCeaeVYzuQwQc/CAhI4/kvz6/i4gB7ms7z6j1aC3p96zRGMqHMOp3YOaLCz1UI
6SUw6n7btHEB2GymqvA/NDVDjZyHD8GBLBg5uTIg7yV2FRDLY0Km7l9Vy+QM7H0y
4CXkwLFosPHTLHVBYKDxt9d7RdQVVjptZwDwb0swk4rkv3o+eaw3dAGWTN5TtiZ3
E4bNf5/XmrZ4l0Aqtqb4yIbaZleCf8w1qJAeIWCGgAUv+s/HJF6l2X0KizOHk5/X
ZgQeQsht/YG79ydWj5QId3o/jvEst3nzo7DcaoJMawnBH+qhjA1Z8rqcsBPEYBDK
es2md82IHXcISjXfpOhLYwJgkqJMkyCj3HS8BQx5bj2VSMcOME9EEIon8+Tfs/3X
1adx+Y7HTYP68M3mbW6Imx4XdVbDfAWOFzfHMghlpV35ALvCEeisS64yrMjnJ8zo
Lf7cQ02wrUjggsiREiVcUH6dDkAYbQZGB/8o2yv3ZDR0X8TN8hsxOTTlMJd+wmQF
Y+7tUc5vhhN2PtHeQi/vEtuGkVx649eoNh1P+RcCox1+07vF8aS3Q7onWj01yUFG
ZiUXNy3QIWJQ/qKS1zAHaALOf7OfiPwhPcw30LsqTVV+StrIx/BwuM4KxV1zAQ8C
AmfbQ5GYkBr1gACZTx8KPche/+hjVWU+3wyDzFaS2AtwJr9YkVysb6ggMf1UsWpN
YOvzxYA9JPW7+iCOBwqGl5LS2fSTE1oK287LpMk2VVd9Y6ENc/4rTKkrWQk7S+wb
PVaoNwFczwpZ5Hjnj05GE9YOlCXJrdRhrt+apA5wByY42IfM5c6lhCT3BIbp8/BV
bYyHYKceEYv44cD3TjJs3rkDWdsQMeb2kIqu53LBtAyka8t3nTT6Vk8xRKvkOfNM
NhqtLWdK4Uw1CeGTwZoPqqYRKgTWkk+qVxdoL9WltlWeO9macUh7h2r3sUKe5K7a
dJyvWhYZvkCJLG6wdNfHUhWPwcjWbpEG/nkqrqsRThHcywGQk3NGQWH4jDenkcov
BjEiqutdUaRISYs5Z88GoG5FKzH9tfTFM5GDyL0BXG2eH/F/wBYD9XRsykfhtcog
9L+f4UK76d2SRXukqETGBUM75+KwG94/ZWzTzWAlCGErQJ5K1Bv7NY8Mi9gYQhRd
Eah7mwmYU7AFZe3bMj0AVJJKbeoEBgoKceL1SLBF4FdhaCmKtuDcb7/6dB7T6FhZ
ldOagyEcPSUZFhoimWz3bfkTP/OrCPjywDddHTxyxoY6H3A9vSzUQWYIfPuFQeEa
12mRJlmcHvkl1++BX0TPUnJ8XhIhtiz7h847XeDBswznb9WqZRPWmy9E/sPTrf/X
7h/Qomb1iwc2EhV1t3wp3oWgJ8rylVIGWuA11pbV8p1A8OjbPuRPuMPrCZGFpIcZ
llINxTrXF9U2webN4hBpR4a0WQdSFPQPnDYfByWXGv8avJqfy7fL9FvmW8xfd4z6
1HEZk/iCnuoYzZuERlj4LE+ItZ33RlEkST5CyIJxGJUUbTuN52wiQ1PWBRckwOmH
Y0zZEVdnazbXhR1tQ/PfEpTdh7bXWXWQwQ40g7f8qQm/cYHGVx+NZJS4MHy7BnI1
ix758rTLgA7Rmpx1y8bwzieUBlHeKvKl4oT+6UGXjqJNuuampUCYO64I73TaK8LW
R1P8rhYztLwUPQ+tPwqh3ZT4WhcvrqCfLbmodOEd/rWlRYomnbj+OeGQMGIj+Dgb
sjMUb4yGqgkcNubUqaLlH0yVotH77WQvJnLhT3jWCgT6pkMra+wdijnq9E2OH60z
02+80LkkDk0YqY56odfxYxHPgmS70qSx7H/o7GDkyY/vR75lownva5n5ZkTyEQQE
cyj16+PAVoQLFnP9DucaLrMDnry9bHLYAzYDxXKZbJ8AK5b5xgGdcUM0Fv5Q68GN
huctxSjyxL1ZejIZsx12L3HRp61E45QOjJXAYyFAzUJZ1TrLxEAiyUFJ10utiHby
J+R+JE8nLs89n1JkaUkaiRJlUZesDhySUZ6G6cMS/DrH2uFibDIPskvYUew7KSxS
yr/8CTr//Ug/Gmvncme2267xdmql3NJx4zyCKdDa9t+L+Uiwe3lZ7XJQ8AdG0JhG
yJvVeT3qC3glkODS0WaCyWjZ9m7KLR3r6vzuMzU8LfYMtHCIpOr++hLRh/insI9e
hbco30gYic1RCz2J70qlbb7kKLvNVqi9Me25JV19k/m0ntf1iMVTp/BukYwRQ7to
IVM7BW1MzLuBJ+ytVlAbr/O87fvZRcVWAjYrBR1z7ULn5Czo/ylUVkOAq61r8XxL
apEHiOxhqNEkG1xjsC4IjQF1CIlKLWXjMlGBjISIUTBiP/I0tM0HGJr1LwuNodL+
dE4ycn9C85aaQa+jE+1ra08wbMM+b8i/obnltahlWnc4SzV6ObWz3tCzbvqN45tv
kBEbKp8jv9sLzuHMEif/P0fnlAIHgLnew3yIVD3qC66JhGf87jLRJtED03hxpz/m
psNfDSjC4GXRc8UcaSilxyXBxQwflyzXmz0YhDKpXVB9w2ld74RE3XRxQV7UbhGt
dLdgVcV4KBWuuWi4/HFg7UJJIDDin5v2KrmOHTtbY/NRBo/xkPytb2KAMEseCS3G
wgbVRZ2kQFrPSaaMLsphYdyumvbJzzIUA6/njqGz7D0k7xFtqYJprPrjiBb2TCOR
JX9xFARkiFZ/9bOPD1s2Tkx1cgOvlcWArispZV7ICY6JSi0IwxIKiq+syHtZh0om
SmrcvVLGmGEz5GxuJ5B6cqBs2AqDveOueDpMSnWJAIbwlfXAK/R6gZHOnYRDNrN3
FBoH8S5wg0Qq/1qj0an9fcQgaC+Zw4aNoNfDwxOd9S3EJu9gTdjWySgxajS7YYM5
t+V7ycyLzI/pxC0cfzHyVA==
`protect END_PROTECTED
