`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7CMy+kanytfMBiysbb3bqisSloYhlff/sPUiAwHD5rvbW50h5H9j3vFY2c6onbX+
T72/Nk0By1ramp3iCuTNBlvQQiK/bU8P8yfiSHF72rkilNObP7PJq1ZT6cFrJ/2j
GsFBwRleWg+sicVKAR1sxDwDwKdrbvxppcCTUf6eOc5egg5mfE1wDDNZQSlLmmT3
wDOYVLzuZl+HNXylbh21OeQWupFbJf5ltfVfQLDMJMWFyxECwdGGVx5GYmq4B4dK
9vJMVp0t7ABlUG8GOF/rdu+4rT5a0vOdeme6eimA8rO6g1CIFkD0IREbJXA+bnOa
QlDw3PQCG7clf5u/0/4YJlv1DcAabTds6bTFGHCv/Vg/m7UNvMop6iXeLLXu4UET
vgxoWEi5SRGPzBCJ5KfiFkJUcWR3lDYAx88zkiMCqqUcD76ZAvrGh8NWDMsJYqS7
TYyhbBrj4YnZ2tKJnFkwBfyvGuXefsx1YqgL6nTzKd35OfVTqPviPmdwnZ/ztX66
1BqGq/OCgJypMuImkwffsMqn/xsQVrsPkHd2CWG/ThlIQdQR9LNeXBCQsn90wKIZ
w/twEnPVmyhXfgvIph5+ucw3e+/r6E8mKrib5Q6M00600cShHxIOX/m7SZS+Ih3k
QORJRJ3+c4Jyvxe9TteyqpHxGWfUhYfKqyBplehUHg8pzntnfU4iRaSRByfWxwiZ
gn8afBzmXbN5bCrWJPhQveydBn+gxUPDXjZHAOksmXMQdEDwNy8WUyEI3DyVk38P
fy3XBodhSshhSdtJtN+F3gBDGn/m4FYWElod8kqxbLeLh5kvZNqgNNC0dRqZrNlf
C2M+OfePWi0nlctEriMFeXf56/nLgpXoD1FeXV9JWtiYeuhLyJVccSmhz+RBirDZ
tgNaKNrNid8BsVbGzpgD5IGVdjndo7i01b1nYWmzPG0vUCCgq11KIeJgOuR0G39e
ItsHo4BBtRbp9oE5qP63MOxenjrPcZNJjsNc+X1lt1v5iFRCuH7/ilniI9naQnuG
ebW4xWVD+3huDyH2TmYQwn2EbhO5qbrD3QCWAhIJLrDKkjhB+OD9CktKx0XuHrkk
j9dpfGLa66QRsuIzleDIB/hBmhiElVLeEFuUsREdy0iAvLARq58Y5YzLK30+k9Vy
Ea6TKze2Sf/twhhw1NDDTIU47pPAwGptG+php6HBCDg9skPGODzenFza1oLrj4dG
jumXqGyztlexAVLBIAf5MhQq8QCAZHmM+640QUnNdXLQvBCygCuqpaEGqb0yJljv
GUpFNPjYy1KuZj0b5mGuif2yHCs82vbSOUrk8klN4uGWiETEaBtlbt3M3MeTu6it
TZXNpbCepLHywu7GicMmhNJ0GrKSLfhxaw53gzYGBYAzjcIgx4pbdNCdYow27s3W
ozK/uutMue7BZl7+dRo1tO3zwN6vCA/XdbtgyXZedHLQL5/jPbz4hQzZ1keU3fcR
jY/cCqhzEbmlLqE3FIVUJPaDEkVo3WfKD5hkR4178NYukwnG5apBA9dZZQftKLR3
E+wacttzfZBIckknOsXUc9lpkDfJlnOvOBf8dBlqjpRiSpUlvQTCnk2zNVxhz/Zs
qCDYz2yFvAZpNx8Udxgbe0GHzmUpA5/a7ExfLrDCwDDX3IvfIZ6DEZ06eJ8lhLxB
+7R4zYxCv/UxP7OSeIocdvlIfJUlbaiiQtKP4S8yzk06FdUOTpPjVPQ+6pyrVu/k
`protect END_PROTECTED
