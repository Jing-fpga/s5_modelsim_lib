`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AYp6N6SYbjPeqf0jkxlpNE/WG4xOKn05EgbdOvFHa039DXEdaRI87/rNvtg8dGNf
xIkYzAjmMtSiCH9lGj6hS27gxd0DGb3Lo9JawjKKriIYb6upCXewhPmFM4CW7BDy
chyQRbmpzU9kmkhgnqCAL8oCFTg2kn2bqpZ/1wLE29lG9GeJ5uiclsWeMFbmduHH
izCIxfamGRktaHP9cfz4QHf/gD0Xy0hP1VrcnhbY1SwOWJxiJzYGtj2fcDslC+Pu
CisawxGPX6vPesk8zJXtpFZ5AERRT/TqcMmnenICXaCKyD+AFlUE4lSGYiENn5DL
q//uoeum/+Xnz344wD8GjJiEb/oue4lyHMRcuZjLBUYKiXVvvkk3K/EF89RVWnlz
kOsYG9YvxG5lKwXTVYo57FA+8LSudDGqLEl5xpHxdk9EE4vmdG1GtzSwecepc0uW
uJEvQ0y4m37+/c2fwFMVcgMpE6SpZDgSsnUuzx1wTEfq8jPiyHnyNnQWWAhF4Mmd
RClhc3xfSON0EfE2p/wMlKUYnDcSPHKVD41ttAL9Zh8lp9+KP50pmMuztgANJE12
06ZKW/p7mSgGELbFHzWXvM4i8oiZJ5Bx9VmxrBBL49qZ+rLSRT7qZYwy/DkNP0YH
IYrmbX5mAnj3Ei1+VN6hsReVqTugMhKqodQ9zOIVFcwiGClcCM4Q2xVUcU1VAOsz
FWfQpJWpN+4YS4giv4XFw+kflbnm71aY1mBhOaRiUQvhSe0fOskbX21FyQI0xjdB
Ii+bheS6th8qlqZSYnjsQnnRAcXOslKFz8pf+P+9PV3UrbrIigXUWDnUnqjlVNSj
D6TtpOmyXrcUrl0SvNkh2I65HAkg0H1eUlHh7nGlRyBhnoB+Q8YoEDdqM49kpzx3
11+QXmy2nITenT6Leef1R/XCp6MiFW/Zez6yopW1cAp76Iiuml5ibqzBlhAjj4FJ
ziyk2M0i9sGF2IzwuFSHOhhmDoCAiJh7eE8l6FtNBkFcBgEKB6nGAJe48bX4rC6J
ZN9x2j8NjS8XDvD/FgRhtCLQTdvhA6mR0UoEBaXtYhlcLCAVVvuEUwFvorq0ferA
4tHLPZz/WDZlRlQuhQqZpb/LzMKX5nb35EFXWQ/4C9A6GdOdKPlFBay+XPPRPkng
Vv8zobbbsbkJa3gaD1WapEqF1r6w9STynMdJ/mAvTngVO0IDlX4ibJgQGJ68HbAg
ZzylzxVzmc4V8b0cSaysZ32WMmv3WhLnk3jpkIBFzMGJkmhEGHi6Px3wWATHLk8q
`protect END_PROTECTED
