`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mn/LO13iusCqkwUaqoRbw44Z1NWRN5n2WU8oSZy9dHcgV+lbiZnHPB6hRcJcl8S4
pyiGR3zzYFJAyIyEpozZ8AC3jef9C3siq+jpg2ZHqMkW0EGskdhzPmeeDCU/rBxH
hHIJNs6RlvMwx6yXPJCC0q37YNXvg4nhJx+1k+KW+6URTVUtQgzz39S1AIhD+1V+
uBV4CDk0v4LZHOsm5R7/t1FeAScu8D6eRZsRej+9QXA4WNsTfxQDSCNFupzeVGUG
fPHwFBsnv/w0C3BXqRVkBgu2OuSSl7+gylW5KkyxKPShTE3WSiYs1MxpmBLCj6V3
ZADW4gdbmTfOrpzaXPVZOyTqbkdAgBYMRyEAfVIazxsw8IZsapPAit2uUge54l/T
1pTCzcNLRjBSE41sjMRmeLBKrJMDmOi70D8Xq6KfSpzhzoqCmTDduaSDoyoDjTYZ
Yft+4C/kYxKNOpvdnTaoxa8++SuDM0yvJYGSnPJytmkpHzY/GpuoWNgidwcIjoVx
JqZ+uTyY0xMlBVbxziZ+J9M4NGh3Fwf35mgRhzA7jKCiIOJl9+rcXAbh0Rmlsd3H
VgOrr7vN28P2VThq27Y3OTfSJGLO9Uc8OZ1wjXIehQB/+KZaZLlAZk0U8og0zZs7
Pw8uRBWSE3VwPR4tMzt97gpStnyEo/FE9nb/28UcmHReUMzJihD2yQUyuYcnnpri
VbOLk12qxq7H1Yy79XB5eLCyZr/VFoRi6nLwThuuKBZsVNJrCR/0OeqQxQ2LtWbg
XpiMRwD1T/49wbJVURAysyKJtT8d4hByVRik3VxTwN0Fs38ZqndDMEpcDYY8iXwh
GuqOoOuy+NnEFakWO7qGxpBnkiueMrlWdJjme7R6kIDmxMYgw90UbLU278XhX3BW
AfN0xXoaXJOyW03Nsqkqs26QAgfzgz5j8bLp8XAYN2cHeaPQTyLi4bOthgVL8IkN
q4VScsSaHQNnIp0r6HItiJPi0mt+Jw7AFrZDNDMgWDY47wVBTJb/B3XEg0e6TY5U
lt0k4ld0ehbM7TBYs/0y/8aRPxVdZllOA+P0+VWh6GrO9UChcKUdJR6DSpZoUH2f
uW39W3LVkMzSxUX/ZNHhnXSD0X08bBQuRpo8TviB4zLWqZyD0x/TpJ2DyJ8mynNl
nHYMwxGZGsU7l6fx33+IFPlizlXCIui4wpbj67nSonjwMUUFa49Dx6OtDjN9bGMv
yQFMtDuoJwwPTOmUPs3XTX1Ntmpm2FyzhynOJNtrzZN90P5p+ef+GF9JWfM2QlQJ
a+EQTxym/gHOxSgRC199ozWONTmI6L831jzvPBo0D2DNtvaavgD2E5nSCImRLjrn
A8y4jiuzGoOO5ksoxiXNBAr83D4nz7EGWyoweuVSKOnjbJxiU8H2fjlSVSEQW2z6
eKeRY7yai6mKhL/NiMjcyplYskYBfQX0m62SuMD6GdD7Eq3WJrMCt3oh7iT7paUE
/hkJNvKMkzHgqBBN70bYXjJ3GpZogV2nMIXjD8qSyLCkURn8pKEt5ldpZiH0Avt/
ycRWM4bMO0Jr+VO8p4HRVDQNTSdDj/Fy2zSSIOpdXV7gk7irlR6i7pvGcD3/iEmR
E06dAmqtwC27NyFVPb7BYNUlb+GceYgxrKfNY30JO8uQYeJgwC+VcbE5LslkP9S+
0HJ5kRFv7Zmx2it9JF6vqSnHZeP2i423UTXq46oyv4UHvpZcQUTvbB/DEVD6mdXI
cNds8X1ErcvWQAMhxFigD1fFUQFb085+RTlLc0elVLFvD/ompFsffK8vFy8JMxKA
PfmmJpe1DwEiHEg8mnS4OF55E0E+zrzU3aW7BFyNQrWayOh8dbUPHGQNa3QNJTOx
e0//lsAEVpYPrd+81YOALHlP9y28YpbVJjUxWibGkRLgN3zt7QPwvtjd8rDI1jAC
1WUGnHU0J/2gTkBzUcdw3PFI+R1Ud9TeI8qfMiSxqGo38Et9uZnRoK1T95sSzxPe
Xyxbt4O6gdQmnALyE9nBJuXhpeKEup/ejeVclHHfeTgfLgiLfH8fXvBuINF7WvCo
Fo3a787SMnpBkGHedQM2KLv8h75bk5j0vJhb4udsU4rkJdCZhHkJgrufArbOHq6i
TMuvW/tS5sWTu0F2Wq0ZPGPIv+ymydEu6WDPTtIRsr0AmGdHO20XVJsBHaHwGVHC
BaVKP6QkYuNARqzaQFt4cSNnLrlidJL9buOaVpkRsU/Feaq3HlrloJv8umhImLTS
nwkK9qR3LiM+liJYUBVtwWrWY7ZIiX9mazfM1Ru+QSwV/Yl5rXrMJDKo+eWAr4yB
`protect END_PROTECTED
