`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OC/xqNbXgekTlP4e4haquiHbsFMn8P/RDhtlVOyIIML15eHC005NuJURaPcGDr/P
2goOwZq8RM/R1Z0XoDmLPDbit9Cz4nSLqi8AVY0qiBGsKoMUSmTLxhhuHrqG9DmR
kpEgyHO8PUPjOPswqYF5C+t2PyiAH7YGNIalBzS1w98t4/xnXAVGPeXSwbmiiSCs
yz84OyZpTHSwrndZ1ymikf5xBjSCMliYtuL5aQDxzMQtrW/ZVX2h/Wmo6sh6rOJm
3v84L11FTkLRJMDKAF3LWW7E13hs3m3oMAK87rE8q6edbOqKRytMbw2vhppBseu2
ylzUr4MyoCSBDMVfUHa64jCYNmcrsjYjGW90JtHHDR4wBqhyfro7cZwssg02Xw3u
yQrKKlWwU11bM76lJE9vSIt6++N1EYrICTtEugpAhCHg9QJZ2m5R6I4B8A/Bl/JY
RVLJucFtsiY4puys7EJPy72Gold1FcZBTJmOqSsP2gh0t2eZu/XTsjhPxdD4o1DA
hj3HO9ZNxCJWlUoL1uRxfMJe/MpGG+9xwpmtsoCY+DDufMeRuS0OCy+M5c88AGvH
n6HTu5u8WDow2iZSkHdzFHsdJ6TtjoFjOWl/OH3ZsmWj9ZFWZg8nmgwHLdeyIZxt
Qy/76BnP4xhA//KF4iVZNE9R+EAsHrguhcmlLcm4yB/V5Ugjn3AJ05f0CRUG+nZH
aLd2oajewOaoKZOaNCWJMfRz4p4wrbax8Vq2nvAa0Vb7dZPBdEh1zRWkW3Rz+CSG
1HJ8S2wXd9IF6I59k9xXeUAOO648E3B9QiwbkbCjvhYJR0E8bzcTAiMbp4K0n4i4
DvkGdHA299B3Xq891/gcR4JHZDY/aN16MhWQht3+Hf63wF/0+pnZqouzkqQ3At6I
h7Lgutf4CSw5gshwwUev1rQRVPU4i1BU1MCJtxBCm1M82XUqwK+qFKAcqIKudhB7
P3CSB1JlSl4pXD4ewx70M3vzwZ/4N0ng5NR9Hl0NaISmeZIhtcO1adUHwzc1xJR7
HVQODVnPABBwosYZI7it2+g4E+Vu/HoiagmV5IpAzbZu1AK8JKGo6bjc97QnKn0b
BA/0Pr1ynMI/TUIhZU22Qq28/dle3FvrWLpyvAIoQG/rwF7NIga3bOfbN+PPapSk
RWB1tflOHKji3yXRAWkmec/a8FuX58Tv4lIJRV/MimtFitFIeDqvyALcFVBwIqxK
nu8FmPluMxkLxiiJFQM9ZwTzw1JWQxLdq4rWaBbT+c/94sKVVC1+NJIJ6BTHwLo4
NKPEFeuMwzDTnPecL//SJdELF9xrtuV6/QYVbKs6wyPdzcIIOdiygY688mj0v+uF
HxlwJc9qCjVLYbNYzHEjsDE7fgAo/XA9itVBK/7MPbhS9OFEKJd40UcmO9IhWT42
fhutv1oi1YD3P35oI22SZCj3O9EW4X1Zsp7B6qJbCE42UC7h0rgTo3QJNhcuZavl
u8WxYxGV7eT4oN8+uwbNbsL6Xj/X9C1QbeU5Z82qoGrR7Ltw5tH11yOLJy4Rkx5T
sbdVFeq3C0emMtRUyDDRh6px0sSpkbOYOjcdy+D5siYCgI0/Gjz6IIWaiFdZKPVX
VOlH5V2znveDCLTwb7OvoGQiz0Yl23iFeuxklDmYl66I9fV85QZZRSHtGitldeAc
nU+TTlMvc6BRmCJ9TsqCDObmgtK05S419Haptj8a22teM7oVyoPRh6A+F+0+3CvN
nBycqHRxiuIVoH+XBsu4VmGFxva9S+X6Ra1vSRqQ353YUiPNRanPgpJ/92g2lgz7
5LXfaO/IM7z74DiD7XZPqQ==
`protect END_PROTECTED
