`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cQijEx6ct44Y4khvOM2tSuIEAZlsCVJfiCGxZQtCuLiAKp71jEZNIyW+Khqd+6+b
1g0+9m2CPafDRLuNrmnAB5S596mD8gSHUQfXuvQi0vNT4L+u55dh9vqREadbVRj2
Bu+vMJZ21kVftrJ7UtmRQSqNn5Ydy/hyM23mhVSzykgSzhfN/sdA3cCeYC13CWDe
91ChGCv0EUVWdJQyp+23YNdBKjFjNBcsBOoWDy+bqaFrYmRtiOud77qaA9PWE+T9
RUi5eR49g3uiSN+gIFow2LUGY86cWBJdGqCifCMiZeedGHKHW/OCIHDETlOhmruc
n9a3Mc/poSQfw+8ejpZx0fePs/ii8/99nB5QlMPKYCo1iIMy/eZxRlbLPtxSP9DX
lTSOrYn+lF5nHkzmACCodAuT5XC2f+OI+DfDYXzkbPBH3I30r3CRuh6IVnTG6Z3R
QJQQu85tujNavALpB8WJWxmhx4/gURUOyy2pr6oWDN7j06yOlRG3ox+5KZyTTHI4
aXNopneEEI92uqCrz8Slw1JBgtBikUCCM9qozx/4cyZMvVUdia3hZFIW4M5iSr/D
uufUxBK4YxHHGFjTV7S2effMJRZX+oLkLX6li9ABSjhTOF0fv/1GsLCa76bLlP29
1qM/89xdv5RSByqoHn8wPwDGynRW8nPRbxfjlUb+UyuJTLVZbkpl+hbSuUMcb7Jy
fO6nw1iTSnHkQBubNW97H56QO4jZq1vErLX5p9jFjgSvJC57dYH3WB1ibCVOab4U
CVZdc5sm+UeCwtm8TMQ+/p5sFFxEZB+pVHZ91Iwxd8LKs814FasmxNfJsiTZJ3NU
VgJ+UnCvg01EpW7NgLI7y2pBZf/HOT4tp4xsTcEe/PMow1HzHbqq6xsHMu3ds9Yw
boss02t1IoG5zFm5a+LaZjhD5mkS8/F8Fs9kwW6rR20hoyuoXIPWePvn1zorR1Iu
WJqYWFPvfr1OvqSd20y+HuGKDDWQieL1GtGNoexn2xMIn+xSyzTwG4N4Wbzmt/v6
ZymHt1851fZs7+QzPTDtdY+Dwz4FDNCvjfQE82MHSXX7sutDxvhHQL99W1StdIjv
d9d/n/3HAldeKbggy1j49wZvvy68XHxDdTfrOOkTurB0TUm8NokrbrN6wJk8OaOF
W6zgjnFNHuTnrztwcpeRflXcrzgDzQPJterxNRgqq3biU+Wk/ixDG/nPiU7KonBD
Waw01TjbgbI/C87BF9XoXxrqnq48C/I6l3UJmzmQ+sg4tvi78Q15q7aRKn0ilp7/
GKd9DxiadLhv2dPtxQhIU8o4obSHeBmpKH9ZGUuLAgknqCQ5y7nwV/N5tdSD6dgX
+iBPoTh9WFlrRTOOvbJxM1+7S3GOg8rTH0muG5gLKveHpbPb8NCn4JGXTmxi4toV
sp5C1V9FXx3bdMUUh4M9iiXstPdPGHQtv4NW02LPZjkRdDC0Ax8mkIBMGG4phtgq
v626+/Oq0m5//Sii/otehsx0z08PPMx/5dkjJeC3Y+zm9vUFusTKdL8uaj3qviaV
au1f/bWP/bOmNsHBeB6hfJtVacjHQ5m6RdQgOScX1UztLYmUgIQIv///NjnIQ4lY
KDcTSmhCC3/Zv+31r0OEqbYLx5dHwyvu533hOWYwsPYEWiWDzK9GTGZ07IPcaqSC
CFall4SlDnvLL19wHOSU7DTwQ0u6ii1zUaZri/ZpwqhQut/A71LTUU5ui13jcUEd
seDgaoJvea5zB+l1llvwGL3asr2m5NQud9ILlB9irkCCJ5c0/u2LqRGXnQ7IWpfU
kxJGTXpo3viGWtaySQDaCLlkI+t72xFQ21Q8IgaK7iZeGtgonqMOb8AegBZQBsoJ
AzHZZ+D09G8nMQgdFcljxAvgS1RGntd4iX3Mf5U5Xw9h6olMDh7nRp9vMFOqFirJ
P8xJsJfyMecXdWcbgZoGFmUWNxFtru25XJq3iaOldb5VKDgNCSo4qPmZUjNn3yCy
m7Fdi8UvSuQuUVL8dA5aR/CE2lBNHEzljnoWgQdio+RzzjRnBO7//E/Ys5FRZs/P
vs7l026w6LGqicqNCM8h8gzL+GcinVs+zXdKn8lf5WgiFSeHGfLVd6SQunN7IZ1w
UDzndFsrqqV3MWWa7pCYZlDlfNmCmminjtXjW4j6Yt5xBOxWVekflKE4GgrVsGbU
2K0m0KWCkU1xguM2Up5WNmcHZkBqIpdpMfk5WyUP1CMiT2/wWYUwHpaaKK/p5HhS
9VvUguRt/D4ia1GkapWQHLgGAsmnOtLTjXLu7hkwqV+sedRnqD74Acn/5tGL4lT/
5N2hSkJEJ02JVY/jH7MUrT9J+Zdb6hOmUeY4AVE9PTftO968B+ix9S5mR+lm0Sd1
yEDzJe0XS9H+7l8oIrMAHIAKG2QOz+xi/niFg0U0DY3QDVbjPaF2IFU+20uJemah
CvFEydd2sYlYaTS21GeiowCahJRD3C1yfxX8ZPMsCvAu8MvLRhTC1cF0x2gsJe/P
CekmY/JPPJsZwuolfSGQq+nOghCPI7HOkMBIf5uNy9cMfsH2jE96Cl94qD4nuEK4
/PGBWjPPAhkhRIxjylRkWxvYVhwz+k1fzh5pWjUyxMTtp7FD5uukOtZbu/uEM3bI
x5C4+q9Ne7DpaZWigCE0ftVQaRnzMq/iA2BvnJaaqNe8cufS+SBjjIcKe/rTYEdm
dz6QNMN2cILmyaSYvtLYExFNJ2LEW+8R+oK6AauoHE8ZVB5VWCrLEpjz26hltqEe
JNtHxi/1QCYe2FtOVTwm1uAXR9SRm5L3RvVGIpNaY+dpVUPOJnLv7b+zzEAlk7iJ
BvW16N4Wr3DBw9f7OCTgTruIYjr8GYk9mY0xAGhy9WX3SaKtK1okwfYzsYy7AqW+
xOoVgls0FibOHxfm8+NdbY+UzpIEyB3/Dnw3kBDgMmSPquHbxv9jM1kNb69+bQOm
pkymi43V51w/1tYLZGdtAJ7W14NI1xnRsQXffdHXcFtz+OSKPOljtVwBtuw+Sg1F
zXRrF4fbGqoN+7ihyLkPIH8DvsSjQQhoX0PQvsfN7wr9xxtNwxt22WKaiOTSNG2k
9ygrE5jB1i1V329XWP/u6HOQdV9IstjA9Mrq+QS4zkpmEJyArrtMvZCeQA6dZtNJ
kcI/gr9dOFbHGzy2VpNlABawzbRFOKcJeROzRrI62TOz9+gHSyVbmrbj1dYLHIjh
qTv/TxYT5JERlSQssl+FDsHwyohPXZNm6kw297lyYY4vPCLSRXkQDvJoy0HtWAbY
HRcbzkO8OnJaNOY+vX9vROxRscEaPFxFypPawtSSkzu5j9abBr8hb//e/pmqrVaw
/LL7L2/Eq9LuSslaD6+UWjuW1aVVFe91QWnOflggatvIrnIuWdBHMXGcahbeyvB8
350Smdof7l+rB9LnoG9Z4sYg8xo7TATkHGgdGhY5G1ROxtknYVYOKw6WWJPpY3hK
5rEEU3Ryd11hcPKOSh1BrPSuXyRiwEvNXnyDfXBOV4vVyNFIqIdAn/QYZb9HDecT
tuLYQ15CZmbJboX2gPem5T3oC93VeHysK1UbFjatMKR3MY6c5XhW1dZvg3Hw5/A0
Ecd7gpyNa1+G6F82qylam9psog/lYvjE0/4Kk2ATCRuoBLVBppw+OXEXXQyaNBEN
xXEFVJ+cairX7f7Wu4g2DkBzqwiHDBVOgF6II24gTIXP+ktxgz8YYbDfv+In/E+m
Uic0xBhfdZJ8L231SyZAsvt/RqRCYRD4/7HH79cBgT7ubR7YzojulMCOmrS3mfZC
UGMZYq1CMtePjPoZ1fL16LFLJKcZadBdYzI837qbpdkWN1S9zcS0MgzmTruRmMs1
OAoUwqZhyxB/9e5tlBsfzw==
`protect END_PROTECTED
