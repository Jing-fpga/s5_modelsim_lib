`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YXwuUQr7YEWn3c7ilHiI2Mpvg/Q7YhxK7919WWLbuZZnGRNvxt2rxbAwhCcIboOF
VjAETsAxu39dOAXA8kB6PqLy2n0Box6/o25BxUFdusf5e7WVwkAz/5hhsryv9cvC
pQeHhCXZZHLgOO0uVq3H7ay3nXHcOr1sHu3rzwEpCcoF8rxlg5TlyXceth+wm8F1
Z5LlyebCi3lEbt1QanHO9jA67vq90JefAKUWHhJxkSANpYSKlRqHcGwCVvgYEIOO
35uYqbchqgy5W4wDSRr/tigc5KOZ1m/RhZH5d/1+A22alvHPEt5GFl5jeREO/by2
4/WWathxz821aywSeySYLtUsD62AA01VFGEH+tNn8QKbNK3PQgB15H6PkfvR8AyI
NEmoBvoyop1/qgPglJnAuIjSkjj4Y4mjb4eijBlnTZNbFW+s+FhS3Z0HzqRlS5ih
bdEWIpQ9gpMaD33fQtPrBUyGuWlTC6Ne95h+w/ucYUmvcjz+1CHlN5ZURcZHzJxn
z53AGDYqaQqQWflt1FX0EBkSCKgZp2h5M26rJSSIEEGWxM7c5Dc15XrugvjPJEcU
XzBJaNglGeVbojb5x6Man52Xn+WzszL35Gqglp5UrxHG40ICzgH/2huhsdJoOcYn
UALSsRdRZRxJU1aG1QlTDLGwRzteMspHwrLD/UVq9BdJ9yqj+ycu+8hWSCbiqWts
xqhaWXKaLzAb+mbubA3Xsh9pKfXkalXPdxxjfU03od6C+/5j9vt7M/kVw/hLxZcX
0QA22LUhcnhS2jcQSH6bSj79PrBKj8jtWMNfs6srukxIcDFAT4t2SZ20M6SYSWee
ow3Ab7/UGstNQ0u2QgASJUwoBSFdTmOjo3A+N2+uAUVGup0RlZeeam9rBZAHBY26
Ci2m6Usr6Z48u2Mzd7wyqEF5bRgQ3UviqG8A5PuS6sGUtoIDdv1kT7mjNqeSyZNo
40sTJEhqTZVkye15M8BZIYxu2DCX+/ysNeYlRzLb2s5SrBqTFkkWr8tnasRGVMUd
UqYzDhheScBDpE0Y/os8Np+O0KUfmOnySfdK3IwZrq1KMngrwhQyNxse4R2S8TBY
Ekg5VBe5U1phKwqBhVSz9buw95fOrqfEaKMJWCMRAYN67k2lHBBr8sHucbLAjZTL
et67DyK7epxBj/QRgp5cQN+rCCN0x8j09ACVHXIER4v/lwG2Hw8Wtgl8FhGVlImk
LRHT2XUlyGetYKMj/jEF/qgwi5xmoQFtWwJZWJtN41S3ABC/npbtELO6+sOnaorv
TYMOLVNuj8GyWOUIJCqXWMj3BfSEqN2IvWkQe+fRtctFLGBt+aQa97C1ckPN61wu
saqOJXvnULROz6UdMVvHjMqb14xPrUaRE0EB9eBbvd6kcJ9LnqmIG2FWxLyzFQe5
V4b9hN+pKUyzQyDlipYPqeA236kdfFfDPhOIvMqK2AKaM1JgVncg7IV5WhCYjNmF
bD6SHpDarAKGjoYTGnWnD4SjtVQwZN7VABa4+Aa//1ONtKGPsBjmGp3k2TL9R4zU
E0TIZNE48KGZ9n63O10HUyeNaPDrHjIb/y1fP/RR7YgajZVaJMpDUuvvCJY2wL8M
O7nAm4AWex3ZuQ5n31DROLGo9Z2M/INdSJ0i90kGCCIEv9jdKUCVeKNxg6G0W5Pc
M1N3xzgPm/rt9+/PbwRBpFZmQUL1k32Epur+ctn2sOny66lQnbB4RrHodAKlXJUx
Uk48VUjb7Eq0LkS0smyeFREMsywuMGfg3HzCvEUNfUsWMqYKbpQ9Q/FUl4M/fHvB
ZiJwYK20yVv6UmKJV+8DbbU0jkftOaIBk66lExa4StDdPxAVDNR7m6QlnHkDxJTA
cDEIPwJkdnz3WDjuKcSUbxz1bN6olBAlZYqaXm3mq0x0nml9lH9aNWOaMGK1oztj
Ur0R2FF143KySMVRdTEj8X3lyz7FzlNvjmwdLGbS6hb/oIeJZlPQ5dbSmwZ9MH0V
GfPTg9EMW5BAEZ0rhD1RhonYb0EWsJlTWcm8vJG2ID6qKu3Rjc/mFfk2PlHSnFkQ
+iijGsp6ouY0HJGorPDfGBOw/78EDk73wZ5zoKVb29089Jh50slLOdYkZPh2QqTC
Oeo932bzUjZa1SWux5x/LDVdoVZR4dBF/fzOWwdd1wc=
`protect END_PROTECTED
