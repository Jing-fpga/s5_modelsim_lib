`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B+uqcEsdDqYC9t04eKAZEilo4O7oYUqIhbdH75rmIpxYy+PmIFnlIWP0L6qJq/ke
WbjAfmmVEu5IlozBMxljLa7tUK0ap6sk/Q7FJ5syMv/I6XTvjrfQ12uRVR00P7GQ
AMfkRGe2eS2247ryUbSptI/Ihy9dRcRNIACKFXkkesN9xUsCtYO8uzjv7hCfgy6i
tRwXu9d/ALzSAU0htk+MkF0314kqIwh76GWB0fZkTq1jTtAhPnReSdtWGDMsUI3r
QuBdMB6nn6aD8Fjuk8m3EiPc4uN3hNQ1FsQRYzztO9aXRaQF80cZpvp0boKLHcHZ
PRnXNHaZn8T2qqmej69FBmHGha7jg/UyqSGjcaFbOpGKHumE6PkhJ946mq/XH+Pf
Xx/cYCmxDM+dDCoHIV1q93C4xQJ+MnVseKU9IoF33RS3lr85UWIZZYPNhqAgwTAW
+S1/DQZA1BoTux7cuNOQu8jP7jDGSqw4WTKXfFTVHTgL1d1esByXeaR0Sn/zXc0n
ZCAtb2THSf0aPfE46Ue9j7aYILvtBULpSwxIPcQfKgeYvzsbQtcFeTdqqS1VeU7N
eKq3ezCAnqsIZO8m1AQ8naBx20jCkStKaJgXFpaO6u8RJzoXvK3kZzYrG3hgTHSq
fyI8BSzuyTzD9xCD/KveZc6XPNLMDDpoch2SGfzWa3QO+a0EWq2suTfOHfhR9l13
9c259N/Bt5uxQcVvy3y5Q1s6XSbFLFgg+ex3X5MEw9Fs7NBNO8WppW5kUpV/q1PG
gKjrx7QT557ystoDgPn60A==
`protect END_PROTECTED
