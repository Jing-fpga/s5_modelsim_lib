`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MsSOfA9bCBOvjvjzrq6wvUWgJFzdh9v22JOJ9I8L+JR5/8O2VU0r45vef9h7tx56
YQ37XBp7I8zPKRSSeRDyDahycDESjF9bZWkE3UsENGx5S1NgKgg77B6WXxKXEtM7
s0LTgW5XOJafP84PDpXi2Ig4OtSYxel0XetdOa4SXvGklzh8Q5KFRR3ldbxO25QX
hfJVLyvy2Ojc5wDOylRbRBMBULDnd8GKX90weiacvW9jWilPAUQUo8cNowlcUt1m
qv487qrxhiJcaGyVnalhussu6EHAuNiNHc2fYBrcIvET59VKAc8/IBcI8XRqZ3ig
b6ij3bUborXrr4UiA3LpxARpf44GV4uKS2hf0jvN9UozRNARheIb6oxvhjKcgjhW
iAFpFl8zeYGjlt1bM3ts3ICHur2fa7XgyF/S6jcde5FkgDoavmZtUPnm5BrZT5k0
Vig1gtVntma8u5QUJBH388pWVSl5NC5vaSHN6ruOZT94RG7ubWcSBWJJKdgsfIuS
VCP/lvbgmOUdoE9eKMRwEHnCXnfsUaT0po7jDm7dMAFr8Zem0+WlVghPrvUo0IPc
eB+XPDhkWmdM3Nl/3wyoXz2UhIYtnCVFMpp7ZnUdD2jmRJdZHoOQ56GRqLlFxDeR
FJQNGvsOo/P1Uzzo26SxGReV6bq5TPRCoTbIejG7hRz4fqmtw5Tc6ZPs5XMEGTuZ
OQmfNHwxCJcXLizMdPRnR6+7gaeKdgDI8NpMB6l4EmTpMZWFne4+nq1UbDSIvNDC
gb5GaFbC38dIsTX7T3z6IcEWBu072x5naHXSeNcJkzxu+pZwIWZcgFd97DDe++BH
pfOsMFWST7qQUrZbeSNMkUE4eXsAeE1OwKTRTHchXzRBwW9g4wK/4N9dm1EGJfVV
mx4UNs/L1CpY36P/6sSHZOk0jBgoBaW0vC6ys63KeUiM5WuFjM8nTEpeis+HiMK5
VlLqt3DaBg3Q6NkkY+B+soJv7ZhQJx4TVJGPEB9V7JvHfHXF/lpGPnhnRbTTYT4w
Imv3dIdcg5SxzZAwc4QDjhtHrxtjjoi3z8oV3FdJ4f8Xq4dEiOhxBjEEj5cbdam7
6JJf0LUtDK+sKlDQ1DLTcesclS2il3RZmXSXbHiv+aISi1U47wc4mmpitELwHgOY
jkjWMx1pfIxcbOUAW1ano5o8Go7IBiC4L6P2NkLyH7p/X/5Y6gpjV+MdplHRCP+3
qbg3EGQWpYiH6RWJYRuURnR/TZFRsK+m71/DpeHFJXjuZYk8cMMjAQilRUd65UGJ
dBEInykXqQEDevYgKqrLDe/Sfl+HSwWOhunLMDmOaOXh0e/v2vH+l2VT15+JMuu+
BShlJX560uBkL9aYV2Z/pxML3Caa46ZorPjYQYrCy0ly5T53jLZiEbOSwvE+C3bI
AC+rspza+i0xQBONeFtAO4sJpYexgcO0IeUyB1BMaBM3pjYqOIEFQWta4VHJCO+4
i6o+oiSLkwsbIgDxPpPqFmdvVr3yviw1mO3K0c6i9v0OQBWPf8es4CGVNKZniHvK
yLppgkahTULA71lH5atBnvSL+yEJFnTVLnQ4kew6iam+6jGcLNIuKAouNX1uVWGa
LGWf6uFpC01e48bi8OSpuGBJziH3NCXdIKjiNjADZW/UwH7sf82SQZL00lDoJrcv
sB/YifnZwuASknVZ4YVD758sdqyRsRd7Wb/Qj6NtSCXdz82Es+84yOspMHiHV4XS
jCAzDpiKGF7DPJZD9squ9JibzzjmsarrQV11yvrzcwZo8ABWhiKd7oEBXk7uCJZ7
mmvQFQ3yGQBFKpW61wcq+2ddswJyWeU0wUGPlM+O3KSFOH+bUuRCHphZ3vqieGyt
QhXt7gNLSminrh7WeYmvpJHJbKvhZesJGLJylIevWb006UKyUCo0IxKAm+3BovwS
pVz9ilFasAT5YZhqM2hECagvzAB4B+DCD9r+QxMjQpGnBiSf3e30QcG6eLMjJ6Iz
cCqlAd0B6ifBRFn/AbTAxMxd6UlL/okp5QnfLbDcm2YPxAm1XKEoUuUKMfByPv1R
t8Fh7nZIB9jZ9IjdVUJhEBmYUglHBsA9xLHGuBdtEtzOJnSGQY75dEstVMEWjPTZ
V671G1ncWKHrZp0QZ8NuxhC0fzXtoEYRxHtzAP0ZEydnVyMCmIoQU5bvKWd8JU0f
GW1fDWRYVECDamNMqUAo62wVAwbX2HAVQxP3iBDmjMzlin09xHIQX0VEX28XbC5N
t+kO1eI2kYKV18gTGGSwDrbCj5g26e9g2Igqgi9A4HtvgUtnQA8luzByAOYEis9a
lXd9GAyK8w1QawWlz0SL1OhBzM0tlGZ67ESAwsF1pdP3VdPj/TFyOwsqnx8wd5Zg
B0Fu+aVMqP+N32kkSITzYTJSJEjiUyUHSjGa37sz3tghMsGIM5Hgw/6PnUjqgddz
RzqJ5WaJUuhIt260lFMGfCyk6Zh/HvctHLOmZ0bCc6ZiaHoWdcGfrR0CcRrT6Ry9
UyqZdrJBoZJIKe35hrCNXzhpLQik0Japi14DjAVxXPXgNbipcvwIcuk3P3pK4lKT
1XKvdB+hEH2UKto7Cv9T7nlqY6iHUeH0AAgQUJWMDbAqDWFWdGuyXo9/ET4xaSzR
v/P9ttxwAi2jtu0iQ/ztJlsGiZ3TdTWzxuFR62NyEJuP8HTdmKL87EGah6eVjihI
G3HdDvk83trKeb42FVqE51HKdbfaChavUIVBXiLBJNI=
`protect END_PROTECTED
